library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs: in std_logic_vector(1023 downto 0);
        outputs: out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs: std_logic_vector(10239 downto 0);
    signal layer1_outputs: std_logic_vector(10239 downto 0);
    signal layer2_outputs: std_logic_vector(10239 downto 0);
    signal layer3_outputs: std_logic_vector(10239 downto 0);
    signal layer4_outputs: std_logic_vector(10239 downto 0);
    signal layer5_outputs: std_logic_vector(10239 downto 0);
    signal layer6_outputs: std_logic_vector(10239 downto 0);

begin
    layer0_outputs(0) <= b;
    layer0_outputs(1) <= '0';
    layer0_outputs(2) <= a and not b;
    layer0_outputs(3) <= a xor b;
    layer0_outputs(4) <= not b or a;
    layer0_outputs(5) <= not b or a;
    layer0_outputs(6) <= not a or b;
    layer0_outputs(7) <= a and not b;
    layer0_outputs(8) <= not b;
    layer0_outputs(9) <= not b or a;
    layer0_outputs(10) <= not b or a;
    layer0_outputs(11) <= not (a xor b);
    layer0_outputs(12) <= not (a or b);
    layer0_outputs(13) <= '0';
    layer0_outputs(14) <= not b or a;
    layer0_outputs(15) <= a xor b;
    layer0_outputs(16) <= not (a xor b);
    layer0_outputs(17) <= not (a and b);
    layer0_outputs(18) <= '0';
    layer0_outputs(19) <= a or b;
    layer0_outputs(20) <= b;
    layer0_outputs(21) <= not a or b;
    layer0_outputs(22) <= a and b;
    layer0_outputs(23) <= '1';
    layer0_outputs(24) <= a or b;
    layer0_outputs(25) <= b and not a;
    layer0_outputs(26) <= b;
    layer0_outputs(27) <= not (a or b);
    layer0_outputs(28) <= not b;
    layer0_outputs(29) <= not a;
    layer0_outputs(30) <= a or b;
    layer0_outputs(31) <= b;
    layer0_outputs(32) <= b;
    layer0_outputs(33) <= not b;
    layer0_outputs(34) <= not (a and b);
    layer0_outputs(35) <= '0';
    layer0_outputs(36) <= not b or a;
    layer0_outputs(37) <= b;
    layer0_outputs(38) <= not b;
    layer0_outputs(39) <= '0';
    layer0_outputs(40) <= not b or a;
    layer0_outputs(41) <= '0';
    layer0_outputs(42) <= b and not a;
    layer0_outputs(43) <= '0';
    layer0_outputs(44) <= not (a or b);
    layer0_outputs(45) <= not (a and b);
    layer0_outputs(46) <= a and not b;
    layer0_outputs(47) <= a and b;
    layer0_outputs(48) <= a and not b;
    layer0_outputs(49) <= a and b;
    layer0_outputs(50) <= a;
    layer0_outputs(51) <= a;
    layer0_outputs(52) <= a or b;
    layer0_outputs(53) <= not (a and b);
    layer0_outputs(54) <= a and not b;
    layer0_outputs(55) <= not a;
    layer0_outputs(56) <= b;
    layer0_outputs(57) <= a;
    layer0_outputs(58) <= '0';
    layer0_outputs(59) <= '1';
    layer0_outputs(60) <= a xor b;
    layer0_outputs(61) <= a or b;
    layer0_outputs(62) <= not b or a;
    layer0_outputs(63) <= not a;
    layer0_outputs(64) <= b and not a;
    layer0_outputs(65) <= b and not a;
    layer0_outputs(66) <= a or b;
    layer0_outputs(67) <= a and not b;
    layer0_outputs(68) <= b and not a;
    layer0_outputs(69) <= not (a xor b);
    layer0_outputs(70) <= not b;
    layer0_outputs(71) <= a xor b;
    layer0_outputs(72) <= not b;
    layer0_outputs(73) <= a or b;
    layer0_outputs(74) <= not a or b;
    layer0_outputs(75) <= a and b;
    layer0_outputs(76) <= not (a or b);
    layer0_outputs(77) <= b and not a;
    layer0_outputs(78) <= not (a xor b);
    layer0_outputs(79) <= not a or b;
    layer0_outputs(80) <= a or b;
    layer0_outputs(81) <= not b;
    layer0_outputs(82) <= not (a and b);
    layer0_outputs(83) <= a and not b;
    layer0_outputs(84) <= a and not b;
    layer0_outputs(85) <= a and not b;
    layer0_outputs(86) <= not a or b;
    layer0_outputs(87) <= a and b;
    layer0_outputs(88) <= a or b;
    layer0_outputs(89) <= not (a or b);
    layer0_outputs(90) <= a or b;
    layer0_outputs(91) <= a and b;
    layer0_outputs(92) <= not (a and b);
    layer0_outputs(93) <= a or b;
    layer0_outputs(94) <= not a;
    layer0_outputs(95) <= not a;
    layer0_outputs(96) <= a and b;
    layer0_outputs(97) <= b;
    layer0_outputs(98) <= not a;
    layer0_outputs(99) <= '0';
    layer0_outputs(100) <= not (a xor b);
    layer0_outputs(101) <= b;
    layer0_outputs(102) <= a or b;
    layer0_outputs(103) <= not b;
    layer0_outputs(104) <= not a or b;
    layer0_outputs(105) <= '0';
    layer0_outputs(106) <= not (a and b);
    layer0_outputs(107) <= not (a or b);
    layer0_outputs(108) <= a and not b;
    layer0_outputs(109) <= a and b;
    layer0_outputs(110) <= not b or a;
    layer0_outputs(111) <= a;
    layer0_outputs(112) <= not (a or b);
    layer0_outputs(113) <= b;
    layer0_outputs(114) <= a;
    layer0_outputs(115) <= not a or b;
    layer0_outputs(116) <= not (a and b);
    layer0_outputs(117) <= not b or a;
    layer0_outputs(118) <= a;
    layer0_outputs(119) <= not (a xor b);
    layer0_outputs(120) <= a or b;
    layer0_outputs(121) <= a and b;
    layer0_outputs(122) <= not (a or b);
    layer0_outputs(123) <= not a;
    layer0_outputs(124) <= a and b;
    layer0_outputs(125) <= not a or b;
    layer0_outputs(126) <= not b;
    layer0_outputs(127) <= b;
    layer0_outputs(128) <= a and not b;
    layer0_outputs(129) <= not b or a;
    layer0_outputs(130) <= a or b;
    layer0_outputs(131) <= '1';
    layer0_outputs(132) <= a xor b;
    layer0_outputs(133) <= a and not b;
    layer0_outputs(134) <= a and b;
    layer0_outputs(135) <= b;
    layer0_outputs(136) <= not a;
    layer0_outputs(137) <= not (a xor b);
    layer0_outputs(138) <= b;
    layer0_outputs(139) <= not (a or b);
    layer0_outputs(140) <= not (a or b);
    layer0_outputs(141) <= a and b;
    layer0_outputs(142) <= a xor b;
    layer0_outputs(143) <= not a;
    layer0_outputs(144) <= a;
    layer0_outputs(145) <= a or b;
    layer0_outputs(146) <= not (a xor b);
    layer0_outputs(147) <= a or b;
    layer0_outputs(148) <= not b;
    layer0_outputs(149) <= a or b;
    layer0_outputs(150) <= a and b;
    layer0_outputs(151) <= a and not b;
    layer0_outputs(152) <= not b;
    layer0_outputs(153) <= b and not a;
    layer0_outputs(154) <= '0';
    layer0_outputs(155) <= b;
    layer0_outputs(156) <= a and b;
    layer0_outputs(157) <= not a;
    layer0_outputs(158) <= not a or b;
    layer0_outputs(159) <= not b;
    layer0_outputs(160) <= not a or b;
    layer0_outputs(161) <= not a;
    layer0_outputs(162) <= a;
    layer0_outputs(163) <= '0';
    layer0_outputs(164) <= not (a xor b);
    layer0_outputs(165) <= b;
    layer0_outputs(166) <= a;
    layer0_outputs(167) <= not (a or b);
    layer0_outputs(168) <= a and not b;
    layer0_outputs(169) <= a;
    layer0_outputs(170) <= a and not b;
    layer0_outputs(171) <= not (a or b);
    layer0_outputs(172) <= not a;
    layer0_outputs(173) <= '1';
    layer0_outputs(174) <= a;
    layer0_outputs(175) <= a;
    layer0_outputs(176) <= not (a and b);
    layer0_outputs(177) <= a;
    layer0_outputs(178) <= b;
    layer0_outputs(179) <= not a;
    layer0_outputs(180) <= a xor b;
    layer0_outputs(181) <= not b or a;
    layer0_outputs(182) <= not (a or b);
    layer0_outputs(183) <= a and not b;
    layer0_outputs(184) <= '0';
    layer0_outputs(185) <= not b;
    layer0_outputs(186) <= a;
    layer0_outputs(187) <= not b;
    layer0_outputs(188) <= not (a xor b);
    layer0_outputs(189) <= b and not a;
    layer0_outputs(190) <= not b;
    layer0_outputs(191) <= a or b;
    layer0_outputs(192) <= a or b;
    layer0_outputs(193) <= not (a and b);
    layer0_outputs(194) <= a xor b;
    layer0_outputs(195) <= b and not a;
    layer0_outputs(196) <= a xor b;
    layer0_outputs(197) <= not (a or b);
    layer0_outputs(198) <= not (a or b);
    layer0_outputs(199) <= a;
    layer0_outputs(200) <= not a;
    layer0_outputs(201) <= not b or a;
    layer0_outputs(202) <= not b;
    layer0_outputs(203) <= not a or b;
    layer0_outputs(204) <= b;
    layer0_outputs(205) <= b and not a;
    layer0_outputs(206) <= b and not a;
    layer0_outputs(207) <= not (a or b);
    layer0_outputs(208) <= not a or b;
    layer0_outputs(209) <= a xor b;
    layer0_outputs(210) <= not (a or b);
    layer0_outputs(211) <= not a;
    layer0_outputs(212) <= '0';
    layer0_outputs(213) <= a and b;
    layer0_outputs(214) <= not (a or b);
    layer0_outputs(215) <= a or b;
    layer0_outputs(216) <= a and not b;
    layer0_outputs(217) <= '0';
    layer0_outputs(218) <= a xor b;
    layer0_outputs(219) <= not a;
    layer0_outputs(220) <= not a or b;
    layer0_outputs(221) <= a or b;
    layer0_outputs(222) <= not a or b;
    layer0_outputs(223) <= a and not b;
    layer0_outputs(224) <= a or b;
    layer0_outputs(225) <= not a or b;
    layer0_outputs(226) <= a;
    layer0_outputs(227) <= not a or b;
    layer0_outputs(228) <= not (a xor b);
    layer0_outputs(229) <= not (a or b);
    layer0_outputs(230) <= '1';
    layer0_outputs(231) <= a;
    layer0_outputs(232) <= '1';
    layer0_outputs(233) <= '0';
    layer0_outputs(234) <= not (a and b);
    layer0_outputs(235) <= b;
    layer0_outputs(236) <= a or b;
    layer0_outputs(237) <= a;
    layer0_outputs(238) <= not (a or b);
    layer0_outputs(239) <= '0';
    layer0_outputs(240) <= not (a or b);
    layer0_outputs(241) <= a;
    layer0_outputs(242) <= not b;
    layer0_outputs(243) <= not b or a;
    layer0_outputs(244) <= b;
    layer0_outputs(245) <= '1';
    layer0_outputs(246) <= not b;
    layer0_outputs(247) <= '1';
    layer0_outputs(248) <= '0';
    layer0_outputs(249) <= a and not b;
    layer0_outputs(250) <= not b;
    layer0_outputs(251) <= b;
    layer0_outputs(252) <= b and not a;
    layer0_outputs(253) <= '1';
    layer0_outputs(254) <= not a or b;
    layer0_outputs(255) <= not b;
    layer0_outputs(256) <= b;
    layer0_outputs(257) <= a and not b;
    layer0_outputs(258) <= not a or b;
    layer0_outputs(259) <= a or b;
    layer0_outputs(260) <= not b;
    layer0_outputs(261) <= a xor b;
    layer0_outputs(262) <= a and not b;
    layer0_outputs(263) <= not b or a;
    layer0_outputs(264) <= not (a or b);
    layer0_outputs(265) <= not b;
    layer0_outputs(266) <= a;
    layer0_outputs(267) <= not a or b;
    layer0_outputs(268) <= '1';
    layer0_outputs(269) <= b;
    layer0_outputs(270) <= not a or b;
    layer0_outputs(271) <= b and not a;
    layer0_outputs(272) <= not a or b;
    layer0_outputs(273) <= b and not a;
    layer0_outputs(274) <= a or b;
    layer0_outputs(275) <= not b;
    layer0_outputs(276) <= a and not b;
    layer0_outputs(277) <= a and not b;
    layer0_outputs(278) <= not b;
    layer0_outputs(279) <= not a;
    layer0_outputs(280) <= not (a xor b);
    layer0_outputs(281) <= a;
    layer0_outputs(282) <= a or b;
    layer0_outputs(283) <= b;
    layer0_outputs(284) <= not b or a;
    layer0_outputs(285) <= a or b;
    layer0_outputs(286) <= not a;
    layer0_outputs(287) <= '0';
    layer0_outputs(288) <= not b;
    layer0_outputs(289) <= '0';
    layer0_outputs(290) <= not a or b;
    layer0_outputs(291) <= b;
    layer0_outputs(292) <= '1';
    layer0_outputs(293) <= not (a xor b);
    layer0_outputs(294) <= a;
    layer0_outputs(295) <= not b;
    layer0_outputs(296) <= not b;
    layer0_outputs(297) <= b and not a;
    layer0_outputs(298) <= not (a or b);
    layer0_outputs(299) <= not (a or b);
    layer0_outputs(300) <= not b;
    layer0_outputs(301) <= not a or b;
    layer0_outputs(302) <= a and not b;
    layer0_outputs(303) <= not a or b;
    layer0_outputs(304) <= a;
    layer0_outputs(305) <= a xor b;
    layer0_outputs(306) <= not a or b;
    layer0_outputs(307) <= b and not a;
    layer0_outputs(308) <= not a;
    layer0_outputs(309) <= not b;
    layer0_outputs(310) <= not b;
    layer0_outputs(311) <= not (a and b);
    layer0_outputs(312) <= not (a xor b);
    layer0_outputs(313) <= not b;
    layer0_outputs(314) <= b;
    layer0_outputs(315) <= a xor b;
    layer0_outputs(316) <= b;
    layer0_outputs(317) <= not (a or b);
    layer0_outputs(318) <= '0';
    layer0_outputs(319) <= a xor b;
    layer0_outputs(320) <= a or b;
    layer0_outputs(321) <= not a;
    layer0_outputs(322) <= '0';
    layer0_outputs(323) <= not (a or b);
    layer0_outputs(324) <= a;
    layer0_outputs(325) <= a;
    layer0_outputs(326) <= not (a or b);
    layer0_outputs(327) <= not (a xor b);
    layer0_outputs(328) <= not b;
    layer0_outputs(329) <= not b or a;
    layer0_outputs(330) <= a xor b;
    layer0_outputs(331) <= a or b;
    layer0_outputs(332) <= b;
    layer0_outputs(333) <= not b;
    layer0_outputs(334) <= not (a or b);
    layer0_outputs(335) <= not b or a;
    layer0_outputs(336) <= not (a and b);
    layer0_outputs(337) <= '1';
    layer0_outputs(338) <= not (a or b);
    layer0_outputs(339) <= not b or a;
    layer0_outputs(340) <= not (a xor b);
    layer0_outputs(341) <= a and b;
    layer0_outputs(342) <= not (a xor b);
    layer0_outputs(343) <= a or b;
    layer0_outputs(344) <= not b or a;
    layer0_outputs(345) <= not b or a;
    layer0_outputs(346) <= b;
    layer0_outputs(347) <= not a or b;
    layer0_outputs(348) <= not (a xor b);
    layer0_outputs(349) <= a or b;
    layer0_outputs(350) <= a and b;
    layer0_outputs(351) <= not (a or b);
    layer0_outputs(352) <= '0';
    layer0_outputs(353) <= a xor b;
    layer0_outputs(354) <= '1';
    layer0_outputs(355) <= a;
    layer0_outputs(356) <= not b;
    layer0_outputs(357) <= not (a or b);
    layer0_outputs(358) <= not a or b;
    layer0_outputs(359) <= a or b;
    layer0_outputs(360) <= not (a and b);
    layer0_outputs(361) <= not (a and b);
    layer0_outputs(362) <= b and not a;
    layer0_outputs(363) <= not b;
    layer0_outputs(364) <= a;
    layer0_outputs(365) <= '0';
    layer0_outputs(366) <= not (a and b);
    layer0_outputs(367) <= '0';
    layer0_outputs(368) <= a and b;
    layer0_outputs(369) <= not b;
    layer0_outputs(370) <= b;
    layer0_outputs(371) <= not (a or b);
    layer0_outputs(372) <= not (a xor b);
    layer0_outputs(373) <= not (a xor b);
    layer0_outputs(374) <= not (a or b);
    layer0_outputs(375) <= '0';
    layer0_outputs(376) <= a and not b;
    layer0_outputs(377) <= not a;
    layer0_outputs(378) <= not (a and b);
    layer0_outputs(379) <= a or b;
    layer0_outputs(380) <= a xor b;
    layer0_outputs(381) <= not (a and b);
    layer0_outputs(382) <= a;
    layer0_outputs(383) <= not b or a;
    layer0_outputs(384) <= not b;
    layer0_outputs(385) <= a;
    layer0_outputs(386) <= not (a or b);
    layer0_outputs(387) <= not a;
    layer0_outputs(388) <= not (a and b);
    layer0_outputs(389) <= not (a or b);
    layer0_outputs(390) <= a xor b;
    layer0_outputs(391) <= not (a or b);
    layer0_outputs(392) <= b and not a;
    layer0_outputs(393) <= b and not a;
    layer0_outputs(394) <= not b;
    layer0_outputs(395) <= not (a xor b);
    layer0_outputs(396) <= not (a and b);
    layer0_outputs(397) <= a and b;
    layer0_outputs(398) <= '1';
    layer0_outputs(399) <= not a or b;
    layer0_outputs(400) <= not b or a;
    layer0_outputs(401) <= a and b;
    layer0_outputs(402) <= a xor b;
    layer0_outputs(403) <= a;
    layer0_outputs(404) <= not b or a;
    layer0_outputs(405) <= not (a xor b);
    layer0_outputs(406) <= b and not a;
    layer0_outputs(407) <= b;
    layer0_outputs(408) <= not a;
    layer0_outputs(409) <= b and not a;
    layer0_outputs(410) <= a and b;
    layer0_outputs(411) <= not a or b;
    layer0_outputs(412) <= not b or a;
    layer0_outputs(413) <= a xor b;
    layer0_outputs(414) <= a and not b;
    layer0_outputs(415) <= '1';
    layer0_outputs(416) <= a or b;
    layer0_outputs(417) <= a and not b;
    layer0_outputs(418) <= not a;
    layer0_outputs(419) <= a and b;
    layer0_outputs(420) <= a xor b;
    layer0_outputs(421) <= not (a or b);
    layer0_outputs(422) <= '1';
    layer0_outputs(423) <= not (a or b);
    layer0_outputs(424) <= not a;
    layer0_outputs(425) <= b;
    layer0_outputs(426) <= a and b;
    layer0_outputs(427) <= not a or b;
    layer0_outputs(428) <= not (a or b);
    layer0_outputs(429) <= not a;
    layer0_outputs(430) <= not b or a;
    layer0_outputs(431) <= not (a or b);
    layer0_outputs(432) <= not b;
    layer0_outputs(433) <= not a;
    layer0_outputs(434) <= not (a xor b);
    layer0_outputs(435) <= b;
    layer0_outputs(436) <= a and b;
    layer0_outputs(437) <= a and not b;
    layer0_outputs(438) <= b;
    layer0_outputs(439) <= not b or a;
    layer0_outputs(440) <= not (a or b);
    layer0_outputs(441) <= b;
    layer0_outputs(442) <= not b;
    layer0_outputs(443) <= not a or b;
    layer0_outputs(444) <= a;
    layer0_outputs(445) <= a xor b;
    layer0_outputs(446) <= not a;
    layer0_outputs(447) <= b;
    layer0_outputs(448) <= not a;
    layer0_outputs(449) <= not (a or b);
    layer0_outputs(450) <= a and not b;
    layer0_outputs(451) <= b;
    layer0_outputs(452) <= not (a and b);
    layer0_outputs(453) <= '1';
    layer0_outputs(454) <= not (a or b);
    layer0_outputs(455) <= not (a or b);
    layer0_outputs(456) <= b and not a;
    layer0_outputs(457) <= b;
    layer0_outputs(458) <= a and b;
    layer0_outputs(459) <= b and not a;
    layer0_outputs(460) <= not (a and b);
    layer0_outputs(461) <= not (a or b);
    layer0_outputs(462) <= a;
    layer0_outputs(463) <= b;
    layer0_outputs(464) <= a and b;
    layer0_outputs(465) <= a and b;
    layer0_outputs(466) <= not a or b;
    layer0_outputs(467) <= a xor b;
    layer0_outputs(468) <= a and b;
    layer0_outputs(469) <= a and not b;
    layer0_outputs(470) <= b and not a;
    layer0_outputs(471) <= not a or b;
    layer0_outputs(472) <= not (a and b);
    layer0_outputs(473) <= not b;
    layer0_outputs(474) <= a;
    layer0_outputs(475) <= b;
    layer0_outputs(476) <= a;
    layer0_outputs(477) <= a;
    layer0_outputs(478) <= a xor b;
    layer0_outputs(479) <= '1';
    layer0_outputs(480) <= not a;
    layer0_outputs(481) <= a or b;
    layer0_outputs(482) <= not (a or b);
    layer0_outputs(483) <= a or b;
    layer0_outputs(484) <= not b or a;
    layer0_outputs(485) <= not a;
    layer0_outputs(486) <= a and b;
    layer0_outputs(487) <= a;
    layer0_outputs(488) <= b;
    layer0_outputs(489) <= '0';
    layer0_outputs(490) <= '1';
    layer0_outputs(491) <= not b or a;
    layer0_outputs(492) <= not a;
    layer0_outputs(493) <= not a;
    layer0_outputs(494) <= not (a or b);
    layer0_outputs(495) <= b and not a;
    layer0_outputs(496) <= b;
    layer0_outputs(497) <= not b or a;
    layer0_outputs(498) <= b;
    layer0_outputs(499) <= a;
    layer0_outputs(500) <= not a;
    layer0_outputs(501) <= '0';
    layer0_outputs(502) <= not a;
    layer0_outputs(503) <= not (a xor b);
    layer0_outputs(504) <= not a or b;
    layer0_outputs(505) <= a or b;
    layer0_outputs(506) <= not (a or b);
    layer0_outputs(507) <= not b or a;
    layer0_outputs(508) <= not a or b;
    layer0_outputs(509) <= '0';
    layer0_outputs(510) <= '0';
    layer0_outputs(511) <= a and not b;
    layer0_outputs(512) <= a;
    layer0_outputs(513) <= '0';
    layer0_outputs(514) <= '0';
    layer0_outputs(515) <= not (a or b);
    layer0_outputs(516) <= not (a or b);
    layer0_outputs(517) <= not (a or b);
    layer0_outputs(518) <= not a;
    layer0_outputs(519) <= a and b;
    layer0_outputs(520) <= b;
    layer0_outputs(521) <= '0';
    layer0_outputs(522) <= b;
    layer0_outputs(523) <= a or b;
    layer0_outputs(524) <= b;
    layer0_outputs(525) <= b;
    layer0_outputs(526) <= a or b;
    layer0_outputs(527) <= not a or b;
    layer0_outputs(528) <= a or b;
    layer0_outputs(529) <= b;
    layer0_outputs(530) <= a and b;
    layer0_outputs(531) <= '0';
    layer0_outputs(532) <= a;
    layer0_outputs(533) <= not (a or b);
    layer0_outputs(534) <= a;
    layer0_outputs(535) <= not (a or b);
    layer0_outputs(536) <= b;
    layer0_outputs(537) <= a;
    layer0_outputs(538) <= a or b;
    layer0_outputs(539) <= a and b;
    layer0_outputs(540) <= a xor b;
    layer0_outputs(541) <= '0';
    layer0_outputs(542) <= '1';
    layer0_outputs(543) <= '0';
    layer0_outputs(544) <= a or b;
    layer0_outputs(545) <= not a;
    layer0_outputs(546) <= a and b;
    layer0_outputs(547) <= '0';
    layer0_outputs(548) <= b and not a;
    layer0_outputs(549) <= b and not a;
    layer0_outputs(550) <= a xor b;
    layer0_outputs(551) <= b and not a;
    layer0_outputs(552) <= '0';
    layer0_outputs(553) <= not (a and b);
    layer0_outputs(554) <= not a or b;
    layer0_outputs(555) <= not a or b;
    layer0_outputs(556) <= a xor b;
    layer0_outputs(557) <= a;
    layer0_outputs(558) <= not b or a;
    layer0_outputs(559) <= '0';
    layer0_outputs(560) <= not (a or b);
    layer0_outputs(561) <= not a;
    layer0_outputs(562) <= not a or b;
    layer0_outputs(563) <= a;
    layer0_outputs(564) <= b and not a;
    layer0_outputs(565) <= '1';
    layer0_outputs(566) <= not b;
    layer0_outputs(567) <= a or b;
    layer0_outputs(568) <= not (a or b);
    layer0_outputs(569) <= a;
    layer0_outputs(570) <= not b;
    layer0_outputs(571) <= not (a and b);
    layer0_outputs(572) <= not b or a;
    layer0_outputs(573) <= a and not b;
    layer0_outputs(574) <= a;
    layer0_outputs(575) <= '1';
    layer0_outputs(576) <= a or b;
    layer0_outputs(577) <= b;
    layer0_outputs(578) <= a or b;
    layer0_outputs(579) <= not b or a;
    layer0_outputs(580) <= not (a and b);
    layer0_outputs(581) <= '0';
    layer0_outputs(582) <= not b or a;
    layer0_outputs(583) <= a;
    layer0_outputs(584) <= a or b;
    layer0_outputs(585) <= b and not a;
    layer0_outputs(586) <= '1';
    layer0_outputs(587) <= not b;
    layer0_outputs(588) <= '0';
    layer0_outputs(589) <= a and not b;
    layer0_outputs(590) <= a xor b;
    layer0_outputs(591) <= a xor b;
    layer0_outputs(592) <= '0';
    layer0_outputs(593) <= not b;
    layer0_outputs(594) <= a and b;
    layer0_outputs(595) <= a or b;
    layer0_outputs(596) <= not (a xor b);
    layer0_outputs(597) <= a or b;
    layer0_outputs(598) <= a or b;
    layer0_outputs(599) <= not (a or b);
    layer0_outputs(600) <= a and not b;
    layer0_outputs(601) <= b and not a;
    layer0_outputs(602) <= a and not b;
    layer0_outputs(603) <= not a or b;
    layer0_outputs(604) <= a and b;
    layer0_outputs(605) <= not (a xor b);
    layer0_outputs(606) <= a;
    layer0_outputs(607) <= not a;
    layer0_outputs(608) <= '0';
    layer0_outputs(609) <= not (a and b);
    layer0_outputs(610) <= not a or b;
    layer0_outputs(611) <= a and b;
    layer0_outputs(612) <= b;
    layer0_outputs(613) <= a xor b;
    layer0_outputs(614) <= '0';
    layer0_outputs(615) <= not a or b;
    layer0_outputs(616) <= not a or b;
    layer0_outputs(617) <= '1';
    layer0_outputs(618) <= a or b;
    layer0_outputs(619) <= not b or a;
    layer0_outputs(620) <= b and not a;
    layer0_outputs(621) <= not b or a;
    layer0_outputs(622) <= '1';
    layer0_outputs(623) <= not a;
    layer0_outputs(624) <= a;
    layer0_outputs(625) <= a;
    layer0_outputs(626) <= a and b;
    layer0_outputs(627) <= not (a or b);
    layer0_outputs(628) <= not (a or b);
    layer0_outputs(629) <= a and not b;
    layer0_outputs(630) <= a or b;
    layer0_outputs(631) <= b;
    layer0_outputs(632) <= not (a xor b);
    layer0_outputs(633) <= a and b;
    layer0_outputs(634) <= not a or b;
    layer0_outputs(635) <= a and not b;
    layer0_outputs(636) <= not (a and b);
    layer0_outputs(637) <= a;
    layer0_outputs(638) <= not b;
    layer0_outputs(639) <= not (a and b);
    layer0_outputs(640) <= a;
    layer0_outputs(641) <= a and not b;
    layer0_outputs(642) <= b;
    layer0_outputs(643) <= not (a xor b);
    layer0_outputs(644) <= b and not a;
    layer0_outputs(645) <= not (a and b);
    layer0_outputs(646) <= not (a xor b);
    layer0_outputs(647) <= not a or b;
    layer0_outputs(648) <= not (a or b);
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= not a or b;
    layer0_outputs(651) <= b and not a;
    layer0_outputs(652) <= b;
    layer0_outputs(653) <= a and not b;
    layer0_outputs(654) <= not b;
    layer0_outputs(655) <= b and not a;
    layer0_outputs(656) <= not b or a;
    layer0_outputs(657) <= a and b;
    layer0_outputs(658) <= not (a and b);
    layer0_outputs(659) <= a;
    layer0_outputs(660) <= not a or b;
    layer0_outputs(661) <= not a;
    layer0_outputs(662) <= a and b;
    layer0_outputs(663) <= not (a or b);
    layer0_outputs(664) <= a;
    layer0_outputs(665) <= not a or b;
    layer0_outputs(666) <= not (a or b);
    layer0_outputs(667) <= not (a xor b);
    layer0_outputs(668) <= a and not b;
    layer0_outputs(669) <= b;
    layer0_outputs(670) <= '1';
    layer0_outputs(671) <= not b;
    layer0_outputs(672) <= a xor b;
    layer0_outputs(673) <= not (a or b);
    layer0_outputs(674) <= not (a or b);
    layer0_outputs(675) <= a;
    layer0_outputs(676) <= b;
    layer0_outputs(677) <= a and not b;
    layer0_outputs(678) <= not (a or b);
    layer0_outputs(679) <= a xor b;
    layer0_outputs(680) <= a xor b;
    layer0_outputs(681) <= not a;
    layer0_outputs(682) <= a and b;
    layer0_outputs(683) <= '1';
    layer0_outputs(684) <= a xor b;
    layer0_outputs(685) <= not (a xor b);
    layer0_outputs(686) <= a or b;
    layer0_outputs(687) <= '0';
    layer0_outputs(688) <= '0';
    layer0_outputs(689) <= not b;
    layer0_outputs(690) <= a or b;
    layer0_outputs(691) <= '1';
    layer0_outputs(692) <= b and not a;
    layer0_outputs(693) <= b;
    layer0_outputs(694) <= a or b;
    layer0_outputs(695) <= a and not b;
    layer0_outputs(696) <= not (a xor b);
    layer0_outputs(697) <= not b or a;
    layer0_outputs(698) <= b;
    layer0_outputs(699) <= b;
    layer0_outputs(700) <= a xor b;
    layer0_outputs(701) <= not b;
    layer0_outputs(702) <= not a or b;
    layer0_outputs(703) <= b;
    layer0_outputs(704) <= b;
    layer0_outputs(705) <= not a or b;
    layer0_outputs(706) <= not a;
    layer0_outputs(707) <= b and not a;
    layer0_outputs(708) <= not a or b;
    layer0_outputs(709) <= '1';
    layer0_outputs(710) <= b and not a;
    layer0_outputs(711) <= a or b;
    layer0_outputs(712) <= not (a or b);
    layer0_outputs(713) <= a xor b;
    layer0_outputs(714) <= a;
    layer0_outputs(715) <= a xor b;
    layer0_outputs(716) <= not b or a;
    layer0_outputs(717) <= not b;
    layer0_outputs(718) <= not a;
    layer0_outputs(719) <= not (a and b);
    layer0_outputs(720) <= a or b;
    layer0_outputs(721) <= not a;
    layer0_outputs(722) <= a and not b;
    layer0_outputs(723) <= a or b;
    layer0_outputs(724) <= not b or a;
    layer0_outputs(725) <= '1';
    layer0_outputs(726) <= not b or a;
    layer0_outputs(727) <= a or b;
    layer0_outputs(728) <= not (a or b);
    layer0_outputs(729) <= not (a and b);
    layer0_outputs(730) <= not a or b;
    layer0_outputs(731) <= not (a or b);
    layer0_outputs(732) <= not (a and b);
    layer0_outputs(733) <= not b;
    layer0_outputs(734) <= not (a xor b);
    layer0_outputs(735) <= a or b;
    layer0_outputs(736) <= a xor b;
    layer0_outputs(737) <= b;
    layer0_outputs(738) <= a;
    layer0_outputs(739) <= a and b;
    layer0_outputs(740) <= '0';
    layer0_outputs(741) <= a;
    layer0_outputs(742) <= a and not b;
    layer0_outputs(743) <= a or b;
    layer0_outputs(744) <= not a or b;
    layer0_outputs(745) <= a;
    layer0_outputs(746) <= a xor b;
    layer0_outputs(747) <= not a;
    layer0_outputs(748) <= not a or b;
    layer0_outputs(749) <= a;
    layer0_outputs(750) <= not (a xor b);
    layer0_outputs(751) <= a xor b;
    layer0_outputs(752) <= not b;
    layer0_outputs(753) <= a or b;
    layer0_outputs(754) <= a and b;
    layer0_outputs(755) <= '1';
    layer0_outputs(756) <= not b or a;
    layer0_outputs(757) <= '1';
    layer0_outputs(758) <= a or b;
    layer0_outputs(759) <= not (a or b);
    layer0_outputs(760) <= not b;
    layer0_outputs(761) <= '1';
    layer0_outputs(762) <= b;
    layer0_outputs(763) <= not (a or b);
    layer0_outputs(764) <= b;
    layer0_outputs(765) <= '0';
    layer0_outputs(766) <= a xor b;
    layer0_outputs(767) <= not (a xor b);
    layer0_outputs(768) <= a or b;
    layer0_outputs(769) <= not b or a;
    layer0_outputs(770) <= not (a or b);
    layer0_outputs(771) <= not (a xor b);
    layer0_outputs(772) <= b and not a;
    layer0_outputs(773) <= not b or a;
    layer0_outputs(774) <= b;
    layer0_outputs(775) <= a xor b;
    layer0_outputs(776) <= not (a and b);
    layer0_outputs(777) <= b and not a;
    layer0_outputs(778) <= '1';
    layer0_outputs(779) <= not (a and b);
    layer0_outputs(780) <= not (a or b);
    layer0_outputs(781) <= b;
    layer0_outputs(782) <= '0';
    layer0_outputs(783) <= not b;
    layer0_outputs(784) <= a and not b;
    layer0_outputs(785) <= a and b;
    layer0_outputs(786) <= '1';
    layer0_outputs(787) <= a;
    layer0_outputs(788) <= not b;
    layer0_outputs(789) <= not (a xor b);
    layer0_outputs(790) <= not b;
    layer0_outputs(791) <= b;
    layer0_outputs(792) <= not (a xor b);
    layer0_outputs(793) <= a or b;
    layer0_outputs(794) <= b and not a;
    layer0_outputs(795) <= a or b;
    layer0_outputs(796) <= not (a or b);
    layer0_outputs(797) <= not (a and b);
    layer0_outputs(798) <= not a;
    layer0_outputs(799) <= b and not a;
    layer0_outputs(800) <= '0';
    layer0_outputs(801) <= not (a xor b);
    layer0_outputs(802) <= not (a or b);
    layer0_outputs(803) <= not (a xor b);
    layer0_outputs(804) <= not (a xor b);
    layer0_outputs(805) <= a and not b;
    layer0_outputs(806) <= a or b;
    layer0_outputs(807) <= a;
    layer0_outputs(808) <= b and not a;
    layer0_outputs(809) <= a or b;
    layer0_outputs(810) <= not (a xor b);
    layer0_outputs(811) <= a and b;
    layer0_outputs(812) <= not a or b;
    layer0_outputs(813) <= not (a xor b);
    layer0_outputs(814) <= a;
    layer0_outputs(815) <= not b;
    layer0_outputs(816) <= not b or a;
    layer0_outputs(817) <= b and not a;
    layer0_outputs(818) <= not a or b;
    layer0_outputs(819) <= not (a or b);
    layer0_outputs(820) <= a and not b;
    layer0_outputs(821) <= not b;
    layer0_outputs(822) <= a or b;
    layer0_outputs(823) <= not (a xor b);
    layer0_outputs(824) <= a;
    layer0_outputs(825) <= a or b;
    layer0_outputs(826) <= a or b;
    layer0_outputs(827) <= '0';
    layer0_outputs(828) <= a or b;
    layer0_outputs(829) <= not (a or b);
    layer0_outputs(830) <= not (a xor b);
    layer0_outputs(831) <= b;
    layer0_outputs(832) <= a or b;
    layer0_outputs(833) <= '0';
    layer0_outputs(834) <= a or b;
    layer0_outputs(835) <= not (a xor b);
    layer0_outputs(836) <= not b;
    layer0_outputs(837) <= a;
    layer0_outputs(838) <= not b;
    layer0_outputs(839) <= b;
    layer0_outputs(840) <= not a;
    layer0_outputs(841) <= b and not a;
    layer0_outputs(842) <= not (a or b);
    layer0_outputs(843) <= a or b;
    layer0_outputs(844) <= a xor b;
    layer0_outputs(845) <= a and not b;
    layer0_outputs(846) <= a and b;
    layer0_outputs(847) <= a and not b;
    layer0_outputs(848) <= a or b;
    layer0_outputs(849) <= '0';
    layer0_outputs(850) <= a and not b;
    layer0_outputs(851) <= a;
    layer0_outputs(852) <= not b;
    layer0_outputs(853) <= '0';
    layer0_outputs(854) <= not b or a;
    layer0_outputs(855) <= b and not a;
    layer0_outputs(856) <= '0';
    layer0_outputs(857) <= b;
    layer0_outputs(858) <= not a or b;
    layer0_outputs(859) <= not (a xor b);
    layer0_outputs(860) <= not b or a;
    layer0_outputs(861) <= a or b;
    layer0_outputs(862) <= a and b;
    layer0_outputs(863) <= b;
    layer0_outputs(864) <= not (a or b);
    layer0_outputs(865) <= a xor b;
    layer0_outputs(866) <= not (a xor b);
    layer0_outputs(867) <= not (a and b);
    layer0_outputs(868) <= b;
    layer0_outputs(869) <= a or b;
    layer0_outputs(870) <= not a;
    layer0_outputs(871) <= not b or a;
    layer0_outputs(872) <= not b or a;
    layer0_outputs(873) <= not a;
    layer0_outputs(874) <= not (a xor b);
    layer0_outputs(875) <= not a;
    layer0_outputs(876) <= a xor b;
    layer0_outputs(877) <= not (a and b);
    layer0_outputs(878) <= a;
    layer0_outputs(879) <= not a or b;
    layer0_outputs(880) <= not b or a;
    layer0_outputs(881) <= b;
    layer0_outputs(882) <= a;
    layer0_outputs(883) <= a;
    layer0_outputs(884) <= a and not b;
    layer0_outputs(885) <= b and not a;
    layer0_outputs(886) <= not (a xor b);
    layer0_outputs(887) <= not a;
    layer0_outputs(888) <= '0';
    layer0_outputs(889) <= a;
    layer0_outputs(890) <= not (a xor b);
    layer0_outputs(891) <= a or b;
    layer0_outputs(892) <= not a or b;
    layer0_outputs(893) <= a or b;
    layer0_outputs(894) <= '0';
    layer0_outputs(895) <= not b;
    layer0_outputs(896) <= not (a and b);
    layer0_outputs(897) <= a and not b;
    layer0_outputs(898) <= '0';
    layer0_outputs(899) <= not (a and b);
    layer0_outputs(900) <= '0';
    layer0_outputs(901) <= b and not a;
    layer0_outputs(902) <= a or b;
    layer0_outputs(903) <= a or b;
    layer0_outputs(904) <= a or b;
    layer0_outputs(905) <= not (a xor b);
    layer0_outputs(906) <= not a;
    layer0_outputs(907) <= not (a and b);
    layer0_outputs(908) <= a and not b;
    layer0_outputs(909) <= not b;
    layer0_outputs(910) <= b and not a;
    layer0_outputs(911) <= a and not b;
    layer0_outputs(912) <= not a or b;
    layer0_outputs(913) <= not (a and b);
    layer0_outputs(914) <= not (a or b);
    layer0_outputs(915) <= not b;
    layer0_outputs(916) <= not a;
    layer0_outputs(917) <= b and not a;
    layer0_outputs(918) <= '0';
    layer0_outputs(919) <= a and b;
    layer0_outputs(920) <= not b or a;
    layer0_outputs(921) <= a xor b;
    layer0_outputs(922) <= a and b;
    layer0_outputs(923) <= a or b;
    layer0_outputs(924) <= not (a and b);
    layer0_outputs(925) <= not (a or b);
    layer0_outputs(926) <= not a;
    layer0_outputs(927) <= not (a and b);
    layer0_outputs(928) <= not a;
    layer0_outputs(929) <= b;
    layer0_outputs(930) <= not b;
    layer0_outputs(931) <= not (a or b);
    layer0_outputs(932) <= a xor b;
    layer0_outputs(933) <= b;
    layer0_outputs(934) <= a and not b;
    layer0_outputs(935) <= a and b;
    layer0_outputs(936) <= b and not a;
    layer0_outputs(937) <= not a;
    layer0_outputs(938) <= a or b;
    layer0_outputs(939) <= not a;
    layer0_outputs(940) <= a xor b;
    layer0_outputs(941) <= a and b;
    layer0_outputs(942) <= b;
    layer0_outputs(943) <= b;
    layer0_outputs(944) <= not (a and b);
    layer0_outputs(945) <= not b or a;
    layer0_outputs(946) <= not b;
    layer0_outputs(947) <= b;
    layer0_outputs(948) <= b;
    layer0_outputs(949) <= b;
    layer0_outputs(950) <= not b;
    layer0_outputs(951) <= a or b;
    layer0_outputs(952) <= a xor b;
    layer0_outputs(953) <= not (a or b);
    layer0_outputs(954) <= not (a xor b);
    layer0_outputs(955) <= not a or b;
    layer0_outputs(956) <= not b;
    layer0_outputs(957) <= '1';
    layer0_outputs(958) <= a or b;
    layer0_outputs(959) <= b and not a;
    layer0_outputs(960) <= not (a or b);
    layer0_outputs(961) <= not b;
    layer0_outputs(962) <= a and b;
    layer0_outputs(963) <= b and not a;
    layer0_outputs(964) <= not (a xor b);
    layer0_outputs(965) <= not a;
    layer0_outputs(966) <= not (a xor b);
    layer0_outputs(967) <= not a or b;
    layer0_outputs(968) <= a;
    layer0_outputs(969) <= not a;
    layer0_outputs(970) <= a or b;
    layer0_outputs(971) <= '1';
    layer0_outputs(972) <= a or b;
    layer0_outputs(973) <= not a;
    layer0_outputs(974) <= not (a or b);
    layer0_outputs(975) <= a xor b;
    layer0_outputs(976) <= b and not a;
    layer0_outputs(977) <= not b;
    layer0_outputs(978) <= not (a or b);
    layer0_outputs(979) <= a or b;
    layer0_outputs(980) <= not (a xor b);
    layer0_outputs(981) <= not b or a;
    layer0_outputs(982) <= not a;
    layer0_outputs(983) <= not (a xor b);
    layer0_outputs(984) <= b;
    layer0_outputs(985) <= not (a xor b);
    layer0_outputs(986) <= a and b;
    layer0_outputs(987) <= '1';
    layer0_outputs(988) <= not b;
    layer0_outputs(989) <= not b or a;
    layer0_outputs(990) <= not (a xor b);
    layer0_outputs(991) <= a and b;
    layer0_outputs(992) <= a and not b;
    layer0_outputs(993) <= '1';
    layer0_outputs(994) <= a;
    layer0_outputs(995) <= '1';
    layer0_outputs(996) <= not a or b;
    layer0_outputs(997) <= '1';
    layer0_outputs(998) <= not a;
    layer0_outputs(999) <= not a;
    layer0_outputs(1000) <= not b;
    layer0_outputs(1001) <= '1';
    layer0_outputs(1002) <= '0';
    layer0_outputs(1003) <= not (a or b);
    layer0_outputs(1004) <= a or b;
    layer0_outputs(1005) <= a;
    layer0_outputs(1006) <= not a;
    layer0_outputs(1007) <= a or b;
    layer0_outputs(1008) <= a and not b;
    layer0_outputs(1009) <= a and b;
    layer0_outputs(1010) <= not a;
    layer0_outputs(1011) <= a xor b;
    layer0_outputs(1012) <= not (a and b);
    layer0_outputs(1013) <= not (a or b);
    layer0_outputs(1014) <= not (a or b);
    layer0_outputs(1015) <= '0';
    layer0_outputs(1016) <= b and not a;
    layer0_outputs(1017) <= not a;
    layer0_outputs(1018) <= a and b;
    layer0_outputs(1019) <= a and not b;
    layer0_outputs(1020) <= not (a xor b);
    layer0_outputs(1021) <= not a or b;
    layer0_outputs(1022) <= not (a and b);
    layer0_outputs(1023) <= not (a and b);
    layer0_outputs(1024) <= b and not a;
    layer0_outputs(1025) <= not b or a;
    layer0_outputs(1026) <= not a or b;
    layer0_outputs(1027) <= not b or a;
    layer0_outputs(1028) <= '0';
    layer0_outputs(1029) <= b and not a;
    layer0_outputs(1030) <= not (a or b);
    layer0_outputs(1031) <= a xor b;
    layer0_outputs(1032) <= b;
    layer0_outputs(1033) <= a or b;
    layer0_outputs(1034) <= a xor b;
    layer0_outputs(1035) <= not a or b;
    layer0_outputs(1036) <= not (a or b);
    layer0_outputs(1037) <= not a or b;
    layer0_outputs(1038) <= a xor b;
    layer0_outputs(1039) <= not (a xor b);
    layer0_outputs(1040) <= a;
    layer0_outputs(1041) <= a or b;
    layer0_outputs(1042) <= a xor b;
    layer0_outputs(1043) <= a or b;
    layer0_outputs(1044) <= a xor b;
    layer0_outputs(1045) <= not (a or b);
    layer0_outputs(1046) <= not b or a;
    layer0_outputs(1047) <= a and not b;
    layer0_outputs(1048) <= not (a and b);
    layer0_outputs(1049) <= a xor b;
    layer0_outputs(1050) <= a and not b;
    layer0_outputs(1051) <= b;
    layer0_outputs(1052) <= not b;
    layer0_outputs(1053) <= not (a xor b);
    layer0_outputs(1054) <= b;
    layer0_outputs(1055) <= '0';
    layer0_outputs(1056) <= a and not b;
    layer0_outputs(1057) <= not a or b;
    layer0_outputs(1058) <= not (a or b);
    layer0_outputs(1059) <= not a;
    layer0_outputs(1060) <= a;
    layer0_outputs(1061) <= a and not b;
    layer0_outputs(1062) <= a and not b;
    layer0_outputs(1063) <= b;
    layer0_outputs(1064) <= b;
    layer0_outputs(1065) <= not (a or b);
    layer0_outputs(1066) <= not b or a;
    layer0_outputs(1067) <= not a;
    layer0_outputs(1068) <= not (a xor b);
    layer0_outputs(1069) <= b and not a;
    layer0_outputs(1070) <= b and not a;
    layer0_outputs(1071) <= not b or a;
    layer0_outputs(1072) <= not b or a;
    layer0_outputs(1073) <= a;
    layer0_outputs(1074) <= not b;
    layer0_outputs(1075) <= not a or b;
    layer0_outputs(1076) <= not (a or b);
    layer0_outputs(1077) <= a and b;
    layer0_outputs(1078) <= not b;
    layer0_outputs(1079) <= a or b;
    layer0_outputs(1080) <= a and b;
    layer0_outputs(1081) <= b;
    layer0_outputs(1082) <= a;
    layer0_outputs(1083) <= not b or a;
    layer0_outputs(1084) <= not (a or b);
    layer0_outputs(1085) <= b and not a;
    layer0_outputs(1086) <= not (a and b);
    layer0_outputs(1087) <= b;
    layer0_outputs(1088) <= '1';
    layer0_outputs(1089) <= not (a and b);
    layer0_outputs(1090) <= a or b;
    layer0_outputs(1091) <= not (a or b);
    layer0_outputs(1092) <= '0';
    layer0_outputs(1093) <= not (a xor b);
    layer0_outputs(1094) <= a xor b;
    layer0_outputs(1095) <= not b;
    layer0_outputs(1096) <= a;
    layer0_outputs(1097) <= not a or b;
    layer0_outputs(1098) <= not a or b;
    layer0_outputs(1099) <= not a;
    layer0_outputs(1100) <= a;
    layer0_outputs(1101) <= b and not a;
    layer0_outputs(1102) <= not a or b;
    layer0_outputs(1103) <= not b or a;
    layer0_outputs(1104) <= not (a and b);
    layer0_outputs(1105) <= not a;
    layer0_outputs(1106) <= a;
    layer0_outputs(1107) <= a;
    layer0_outputs(1108) <= not b or a;
    layer0_outputs(1109) <= not (a xor b);
    layer0_outputs(1110) <= a xor b;
    layer0_outputs(1111) <= '0';
    layer0_outputs(1112) <= not a;
    layer0_outputs(1113) <= '1';
    layer0_outputs(1114) <= not b;
    layer0_outputs(1115) <= a or b;
    layer0_outputs(1116) <= b;
    layer0_outputs(1117) <= not (a xor b);
    layer0_outputs(1118) <= not (a or b);
    layer0_outputs(1119) <= not a;
    layer0_outputs(1120) <= not b or a;
    layer0_outputs(1121) <= '0';
    layer0_outputs(1122) <= a and b;
    layer0_outputs(1123) <= not a;
    layer0_outputs(1124) <= not a;
    layer0_outputs(1125) <= b and not a;
    layer0_outputs(1126) <= a and not b;
    layer0_outputs(1127) <= not (a and b);
    layer0_outputs(1128) <= not (a or b);
    layer0_outputs(1129) <= not a;
    layer0_outputs(1130) <= not a or b;
    layer0_outputs(1131) <= b and not a;
    layer0_outputs(1132) <= b;
    layer0_outputs(1133) <= not (a or b);
    layer0_outputs(1134) <= a;
    layer0_outputs(1135) <= b;
    layer0_outputs(1136) <= a and b;
    layer0_outputs(1137) <= '1';
    layer0_outputs(1138) <= a and b;
    layer0_outputs(1139) <= not (a xor b);
    layer0_outputs(1140) <= not (a and b);
    layer0_outputs(1141) <= not (a xor b);
    layer0_outputs(1142) <= not (a or b);
    layer0_outputs(1143) <= a and not b;
    layer0_outputs(1144) <= not a;
    layer0_outputs(1145) <= b;
    layer0_outputs(1146) <= not a or b;
    layer0_outputs(1147) <= not a or b;
    layer0_outputs(1148) <= not a or b;
    layer0_outputs(1149) <= not a or b;
    layer0_outputs(1150) <= not a or b;
    layer0_outputs(1151) <= b and not a;
    layer0_outputs(1152) <= a and not b;
    layer0_outputs(1153) <= b;
    layer0_outputs(1154) <= a xor b;
    layer0_outputs(1155) <= b;
    layer0_outputs(1156) <= a and not b;
    layer0_outputs(1157) <= a;
    layer0_outputs(1158) <= not a;
    layer0_outputs(1159) <= a;
    layer0_outputs(1160) <= not b or a;
    layer0_outputs(1161) <= a and not b;
    layer0_outputs(1162) <= a;
    layer0_outputs(1163) <= not a;
    layer0_outputs(1164) <= not a or b;
    layer0_outputs(1165) <= not a;
    layer0_outputs(1166) <= '0';
    layer0_outputs(1167) <= not (a xor b);
    layer0_outputs(1168) <= not (a xor b);
    layer0_outputs(1169) <= not (a or b);
    layer0_outputs(1170) <= '0';
    layer0_outputs(1171) <= '1';
    layer0_outputs(1172) <= not b;
    layer0_outputs(1173) <= a or b;
    layer0_outputs(1174) <= not (a or b);
    layer0_outputs(1175) <= not a;
    layer0_outputs(1176) <= not (a xor b);
    layer0_outputs(1177) <= b and not a;
    layer0_outputs(1178) <= a xor b;
    layer0_outputs(1179) <= not a;
    layer0_outputs(1180) <= a and not b;
    layer0_outputs(1181) <= a or b;
    layer0_outputs(1182) <= '1';
    layer0_outputs(1183) <= b and not a;
    layer0_outputs(1184) <= b and not a;
    layer0_outputs(1185) <= a;
    layer0_outputs(1186) <= not (a and b);
    layer0_outputs(1187) <= not (a xor b);
    layer0_outputs(1188) <= not (a and b);
    layer0_outputs(1189) <= a or b;
    layer0_outputs(1190) <= b;
    layer0_outputs(1191) <= not (a or b);
    layer0_outputs(1192) <= not b or a;
    layer0_outputs(1193) <= a or b;
    layer0_outputs(1194) <= not b or a;
    layer0_outputs(1195) <= not a or b;
    layer0_outputs(1196) <= not b or a;
    layer0_outputs(1197) <= b and not a;
    layer0_outputs(1198) <= not b or a;
    layer0_outputs(1199) <= a or b;
    layer0_outputs(1200) <= '0';
    layer0_outputs(1201) <= a and not b;
    layer0_outputs(1202) <= not (a xor b);
    layer0_outputs(1203) <= a and b;
    layer0_outputs(1204) <= a xor b;
    layer0_outputs(1205) <= not a or b;
    layer0_outputs(1206) <= not (a or b);
    layer0_outputs(1207) <= a or b;
    layer0_outputs(1208) <= not (a xor b);
    layer0_outputs(1209) <= not (a and b);
    layer0_outputs(1210) <= b and not a;
    layer0_outputs(1211) <= not (a xor b);
    layer0_outputs(1212) <= not a or b;
    layer0_outputs(1213) <= not (a or b);
    layer0_outputs(1214) <= '0';
    layer0_outputs(1215) <= not b;
    layer0_outputs(1216) <= a;
    layer0_outputs(1217) <= not (a or b);
    layer0_outputs(1218) <= not b;
    layer0_outputs(1219) <= not a or b;
    layer0_outputs(1220) <= a;
    layer0_outputs(1221) <= a;
    layer0_outputs(1222) <= '1';
    layer0_outputs(1223) <= b;
    layer0_outputs(1224) <= a;
    layer0_outputs(1225) <= not b;
    layer0_outputs(1226) <= a and b;
    layer0_outputs(1227) <= a;
    layer0_outputs(1228) <= a;
    layer0_outputs(1229) <= not b or a;
    layer0_outputs(1230) <= not b;
    layer0_outputs(1231) <= not (a or b);
    layer0_outputs(1232) <= not b or a;
    layer0_outputs(1233) <= a or b;
    layer0_outputs(1234) <= a and b;
    layer0_outputs(1235) <= not (a and b);
    layer0_outputs(1236) <= '1';
    layer0_outputs(1237) <= not b;
    layer0_outputs(1238) <= not b;
    layer0_outputs(1239) <= a and b;
    layer0_outputs(1240) <= not (a or b);
    layer0_outputs(1241) <= b and not a;
    layer0_outputs(1242) <= a xor b;
    layer0_outputs(1243) <= a and not b;
    layer0_outputs(1244) <= a or b;
    layer0_outputs(1245) <= a and b;
    layer0_outputs(1246) <= not a;
    layer0_outputs(1247) <= a and b;
    layer0_outputs(1248) <= not a;
    layer0_outputs(1249) <= not a;
    layer0_outputs(1250) <= not (a and b);
    layer0_outputs(1251) <= a;
    layer0_outputs(1252) <= not (a or b);
    layer0_outputs(1253) <= not (a and b);
    layer0_outputs(1254) <= not (a xor b);
    layer0_outputs(1255) <= a or b;
    layer0_outputs(1256) <= a;
    layer0_outputs(1257) <= a xor b;
    layer0_outputs(1258) <= a xor b;
    layer0_outputs(1259) <= not a;
    layer0_outputs(1260) <= '1';
    layer0_outputs(1261) <= not b;
    layer0_outputs(1262) <= b;
    layer0_outputs(1263) <= not a;
    layer0_outputs(1264) <= not a;
    layer0_outputs(1265) <= b and not a;
    layer0_outputs(1266) <= not b or a;
    layer0_outputs(1267) <= a and b;
    layer0_outputs(1268) <= not a;
    layer0_outputs(1269) <= not b;
    layer0_outputs(1270) <= not (a xor b);
    layer0_outputs(1271) <= not b;
    layer0_outputs(1272) <= not b or a;
    layer0_outputs(1273) <= not (a xor b);
    layer0_outputs(1274) <= not (a or b);
    layer0_outputs(1275) <= a and not b;
    layer0_outputs(1276) <= a;
    layer0_outputs(1277) <= '0';
    layer0_outputs(1278) <= not a or b;
    layer0_outputs(1279) <= not b;
    layer0_outputs(1280) <= not b or a;
    layer0_outputs(1281) <= not a or b;
    layer0_outputs(1282) <= not (a xor b);
    layer0_outputs(1283) <= not (a or b);
    layer0_outputs(1284) <= a and b;
    layer0_outputs(1285) <= not a or b;
    layer0_outputs(1286) <= not (a and b);
    layer0_outputs(1287) <= not a;
    layer0_outputs(1288) <= '1';
    layer0_outputs(1289) <= b;
    layer0_outputs(1290) <= not b;
    layer0_outputs(1291) <= not (a xor b);
    layer0_outputs(1292) <= not b or a;
    layer0_outputs(1293) <= a or b;
    layer0_outputs(1294) <= not a or b;
    layer0_outputs(1295) <= not (a xor b);
    layer0_outputs(1296) <= not (a or b);
    layer0_outputs(1297) <= not a or b;
    layer0_outputs(1298) <= not b;
    layer0_outputs(1299) <= a;
    layer0_outputs(1300) <= a xor b;
    layer0_outputs(1301) <= not a;
    layer0_outputs(1302) <= not a;
    layer0_outputs(1303) <= a xor b;
    layer0_outputs(1304) <= a and not b;
    layer0_outputs(1305) <= a or b;
    layer0_outputs(1306) <= not b or a;
    layer0_outputs(1307) <= '0';
    layer0_outputs(1308) <= b;
    layer0_outputs(1309) <= '0';
    layer0_outputs(1310) <= not a;
    layer0_outputs(1311) <= '1';
    layer0_outputs(1312) <= not (a and b);
    layer0_outputs(1313) <= not a;
    layer0_outputs(1314) <= '1';
    layer0_outputs(1315) <= not a;
    layer0_outputs(1316) <= not (a xor b);
    layer0_outputs(1317) <= a and b;
    layer0_outputs(1318) <= b and not a;
    layer0_outputs(1319) <= not b;
    layer0_outputs(1320) <= b and not a;
    layer0_outputs(1321) <= not a or b;
    layer0_outputs(1322) <= not a;
    layer0_outputs(1323) <= not (a xor b);
    layer0_outputs(1324) <= '1';
    layer0_outputs(1325) <= not a or b;
    layer0_outputs(1326) <= '1';
    layer0_outputs(1327) <= not a or b;
    layer0_outputs(1328) <= not b;
    layer0_outputs(1329) <= a or b;
    layer0_outputs(1330) <= not (a or b);
    layer0_outputs(1331) <= not (a and b);
    layer0_outputs(1332) <= a xor b;
    layer0_outputs(1333) <= '1';
    layer0_outputs(1334) <= b and not a;
    layer0_outputs(1335) <= b;
    layer0_outputs(1336) <= not (a and b);
    layer0_outputs(1337) <= b and not a;
    layer0_outputs(1338) <= a;
    layer0_outputs(1339) <= not a or b;
    layer0_outputs(1340) <= not b;
    layer0_outputs(1341) <= not a;
    layer0_outputs(1342) <= not (a xor b);
    layer0_outputs(1343) <= not b or a;
    layer0_outputs(1344) <= not a or b;
    layer0_outputs(1345) <= not (a or b);
    layer0_outputs(1346) <= not a or b;
    layer0_outputs(1347) <= b and not a;
    layer0_outputs(1348) <= a or b;
    layer0_outputs(1349) <= not (a or b);
    layer0_outputs(1350) <= a and b;
    layer0_outputs(1351) <= not (a xor b);
    layer0_outputs(1352) <= b;
    layer0_outputs(1353) <= not a;
    layer0_outputs(1354) <= '1';
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= b;
    layer0_outputs(1357) <= a;
    layer0_outputs(1358) <= a and not b;
    layer0_outputs(1359) <= '1';
    layer0_outputs(1360) <= not (a or b);
    layer0_outputs(1361) <= a or b;
    layer0_outputs(1362) <= not a or b;
    layer0_outputs(1363) <= not a;
    layer0_outputs(1364) <= not (a xor b);
    layer0_outputs(1365) <= not a;
    layer0_outputs(1366) <= not a or b;
    layer0_outputs(1367) <= a xor b;
    layer0_outputs(1368) <= b and not a;
    layer0_outputs(1369) <= not a;
    layer0_outputs(1370) <= '1';
    layer0_outputs(1371) <= not (a or b);
    layer0_outputs(1372) <= b and not a;
    layer0_outputs(1373) <= b;
    layer0_outputs(1374) <= '1';
    layer0_outputs(1375) <= a xor b;
    layer0_outputs(1376) <= not b;
    layer0_outputs(1377) <= not (a or b);
    layer0_outputs(1378) <= not a;
    layer0_outputs(1379) <= b;
    layer0_outputs(1380) <= not (a or b);
    layer0_outputs(1381) <= not a;
    layer0_outputs(1382) <= b;
    layer0_outputs(1383) <= not b or a;
    layer0_outputs(1384) <= a xor b;
    layer0_outputs(1385) <= '0';
    layer0_outputs(1386) <= not (a and b);
    layer0_outputs(1387) <= not b;
    layer0_outputs(1388) <= not b;
    layer0_outputs(1389) <= not (a and b);
    layer0_outputs(1390) <= b and not a;
    layer0_outputs(1391) <= a xor b;
    layer0_outputs(1392) <= '1';
    layer0_outputs(1393) <= not (a or b);
    layer0_outputs(1394) <= not b or a;
    layer0_outputs(1395) <= b;
    layer0_outputs(1396) <= '0';
    layer0_outputs(1397) <= b and not a;
    layer0_outputs(1398) <= a or b;
    layer0_outputs(1399) <= not (a xor b);
    layer0_outputs(1400) <= not a or b;
    layer0_outputs(1401) <= a xor b;
    layer0_outputs(1402) <= not a;
    layer0_outputs(1403) <= not (a and b);
    layer0_outputs(1404) <= a and b;
    layer0_outputs(1405) <= not b;
    layer0_outputs(1406) <= a and b;
    layer0_outputs(1407) <= a and not b;
    layer0_outputs(1408) <= a and not b;
    layer0_outputs(1409) <= a or b;
    layer0_outputs(1410) <= not (a or b);
    layer0_outputs(1411) <= not b or a;
    layer0_outputs(1412) <= '0';
    layer0_outputs(1413) <= '0';
    layer0_outputs(1414) <= not (a or b);
    layer0_outputs(1415) <= not a or b;
    layer0_outputs(1416) <= not b or a;
    layer0_outputs(1417) <= not a;
    layer0_outputs(1418) <= not b;
    layer0_outputs(1419) <= a or b;
    layer0_outputs(1420) <= b;
    layer0_outputs(1421) <= not b;
    layer0_outputs(1422) <= not (a or b);
    layer0_outputs(1423) <= a or b;
    layer0_outputs(1424) <= b;
    layer0_outputs(1425) <= not (a or b);
    layer0_outputs(1426) <= a and not b;
    layer0_outputs(1427) <= a and not b;
    layer0_outputs(1428) <= a and not b;
    layer0_outputs(1429) <= '0';
    layer0_outputs(1430) <= not a or b;
    layer0_outputs(1431) <= a or b;
    layer0_outputs(1432) <= not b or a;
    layer0_outputs(1433) <= b;
    layer0_outputs(1434) <= b and not a;
    layer0_outputs(1435) <= not b;
    layer0_outputs(1436) <= not (a and b);
    layer0_outputs(1437) <= b and not a;
    layer0_outputs(1438) <= not a or b;
    layer0_outputs(1439) <= b and not a;
    layer0_outputs(1440) <= a;
    layer0_outputs(1441) <= a xor b;
    layer0_outputs(1442) <= a xor b;
    layer0_outputs(1443) <= a or b;
    layer0_outputs(1444) <= a or b;
    layer0_outputs(1445) <= '0';
    layer0_outputs(1446) <= a;
    layer0_outputs(1447) <= b and not a;
    layer0_outputs(1448) <= '1';
    layer0_outputs(1449) <= a and not b;
    layer0_outputs(1450) <= '0';
    layer0_outputs(1451) <= not b;
    layer0_outputs(1452) <= not a or b;
    layer0_outputs(1453) <= '1';
    layer0_outputs(1454) <= b;
    layer0_outputs(1455) <= a xor b;
    layer0_outputs(1456) <= '0';
    layer0_outputs(1457) <= not b;
    layer0_outputs(1458) <= a xor b;
    layer0_outputs(1459) <= not b or a;
    layer0_outputs(1460) <= not a;
    layer0_outputs(1461) <= a and not b;
    layer0_outputs(1462) <= not (a or b);
    layer0_outputs(1463) <= b;
    layer0_outputs(1464) <= not (a and b);
    layer0_outputs(1465) <= not (a xor b);
    layer0_outputs(1466) <= not (a or b);
    layer0_outputs(1467) <= '0';
    layer0_outputs(1468) <= a xor b;
    layer0_outputs(1469) <= not a;
    layer0_outputs(1470) <= not b;
    layer0_outputs(1471) <= b;
    layer0_outputs(1472) <= a and b;
    layer0_outputs(1473) <= a or b;
    layer0_outputs(1474) <= not b or a;
    layer0_outputs(1475) <= not b;
    layer0_outputs(1476) <= not (a xor b);
    layer0_outputs(1477) <= a;
    layer0_outputs(1478) <= a xor b;
    layer0_outputs(1479) <= not b or a;
    layer0_outputs(1480) <= a;
    layer0_outputs(1481) <= not (a xor b);
    layer0_outputs(1482) <= not b;
    layer0_outputs(1483) <= a and b;
    layer0_outputs(1484) <= not (a and b);
    layer0_outputs(1485) <= a and b;
    layer0_outputs(1486) <= a xor b;
    layer0_outputs(1487) <= a and b;
    layer0_outputs(1488) <= not b or a;
    layer0_outputs(1489) <= not a;
    layer0_outputs(1490) <= a and b;
    layer0_outputs(1491) <= not a;
    layer0_outputs(1492) <= a and b;
    layer0_outputs(1493) <= a and b;
    layer0_outputs(1494) <= '1';
    layer0_outputs(1495) <= not b or a;
    layer0_outputs(1496) <= a or b;
    layer0_outputs(1497) <= '0';
    layer0_outputs(1498) <= not (a or b);
    layer0_outputs(1499) <= not b or a;
    layer0_outputs(1500) <= a;
    layer0_outputs(1501) <= not b;
    layer0_outputs(1502) <= a;
    layer0_outputs(1503) <= not b;
    layer0_outputs(1504) <= a;
    layer0_outputs(1505) <= not b or a;
    layer0_outputs(1506) <= a and b;
    layer0_outputs(1507) <= not (a and b);
    layer0_outputs(1508) <= b;
    layer0_outputs(1509) <= not (a and b);
    layer0_outputs(1510) <= not b;
    layer0_outputs(1511) <= not (a xor b);
    layer0_outputs(1512) <= not (a and b);
    layer0_outputs(1513) <= not (a or b);
    layer0_outputs(1514) <= a or b;
    layer0_outputs(1515) <= b;
    layer0_outputs(1516) <= not (a xor b);
    layer0_outputs(1517) <= not (a xor b);
    layer0_outputs(1518) <= '1';
    layer0_outputs(1519) <= '0';
    layer0_outputs(1520) <= a xor b;
    layer0_outputs(1521) <= b;
    layer0_outputs(1522) <= not (a or b);
    layer0_outputs(1523) <= '0';
    layer0_outputs(1524) <= a or b;
    layer0_outputs(1525) <= b;
    layer0_outputs(1526) <= not a or b;
    layer0_outputs(1527) <= '0';
    layer0_outputs(1528) <= a and b;
    layer0_outputs(1529) <= a xor b;
    layer0_outputs(1530) <= a;
    layer0_outputs(1531) <= not b;
    layer0_outputs(1532) <= not b;
    layer0_outputs(1533) <= a or b;
    layer0_outputs(1534) <= not b;
    layer0_outputs(1535) <= not b;
    layer0_outputs(1536) <= a or b;
    layer0_outputs(1537) <= '0';
    layer0_outputs(1538) <= a;
    layer0_outputs(1539) <= not b;
    layer0_outputs(1540) <= not (a xor b);
    layer0_outputs(1541) <= b and not a;
    layer0_outputs(1542) <= b and not a;
    layer0_outputs(1543) <= a;
    layer0_outputs(1544) <= not (a or b);
    layer0_outputs(1545) <= not (a xor b);
    layer0_outputs(1546) <= a;
    layer0_outputs(1547) <= a xor b;
    layer0_outputs(1548) <= not a or b;
    layer0_outputs(1549) <= a;
    layer0_outputs(1550) <= a or b;
    layer0_outputs(1551) <= b;
    layer0_outputs(1552) <= a or b;
    layer0_outputs(1553) <= not b;
    layer0_outputs(1554) <= a;
    layer0_outputs(1555) <= a or b;
    layer0_outputs(1556) <= a;
    layer0_outputs(1557) <= not a;
    layer0_outputs(1558) <= not a;
    layer0_outputs(1559) <= not (a or b);
    layer0_outputs(1560) <= not b or a;
    layer0_outputs(1561) <= not b;
    layer0_outputs(1562) <= not a or b;
    layer0_outputs(1563) <= a and b;
    layer0_outputs(1564) <= not (a and b);
    layer0_outputs(1565) <= a;
    layer0_outputs(1566) <= a and b;
    layer0_outputs(1567) <= b;
    layer0_outputs(1568) <= b;
    layer0_outputs(1569) <= '1';
    layer0_outputs(1570) <= not (a xor b);
    layer0_outputs(1571) <= not b;
    layer0_outputs(1572) <= a and not b;
    layer0_outputs(1573) <= not (a and b);
    layer0_outputs(1574) <= a and not b;
    layer0_outputs(1575) <= not b or a;
    layer0_outputs(1576) <= a;
    layer0_outputs(1577) <= not a;
    layer0_outputs(1578) <= not a or b;
    layer0_outputs(1579) <= a;
    layer0_outputs(1580) <= '1';
    layer0_outputs(1581) <= a xor b;
    layer0_outputs(1582) <= b;
    layer0_outputs(1583) <= a;
    layer0_outputs(1584) <= a or b;
    layer0_outputs(1585) <= not b;
    layer0_outputs(1586) <= not (a xor b);
    layer0_outputs(1587) <= '1';
    layer0_outputs(1588) <= not b;
    layer0_outputs(1589) <= '1';
    layer0_outputs(1590) <= not b;
    layer0_outputs(1591) <= a xor b;
    layer0_outputs(1592) <= not (a and b);
    layer0_outputs(1593) <= '1';
    layer0_outputs(1594) <= b;
    layer0_outputs(1595) <= not (a and b);
    layer0_outputs(1596) <= not (a or b);
    layer0_outputs(1597) <= a xor b;
    layer0_outputs(1598) <= not (a and b);
    layer0_outputs(1599) <= '0';
    layer0_outputs(1600) <= b and not a;
    layer0_outputs(1601) <= '0';
    layer0_outputs(1602) <= not (a or b);
    layer0_outputs(1603) <= not (a xor b);
    layer0_outputs(1604) <= a and not b;
    layer0_outputs(1605) <= a xor b;
    layer0_outputs(1606) <= a;
    layer0_outputs(1607) <= not b;
    layer0_outputs(1608) <= not (a or b);
    layer0_outputs(1609) <= b;
    layer0_outputs(1610) <= b and not a;
    layer0_outputs(1611) <= not b or a;
    layer0_outputs(1612) <= a and not b;
    layer0_outputs(1613) <= not (a and b);
    layer0_outputs(1614) <= a and b;
    layer0_outputs(1615) <= a;
    layer0_outputs(1616) <= b;
    layer0_outputs(1617) <= '1';
    layer0_outputs(1618) <= not b;
    layer0_outputs(1619) <= not a;
    layer0_outputs(1620) <= not b;
    layer0_outputs(1621) <= not (a and b);
    layer0_outputs(1622) <= not (a xor b);
    layer0_outputs(1623) <= not b or a;
    layer0_outputs(1624) <= not b or a;
    layer0_outputs(1625) <= a;
    layer0_outputs(1626) <= not b or a;
    layer0_outputs(1627) <= '0';
    layer0_outputs(1628) <= not a or b;
    layer0_outputs(1629) <= not a;
    layer0_outputs(1630) <= b;
    layer0_outputs(1631) <= a or b;
    layer0_outputs(1632) <= not (a or b);
    layer0_outputs(1633) <= a xor b;
    layer0_outputs(1634) <= '0';
    layer0_outputs(1635) <= not b;
    layer0_outputs(1636) <= not (a or b);
    layer0_outputs(1637) <= '1';
    layer0_outputs(1638) <= a xor b;
    layer0_outputs(1639) <= b and not a;
    layer0_outputs(1640) <= a xor b;
    layer0_outputs(1641) <= a or b;
    layer0_outputs(1642) <= a or b;
    layer0_outputs(1643) <= not b;
    layer0_outputs(1644) <= a;
    layer0_outputs(1645) <= a xor b;
    layer0_outputs(1646) <= '0';
    layer0_outputs(1647) <= not a or b;
    layer0_outputs(1648) <= not (a or b);
    layer0_outputs(1649) <= not b or a;
    layer0_outputs(1650) <= not b;
    layer0_outputs(1651) <= not b;
    layer0_outputs(1652) <= a and b;
    layer0_outputs(1653) <= a and not b;
    layer0_outputs(1654) <= a and not b;
    layer0_outputs(1655) <= a xor b;
    layer0_outputs(1656) <= not (a and b);
    layer0_outputs(1657) <= not (a or b);
    layer0_outputs(1658) <= not b or a;
    layer0_outputs(1659) <= a and b;
    layer0_outputs(1660) <= not b or a;
    layer0_outputs(1661) <= not b or a;
    layer0_outputs(1662) <= b;
    layer0_outputs(1663) <= not a or b;
    layer0_outputs(1664) <= not (a or b);
    layer0_outputs(1665) <= '0';
    layer0_outputs(1666) <= a or b;
    layer0_outputs(1667) <= a and not b;
    layer0_outputs(1668) <= a or b;
    layer0_outputs(1669) <= a xor b;
    layer0_outputs(1670) <= b and not a;
    layer0_outputs(1671) <= not (a or b);
    layer0_outputs(1672) <= not (a xor b);
    layer0_outputs(1673) <= b and not a;
    layer0_outputs(1674) <= not a;
    layer0_outputs(1675) <= not (a or b);
    layer0_outputs(1676) <= not b or a;
    layer0_outputs(1677) <= '1';
    layer0_outputs(1678) <= not a;
    layer0_outputs(1679) <= not (a or b);
    layer0_outputs(1680) <= not b or a;
    layer0_outputs(1681) <= not (a and b);
    layer0_outputs(1682) <= a or b;
    layer0_outputs(1683) <= not b;
    layer0_outputs(1684) <= '0';
    layer0_outputs(1685) <= not (a xor b);
    layer0_outputs(1686) <= not a;
    layer0_outputs(1687) <= b;
    layer0_outputs(1688) <= '0';
    layer0_outputs(1689) <= a xor b;
    layer0_outputs(1690) <= not b or a;
    layer0_outputs(1691) <= not b or a;
    layer0_outputs(1692) <= not b or a;
    layer0_outputs(1693) <= b;
    layer0_outputs(1694) <= not a or b;
    layer0_outputs(1695) <= not b or a;
    layer0_outputs(1696) <= not (a and b);
    layer0_outputs(1697) <= '0';
    layer0_outputs(1698) <= a;
    layer0_outputs(1699) <= '1';
    layer0_outputs(1700) <= not (a xor b);
    layer0_outputs(1701) <= not a;
    layer0_outputs(1702) <= not (a or b);
    layer0_outputs(1703) <= a xor b;
    layer0_outputs(1704) <= b;
    layer0_outputs(1705) <= not (a or b);
    layer0_outputs(1706) <= a and not b;
    layer0_outputs(1707) <= not b or a;
    layer0_outputs(1708) <= a xor b;
    layer0_outputs(1709) <= not b;
    layer0_outputs(1710) <= a and not b;
    layer0_outputs(1711) <= not a or b;
    layer0_outputs(1712) <= not a or b;
    layer0_outputs(1713) <= '0';
    layer0_outputs(1714) <= a xor b;
    layer0_outputs(1715) <= not b or a;
    layer0_outputs(1716) <= not (a or b);
    layer0_outputs(1717) <= b and not a;
    layer0_outputs(1718) <= not b or a;
    layer0_outputs(1719) <= not (a and b);
    layer0_outputs(1720) <= not (a and b);
    layer0_outputs(1721) <= a xor b;
    layer0_outputs(1722) <= not (a or b);
    layer0_outputs(1723) <= not a;
    layer0_outputs(1724) <= b and not a;
    layer0_outputs(1725) <= a and not b;
    layer0_outputs(1726) <= not b or a;
    layer0_outputs(1727) <= not b or a;
    layer0_outputs(1728) <= not (a or b);
    layer0_outputs(1729) <= not a;
    layer0_outputs(1730) <= '0';
    layer0_outputs(1731) <= a and b;
    layer0_outputs(1732) <= a and not b;
    layer0_outputs(1733) <= not b or a;
    layer0_outputs(1734) <= '1';
    layer0_outputs(1735) <= not b;
    layer0_outputs(1736) <= not (a or b);
    layer0_outputs(1737) <= '0';
    layer0_outputs(1738) <= not b or a;
    layer0_outputs(1739) <= not a or b;
    layer0_outputs(1740) <= b and not a;
    layer0_outputs(1741) <= a xor b;
    layer0_outputs(1742) <= not (a xor b);
    layer0_outputs(1743) <= not a;
    layer0_outputs(1744) <= not (a xor b);
    layer0_outputs(1745) <= not (a and b);
    layer0_outputs(1746) <= not (a or b);
    layer0_outputs(1747) <= not a;
    layer0_outputs(1748) <= a or b;
    layer0_outputs(1749) <= a and not b;
    layer0_outputs(1750) <= '0';
    layer0_outputs(1751) <= a;
    layer0_outputs(1752) <= not a or b;
    layer0_outputs(1753) <= not a or b;
    layer0_outputs(1754) <= b;
    layer0_outputs(1755) <= not (a or b);
    layer0_outputs(1756) <= not b or a;
    layer0_outputs(1757) <= not (a and b);
    layer0_outputs(1758) <= a;
    layer0_outputs(1759) <= a xor b;
    layer0_outputs(1760) <= not b or a;
    layer0_outputs(1761) <= not (a xor b);
    layer0_outputs(1762) <= a xor b;
    layer0_outputs(1763) <= not a or b;
    layer0_outputs(1764) <= '1';
    layer0_outputs(1765) <= a and not b;
    layer0_outputs(1766) <= b;
    layer0_outputs(1767) <= not (a and b);
    layer0_outputs(1768) <= a xor b;
    layer0_outputs(1769) <= b;
    layer0_outputs(1770) <= not a;
    layer0_outputs(1771) <= not a or b;
    layer0_outputs(1772) <= a or b;
    layer0_outputs(1773) <= not a;
    layer0_outputs(1774) <= a and b;
    layer0_outputs(1775) <= a;
    layer0_outputs(1776) <= a and not b;
    layer0_outputs(1777) <= a or b;
    layer0_outputs(1778) <= a;
    layer0_outputs(1779) <= a and not b;
    layer0_outputs(1780) <= not (a xor b);
    layer0_outputs(1781) <= not b;
    layer0_outputs(1782) <= not (a xor b);
    layer0_outputs(1783) <= b and not a;
    layer0_outputs(1784) <= not (a and b);
    layer0_outputs(1785) <= not a;
    layer0_outputs(1786) <= b and not a;
    layer0_outputs(1787) <= not (a or b);
    layer0_outputs(1788) <= b and not a;
    layer0_outputs(1789) <= a and not b;
    layer0_outputs(1790) <= a;
    layer0_outputs(1791) <= b;
    layer0_outputs(1792) <= a or b;
    layer0_outputs(1793) <= not b or a;
    layer0_outputs(1794) <= not b;
    layer0_outputs(1795) <= a;
    layer0_outputs(1796) <= a and b;
    layer0_outputs(1797) <= a or b;
    layer0_outputs(1798) <= not (a or b);
    layer0_outputs(1799) <= '1';
    layer0_outputs(1800) <= a or b;
    layer0_outputs(1801) <= b;
    layer0_outputs(1802) <= '0';
    layer0_outputs(1803) <= a xor b;
    layer0_outputs(1804) <= b;
    layer0_outputs(1805) <= a xor b;
    layer0_outputs(1806) <= a;
    layer0_outputs(1807) <= not b;
    layer0_outputs(1808) <= b and not a;
    layer0_outputs(1809) <= '1';
    layer0_outputs(1810) <= a and b;
    layer0_outputs(1811) <= a or b;
    layer0_outputs(1812) <= not b;
    layer0_outputs(1813) <= not b or a;
    layer0_outputs(1814) <= a xor b;
    layer0_outputs(1815) <= not (a xor b);
    layer0_outputs(1816) <= not a;
    layer0_outputs(1817) <= '1';
    layer0_outputs(1818) <= not (a or b);
    layer0_outputs(1819) <= not (a xor b);
    layer0_outputs(1820) <= not (a or b);
    layer0_outputs(1821) <= not (a and b);
    layer0_outputs(1822) <= not a or b;
    layer0_outputs(1823) <= '0';
    layer0_outputs(1824) <= not a or b;
    layer0_outputs(1825) <= '0';
    layer0_outputs(1826) <= not (a or b);
    layer0_outputs(1827) <= a and not b;
    layer0_outputs(1828) <= a;
    layer0_outputs(1829) <= not b or a;
    layer0_outputs(1830) <= not (a and b);
    layer0_outputs(1831) <= b and not a;
    layer0_outputs(1832) <= '0';
    layer0_outputs(1833) <= not b or a;
    layer0_outputs(1834) <= b;
    layer0_outputs(1835) <= b;
    layer0_outputs(1836) <= not (a or b);
    layer0_outputs(1837) <= not a;
    layer0_outputs(1838) <= a or b;
    layer0_outputs(1839) <= not a or b;
    layer0_outputs(1840) <= b and not a;
    layer0_outputs(1841) <= b and not a;
    layer0_outputs(1842) <= a or b;
    layer0_outputs(1843) <= not (a xor b);
    layer0_outputs(1844) <= not (a and b);
    layer0_outputs(1845) <= a or b;
    layer0_outputs(1846) <= not (a or b);
    layer0_outputs(1847) <= not (a or b);
    layer0_outputs(1848) <= b;
    layer0_outputs(1849) <= a and not b;
    layer0_outputs(1850) <= a xor b;
    layer0_outputs(1851) <= not a;
    layer0_outputs(1852) <= b;
    layer0_outputs(1853) <= b;
    layer0_outputs(1854) <= '0';
    layer0_outputs(1855) <= b;
    layer0_outputs(1856) <= not a;
    layer0_outputs(1857) <= a or b;
    layer0_outputs(1858) <= b and not a;
    layer0_outputs(1859) <= b and not a;
    layer0_outputs(1860) <= '0';
    layer0_outputs(1861) <= b and not a;
    layer0_outputs(1862) <= b and not a;
    layer0_outputs(1863) <= a and not b;
    layer0_outputs(1864) <= b;
    layer0_outputs(1865) <= not a or b;
    layer0_outputs(1866) <= b;
    layer0_outputs(1867) <= not b or a;
    layer0_outputs(1868) <= not a or b;
    layer0_outputs(1869) <= a and b;
    layer0_outputs(1870) <= a xor b;
    layer0_outputs(1871) <= '1';
    layer0_outputs(1872) <= a or b;
    layer0_outputs(1873) <= b and not a;
    layer0_outputs(1874) <= not b or a;
    layer0_outputs(1875) <= not (a and b);
    layer0_outputs(1876) <= not b;
    layer0_outputs(1877) <= a and b;
    layer0_outputs(1878) <= a xor b;
    layer0_outputs(1879) <= a or b;
    layer0_outputs(1880) <= a and b;
    layer0_outputs(1881) <= not (a and b);
    layer0_outputs(1882) <= a and b;
    layer0_outputs(1883) <= b and not a;
    layer0_outputs(1884) <= a xor b;
    layer0_outputs(1885) <= not a or b;
    layer0_outputs(1886) <= '1';
    layer0_outputs(1887) <= a and not b;
    layer0_outputs(1888) <= a;
    layer0_outputs(1889) <= a;
    layer0_outputs(1890) <= '0';
    layer0_outputs(1891) <= not a or b;
    layer0_outputs(1892) <= a;
    layer0_outputs(1893) <= a and not b;
    layer0_outputs(1894) <= not a;
    layer0_outputs(1895) <= a and not b;
    layer0_outputs(1896) <= a and b;
    layer0_outputs(1897) <= '0';
    layer0_outputs(1898) <= not (a or b);
    layer0_outputs(1899) <= a;
    layer0_outputs(1900) <= not a or b;
    layer0_outputs(1901) <= '1';
    layer0_outputs(1902) <= not a;
    layer0_outputs(1903) <= a xor b;
    layer0_outputs(1904) <= not (a xor b);
    layer0_outputs(1905) <= b;
    layer0_outputs(1906) <= not (a xor b);
    layer0_outputs(1907) <= '1';
    layer0_outputs(1908) <= a;
    layer0_outputs(1909) <= b;
    layer0_outputs(1910) <= not b or a;
    layer0_outputs(1911) <= b;
    layer0_outputs(1912) <= a or b;
    layer0_outputs(1913) <= not b or a;
    layer0_outputs(1914) <= not (a or b);
    layer0_outputs(1915) <= a or b;
    layer0_outputs(1916) <= not a or b;
    layer0_outputs(1917) <= not b;
    layer0_outputs(1918) <= not a or b;
    layer0_outputs(1919) <= a;
    layer0_outputs(1920) <= not (a or b);
    layer0_outputs(1921) <= not a;
    layer0_outputs(1922) <= a or b;
    layer0_outputs(1923) <= '1';
    layer0_outputs(1924) <= not b;
    layer0_outputs(1925) <= not (a or b);
    layer0_outputs(1926) <= a or b;
    layer0_outputs(1927) <= not (a xor b);
    layer0_outputs(1928) <= not (a xor b);
    layer0_outputs(1929) <= not b;
    layer0_outputs(1930) <= a;
    layer0_outputs(1931) <= a or b;
    layer0_outputs(1932) <= not b;
    layer0_outputs(1933) <= not a or b;
    layer0_outputs(1934) <= b and not a;
    layer0_outputs(1935) <= '1';
    layer0_outputs(1936) <= a;
    layer0_outputs(1937) <= not (a xor b);
    layer0_outputs(1938) <= '1';
    layer0_outputs(1939) <= a;
    layer0_outputs(1940) <= not a;
    layer0_outputs(1941) <= not b;
    layer0_outputs(1942) <= '1';
    layer0_outputs(1943) <= not b or a;
    layer0_outputs(1944) <= '1';
    layer0_outputs(1945) <= not a or b;
    layer0_outputs(1946) <= not b or a;
    layer0_outputs(1947) <= a xor b;
    layer0_outputs(1948) <= not a or b;
    layer0_outputs(1949) <= a and not b;
    layer0_outputs(1950) <= b and not a;
    layer0_outputs(1951) <= a xor b;
    layer0_outputs(1952) <= not a;
    layer0_outputs(1953) <= not (a or b);
    layer0_outputs(1954) <= a or b;
    layer0_outputs(1955) <= not (a or b);
    layer0_outputs(1956) <= '0';
    layer0_outputs(1957) <= a and b;
    layer0_outputs(1958) <= not b or a;
    layer0_outputs(1959) <= a and not b;
    layer0_outputs(1960) <= a;
    layer0_outputs(1961) <= b and not a;
    layer0_outputs(1962) <= b;
    layer0_outputs(1963) <= b and not a;
    layer0_outputs(1964) <= not a;
    layer0_outputs(1965) <= not b;
    layer0_outputs(1966) <= not a or b;
    layer0_outputs(1967) <= '1';
    layer0_outputs(1968) <= a;
    layer0_outputs(1969) <= a or b;
    layer0_outputs(1970) <= b;
    layer0_outputs(1971) <= not b or a;
    layer0_outputs(1972) <= a xor b;
    layer0_outputs(1973) <= '1';
    layer0_outputs(1974) <= '1';
    layer0_outputs(1975) <= not (a or b);
    layer0_outputs(1976) <= not (a xor b);
    layer0_outputs(1977) <= not (a xor b);
    layer0_outputs(1978) <= b;
    layer0_outputs(1979) <= not (a or b);
    layer0_outputs(1980) <= a xor b;
    layer0_outputs(1981) <= a or b;
    layer0_outputs(1982) <= not a or b;
    layer0_outputs(1983) <= not (a or b);
    layer0_outputs(1984) <= a xor b;
    layer0_outputs(1985) <= '1';
    layer0_outputs(1986) <= a;
    layer0_outputs(1987) <= not a;
    layer0_outputs(1988) <= not (a or b);
    layer0_outputs(1989) <= a xor b;
    layer0_outputs(1990) <= b;
    layer0_outputs(1991) <= b and not a;
    layer0_outputs(1992) <= not (a xor b);
    layer0_outputs(1993) <= a or b;
    layer0_outputs(1994) <= b and not a;
    layer0_outputs(1995) <= not b;
    layer0_outputs(1996) <= '1';
    layer0_outputs(1997) <= not (a xor b);
    layer0_outputs(1998) <= not (a or b);
    layer0_outputs(1999) <= not (a or b);
    layer0_outputs(2000) <= a;
    layer0_outputs(2001) <= a xor b;
    layer0_outputs(2002) <= not a;
    layer0_outputs(2003) <= a;
    layer0_outputs(2004) <= not b;
    layer0_outputs(2005) <= a;
    layer0_outputs(2006) <= not b or a;
    layer0_outputs(2007) <= a or b;
    layer0_outputs(2008) <= a;
    layer0_outputs(2009) <= not b or a;
    layer0_outputs(2010) <= b;
    layer0_outputs(2011) <= b;
    layer0_outputs(2012) <= b and not a;
    layer0_outputs(2013) <= not (a or b);
    layer0_outputs(2014) <= b;
    layer0_outputs(2015) <= a xor b;
    layer0_outputs(2016) <= not a;
    layer0_outputs(2017) <= not a or b;
    layer0_outputs(2018) <= not b;
    layer0_outputs(2019) <= not a or b;
    layer0_outputs(2020) <= not b;
    layer0_outputs(2021) <= not (a or b);
    layer0_outputs(2022) <= a xor b;
    layer0_outputs(2023) <= not (a xor b);
    layer0_outputs(2024) <= b;
    layer0_outputs(2025) <= not a or b;
    layer0_outputs(2026) <= a and not b;
    layer0_outputs(2027) <= b;
    layer0_outputs(2028) <= not a or b;
    layer0_outputs(2029) <= '1';
    layer0_outputs(2030) <= not b or a;
    layer0_outputs(2031) <= a xor b;
    layer0_outputs(2032) <= a;
    layer0_outputs(2033) <= not b;
    layer0_outputs(2034) <= b;
    layer0_outputs(2035) <= a or b;
    layer0_outputs(2036) <= '1';
    layer0_outputs(2037) <= a or b;
    layer0_outputs(2038) <= b and not a;
    layer0_outputs(2039) <= not a or b;
    layer0_outputs(2040) <= a and b;
    layer0_outputs(2041) <= not a;
    layer0_outputs(2042) <= not b or a;
    layer0_outputs(2043) <= '1';
    layer0_outputs(2044) <= not b;
    layer0_outputs(2045) <= '1';
    layer0_outputs(2046) <= not (a xor b);
    layer0_outputs(2047) <= b and not a;
    layer0_outputs(2048) <= a and b;
    layer0_outputs(2049) <= not a or b;
    layer0_outputs(2050) <= b;
    layer0_outputs(2051) <= not a or b;
    layer0_outputs(2052) <= not (a or b);
    layer0_outputs(2053) <= b;
    layer0_outputs(2054) <= not (a xor b);
    layer0_outputs(2055) <= '0';
    layer0_outputs(2056) <= not (a xor b);
    layer0_outputs(2057) <= not b or a;
    layer0_outputs(2058) <= not (a or b);
    layer0_outputs(2059) <= a xor b;
    layer0_outputs(2060) <= not (a and b);
    layer0_outputs(2061) <= not (a or b);
    layer0_outputs(2062) <= not a or b;
    layer0_outputs(2063) <= not (a xor b);
    layer0_outputs(2064) <= a or b;
    layer0_outputs(2065) <= not (a xor b);
    layer0_outputs(2066) <= not a or b;
    layer0_outputs(2067) <= not (a or b);
    layer0_outputs(2068) <= b;
    layer0_outputs(2069) <= not (a xor b);
    layer0_outputs(2070) <= not a;
    layer0_outputs(2071) <= b and not a;
    layer0_outputs(2072) <= a;
    layer0_outputs(2073) <= not (a xor b);
    layer0_outputs(2074) <= '0';
    layer0_outputs(2075) <= not a;
    layer0_outputs(2076) <= not b;
    layer0_outputs(2077) <= a or b;
    layer0_outputs(2078) <= a and b;
    layer0_outputs(2079) <= '1';
    layer0_outputs(2080) <= a and not b;
    layer0_outputs(2081) <= '0';
    layer0_outputs(2082) <= '1';
    layer0_outputs(2083) <= '1';
    layer0_outputs(2084) <= a and not b;
    layer0_outputs(2085) <= a and b;
    layer0_outputs(2086) <= a and b;
    layer0_outputs(2087) <= a xor b;
    layer0_outputs(2088) <= not (a or b);
    layer0_outputs(2089) <= a;
    layer0_outputs(2090) <= a and not b;
    layer0_outputs(2091) <= not (a or b);
    layer0_outputs(2092) <= not a;
    layer0_outputs(2093) <= not b or a;
    layer0_outputs(2094) <= a xor b;
    layer0_outputs(2095) <= not (a xor b);
    layer0_outputs(2096) <= '1';
    layer0_outputs(2097) <= a and not b;
    layer0_outputs(2098) <= not a;
    layer0_outputs(2099) <= b;
    layer0_outputs(2100) <= not b or a;
    layer0_outputs(2101) <= a xor b;
    layer0_outputs(2102) <= not a or b;
    layer0_outputs(2103) <= a and not b;
    layer0_outputs(2104) <= a or b;
    layer0_outputs(2105) <= '0';
    layer0_outputs(2106) <= not a or b;
    layer0_outputs(2107) <= a and b;
    layer0_outputs(2108) <= not (a and b);
    layer0_outputs(2109) <= a and b;
    layer0_outputs(2110) <= not (a and b);
    layer0_outputs(2111) <= not (a and b);
    layer0_outputs(2112) <= not b;
    layer0_outputs(2113) <= '1';
    layer0_outputs(2114) <= not (a xor b);
    layer0_outputs(2115) <= a xor b;
    layer0_outputs(2116) <= a and b;
    layer0_outputs(2117) <= not (a or b);
    layer0_outputs(2118) <= not a or b;
    layer0_outputs(2119) <= a xor b;
    layer0_outputs(2120) <= not b;
    layer0_outputs(2121) <= a;
    layer0_outputs(2122) <= not b;
    layer0_outputs(2123) <= a and b;
    layer0_outputs(2124) <= a and b;
    layer0_outputs(2125) <= not (a xor b);
    layer0_outputs(2126) <= a and b;
    layer0_outputs(2127) <= '1';
    layer0_outputs(2128) <= '1';
    layer0_outputs(2129) <= b and not a;
    layer0_outputs(2130) <= b;
    layer0_outputs(2131) <= a and b;
    layer0_outputs(2132) <= not (a or b);
    layer0_outputs(2133) <= '1';
    layer0_outputs(2134) <= not a or b;
    layer0_outputs(2135) <= a xor b;
    layer0_outputs(2136) <= b and not a;
    layer0_outputs(2137) <= not b or a;
    layer0_outputs(2138) <= not (a xor b);
    layer0_outputs(2139) <= b and not a;
    layer0_outputs(2140) <= not (a or b);
    layer0_outputs(2141) <= not (a or b);
    layer0_outputs(2142) <= not (a or b);
    layer0_outputs(2143) <= b;
    layer0_outputs(2144) <= not (a or b);
    layer0_outputs(2145) <= '1';
    layer0_outputs(2146) <= a or b;
    layer0_outputs(2147) <= not (a and b);
    layer0_outputs(2148) <= not a;
    layer0_outputs(2149) <= b and not a;
    layer0_outputs(2150) <= b;
    layer0_outputs(2151) <= b;
    layer0_outputs(2152) <= a;
    layer0_outputs(2153) <= a;
    layer0_outputs(2154) <= a and not b;
    layer0_outputs(2155) <= not a or b;
    layer0_outputs(2156) <= a and not b;
    layer0_outputs(2157) <= '1';
    layer0_outputs(2158) <= b;
    layer0_outputs(2159) <= not a or b;
    layer0_outputs(2160) <= a;
    layer0_outputs(2161) <= a and b;
    layer0_outputs(2162) <= not (a or b);
    layer0_outputs(2163) <= '0';
    layer0_outputs(2164) <= a and not b;
    layer0_outputs(2165) <= a and not b;
    layer0_outputs(2166) <= not a;
    layer0_outputs(2167) <= not (a xor b);
    layer0_outputs(2168) <= not (a and b);
    layer0_outputs(2169) <= a xor b;
    layer0_outputs(2170) <= b and not a;
    layer0_outputs(2171) <= not b;
    layer0_outputs(2172) <= b and not a;
    layer0_outputs(2173) <= b and not a;
    layer0_outputs(2174) <= '1';
    layer0_outputs(2175) <= not (a or b);
    layer0_outputs(2176) <= not a or b;
    layer0_outputs(2177) <= not (a or b);
    layer0_outputs(2178) <= a or b;
    layer0_outputs(2179) <= a and b;
    layer0_outputs(2180) <= a xor b;
    layer0_outputs(2181) <= a;
    layer0_outputs(2182) <= '1';
    layer0_outputs(2183) <= b;
    layer0_outputs(2184) <= '0';
    layer0_outputs(2185) <= a xor b;
    layer0_outputs(2186) <= '0';
    layer0_outputs(2187) <= not b or a;
    layer0_outputs(2188) <= not (a or b);
    layer0_outputs(2189) <= b;
    layer0_outputs(2190) <= '0';
    layer0_outputs(2191) <= not a or b;
    layer0_outputs(2192) <= not (a and b);
    layer0_outputs(2193) <= b and not a;
    layer0_outputs(2194) <= '1';
    layer0_outputs(2195) <= not (a or b);
    layer0_outputs(2196) <= not (a or b);
    layer0_outputs(2197) <= not (a or b);
    layer0_outputs(2198) <= a and b;
    layer0_outputs(2199) <= a xor b;
    layer0_outputs(2200) <= a or b;
    layer0_outputs(2201) <= not b or a;
    layer0_outputs(2202) <= a;
    layer0_outputs(2203) <= a and not b;
    layer0_outputs(2204) <= a;
    layer0_outputs(2205) <= a and not b;
    layer0_outputs(2206) <= a;
    layer0_outputs(2207) <= not (a xor b);
    layer0_outputs(2208) <= a and not b;
    layer0_outputs(2209) <= a or b;
    layer0_outputs(2210) <= a;
    layer0_outputs(2211) <= a or b;
    layer0_outputs(2212) <= not (a or b);
    layer0_outputs(2213) <= a or b;
    layer0_outputs(2214) <= not (a xor b);
    layer0_outputs(2215) <= not b or a;
    layer0_outputs(2216) <= a;
    layer0_outputs(2217) <= not (a or b);
    layer0_outputs(2218) <= a and not b;
    layer0_outputs(2219) <= a xor b;
    layer0_outputs(2220) <= not (a xor b);
    layer0_outputs(2221) <= not a;
    layer0_outputs(2222) <= not (a or b);
    layer0_outputs(2223) <= not b or a;
    layer0_outputs(2224) <= a or b;
    layer0_outputs(2225) <= not (a or b);
    layer0_outputs(2226) <= not (a or b);
    layer0_outputs(2227) <= a and not b;
    layer0_outputs(2228) <= not (a xor b);
    layer0_outputs(2229) <= '0';
    layer0_outputs(2230) <= a and b;
    layer0_outputs(2231) <= a and not b;
    layer0_outputs(2232) <= b;
    layer0_outputs(2233) <= b;
    layer0_outputs(2234) <= not a or b;
    layer0_outputs(2235) <= a and b;
    layer0_outputs(2236) <= a xor b;
    layer0_outputs(2237) <= not b or a;
    layer0_outputs(2238) <= not a or b;
    layer0_outputs(2239) <= not (a and b);
    layer0_outputs(2240) <= b and not a;
    layer0_outputs(2241) <= b;
    layer0_outputs(2242) <= a and b;
    layer0_outputs(2243) <= not a or b;
    layer0_outputs(2244) <= not a or b;
    layer0_outputs(2245) <= not (a and b);
    layer0_outputs(2246) <= b;
    layer0_outputs(2247) <= not b or a;
    layer0_outputs(2248) <= not a;
    layer0_outputs(2249) <= b;
    layer0_outputs(2250) <= not (a and b);
    layer0_outputs(2251) <= a xor b;
    layer0_outputs(2252) <= a or b;
    layer0_outputs(2253) <= not b or a;
    layer0_outputs(2254) <= b;
    layer0_outputs(2255) <= '1';
    layer0_outputs(2256) <= a or b;
    layer0_outputs(2257) <= b;
    layer0_outputs(2258) <= not (a and b);
    layer0_outputs(2259) <= '0';
    layer0_outputs(2260) <= not b or a;
    layer0_outputs(2261) <= '0';
    layer0_outputs(2262) <= not (a xor b);
    layer0_outputs(2263) <= '0';
    layer0_outputs(2264) <= not a;
    layer0_outputs(2265) <= not a or b;
    layer0_outputs(2266) <= '0';
    layer0_outputs(2267) <= b;
    layer0_outputs(2268) <= not b;
    layer0_outputs(2269) <= b;
    layer0_outputs(2270) <= a xor b;
    layer0_outputs(2271) <= not b or a;
    layer0_outputs(2272) <= b;
    layer0_outputs(2273) <= '0';
    layer0_outputs(2274) <= not b;
    layer0_outputs(2275) <= a or b;
    layer0_outputs(2276) <= not (a xor b);
    layer0_outputs(2277) <= not b;
    layer0_outputs(2278) <= not (a and b);
    layer0_outputs(2279) <= not (a or b);
    layer0_outputs(2280) <= a or b;
    layer0_outputs(2281) <= b and not a;
    layer0_outputs(2282) <= a;
    layer0_outputs(2283) <= not b or a;
    layer0_outputs(2284) <= not (a or b);
    layer0_outputs(2285) <= not b;
    layer0_outputs(2286) <= a;
    layer0_outputs(2287) <= b;
    layer0_outputs(2288) <= not (a xor b);
    layer0_outputs(2289) <= b;
    layer0_outputs(2290) <= a or b;
    layer0_outputs(2291) <= not (a or b);
    layer0_outputs(2292) <= not (a or b);
    layer0_outputs(2293) <= '0';
    layer0_outputs(2294) <= not (a xor b);
    layer0_outputs(2295) <= '1';
    layer0_outputs(2296) <= not (a or b);
    layer0_outputs(2297) <= '0';
    layer0_outputs(2298) <= not a or b;
    layer0_outputs(2299) <= b;
    layer0_outputs(2300) <= not b;
    layer0_outputs(2301) <= not b;
    layer0_outputs(2302) <= '0';
    layer0_outputs(2303) <= b and not a;
    layer0_outputs(2304) <= not b;
    layer0_outputs(2305) <= b;
    layer0_outputs(2306) <= not a;
    layer0_outputs(2307) <= not b;
    layer0_outputs(2308) <= not a or b;
    layer0_outputs(2309) <= '1';
    layer0_outputs(2310) <= not b;
    layer0_outputs(2311) <= a;
    layer0_outputs(2312) <= not b;
    layer0_outputs(2313) <= not (a xor b);
    layer0_outputs(2314) <= a xor b;
    layer0_outputs(2315) <= not (a xor b);
    layer0_outputs(2316) <= b;
    layer0_outputs(2317) <= not a or b;
    layer0_outputs(2318) <= not a or b;
    layer0_outputs(2319) <= b;
    layer0_outputs(2320) <= b and not a;
    layer0_outputs(2321) <= a xor b;
    layer0_outputs(2322) <= not (a and b);
    layer0_outputs(2323) <= '0';
    layer0_outputs(2324) <= not b or a;
    layer0_outputs(2325) <= not a or b;
    layer0_outputs(2326) <= b;
    layer0_outputs(2327) <= b;
    layer0_outputs(2328) <= not (a xor b);
    layer0_outputs(2329) <= a xor b;
    layer0_outputs(2330) <= not b;
    layer0_outputs(2331) <= b;
    layer0_outputs(2332) <= a;
    layer0_outputs(2333) <= a and not b;
    layer0_outputs(2334) <= '1';
    layer0_outputs(2335) <= not (a and b);
    layer0_outputs(2336) <= not b or a;
    layer0_outputs(2337) <= not a or b;
    layer0_outputs(2338) <= not (a xor b);
    layer0_outputs(2339) <= a and b;
    layer0_outputs(2340) <= '0';
    layer0_outputs(2341) <= not a or b;
    layer0_outputs(2342) <= not (a or b);
    layer0_outputs(2343) <= b;
    layer0_outputs(2344) <= not (a xor b);
    layer0_outputs(2345) <= not b or a;
    layer0_outputs(2346) <= b;
    layer0_outputs(2347) <= a;
    layer0_outputs(2348) <= b and not a;
    layer0_outputs(2349) <= a;
    layer0_outputs(2350) <= b;
    layer0_outputs(2351) <= a and not b;
    layer0_outputs(2352) <= a;
    layer0_outputs(2353) <= not (a and b);
    layer0_outputs(2354) <= not a or b;
    layer0_outputs(2355) <= a and b;
    layer0_outputs(2356) <= not (a xor b);
    layer0_outputs(2357) <= not (a or b);
    layer0_outputs(2358) <= not b;
    layer0_outputs(2359) <= not b;
    layer0_outputs(2360) <= not (a and b);
    layer0_outputs(2361) <= not (a or b);
    layer0_outputs(2362) <= a or b;
    layer0_outputs(2363) <= not a or b;
    layer0_outputs(2364) <= not (a and b);
    layer0_outputs(2365) <= a and b;
    layer0_outputs(2366) <= not (a or b);
    layer0_outputs(2367) <= '0';
    layer0_outputs(2368) <= a or b;
    layer0_outputs(2369) <= '1';
    layer0_outputs(2370) <= not (a or b);
    layer0_outputs(2371) <= b;
    layer0_outputs(2372) <= not b;
    layer0_outputs(2373) <= not (a xor b);
    layer0_outputs(2374) <= a xor b;
    layer0_outputs(2375) <= not (a xor b);
    layer0_outputs(2376) <= a;
    layer0_outputs(2377) <= not (a xor b);
    layer0_outputs(2378) <= not a;
    layer0_outputs(2379) <= not (a and b);
    layer0_outputs(2380) <= not (a xor b);
    layer0_outputs(2381) <= a xor b;
    layer0_outputs(2382) <= not a;
    layer0_outputs(2383) <= not b or a;
    layer0_outputs(2384) <= a or b;
    layer0_outputs(2385) <= a or b;
    layer0_outputs(2386) <= a or b;
    layer0_outputs(2387) <= b;
    layer0_outputs(2388) <= not (a xor b);
    layer0_outputs(2389) <= not b;
    layer0_outputs(2390) <= a or b;
    layer0_outputs(2391) <= '0';
    layer0_outputs(2392) <= not b;
    layer0_outputs(2393) <= not b or a;
    layer0_outputs(2394) <= b and not a;
    layer0_outputs(2395) <= not b;
    layer0_outputs(2396) <= b;
    layer0_outputs(2397) <= a xor b;
    layer0_outputs(2398) <= not (a and b);
    layer0_outputs(2399) <= a and not b;
    layer0_outputs(2400) <= not (a or b);
    layer0_outputs(2401) <= a xor b;
    layer0_outputs(2402) <= a;
    layer0_outputs(2403) <= not b or a;
    layer0_outputs(2404) <= b and not a;
    layer0_outputs(2405) <= a and not b;
    layer0_outputs(2406) <= a xor b;
    layer0_outputs(2407) <= not b;
    layer0_outputs(2408) <= not b or a;
    layer0_outputs(2409) <= not a or b;
    layer0_outputs(2410) <= a;
    layer0_outputs(2411) <= '1';
    layer0_outputs(2412) <= not b;
    layer0_outputs(2413) <= '0';
    layer0_outputs(2414) <= a or b;
    layer0_outputs(2415) <= not (a or b);
    layer0_outputs(2416) <= b;
    layer0_outputs(2417) <= a;
    layer0_outputs(2418) <= b and not a;
    layer0_outputs(2419) <= b and not a;
    layer0_outputs(2420) <= not b or a;
    layer0_outputs(2421) <= not a;
    layer0_outputs(2422) <= a or b;
    layer0_outputs(2423) <= not b or a;
    layer0_outputs(2424) <= a and not b;
    layer0_outputs(2425) <= b and not a;
    layer0_outputs(2426) <= not b;
    layer0_outputs(2427) <= not (a and b);
    layer0_outputs(2428) <= a;
    layer0_outputs(2429) <= a or b;
    layer0_outputs(2430) <= a;
    layer0_outputs(2431) <= b;
    layer0_outputs(2432) <= a;
    layer0_outputs(2433) <= not (a and b);
    layer0_outputs(2434) <= a or b;
    layer0_outputs(2435) <= not b or a;
    layer0_outputs(2436) <= a and b;
    layer0_outputs(2437) <= b;
    layer0_outputs(2438) <= a;
    layer0_outputs(2439) <= a or b;
    layer0_outputs(2440) <= not (a or b);
    layer0_outputs(2441) <= a and not b;
    layer0_outputs(2442) <= not a or b;
    layer0_outputs(2443) <= '1';
    layer0_outputs(2444) <= b;
    layer0_outputs(2445) <= a;
    layer0_outputs(2446) <= not (a xor b);
    layer0_outputs(2447) <= not b;
    layer0_outputs(2448) <= not a;
    layer0_outputs(2449) <= not (a xor b);
    layer0_outputs(2450) <= not b or a;
    layer0_outputs(2451) <= not a;
    layer0_outputs(2452) <= a;
    layer0_outputs(2453) <= '0';
    layer0_outputs(2454) <= b and not a;
    layer0_outputs(2455) <= not (a or b);
    layer0_outputs(2456) <= a and b;
    layer0_outputs(2457) <= a;
    layer0_outputs(2458) <= not b;
    layer0_outputs(2459) <= not (a or b);
    layer0_outputs(2460) <= a or b;
    layer0_outputs(2461) <= a and b;
    layer0_outputs(2462) <= a or b;
    layer0_outputs(2463) <= a xor b;
    layer0_outputs(2464) <= not a or b;
    layer0_outputs(2465) <= a and b;
    layer0_outputs(2466) <= b and not a;
    layer0_outputs(2467) <= not a or b;
    layer0_outputs(2468) <= not (a or b);
    layer0_outputs(2469) <= not (a or b);
    layer0_outputs(2470) <= b;
    layer0_outputs(2471) <= a and b;
    layer0_outputs(2472) <= b and not a;
    layer0_outputs(2473) <= a and b;
    layer0_outputs(2474) <= b;
    layer0_outputs(2475) <= a and not b;
    layer0_outputs(2476) <= a or b;
    layer0_outputs(2477) <= not (a xor b);
    layer0_outputs(2478) <= a and b;
    layer0_outputs(2479) <= a or b;
    layer0_outputs(2480) <= b and not a;
    layer0_outputs(2481) <= not (a or b);
    layer0_outputs(2482) <= b;
    layer0_outputs(2483) <= not (a or b);
    layer0_outputs(2484) <= not (a and b);
    layer0_outputs(2485) <= not (a xor b);
    layer0_outputs(2486) <= a;
    layer0_outputs(2487) <= b and not a;
    layer0_outputs(2488) <= a;
    layer0_outputs(2489) <= not b or a;
    layer0_outputs(2490) <= b and not a;
    layer0_outputs(2491) <= not (a and b);
    layer0_outputs(2492) <= a xor b;
    layer0_outputs(2493) <= a and b;
    layer0_outputs(2494) <= a or b;
    layer0_outputs(2495) <= a or b;
    layer0_outputs(2496) <= a or b;
    layer0_outputs(2497) <= a and b;
    layer0_outputs(2498) <= not a;
    layer0_outputs(2499) <= a and not b;
    layer0_outputs(2500) <= b;
    layer0_outputs(2501) <= not (a and b);
    layer0_outputs(2502) <= b;
    layer0_outputs(2503) <= a;
    layer0_outputs(2504) <= not a;
    layer0_outputs(2505) <= '1';
    layer0_outputs(2506) <= not (a or b);
    layer0_outputs(2507) <= a or b;
    layer0_outputs(2508) <= not b or a;
    layer0_outputs(2509) <= not a;
    layer0_outputs(2510) <= a;
    layer0_outputs(2511) <= not (a or b);
    layer0_outputs(2512) <= a and b;
    layer0_outputs(2513) <= not b;
    layer0_outputs(2514) <= not b;
    layer0_outputs(2515) <= a or b;
    layer0_outputs(2516) <= not b;
    layer0_outputs(2517) <= b and not a;
    layer0_outputs(2518) <= not (a or b);
    layer0_outputs(2519) <= not a;
    layer0_outputs(2520) <= a;
    layer0_outputs(2521) <= a and not b;
    layer0_outputs(2522) <= b;
    layer0_outputs(2523) <= not b;
    layer0_outputs(2524) <= not (a or b);
    layer0_outputs(2525) <= not a or b;
    layer0_outputs(2526) <= not (a or b);
    layer0_outputs(2527) <= b and not a;
    layer0_outputs(2528) <= not a or b;
    layer0_outputs(2529) <= b;
    layer0_outputs(2530) <= not (a and b);
    layer0_outputs(2531) <= b and not a;
    layer0_outputs(2532) <= not (a or b);
    layer0_outputs(2533) <= b and not a;
    layer0_outputs(2534) <= not a or b;
    layer0_outputs(2535) <= not b or a;
    layer0_outputs(2536) <= not (a xor b);
    layer0_outputs(2537) <= a;
    layer0_outputs(2538) <= a xor b;
    layer0_outputs(2539) <= '0';
    layer0_outputs(2540) <= b and not a;
    layer0_outputs(2541) <= not (a xor b);
    layer0_outputs(2542) <= b and not a;
    layer0_outputs(2543) <= a and not b;
    layer0_outputs(2544) <= a or b;
    layer0_outputs(2545) <= a or b;
    layer0_outputs(2546) <= a or b;
    layer0_outputs(2547) <= a xor b;
    layer0_outputs(2548) <= not b;
    layer0_outputs(2549) <= '0';
    layer0_outputs(2550) <= not a;
    layer0_outputs(2551) <= '1';
    layer0_outputs(2552) <= a xor b;
    layer0_outputs(2553) <= a and not b;
    layer0_outputs(2554) <= not (a or b);
    layer0_outputs(2555) <= not (a or b);
    layer0_outputs(2556) <= not (a or b);
    layer0_outputs(2557) <= not b or a;
    layer0_outputs(2558) <= not (a and b);
    layer0_outputs(2559) <= not (a or b);
    layer0_outputs(2560) <= not (a xor b);
    layer0_outputs(2561) <= not a or b;
    layer0_outputs(2562) <= b;
    layer0_outputs(2563) <= not (a xor b);
    layer0_outputs(2564) <= not (a xor b);
    layer0_outputs(2565) <= not b or a;
    layer0_outputs(2566) <= not (a xor b);
    layer0_outputs(2567) <= a and not b;
    layer0_outputs(2568) <= not b;
    layer0_outputs(2569) <= a and b;
    layer0_outputs(2570) <= a and not b;
    layer0_outputs(2571) <= a;
    layer0_outputs(2572) <= not b;
    layer0_outputs(2573) <= a xor b;
    layer0_outputs(2574) <= a xor b;
    layer0_outputs(2575) <= not (a and b);
    layer0_outputs(2576) <= not (a and b);
    layer0_outputs(2577) <= a and not b;
    layer0_outputs(2578) <= not b or a;
    layer0_outputs(2579) <= not a;
    layer0_outputs(2580) <= b;
    layer0_outputs(2581) <= '0';
    layer0_outputs(2582) <= '0';
    layer0_outputs(2583) <= a;
    layer0_outputs(2584) <= not a or b;
    layer0_outputs(2585) <= b and not a;
    layer0_outputs(2586) <= '0';
    layer0_outputs(2587) <= not b or a;
    layer0_outputs(2588) <= a or b;
    layer0_outputs(2589) <= not a or b;
    layer0_outputs(2590) <= not (a or b);
    layer0_outputs(2591) <= not (a or b);
    layer0_outputs(2592) <= not b;
    layer0_outputs(2593) <= not a;
    layer0_outputs(2594) <= not (a xor b);
    layer0_outputs(2595) <= a;
    layer0_outputs(2596) <= not a;
    layer0_outputs(2597) <= not b;
    layer0_outputs(2598) <= a and b;
    layer0_outputs(2599) <= '1';
    layer0_outputs(2600) <= '1';
    layer0_outputs(2601) <= a and not b;
    layer0_outputs(2602) <= not b;
    layer0_outputs(2603) <= a or b;
    layer0_outputs(2604) <= b;
    layer0_outputs(2605) <= not (a xor b);
    layer0_outputs(2606) <= a and not b;
    layer0_outputs(2607) <= not (a or b);
    layer0_outputs(2608) <= a and not b;
    layer0_outputs(2609) <= a and not b;
    layer0_outputs(2610) <= '0';
    layer0_outputs(2611) <= not a;
    layer0_outputs(2612) <= a or b;
    layer0_outputs(2613) <= a;
    layer0_outputs(2614) <= a and b;
    layer0_outputs(2615) <= not (a or b);
    layer0_outputs(2616) <= '0';
    layer0_outputs(2617) <= '1';
    layer0_outputs(2618) <= b;
    layer0_outputs(2619) <= not (a or b);
    layer0_outputs(2620) <= '1';
    layer0_outputs(2621) <= a or b;
    layer0_outputs(2622) <= b and not a;
    layer0_outputs(2623) <= not a;
    layer0_outputs(2624) <= not a;
    layer0_outputs(2625) <= not a;
    layer0_outputs(2626) <= a or b;
    layer0_outputs(2627) <= a or b;
    layer0_outputs(2628) <= not b or a;
    layer0_outputs(2629) <= a xor b;
    layer0_outputs(2630) <= not (a or b);
    layer0_outputs(2631) <= '1';
    layer0_outputs(2632) <= a xor b;
    layer0_outputs(2633) <= not (a and b);
    layer0_outputs(2634) <= a or b;
    layer0_outputs(2635) <= a xor b;
    layer0_outputs(2636) <= not b or a;
    layer0_outputs(2637) <= not (a or b);
    layer0_outputs(2638) <= not (a and b);
    layer0_outputs(2639) <= a or b;
    layer0_outputs(2640) <= not b or a;
    layer0_outputs(2641) <= a and not b;
    layer0_outputs(2642) <= a and b;
    layer0_outputs(2643) <= '0';
    layer0_outputs(2644) <= not b or a;
    layer0_outputs(2645) <= '1';
    layer0_outputs(2646) <= b;
    layer0_outputs(2647) <= not (a xor b);
    layer0_outputs(2648) <= '1';
    layer0_outputs(2649) <= not b or a;
    layer0_outputs(2650) <= not a or b;
    layer0_outputs(2651) <= a;
    layer0_outputs(2652) <= a and not b;
    layer0_outputs(2653) <= '0';
    layer0_outputs(2654) <= a and not b;
    layer0_outputs(2655) <= a;
    layer0_outputs(2656) <= not (a or b);
    layer0_outputs(2657) <= b;
    layer0_outputs(2658) <= a;
    layer0_outputs(2659) <= not a or b;
    layer0_outputs(2660) <= not (a xor b);
    layer0_outputs(2661) <= b;
    layer0_outputs(2662) <= a;
    layer0_outputs(2663) <= a;
    layer0_outputs(2664) <= not (a and b);
    layer0_outputs(2665) <= not a or b;
    layer0_outputs(2666) <= not a;
    layer0_outputs(2667) <= not b;
    layer0_outputs(2668) <= not (a or b);
    layer0_outputs(2669) <= b;
    layer0_outputs(2670) <= not a;
    layer0_outputs(2671) <= a or b;
    layer0_outputs(2672) <= a and not b;
    layer0_outputs(2673) <= a or b;
    layer0_outputs(2674) <= a and not b;
    layer0_outputs(2675) <= b;
    layer0_outputs(2676) <= not (a or b);
    layer0_outputs(2677) <= not (a xor b);
    layer0_outputs(2678) <= b and not a;
    layer0_outputs(2679) <= not (a xor b);
    layer0_outputs(2680) <= b and not a;
    layer0_outputs(2681) <= a;
    layer0_outputs(2682) <= not a or b;
    layer0_outputs(2683) <= not (a xor b);
    layer0_outputs(2684) <= not (a and b);
    layer0_outputs(2685) <= a xor b;
    layer0_outputs(2686) <= not a;
    layer0_outputs(2687) <= not a;
    layer0_outputs(2688) <= b;
    layer0_outputs(2689) <= '0';
    layer0_outputs(2690) <= not a or b;
    layer0_outputs(2691) <= a and not b;
    layer0_outputs(2692) <= not (a or b);
    layer0_outputs(2693) <= b and not a;
    layer0_outputs(2694) <= '1';
    layer0_outputs(2695) <= not a or b;
    layer0_outputs(2696) <= not (a xor b);
    layer0_outputs(2697) <= not b or a;
    layer0_outputs(2698) <= '0';
    layer0_outputs(2699) <= not a;
    layer0_outputs(2700) <= a and b;
    layer0_outputs(2701) <= not b;
    layer0_outputs(2702) <= not a;
    layer0_outputs(2703) <= not (a xor b);
    layer0_outputs(2704) <= '0';
    layer0_outputs(2705) <= a and not b;
    layer0_outputs(2706) <= not b;
    layer0_outputs(2707) <= not a or b;
    layer0_outputs(2708) <= not b;
    layer0_outputs(2709) <= not b or a;
    layer0_outputs(2710) <= not a;
    layer0_outputs(2711) <= a and b;
    layer0_outputs(2712) <= a and b;
    layer0_outputs(2713) <= b and not a;
    layer0_outputs(2714) <= a and b;
    layer0_outputs(2715) <= '1';
    layer0_outputs(2716) <= not (a or b);
    layer0_outputs(2717) <= b and not a;
    layer0_outputs(2718) <= not b;
    layer0_outputs(2719) <= b;
    layer0_outputs(2720) <= not b or a;
    layer0_outputs(2721) <= a or b;
    layer0_outputs(2722) <= not (a or b);
    layer0_outputs(2723) <= not b;
    layer0_outputs(2724) <= a and not b;
    layer0_outputs(2725) <= not a or b;
    layer0_outputs(2726) <= not (a or b);
    layer0_outputs(2727) <= b;
    layer0_outputs(2728) <= a;
    layer0_outputs(2729) <= not (a and b);
    layer0_outputs(2730) <= not b or a;
    layer0_outputs(2731) <= '1';
    layer0_outputs(2732) <= '0';
    layer0_outputs(2733) <= not a or b;
    layer0_outputs(2734) <= not a or b;
    layer0_outputs(2735) <= a xor b;
    layer0_outputs(2736) <= not b or a;
    layer0_outputs(2737) <= '1';
    layer0_outputs(2738) <= not b;
    layer0_outputs(2739) <= not b;
    layer0_outputs(2740) <= not (a or b);
    layer0_outputs(2741) <= not (a or b);
    layer0_outputs(2742) <= a and b;
    layer0_outputs(2743) <= not b or a;
    layer0_outputs(2744) <= a;
    layer0_outputs(2745) <= a;
    layer0_outputs(2746) <= a and not b;
    layer0_outputs(2747) <= a;
    layer0_outputs(2748) <= a and not b;
    layer0_outputs(2749) <= '0';
    layer0_outputs(2750) <= not b or a;
    layer0_outputs(2751) <= not (a or b);
    layer0_outputs(2752) <= b and not a;
    layer0_outputs(2753) <= not a or b;
    layer0_outputs(2754) <= a;
    layer0_outputs(2755) <= not (a or b);
    layer0_outputs(2756) <= not a;
    layer0_outputs(2757) <= not a or b;
    layer0_outputs(2758) <= not b;
    layer0_outputs(2759) <= not (a and b);
    layer0_outputs(2760) <= not b or a;
    layer0_outputs(2761) <= a and not b;
    layer0_outputs(2762) <= a or b;
    layer0_outputs(2763) <= '0';
    layer0_outputs(2764) <= not (a and b);
    layer0_outputs(2765) <= not (a or b);
    layer0_outputs(2766) <= not b or a;
    layer0_outputs(2767) <= not b or a;
    layer0_outputs(2768) <= a and b;
    layer0_outputs(2769) <= a or b;
    layer0_outputs(2770) <= a;
    layer0_outputs(2771) <= '0';
    layer0_outputs(2772) <= not a or b;
    layer0_outputs(2773) <= not (a xor b);
    layer0_outputs(2774) <= not a or b;
    layer0_outputs(2775) <= not (a xor b);
    layer0_outputs(2776) <= b;
    layer0_outputs(2777) <= '0';
    layer0_outputs(2778) <= not a;
    layer0_outputs(2779) <= a;
    layer0_outputs(2780) <= b;
    layer0_outputs(2781) <= '0';
    layer0_outputs(2782) <= b and not a;
    layer0_outputs(2783) <= not b or a;
    layer0_outputs(2784) <= not (a and b);
    layer0_outputs(2785) <= b;
    layer0_outputs(2786) <= a and not b;
    layer0_outputs(2787) <= not (a or b);
    layer0_outputs(2788) <= b;
    layer0_outputs(2789) <= not b;
    layer0_outputs(2790) <= not a or b;
    layer0_outputs(2791) <= '1';
    layer0_outputs(2792) <= a or b;
    layer0_outputs(2793) <= '0';
    layer0_outputs(2794) <= a or b;
    layer0_outputs(2795) <= a xor b;
    layer0_outputs(2796) <= not b or a;
    layer0_outputs(2797) <= a or b;
    layer0_outputs(2798) <= a or b;
    layer0_outputs(2799) <= not b;
    layer0_outputs(2800) <= b and not a;
    layer0_outputs(2801) <= not b or a;
    layer0_outputs(2802) <= not b;
    layer0_outputs(2803) <= a;
    layer0_outputs(2804) <= b;
    layer0_outputs(2805) <= b;
    layer0_outputs(2806) <= b;
    layer0_outputs(2807) <= '0';
    layer0_outputs(2808) <= b;
    layer0_outputs(2809) <= a;
    layer0_outputs(2810) <= '1';
    layer0_outputs(2811) <= not (a or b);
    layer0_outputs(2812) <= not a;
    layer0_outputs(2813) <= not (a xor b);
    layer0_outputs(2814) <= not b or a;
    layer0_outputs(2815) <= '0';
    layer0_outputs(2816) <= not a or b;
    layer0_outputs(2817) <= a;
    layer0_outputs(2818) <= a and not b;
    layer0_outputs(2819) <= not (a xor b);
    layer0_outputs(2820) <= not b;
    layer0_outputs(2821) <= not (a or b);
    layer0_outputs(2822) <= a and not b;
    layer0_outputs(2823) <= not b or a;
    layer0_outputs(2824) <= '0';
    layer0_outputs(2825) <= not (a xor b);
    layer0_outputs(2826) <= a and not b;
    layer0_outputs(2827) <= a xor b;
    layer0_outputs(2828) <= a and not b;
    layer0_outputs(2829) <= a or b;
    layer0_outputs(2830) <= a;
    layer0_outputs(2831) <= '0';
    layer0_outputs(2832) <= b and not a;
    layer0_outputs(2833) <= not a or b;
    layer0_outputs(2834) <= a xor b;
    layer0_outputs(2835) <= not (a xor b);
    layer0_outputs(2836) <= not b;
    layer0_outputs(2837) <= not (a xor b);
    layer0_outputs(2838) <= '1';
    layer0_outputs(2839) <= b;
    layer0_outputs(2840) <= '0';
    layer0_outputs(2841) <= '0';
    layer0_outputs(2842) <= b;
    layer0_outputs(2843) <= '1';
    layer0_outputs(2844) <= a;
    layer0_outputs(2845) <= not (a and b);
    layer0_outputs(2846) <= not b;
    layer0_outputs(2847) <= not b;
    layer0_outputs(2848) <= not b or a;
    layer0_outputs(2849) <= a xor b;
    layer0_outputs(2850) <= a and b;
    layer0_outputs(2851) <= a;
    layer0_outputs(2852) <= not a;
    layer0_outputs(2853) <= not (a or b);
    layer0_outputs(2854) <= a and b;
    layer0_outputs(2855) <= a and not b;
    layer0_outputs(2856) <= b;
    layer0_outputs(2857) <= a;
    layer0_outputs(2858) <= not b;
    layer0_outputs(2859) <= b;
    layer0_outputs(2860) <= '0';
    layer0_outputs(2861) <= not b;
    layer0_outputs(2862) <= a and b;
    layer0_outputs(2863) <= b;
    layer0_outputs(2864) <= a or b;
    layer0_outputs(2865) <= '0';
    layer0_outputs(2866) <= a and not b;
    layer0_outputs(2867) <= a or b;
    layer0_outputs(2868) <= a and b;
    layer0_outputs(2869) <= a and b;
    layer0_outputs(2870) <= not (a xor b);
    layer0_outputs(2871) <= '0';
    layer0_outputs(2872) <= '0';
    layer0_outputs(2873) <= a;
    layer0_outputs(2874) <= not (a xor b);
    layer0_outputs(2875) <= b and not a;
    layer0_outputs(2876) <= a and not b;
    layer0_outputs(2877) <= a xor b;
    layer0_outputs(2878) <= not b;
    layer0_outputs(2879) <= not (a xor b);
    layer0_outputs(2880) <= a or b;
    layer0_outputs(2881) <= not a or b;
    layer0_outputs(2882) <= a or b;
    layer0_outputs(2883) <= a or b;
    layer0_outputs(2884) <= not b or a;
    layer0_outputs(2885) <= not a;
    layer0_outputs(2886) <= not (a or b);
    layer0_outputs(2887) <= not b or a;
    layer0_outputs(2888) <= a or b;
    layer0_outputs(2889) <= not a or b;
    layer0_outputs(2890) <= a;
    layer0_outputs(2891) <= not (a xor b);
    layer0_outputs(2892) <= a;
    layer0_outputs(2893) <= b;
    layer0_outputs(2894) <= a or b;
    layer0_outputs(2895) <= '1';
    layer0_outputs(2896) <= not b;
    layer0_outputs(2897) <= b;
    layer0_outputs(2898) <= not b;
    layer0_outputs(2899) <= '1';
    layer0_outputs(2900) <= a or b;
    layer0_outputs(2901) <= a xor b;
    layer0_outputs(2902) <= not a or b;
    layer0_outputs(2903) <= not b or a;
    layer0_outputs(2904) <= '1';
    layer0_outputs(2905) <= not (a xor b);
    layer0_outputs(2906) <= not b;
    layer0_outputs(2907) <= b;
    layer0_outputs(2908) <= a or b;
    layer0_outputs(2909) <= not a;
    layer0_outputs(2910) <= not b;
    layer0_outputs(2911) <= not a or b;
    layer0_outputs(2912) <= a xor b;
    layer0_outputs(2913) <= not (a xor b);
    layer0_outputs(2914) <= not b;
    layer0_outputs(2915) <= not a or b;
    layer0_outputs(2916) <= not b or a;
    layer0_outputs(2917) <= not b or a;
    layer0_outputs(2918) <= a or b;
    layer0_outputs(2919) <= '0';
    layer0_outputs(2920) <= not (a xor b);
    layer0_outputs(2921) <= '1';
    layer0_outputs(2922) <= not (a and b);
    layer0_outputs(2923) <= not b or a;
    layer0_outputs(2924) <= a and b;
    layer0_outputs(2925) <= a xor b;
    layer0_outputs(2926) <= '1';
    layer0_outputs(2927) <= b and not a;
    layer0_outputs(2928) <= a;
    layer0_outputs(2929) <= a or b;
    layer0_outputs(2930) <= a and not b;
    layer0_outputs(2931) <= not a;
    layer0_outputs(2932) <= '0';
    layer0_outputs(2933) <= b;
    layer0_outputs(2934) <= a;
    layer0_outputs(2935) <= not a or b;
    layer0_outputs(2936) <= '1';
    layer0_outputs(2937) <= b and not a;
    layer0_outputs(2938) <= a or b;
    layer0_outputs(2939) <= b and not a;
    layer0_outputs(2940) <= a and not b;
    layer0_outputs(2941) <= a xor b;
    layer0_outputs(2942) <= '0';
    layer0_outputs(2943) <= '1';
    layer0_outputs(2944) <= not b or a;
    layer0_outputs(2945) <= b;
    layer0_outputs(2946) <= a xor b;
    layer0_outputs(2947) <= not (a xor b);
    layer0_outputs(2948) <= a xor b;
    layer0_outputs(2949) <= not b;
    layer0_outputs(2950) <= '0';
    layer0_outputs(2951) <= not a;
    layer0_outputs(2952) <= not b or a;
    layer0_outputs(2953) <= '1';
    layer0_outputs(2954) <= b and not a;
    layer0_outputs(2955) <= a;
    layer0_outputs(2956) <= not (a or b);
    layer0_outputs(2957) <= not a;
    layer0_outputs(2958) <= not a;
    layer0_outputs(2959) <= a and b;
    layer0_outputs(2960) <= not a or b;
    layer0_outputs(2961) <= '0';
    layer0_outputs(2962) <= not b or a;
    layer0_outputs(2963) <= '1';
    layer0_outputs(2964) <= not b;
    layer0_outputs(2965) <= b;
    layer0_outputs(2966) <= a;
    layer0_outputs(2967) <= not (a xor b);
    layer0_outputs(2968) <= b;
    layer0_outputs(2969) <= not b;
    layer0_outputs(2970) <= not (a and b);
    layer0_outputs(2971) <= '1';
    layer0_outputs(2972) <= not a or b;
    layer0_outputs(2973) <= not (a xor b);
    layer0_outputs(2974) <= not a or b;
    layer0_outputs(2975) <= not a;
    layer0_outputs(2976) <= a xor b;
    layer0_outputs(2977) <= b;
    layer0_outputs(2978) <= not a;
    layer0_outputs(2979) <= not (a xor b);
    layer0_outputs(2980) <= a and b;
    layer0_outputs(2981) <= a;
    layer0_outputs(2982) <= not (a or b);
    layer0_outputs(2983) <= not a;
    layer0_outputs(2984) <= '0';
    layer0_outputs(2985) <= not (a or b);
    layer0_outputs(2986) <= a and b;
    layer0_outputs(2987) <= b;
    layer0_outputs(2988) <= not (a or b);
    layer0_outputs(2989) <= '0';
    layer0_outputs(2990) <= a or b;
    layer0_outputs(2991) <= not (a xor b);
    layer0_outputs(2992) <= not (a xor b);
    layer0_outputs(2993) <= a xor b;
    layer0_outputs(2994) <= b;
    layer0_outputs(2995) <= a xor b;
    layer0_outputs(2996) <= not b;
    layer0_outputs(2997) <= not a or b;
    layer0_outputs(2998) <= not (a or b);
    layer0_outputs(2999) <= b;
    layer0_outputs(3000) <= not b or a;
    layer0_outputs(3001) <= not b;
    layer0_outputs(3002) <= '1';
    layer0_outputs(3003) <= a xor b;
    layer0_outputs(3004) <= not (a xor b);
    layer0_outputs(3005) <= not b;
    layer0_outputs(3006) <= b and not a;
    layer0_outputs(3007) <= not (a or b);
    layer0_outputs(3008) <= a and b;
    layer0_outputs(3009) <= b;
    layer0_outputs(3010) <= '0';
    layer0_outputs(3011) <= a;
    layer0_outputs(3012) <= not (a xor b);
    layer0_outputs(3013) <= a or b;
    layer0_outputs(3014) <= a and not b;
    layer0_outputs(3015) <= a;
    layer0_outputs(3016) <= '1';
    layer0_outputs(3017) <= not (a xor b);
    layer0_outputs(3018) <= not a;
    layer0_outputs(3019) <= not (a xor b);
    layer0_outputs(3020) <= not a;
    layer0_outputs(3021) <= a or b;
    layer0_outputs(3022) <= a xor b;
    layer0_outputs(3023) <= a xor b;
    layer0_outputs(3024) <= a and not b;
    layer0_outputs(3025) <= b;
    layer0_outputs(3026) <= a;
    layer0_outputs(3027) <= a and b;
    layer0_outputs(3028) <= not a or b;
    layer0_outputs(3029) <= a;
    layer0_outputs(3030) <= not a or b;
    layer0_outputs(3031) <= not a;
    layer0_outputs(3032) <= b;
    layer0_outputs(3033) <= a and b;
    layer0_outputs(3034) <= a and not b;
    layer0_outputs(3035) <= not a or b;
    layer0_outputs(3036) <= not b;
    layer0_outputs(3037) <= not (a or b);
    layer0_outputs(3038) <= a xor b;
    layer0_outputs(3039) <= not (a or b);
    layer0_outputs(3040) <= a;
    layer0_outputs(3041) <= not b;
    layer0_outputs(3042) <= a and not b;
    layer0_outputs(3043) <= a;
    layer0_outputs(3044) <= '1';
    layer0_outputs(3045) <= '0';
    layer0_outputs(3046) <= '0';
    layer0_outputs(3047) <= not (a or b);
    layer0_outputs(3048) <= not b or a;
    layer0_outputs(3049) <= not (a or b);
    layer0_outputs(3050) <= not a or b;
    layer0_outputs(3051) <= b;
    layer0_outputs(3052) <= not b;
    layer0_outputs(3053) <= not b or a;
    layer0_outputs(3054) <= not b or a;
    layer0_outputs(3055) <= not a;
    layer0_outputs(3056) <= not (a and b);
    layer0_outputs(3057) <= '1';
    layer0_outputs(3058) <= not b or a;
    layer0_outputs(3059) <= a or b;
    layer0_outputs(3060) <= a and b;
    layer0_outputs(3061) <= b and not a;
    layer0_outputs(3062) <= a;
    layer0_outputs(3063) <= '1';
    layer0_outputs(3064) <= not a;
    layer0_outputs(3065) <= b;
    layer0_outputs(3066) <= '1';
    layer0_outputs(3067) <= a;
    layer0_outputs(3068) <= '1';
    layer0_outputs(3069) <= b and not a;
    layer0_outputs(3070) <= not b;
    layer0_outputs(3071) <= not (a or b);
    layer0_outputs(3072) <= a;
    layer0_outputs(3073) <= not b;
    layer0_outputs(3074) <= not b;
    layer0_outputs(3075) <= not (a xor b);
    layer0_outputs(3076) <= not b or a;
    layer0_outputs(3077) <= a or b;
    layer0_outputs(3078) <= a;
    layer0_outputs(3079) <= not b or a;
    layer0_outputs(3080) <= not (a and b);
    layer0_outputs(3081) <= not b;
    layer0_outputs(3082) <= b and not a;
    layer0_outputs(3083) <= not (a or b);
    layer0_outputs(3084) <= a or b;
    layer0_outputs(3085) <= b;
    layer0_outputs(3086) <= a;
    layer0_outputs(3087) <= a and b;
    layer0_outputs(3088) <= b and not a;
    layer0_outputs(3089) <= not b or a;
    layer0_outputs(3090) <= a and b;
    layer0_outputs(3091) <= not (a or b);
    layer0_outputs(3092) <= a and not b;
    layer0_outputs(3093) <= a and b;
    layer0_outputs(3094) <= b and not a;
    layer0_outputs(3095) <= a or b;
    layer0_outputs(3096) <= not b;
    layer0_outputs(3097) <= b and not a;
    layer0_outputs(3098) <= a and not b;
    layer0_outputs(3099) <= not b;
    layer0_outputs(3100) <= a and not b;
    layer0_outputs(3101) <= a and b;
    layer0_outputs(3102) <= b and not a;
    layer0_outputs(3103) <= not b;
    layer0_outputs(3104) <= b and not a;
    layer0_outputs(3105) <= a and b;
    layer0_outputs(3106) <= not b or a;
    layer0_outputs(3107) <= a or b;
    layer0_outputs(3108) <= a xor b;
    layer0_outputs(3109) <= a or b;
    layer0_outputs(3110) <= a and not b;
    layer0_outputs(3111) <= not a;
    layer0_outputs(3112) <= a;
    layer0_outputs(3113) <= a;
    layer0_outputs(3114) <= a or b;
    layer0_outputs(3115) <= not a;
    layer0_outputs(3116) <= a;
    layer0_outputs(3117) <= '1';
    layer0_outputs(3118) <= a and b;
    layer0_outputs(3119) <= not (a or b);
    layer0_outputs(3120) <= not b;
    layer0_outputs(3121) <= b and not a;
    layer0_outputs(3122) <= b;
    layer0_outputs(3123) <= b;
    layer0_outputs(3124) <= not b;
    layer0_outputs(3125) <= not a;
    layer0_outputs(3126) <= not b;
    layer0_outputs(3127) <= not (a xor b);
    layer0_outputs(3128) <= b and not a;
    layer0_outputs(3129) <= a xor b;
    layer0_outputs(3130) <= a;
    layer0_outputs(3131) <= a;
    layer0_outputs(3132) <= b;
    layer0_outputs(3133) <= a;
    layer0_outputs(3134) <= not (a and b);
    layer0_outputs(3135) <= not a or b;
    layer0_outputs(3136) <= not a or b;
    layer0_outputs(3137) <= not a;
    layer0_outputs(3138) <= a and not b;
    layer0_outputs(3139) <= b;
    layer0_outputs(3140) <= a xor b;
    layer0_outputs(3141) <= b;
    layer0_outputs(3142) <= a xor b;
    layer0_outputs(3143) <= not (a or b);
    layer0_outputs(3144) <= not b or a;
    layer0_outputs(3145) <= not (a or b);
    layer0_outputs(3146) <= a and not b;
    layer0_outputs(3147) <= a or b;
    layer0_outputs(3148) <= a and b;
    layer0_outputs(3149) <= a and b;
    layer0_outputs(3150) <= not b or a;
    layer0_outputs(3151) <= b;
    layer0_outputs(3152) <= a and b;
    layer0_outputs(3153) <= a and not b;
    layer0_outputs(3154) <= not a;
    layer0_outputs(3155) <= '1';
    layer0_outputs(3156) <= not a or b;
    layer0_outputs(3157) <= not b or a;
    layer0_outputs(3158) <= not a;
    layer0_outputs(3159) <= b;
    layer0_outputs(3160) <= not b or a;
    layer0_outputs(3161) <= not b or a;
    layer0_outputs(3162) <= not b;
    layer0_outputs(3163) <= not (a and b);
    layer0_outputs(3164) <= b and not a;
    layer0_outputs(3165) <= a xor b;
    layer0_outputs(3166) <= a or b;
    layer0_outputs(3167) <= not (a xor b);
    layer0_outputs(3168) <= not (a xor b);
    layer0_outputs(3169) <= not (a or b);
    layer0_outputs(3170) <= b;
    layer0_outputs(3171) <= a xor b;
    layer0_outputs(3172) <= not b or a;
    layer0_outputs(3173) <= not a or b;
    layer0_outputs(3174) <= b;
    layer0_outputs(3175) <= not b;
    layer0_outputs(3176) <= b;
    layer0_outputs(3177) <= not (a xor b);
    layer0_outputs(3178) <= a;
    layer0_outputs(3179) <= a or b;
    layer0_outputs(3180) <= not b or a;
    layer0_outputs(3181) <= b and not a;
    layer0_outputs(3182) <= not a;
    layer0_outputs(3183) <= not (a or b);
    layer0_outputs(3184) <= not a or b;
    layer0_outputs(3185) <= not b or a;
    layer0_outputs(3186) <= not (a and b);
    layer0_outputs(3187) <= not (a or b);
    layer0_outputs(3188) <= not a or b;
    layer0_outputs(3189) <= not b;
    layer0_outputs(3190) <= a xor b;
    layer0_outputs(3191) <= not (a or b);
    layer0_outputs(3192) <= a or b;
    layer0_outputs(3193) <= not (a xor b);
    layer0_outputs(3194) <= '0';
    layer0_outputs(3195) <= a and not b;
    layer0_outputs(3196) <= a and b;
    layer0_outputs(3197) <= a and b;
    layer0_outputs(3198) <= not b or a;
    layer0_outputs(3199) <= not (a and b);
    layer0_outputs(3200) <= a and b;
    layer0_outputs(3201) <= a or b;
    layer0_outputs(3202) <= not (a or b);
    layer0_outputs(3203) <= not (a or b);
    layer0_outputs(3204) <= a and not b;
    layer0_outputs(3205) <= '0';
    layer0_outputs(3206) <= b and not a;
    layer0_outputs(3207) <= '1';
    layer0_outputs(3208) <= not (a xor b);
    layer0_outputs(3209) <= a and not b;
    layer0_outputs(3210) <= not a or b;
    layer0_outputs(3211) <= a and not b;
    layer0_outputs(3212) <= '1';
    layer0_outputs(3213) <= a or b;
    layer0_outputs(3214) <= not b or a;
    layer0_outputs(3215) <= not b or a;
    layer0_outputs(3216) <= b and not a;
    layer0_outputs(3217) <= not b;
    layer0_outputs(3218) <= not a or b;
    layer0_outputs(3219) <= a or b;
    layer0_outputs(3220) <= not a;
    layer0_outputs(3221) <= not (a and b);
    layer0_outputs(3222) <= not b;
    layer0_outputs(3223) <= not b or a;
    layer0_outputs(3224) <= not a or b;
    layer0_outputs(3225) <= not (a xor b);
    layer0_outputs(3226) <= not b or a;
    layer0_outputs(3227) <= a;
    layer0_outputs(3228) <= not a or b;
    layer0_outputs(3229) <= not b;
    layer0_outputs(3230) <= not b;
    layer0_outputs(3231) <= a and b;
    layer0_outputs(3232) <= not b or a;
    layer0_outputs(3233) <= a;
    layer0_outputs(3234) <= a xor b;
    layer0_outputs(3235) <= not (a or b);
    layer0_outputs(3236) <= not a or b;
    layer0_outputs(3237) <= not (a and b);
    layer0_outputs(3238) <= b;
    layer0_outputs(3239) <= a and b;
    layer0_outputs(3240) <= b;
    layer0_outputs(3241) <= not b;
    layer0_outputs(3242) <= '1';
    layer0_outputs(3243) <= not (a or b);
    layer0_outputs(3244) <= a;
    layer0_outputs(3245) <= a;
    layer0_outputs(3246) <= not (a or b);
    layer0_outputs(3247) <= b and not a;
    layer0_outputs(3248) <= a;
    layer0_outputs(3249) <= '0';
    layer0_outputs(3250) <= not (a or b);
    layer0_outputs(3251) <= a;
    layer0_outputs(3252) <= a and b;
    layer0_outputs(3253) <= a xor b;
    layer0_outputs(3254) <= a xor b;
    layer0_outputs(3255) <= a xor b;
    layer0_outputs(3256) <= a or b;
    layer0_outputs(3257) <= not (a and b);
    layer0_outputs(3258) <= a or b;
    layer0_outputs(3259) <= not (a xor b);
    layer0_outputs(3260) <= a and b;
    layer0_outputs(3261) <= not a or b;
    layer0_outputs(3262) <= a and b;
    layer0_outputs(3263) <= not a or b;
    layer0_outputs(3264) <= b;
    layer0_outputs(3265) <= '1';
    layer0_outputs(3266) <= b;
    layer0_outputs(3267) <= a or b;
    layer0_outputs(3268) <= '1';
    layer0_outputs(3269) <= not (a xor b);
    layer0_outputs(3270) <= not (a or b);
    layer0_outputs(3271) <= not (a or b);
    layer0_outputs(3272) <= a;
    layer0_outputs(3273) <= not b;
    layer0_outputs(3274) <= not b or a;
    layer0_outputs(3275) <= not a;
    layer0_outputs(3276) <= not b;
    layer0_outputs(3277) <= a;
    layer0_outputs(3278) <= not b or a;
    layer0_outputs(3279) <= not b;
    layer0_outputs(3280) <= not b or a;
    layer0_outputs(3281) <= not a;
    layer0_outputs(3282) <= not a;
    layer0_outputs(3283) <= not (a xor b);
    layer0_outputs(3284) <= a and b;
    layer0_outputs(3285) <= a and not b;
    layer0_outputs(3286) <= a;
    layer0_outputs(3287) <= not b;
    layer0_outputs(3288) <= a;
    layer0_outputs(3289) <= not b;
    layer0_outputs(3290) <= not a;
    layer0_outputs(3291) <= not (a or b);
    layer0_outputs(3292) <= a or b;
    layer0_outputs(3293) <= a and b;
    layer0_outputs(3294) <= a and b;
    layer0_outputs(3295) <= a and b;
    layer0_outputs(3296) <= '1';
    layer0_outputs(3297) <= '0';
    layer0_outputs(3298) <= a and b;
    layer0_outputs(3299) <= a and not b;
    layer0_outputs(3300) <= not a;
    layer0_outputs(3301) <= not (a or b);
    layer0_outputs(3302) <= not b or a;
    layer0_outputs(3303) <= not a;
    layer0_outputs(3304) <= '1';
    layer0_outputs(3305) <= not b;
    layer0_outputs(3306) <= not b;
    layer0_outputs(3307) <= not b;
    layer0_outputs(3308) <= '1';
    layer0_outputs(3309) <= a or b;
    layer0_outputs(3310) <= b;
    layer0_outputs(3311) <= not (a or b);
    layer0_outputs(3312) <= not a;
    layer0_outputs(3313) <= not (a xor b);
    layer0_outputs(3314) <= a;
    layer0_outputs(3315) <= not (a or b);
    layer0_outputs(3316) <= not a;
    layer0_outputs(3317) <= not b;
    layer0_outputs(3318) <= a or b;
    layer0_outputs(3319) <= a xor b;
    layer0_outputs(3320) <= not b or a;
    layer0_outputs(3321) <= not a;
    layer0_outputs(3322) <= '0';
    layer0_outputs(3323) <= a;
    layer0_outputs(3324) <= not b or a;
    layer0_outputs(3325) <= not (a or b);
    layer0_outputs(3326) <= not a;
    layer0_outputs(3327) <= not (a or b);
    layer0_outputs(3328) <= '1';
    layer0_outputs(3329) <= not a or b;
    layer0_outputs(3330) <= b;
    layer0_outputs(3331) <= '1';
    layer0_outputs(3332) <= not a or b;
    layer0_outputs(3333) <= a;
    layer0_outputs(3334) <= not (a xor b);
    layer0_outputs(3335) <= not (a and b);
    layer0_outputs(3336) <= a or b;
    layer0_outputs(3337) <= b;
    layer0_outputs(3338) <= not (a xor b);
    layer0_outputs(3339) <= a and b;
    layer0_outputs(3340) <= not (a or b);
    layer0_outputs(3341) <= b and not a;
    layer0_outputs(3342) <= a;
    layer0_outputs(3343) <= not (a or b);
    layer0_outputs(3344) <= a xor b;
    layer0_outputs(3345) <= not b or a;
    layer0_outputs(3346) <= a and not b;
    layer0_outputs(3347) <= a xor b;
    layer0_outputs(3348) <= not b or a;
    layer0_outputs(3349) <= not (a or b);
    layer0_outputs(3350) <= a and b;
    layer0_outputs(3351) <= not a or b;
    layer0_outputs(3352) <= b and not a;
    layer0_outputs(3353) <= not (a and b);
    layer0_outputs(3354) <= not (a and b);
    layer0_outputs(3355) <= not b;
    layer0_outputs(3356) <= a or b;
    layer0_outputs(3357) <= b and not a;
    layer0_outputs(3358) <= '0';
    layer0_outputs(3359) <= '0';
    layer0_outputs(3360) <= not (a xor b);
    layer0_outputs(3361) <= a and b;
    layer0_outputs(3362) <= '1';
    layer0_outputs(3363) <= a xor b;
    layer0_outputs(3364) <= a;
    layer0_outputs(3365) <= '1';
    layer0_outputs(3366) <= a and not b;
    layer0_outputs(3367) <= '1';
    layer0_outputs(3368) <= '1';
    layer0_outputs(3369) <= not (a xor b);
    layer0_outputs(3370) <= not a;
    layer0_outputs(3371) <= not (a or b);
    layer0_outputs(3372) <= a;
    layer0_outputs(3373) <= '1';
    layer0_outputs(3374) <= not b or a;
    layer0_outputs(3375) <= a and b;
    layer0_outputs(3376) <= not (a or b);
    layer0_outputs(3377) <= '0';
    layer0_outputs(3378) <= not a;
    layer0_outputs(3379) <= a or b;
    layer0_outputs(3380) <= b;
    layer0_outputs(3381) <= not b;
    layer0_outputs(3382) <= a or b;
    layer0_outputs(3383) <= b;
    layer0_outputs(3384) <= a or b;
    layer0_outputs(3385) <= '0';
    layer0_outputs(3386) <= not a;
    layer0_outputs(3387) <= not b;
    layer0_outputs(3388) <= a and not b;
    layer0_outputs(3389) <= not b or a;
    layer0_outputs(3390) <= not b;
    layer0_outputs(3391) <= a and b;
    layer0_outputs(3392) <= a and not b;
    layer0_outputs(3393) <= '1';
    layer0_outputs(3394) <= a or b;
    layer0_outputs(3395) <= not b or a;
    layer0_outputs(3396) <= a and not b;
    layer0_outputs(3397) <= a and not b;
    layer0_outputs(3398) <= a;
    layer0_outputs(3399) <= a and not b;
    layer0_outputs(3400) <= not (a xor b);
    layer0_outputs(3401) <= not (a xor b);
    layer0_outputs(3402) <= not (a and b);
    layer0_outputs(3403) <= a and not b;
    layer0_outputs(3404) <= not a;
    layer0_outputs(3405) <= not b;
    layer0_outputs(3406) <= b and not a;
    layer0_outputs(3407) <= not a or b;
    layer0_outputs(3408) <= not a;
    layer0_outputs(3409) <= not b or a;
    layer0_outputs(3410) <= a and b;
    layer0_outputs(3411) <= a or b;
    layer0_outputs(3412) <= a;
    layer0_outputs(3413) <= a xor b;
    layer0_outputs(3414) <= '0';
    layer0_outputs(3415) <= '1';
    layer0_outputs(3416) <= a;
    layer0_outputs(3417) <= not a or b;
    layer0_outputs(3418) <= not (a or b);
    layer0_outputs(3419) <= not b;
    layer0_outputs(3420) <= not b;
    layer0_outputs(3421) <= b;
    layer0_outputs(3422) <= '0';
    layer0_outputs(3423) <= a;
    layer0_outputs(3424) <= not b;
    layer0_outputs(3425) <= not b or a;
    layer0_outputs(3426) <= a xor b;
    layer0_outputs(3427) <= a;
    layer0_outputs(3428) <= a xor b;
    layer0_outputs(3429) <= not b or a;
    layer0_outputs(3430) <= not b or a;
    layer0_outputs(3431) <= not a;
    layer0_outputs(3432) <= b;
    layer0_outputs(3433) <= not (a or b);
    layer0_outputs(3434) <= not (a or b);
    layer0_outputs(3435) <= not b or a;
    layer0_outputs(3436) <= not a or b;
    layer0_outputs(3437) <= not a or b;
    layer0_outputs(3438) <= a xor b;
    layer0_outputs(3439) <= a;
    layer0_outputs(3440) <= a xor b;
    layer0_outputs(3441) <= a xor b;
    layer0_outputs(3442) <= not a;
    layer0_outputs(3443) <= not (a or b);
    layer0_outputs(3444) <= a xor b;
    layer0_outputs(3445) <= b and not a;
    layer0_outputs(3446) <= a and not b;
    layer0_outputs(3447) <= not b;
    layer0_outputs(3448) <= not a or b;
    layer0_outputs(3449) <= a and not b;
    layer0_outputs(3450) <= a or b;
    layer0_outputs(3451) <= b and not a;
    layer0_outputs(3452) <= not (a or b);
    layer0_outputs(3453) <= a;
    layer0_outputs(3454) <= '0';
    layer0_outputs(3455) <= b;
    layer0_outputs(3456) <= not (a or b);
    layer0_outputs(3457) <= b and not a;
    layer0_outputs(3458) <= a or b;
    layer0_outputs(3459) <= a;
    layer0_outputs(3460) <= not (a and b);
    layer0_outputs(3461) <= b and not a;
    layer0_outputs(3462) <= a or b;
    layer0_outputs(3463) <= not a;
    layer0_outputs(3464) <= '1';
    layer0_outputs(3465) <= not (a or b);
    layer0_outputs(3466) <= not a or b;
    layer0_outputs(3467) <= not (a or b);
    layer0_outputs(3468) <= not a or b;
    layer0_outputs(3469) <= a;
    layer0_outputs(3470) <= not (a or b);
    layer0_outputs(3471) <= a xor b;
    layer0_outputs(3472) <= not (a and b);
    layer0_outputs(3473) <= '1';
    layer0_outputs(3474) <= b;
    layer0_outputs(3475) <= not a or b;
    layer0_outputs(3476) <= a xor b;
    layer0_outputs(3477) <= not a;
    layer0_outputs(3478) <= b and not a;
    layer0_outputs(3479) <= a and b;
    layer0_outputs(3480) <= not a;
    layer0_outputs(3481) <= b and not a;
    layer0_outputs(3482) <= not b or a;
    layer0_outputs(3483) <= not b;
    layer0_outputs(3484) <= not b;
    layer0_outputs(3485) <= a xor b;
    layer0_outputs(3486) <= not a;
    layer0_outputs(3487) <= not a or b;
    layer0_outputs(3488) <= '0';
    layer0_outputs(3489) <= a;
    layer0_outputs(3490) <= not b;
    layer0_outputs(3491) <= not a;
    layer0_outputs(3492) <= a;
    layer0_outputs(3493) <= a or b;
    layer0_outputs(3494) <= not (a xor b);
    layer0_outputs(3495) <= a xor b;
    layer0_outputs(3496) <= not a or b;
    layer0_outputs(3497) <= not b or a;
    layer0_outputs(3498) <= not b or a;
    layer0_outputs(3499) <= not (a and b);
    layer0_outputs(3500) <= not (a xor b);
    layer0_outputs(3501) <= a;
    layer0_outputs(3502) <= not (a or b);
    layer0_outputs(3503) <= '1';
    layer0_outputs(3504) <= '0';
    layer0_outputs(3505) <= a;
    layer0_outputs(3506) <= not (a or b);
    layer0_outputs(3507) <= a and not b;
    layer0_outputs(3508) <= not a;
    layer0_outputs(3509) <= b and not a;
    layer0_outputs(3510) <= '1';
    layer0_outputs(3511) <= not a or b;
    layer0_outputs(3512) <= not b or a;
    layer0_outputs(3513) <= a;
    layer0_outputs(3514) <= a xor b;
    layer0_outputs(3515) <= not b;
    layer0_outputs(3516) <= not a or b;
    layer0_outputs(3517) <= not b or a;
    layer0_outputs(3518) <= not a or b;
    layer0_outputs(3519) <= not b;
    layer0_outputs(3520) <= not (a xor b);
    layer0_outputs(3521) <= a or b;
    layer0_outputs(3522) <= not b or a;
    layer0_outputs(3523) <= not (a or b);
    layer0_outputs(3524) <= a and not b;
    layer0_outputs(3525) <= not b or a;
    layer0_outputs(3526) <= a or b;
    layer0_outputs(3527) <= b and not a;
    layer0_outputs(3528) <= not b;
    layer0_outputs(3529) <= a and not b;
    layer0_outputs(3530) <= a;
    layer0_outputs(3531) <= a xor b;
    layer0_outputs(3532) <= a and not b;
    layer0_outputs(3533) <= not b or a;
    layer0_outputs(3534) <= not a;
    layer0_outputs(3535) <= not a or b;
    layer0_outputs(3536) <= a;
    layer0_outputs(3537) <= '1';
    layer0_outputs(3538) <= not a;
    layer0_outputs(3539) <= b;
    layer0_outputs(3540) <= a and b;
    layer0_outputs(3541) <= '0';
    layer0_outputs(3542) <= not b or a;
    layer0_outputs(3543) <= b;
    layer0_outputs(3544) <= not b;
    layer0_outputs(3545) <= not (a or b);
    layer0_outputs(3546) <= not b or a;
    layer0_outputs(3547) <= not b;
    layer0_outputs(3548) <= a;
    layer0_outputs(3549) <= a xor b;
    layer0_outputs(3550) <= b and not a;
    layer0_outputs(3551) <= not a;
    layer0_outputs(3552) <= not (a or b);
    layer0_outputs(3553) <= not a;
    layer0_outputs(3554) <= not a;
    layer0_outputs(3555) <= a;
    layer0_outputs(3556) <= not b;
    layer0_outputs(3557) <= not b;
    layer0_outputs(3558) <= '0';
    layer0_outputs(3559) <= '1';
    layer0_outputs(3560) <= b;
    layer0_outputs(3561) <= b;
    layer0_outputs(3562) <= not b;
    layer0_outputs(3563) <= a and not b;
    layer0_outputs(3564) <= '0';
    layer0_outputs(3565) <= b and not a;
    layer0_outputs(3566) <= not (a xor b);
    layer0_outputs(3567) <= not b or a;
    layer0_outputs(3568) <= not a or b;
    layer0_outputs(3569) <= not (a or b);
    layer0_outputs(3570) <= a;
    layer0_outputs(3571) <= not a;
    layer0_outputs(3572) <= not (a and b);
    layer0_outputs(3573) <= a and b;
    layer0_outputs(3574) <= a or b;
    layer0_outputs(3575) <= b;
    layer0_outputs(3576) <= not b;
    layer0_outputs(3577) <= not b or a;
    layer0_outputs(3578) <= not (a xor b);
    layer0_outputs(3579) <= '1';
    layer0_outputs(3580) <= not a or b;
    layer0_outputs(3581) <= a and b;
    layer0_outputs(3582) <= not b or a;
    layer0_outputs(3583) <= a or b;
    layer0_outputs(3584) <= b and not a;
    layer0_outputs(3585) <= b;
    layer0_outputs(3586) <= a xor b;
    layer0_outputs(3587) <= '0';
    layer0_outputs(3588) <= not a;
    layer0_outputs(3589) <= not b;
    layer0_outputs(3590) <= a or b;
    layer0_outputs(3591) <= not a;
    layer0_outputs(3592) <= not (a and b);
    layer0_outputs(3593) <= not a;
    layer0_outputs(3594) <= not a or b;
    layer0_outputs(3595) <= not a or b;
    layer0_outputs(3596) <= a or b;
    layer0_outputs(3597) <= a;
    layer0_outputs(3598) <= not b;
    layer0_outputs(3599) <= a or b;
    layer0_outputs(3600) <= a;
    layer0_outputs(3601) <= not b or a;
    layer0_outputs(3602) <= not b or a;
    layer0_outputs(3603) <= not b;
    layer0_outputs(3604) <= a and not b;
    layer0_outputs(3605) <= a;
    layer0_outputs(3606) <= b;
    layer0_outputs(3607) <= b;
    layer0_outputs(3608) <= a;
    layer0_outputs(3609) <= a xor b;
    layer0_outputs(3610) <= b and not a;
    layer0_outputs(3611) <= not (a or b);
    layer0_outputs(3612) <= not b;
    layer0_outputs(3613) <= a xor b;
    layer0_outputs(3614) <= a and not b;
    layer0_outputs(3615) <= not a;
    layer0_outputs(3616) <= not b;
    layer0_outputs(3617) <= '0';
    layer0_outputs(3618) <= not (a or b);
    layer0_outputs(3619) <= not (a and b);
    layer0_outputs(3620) <= a or b;
    layer0_outputs(3621) <= a and b;
    layer0_outputs(3622) <= '1';
    layer0_outputs(3623) <= not a;
    layer0_outputs(3624) <= not (a and b);
    layer0_outputs(3625) <= not a;
    layer0_outputs(3626) <= '1';
    layer0_outputs(3627) <= a xor b;
    layer0_outputs(3628) <= not (a or b);
    layer0_outputs(3629) <= a or b;
    layer0_outputs(3630) <= not a or b;
    layer0_outputs(3631) <= not a;
    layer0_outputs(3632) <= not (a or b);
    layer0_outputs(3633) <= not a;
    layer0_outputs(3634) <= a or b;
    layer0_outputs(3635) <= not a or b;
    layer0_outputs(3636) <= '0';
    layer0_outputs(3637) <= a;
    layer0_outputs(3638) <= a and b;
    layer0_outputs(3639) <= '0';
    layer0_outputs(3640) <= not a or b;
    layer0_outputs(3641) <= not (a or b);
    layer0_outputs(3642) <= not (a xor b);
    layer0_outputs(3643) <= b;
    layer0_outputs(3644) <= not (a xor b);
    layer0_outputs(3645) <= a and b;
    layer0_outputs(3646) <= b;
    layer0_outputs(3647) <= not a;
    layer0_outputs(3648) <= not b or a;
    layer0_outputs(3649) <= a or b;
    layer0_outputs(3650) <= a or b;
    layer0_outputs(3651) <= a and b;
    layer0_outputs(3652) <= b;
    layer0_outputs(3653) <= '0';
    layer0_outputs(3654) <= b and not a;
    layer0_outputs(3655) <= not a;
    layer0_outputs(3656) <= a or b;
    layer0_outputs(3657) <= b and not a;
    layer0_outputs(3658) <= not (a xor b);
    layer0_outputs(3659) <= b and not a;
    layer0_outputs(3660) <= not b;
    layer0_outputs(3661) <= b and not a;
    layer0_outputs(3662) <= not (a xor b);
    layer0_outputs(3663) <= not (a or b);
    layer0_outputs(3664) <= not (a and b);
    layer0_outputs(3665) <= '0';
    layer0_outputs(3666) <= not a or b;
    layer0_outputs(3667) <= not (a or b);
    layer0_outputs(3668) <= a xor b;
    layer0_outputs(3669) <= '0';
    layer0_outputs(3670) <= a;
    layer0_outputs(3671) <= b and not a;
    layer0_outputs(3672) <= not a or b;
    layer0_outputs(3673) <= not (a or b);
    layer0_outputs(3674) <= not (a or b);
    layer0_outputs(3675) <= not a;
    layer0_outputs(3676) <= b;
    layer0_outputs(3677) <= not (a xor b);
    layer0_outputs(3678) <= not b;
    layer0_outputs(3679) <= not b;
    layer0_outputs(3680) <= not b;
    layer0_outputs(3681) <= b;
    layer0_outputs(3682) <= b and not a;
    layer0_outputs(3683) <= b;
    layer0_outputs(3684) <= a or b;
    layer0_outputs(3685) <= not a or b;
    layer0_outputs(3686) <= not a;
    layer0_outputs(3687) <= a and not b;
    layer0_outputs(3688) <= not a or b;
    layer0_outputs(3689) <= not (a and b);
    layer0_outputs(3690) <= not (a and b);
    layer0_outputs(3691) <= a and not b;
    layer0_outputs(3692) <= a and not b;
    layer0_outputs(3693) <= not b;
    layer0_outputs(3694) <= a xor b;
    layer0_outputs(3695) <= not b;
    layer0_outputs(3696) <= '1';
    layer0_outputs(3697) <= b and not a;
    layer0_outputs(3698) <= a and not b;
    layer0_outputs(3699) <= not b or a;
    layer0_outputs(3700) <= not a;
    layer0_outputs(3701) <= a xor b;
    layer0_outputs(3702) <= a or b;
    layer0_outputs(3703) <= a and not b;
    layer0_outputs(3704) <= a xor b;
    layer0_outputs(3705) <= not b;
    layer0_outputs(3706) <= a or b;
    layer0_outputs(3707) <= not (a xor b);
    layer0_outputs(3708) <= a and not b;
    layer0_outputs(3709) <= not (a or b);
    layer0_outputs(3710) <= a;
    layer0_outputs(3711) <= b and not a;
    layer0_outputs(3712) <= a or b;
    layer0_outputs(3713) <= b;
    layer0_outputs(3714) <= a or b;
    layer0_outputs(3715) <= not (a or b);
    layer0_outputs(3716) <= b;
    layer0_outputs(3717) <= not (a or b);
    layer0_outputs(3718) <= a xor b;
    layer0_outputs(3719) <= not (a xor b);
    layer0_outputs(3720) <= not a or b;
    layer0_outputs(3721) <= not (a xor b);
    layer0_outputs(3722) <= not (a or b);
    layer0_outputs(3723) <= not a or b;
    layer0_outputs(3724) <= not (a xor b);
    layer0_outputs(3725) <= a;
    layer0_outputs(3726) <= not b;
    layer0_outputs(3727) <= not a;
    layer0_outputs(3728) <= a or b;
    layer0_outputs(3729) <= not b or a;
    layer0_outputs(3730) <= not (a and b);
    layer0_outputs(3731) <= not a or b;
    layer0_outputs(3732) <= not (a or b);
    layer0_outputs(3733) <= not b or a;
    layer0_outputs(3734) <= b and not a;
    layer0_outputs(3735) <= a and not b;
    layer0_outputs(3736) <= '0';
    layer0_outputs(3737) <= a and not b;
    layer0_outputs(3738) <= a and not b;
    layer0_outputs(3739) <= b and not a;
    layer0_outputs(3740) <= a or b;
    layer0_outputs(3741) <= a xor b;
    layer0_outputs(3742) <= not (a and b);
    layer0_outputs(3743) <= not (a and b);
    layer0_outputs(3744) <= a and b;
    layer0_outputs(3745) <= b and not a;
    layer0_outputs(3746) <= '0';
    layer0_outputs(3747) <= a or b;
    layer0_outputs(3748) <= not b;
    layer0_outputs(3749) <= '0';
    layer0_outputs(3750) <= not a or b;
    layer0_outputs(3751) <= not a;
    layer0_outputs(3752) <= not a or b;
    layer0_outputs(3753) <= a xor b;
    layer0_outputs(3754) <= b;
    layer0_outputs(3755) <= not a or b;
    layer0_outputs(3756) <= not b or a;
    layer0_outputs(3757) <= not a;
    layer0_outputs(3758) <= not b;
    layer0_outputs(3759) <= a;
    layer0_outputs(3760) <= not b or a;
    layer0_outputs(3761) <= not (a and b);
    layer0_outputs(3762) <= not b;
    layer0_outputs(3763) <= not a;
    layer0_outputs(3764) <= not (a or b);
    layer0_outputs(3765) <= not b or a;
    layer0_outputs(3766) <= a and b;
    layer0_outputs(3767) <= not a or b;
    layer0_outputs(3768) <= not a;
    layer0_outputs(3769) <= not b;
    layer0_outputs(3770) <= not (a or b);
    layer0_outputs(3771) <= not b;
    layer0_outputs(3772) <= '0';
    layer0_outputs(3773) <= a and not b;
    layer0_outputs(3774) <= not a or b;
    layer0_outputs(3775) <= not (a xor b);
    layer0_outputs(3776) <= not (a xor b);
    layer0_outputs(3777) <= a or b;
    layer0_outputs(3778) <= '1';
    layer0_outputs(3779) <= a xor b;
    layer0_outputs(3780) <= not b or a;
    layer0_outputs(3781) <= not a;
    layer0_outputs(3782) <= a xor b;
    layer0_outputs(3783) <= not (a or b);
    layer0_outputs(3784) <= a xor b;
    layer0_outputs(3785) <= not a;
    layer0_outputs(3786) <= not b or a;
    layer0_outputs(3787) <= not a;
    layer0_outputs(3788) <= not a or b;
    layer0_outputs(3789) <= not a;
    layer0_outputs(3790) <= not a or b;
    layer0_outputs(3791) <= not (a xor b);
    layer0_outputs(3792) <= not b;
    layer0_outputs(3793) <= not (a or b);
    layer0_outputs(3794) <= '1';
    layer0_outputs(3795) <= a and not b;
    layer0_outputs(3796) <= not (a xor b);
    layer0_outputs(3797) <= a and not b;
    layer0_outputs(3798) <= a;
    layer0_outputs(3799) <= a or b;
    layer0_outputs(3800) <= not b or a;
    layer0_outputs(3801) <= not (a or b);
    layer0_outputs(3802) <= b;
    layer0_outputs(3803) <= b;
    layer0_outputs(3804) <= not b or a;
    layer0_outputs(3805) <= not (a and b);
    layer0_outputs(3806) <= not a;
    layer0_outputs(3807) <= a;
    layer0_outputs(3808) <= a;
    layer0_outputs(3809) <= a and not b;
    layer0_outputs(3810) <= b;
    layer0_outputs(3811) <= not b;
    layer0_outputs(3812) <= '1';
    layer0_outputs(3813) <= b;
    layer0_outputs(3814) <= not b;
    layer0_outputs(3815) <= a;
    layer0_outputs(3816) <= not b or a;
    layer0_outputs(3817) <= not b or a;
    layer0_outputs(3818) <= b and not a;
    layer0_outputs(3819) <= a or b;
    layer0_outputs(3820) <= not b;
    layer0_outputs(3821) <= not a or b;
    layer0_outputs(3822) <= not b;
    layer0_outputs(3823) <= not a;
    layer0_outputs(3824) <= b;
    layer0_outputs(3825) <= not a;
    layer0_outputs(3826) <= not b or a;
    layer0_outputs(3827) <= not (a and b);
    layer0_outputs(3828) <= '1';
    layer0_outputs(3829) <= b;
    layer0_outputs(3830) <= not a or b;
    layer0_outputs(3831) <= a xor b;
    layer0_outputs(3832) <= not b;
    layer0_outputs(3833) <= a or b;
    layer0_outputs(3834) <= not b or a;
    layer0_outputs(3835) <= b;
    layer0_outputs(3836) <= not a;
    layer0_outputs(3837) <= a and not b;
    layer0_outputs(3838) <= a or b;
    layer0_outputs(3839) <= not (a xor b);
    layer0_outputs(3840) <= '1';
    layer0_outputs(3841) <= not a or b;
    layer0_outputs(3842) <= '1';
    layer0_outputs(3843) <= a or b;
    layer0_outputs(3844) <= not a;
    layer0_outputs(3845) <= not (a xor b);
    layer0_outputs(3846) <= not (a and b);
    layer0_outputs(3847) <= a and b;
    layer0_outputs(3848) <= not a or b;
    layer0_outputs(3849) <= not a;
    layer0_outputs(3850) <= not a;
    layer0_outputs(3851) <= b and not a;
    layer0_outputs(3852) <= '0';
    layer0_outputs(3853) <= b;
    layer0_outputs(3854) <= not b or a;
    layer0_outputs(3855) <= not a or b;
    layer0_outputs(3856) <= not (a or b);
    layer0_outputs(3857) <= a and not b;
    layer0_outputs(3858) <= b;
    layer0_outputs(3859) <= not b or a;
    layer0_outputs(3860) <= '0';
    layer0_outputs(3861) <= a xor b;
    layer0_outputs(3862) <= a and b;
    layer0_outputs(3863) <= '0';
    layer0_outputs(3864) <= a and b;
    layer0_outputs(3865) <= a or b;
    layer0_outputs(3866) <= a and b;
    layer0_outputs(3867) <= not a;
    layer0_outputs(3868) <= a and not b;
    layer0_outputs(3869) <= not b;
    layer0_outputs(3870) <= a and not b;
    layer0_outputs(3871) <= a or b;
    layer0_outputs(3872) <= not b;
    layer0_outputs(3873) <= not b;
    layer0_outputs(3874) <= '1';
    layer0_outputs(3875) <= not (a or b);
    layer0_outputs(3876) <= not b;
    layer0_outputs(3877) <= not b or a;
    layer0_outputs(3878) <= '1';
    layer0_outputs(3879) <= not a or b;
    layer0_outputs(3880) <= not (a xor b);
    layer0_outputs(3881) <= not (a or b);
    layer0_outputs(3882) <= a or b;
    layer0_outputs(3883) <= not a;
    layer0_outputs(3884) <= not (a xor b);
    layer0_outputs(3885) <= b and not a;
    layer0_outputs(3886) <= not a;
    layer0_outputs(3887) <= b and not a;
    layer0_outputs(3888) <= not b or a;
    layer0_outputs(3889) <= a and b;
    layer0_outputs(3890) <= not a;
    layer0_outputs(3891) <= a or b;
    layer0_outputs(3892) <= not b or a;
    layer0_outputs(3893) <= not a;
    layer0_outputs(3894) <= not a or b;
    layer0_outputs(3895) <= not a or b;
    layer0_outputs(3896) <= a xor b;
    layer0_outputs(3897) <= a and not b;
    layer0_outputs(3898) <= not b;
    layer0_outputs(3899) <= not (a xor b);
    layer0_outputs(3900) <= not b or a;
    layer0_outputs(3901) <= b and not a;
    layer0_outputs(3902) <= not a or b;
    layer0_outputs(3903) <= not a or b;
    layer0_outputs(3904) <= b and not a;
    layer0_outputs(3905) <= not (a or b);
    layer0_outputs(3906) <= a xor b;
    layer0_outputs(3907) <= not (a and b);
    layer0_outputs(3908) <= a and not b;
    layer0_outputs(3909) <= not b or a;
    layer0_outputs(3910) <= not a or b;
    layer0_outputs(3911) <= b;
    layer0_outputs(3912) <= b;
    layer0_outputs(3913) <= b and not a;
    layer0_outputs(3914) <= not (a and b);
    layer0_outputs(3915) <= '0';
    layer0_outputs(3916) <= not a;
    layer0_outputs(3917) <= a or b;
    layer0_outputs(3918) <= b;
    layer0_outputs(3919) <= a xor b;
    layer0_outputs(3920) <= not a or b;
    layer0_outputs(3921) <= '0';
    layer0_outputs(3922) <= b;
    layer0_outputs(3923) <= a xor b;
    layer0_outputs(3924) <= a xor b;
    layer0_outputs(3925) <= a and b;
    layer0_outputs(3926) <= a xor b;
    layer0_outputs(3927) <= a or b;
    layer0_outputs(3928) <= not a or b;
    layer0_outputs(3929) <= not (a or b);
    layer0_outputs(3930) <= not a or b;
    layer0_outputs(3931) <= not a or b;
    layer0_outputs(3932) <= a or b;
    layer0_outputs(3933) <= a and not b;
    layer0_outputs(3934) <= a and not b;
    layer0_outputs(3935) <= a or b;
    layer0_outputs(3936) <= not b or a;
    layer0_outputs(3937) <= b;
    layer0_outputs(3938) <= '1';
    layer0_outputs(3939) <= a;
    layer0_outputs(3940) <= not a or b;
    layer0_outputs(3941) <= b;
    layer0_outputs(3942) <= a or b;
    layer0_outputs(3943) <= a or b;
    layer0_outputs(3944) <= not a;
    layer0_outputs(3945) <= a or b;
    layer0_outputs(3946) <= '1';
    layer0_outputs(3947) <= not (a or b);
    layer0_outputs(3948) <= a or b;
    layer0_outputs(3949) <= b;
    layer0_outputs(3950) <= not (a xor b);
    layer0_outputs(3951) <= a xor b;
    layer0_outputs(3952) <= not (a and b);
    layer0_outputs(3953) <= a and not b;
    layer0_outputs(3954) <= not (a xor b);
    layer0_outputs(3955) <= a and not b;
    layer0_outputs(3956) <= a;
    layer0_outputs(3957) <= not (a or b);
    layer0_outputs(3958) <= not b or a;
    layer0_outputs(3959) <= a or b;
    layer0_outputs(3960) <= a or b;
    layer0_outputs(3961) <= not (a and b);
    layer0_outputs(3962) <= not a;
    layer0_outputs(3963) <= not b or a;
    layer0_outputs(3964) <= a or b;
    layer0_outputs(3965) <= a or b;
    layer0_outputs(3966) <= '0';
    layer0_outputs(3967) <= a and b;
    layer0_outputs(3968) <= not a or b;
    layer0_outputs(3969) <= not a or b;
    layer0_outputs(3970) <= a xor b;
    layer0_outputs(3971) <= not a;
    layer0_outputs(3972) <= not (a and b);
    layer0_outputs(3973) <= a or b;
    layer0_outputs(3974) <= not (a or b);
    layer0_outputs(3975) <= not a;
    layer0_outputs(3976) <= '0';
    layer0_outputs(3977) <= not b or a;
    layer0_outputs(3978) <= a xor b;
    layer0_outputs(3979) <= a and b;
    layer0_outputs(3980) <= '0';
    layer0_outputs(3981) <= '1';
    layer0_outputs(3982) <= not a;
    layer0_outputs(3983) <= a or b;
    layer0_outputs(3984) <= b;
    layer0_outputs(3985) <= not (a xor b);
    layer0_outputs(3986) <= not (a or b);
    layer0_outputs(3987) <= not b or a;
    layer0_outputs(3988) <= not b or a;
    layer0_outputs(3989) <= b;
    layer0_outputs(3990) <= a and not b;
    layer0_outputs(3991) <= b and not a;
    layer0_outputs(3992) <= a;
    layer0_outputs(3993) <= '1';
    layer0_outputs(3994) <= not a or b;
    layer0_outputs(3995) <= a and not b;
    layer0_outputs(3996) <= '0';
    layer0_outputs(3997) <= b;
    layer0_outputs(3998) <= not (a and b);
    layer0_outputs(3999) <= a and b;
    layer0_outputs(4000) <= a or b;
    layer0_outputs(4001) <= not a or b;
    layer0_outputs(4002) <= b and not a;
    layer0_outputs(4003) <= not b or a;
    layer0_outputs(4004) <= not b or a;
    layer0_outputs(4005) <= a and b;
    layer0_outputs(4006) <= not a or b;
    layer0_outputs(4007) <= not b or a;
    layer0_outputs(4008) <= not a or b;
    layer0_outputs(4009) <= a and b;
    layer0_outputs(4010) <= a or b;
    layer0_outputs(4011) <= not (a and b);
    layer0_outputs(4012) <= not (a or b);
    layer0_outputs(4013) <= b and not a;
    layer0_outputs(4014) <= '1';
    layer0_outputs(4015) <= not a;
    layer0_outputs(4016) <= a or b;
    layer0_outputs(4017) <= not a;
    layer0_outputs(4018) <= a or b;
    layer0_outputs(4019) <= b;
    layer0_outputs(4020) <= not (a xor b);
    layer0_outputs(4021) <= not (a or b);
    layer0_outputs(4022) <= not (a and b);
    layer0_outputs(4023) <= not b;
    layer0_outputs(4024) <= a and b;
    layer0_outputs(4025) <= '0';
    layer0_outputs(4026) <= b and not a;
    layer0_outputs(4027) <= not b or a;
    layer0_outputs(4028) <= a xor b;
    layer0_outputs(4029) <= b and not a;
    layer0_outputs(4030) <= a;
    layer0_outputs(4031) <= not b or a;
    layer0_outputs(4032) <= not (a and b);
    layer0_outputs(4033) <= '1';
    layer0_outputs(4034) <= a;
    layer0_outputs(4035) <= a or b;
    layer0_outputs(4036) <= not (a xor b);
    layer0_outputs(4037) <= '0';
    layer0_outputs(4038) <= a xor b;
    layer0_outputs(4039) <= not b or a;
    layer0_outputs(4040) <= not b or a;
    layer0_outputs(4041) <= b and not a;
    layer0_outputs(4042) <= a and not b;
    layer0_outputs(4043) <= not (a xor b);
    layer0_outputs(4044) <= not b or a;
    layer0_outputs(4045) <= a;
    layer0_outputs(4046) <= a and b;
    layer0_outputs(4047) <= not a or b;
    layer0_outputs(4048) <= a and b;
    layer0_outputs(4049) <= '0';
    layer0_outputs(4050) <= a;
    layer0_outputs(4051) <= a xor b;
    layer0_outputs(4052) <= a and b;
    layer0_outputs(4053) <= not (a or b);
    layer0_outputs(4054) <= b;
    layer0_outputs(4055) <= not b or a;
    layer0_outputs(4056) <= not a;
    layer0_outputs(4057) <= a;
    layer0_outputs(4058) <= not a;
    layer0_outputs(4059) <= not b;
    layer0_outputs(4060) <= '0';
    layer0_outputs(4061) <= b and not a;
    layer0_outputs(4062) <= b and not a;
    layer0_outputs(4063) <= '0';
    layer0_outputs(4064) <= a or b;
    layer0_outputs(4065) <= not (a xor b);
    layer0_outputs(4066) <= not a;
    layer0_outputs(4067) <= not a or b;
    layer0_outputs(4068) <= a and not b;
    layer0_outputs(4069) <= not (a or b);
    layer0_outputs(4070) <= a;
    layer0_outputs(4071) <= b and not a;
    layer0_outputs(4072) <= not a or b;
    layer0_outputs(4073) <= '0';
    layer0_outputs(4074) <= a or b;
    layer0_outputs(4075) <= not b;
    layer0_outputs(4076) <= not (a and b);
    layer0_outputs(4077) <= not (a or b);
    layer0_outputs(4078) <= a or b;
    layer0_outputs(4079) <= a;
    layer0_outputs(4080) <= a and b;
    layer0_outputs(4081) <= not a;
    layer0_outputs(4082) <= '0';
    layer0_outputs(4083) <= '1';
    layer0_outputs(4084) <= b and not a;
    layer0_outputs(4085) <= a and not b;
    layer0_outputs(4086) <= not a;
    layer0_outputs(4087) <= '1';
    layer0_outputs(4088) <= not (a xor b);
    layer0_outputs(4089) <= not (a or b);
    layer0_outputs(4090) <= not (a and b);
    layer0_outputs(4091) <= not (a xor b);
    layer0_outputs(4092) <= b and not a;
    layer0_outputs(4093) <= a or b;
    layer0_outputs(4094) <= b and not a;
    layer0_outputs(4095) <= a and b;
    layer0_outputs(4096) <= a and b;
    layer0_outputs(4097) <= not a;
    layer0_outputs(4098) <= '1';
    layer0_outputs(4099) <= a;
    layer0_outputs(4100) <= not b;
    layer0_outputs(4101) <= a and not b;
    layer0_outputs(4102) <= '0';
    layer0_outputs(4103) <= a or b;
    layer0_outputs(4104) <= not b;
    layer0_outputs(4105) <= not (a or b);
    layer0_outputs(4106) <= not (a and b);
    layer0_outputs(4107) <= a;
    layer0_outputs(4108) <= not (a xor b);
    layer0_outputs(4109) <= not (a and b);
    layer0_outputs(4110) <= b and not a;
    layer0_outputs(4111) <= '1';
    layer0_outputs(4112) <= not b;
    layer0_outputs(4113) <= not b or a;
    layer0_outputs(4114) <= a;
    layer0_outputs(4115) <= not a;
    layer0_outputs(4116) <= '0';
    layer0_outputs(4117) <= a and not b;
    layer0_outputs(4118) <= not (a and b);
    layer0_outputs(4119) <= a and not b;
    layer0_outputs(4120) <= not a;
    layer0_outputs(4121) <= b;
    layer0_outputs(4122) <= not a;
    layer0_outputs(4123) <= a;
    layer0_outputs(4124) <= not b or a;
    layer0_outputs(4125) <= not a or b;
    layer0_outputs(4126) <= not a;
    layer0_outputs(4127) <= not (a and b);
    layer0_outputs(4128) <= a;
    layer0_outputs(4129) <= a and not b;
    layer0_outputs(4130) <= not (a or b);
    layer0_outputs(4131) <= a;
    layer0_outputs(4132) <= a;
    layer0_outputs(4133) <= not b or a;
    layer0_outputs(4134) <= a or b;
    layer0_outputs(4135) <= not b;
    layer0_outputs(4136) <= not a or b;
    layer0_outputs(4137) <= not b or a;
    layer0_outputs(4138) <= b and not a;
    layer0_outputs(4139) <= a and not b;
    layer0_outputs(4140) <= not b;
    layer0_outputs(4141) <= not (a or b);
    layer0_outputs(4142) <= b;
    layer0_outputs(4143) <= a or b;
    layer0_outputs(4144) <= a or b;
    layer0_outputs(4145) <= b;
    layer0_outputs(4146) <= not (a and b);
    layer0_outputs(4147) <= a or b;
    layer0_outputs(4148) <= not (a or b);
    layer0_outputs(4149) <= not (a or b);
    layer0_outputs(4150) <= '1';
    layer0_outputs(4151) <= a;
    layer0_outputs(4152) <= not (a or b);
    layer0_outputs(4153) <= a xor b;
    layer0_outputs(4154) <= a or b;
    layer0_outputs(4155) <= not (a or b);
    layer0_outputs(4156) <= not (a or b);
    layer0_outputs(4157) <= not (a xor b);
    layer0_outputs(4158) <= not a;
    layer0_outputs(4159) <= a and b;
    layer0_outputs(4160) <= not a or b;
    layer0_outputs(4161) <= not (a and b);
    layer0_outputs(4162) <= not (a xor b);
    layer0_outputs(4163) <= not (a xor b);
    layer0_outputs(4164) <= not a;
    layer0_outputs(4165) <= a or b;
    layer0_outputs(4166) <= not (a or b);
    layer0_outputs(4167) <= not (a and b);
    layer0_outputs(4168) <= b;
    layer0_outputs(4169) <= not (a and b);
    layer0_outputs(4170) <= a or b;
    layer0_outputs(4171) <= a or b;
    layer0_outputs(4172) <= b and not a;
    layer0_outputs(4173) <= '1';
    layer0_outputs(4174) <= a;
    layer0_outputs(4175) <= not (a and b);
    layer0_outputs(4176) <= a and b;
    layer0_outputs(4177) <= a or b;
    layer0_outputs(4178) <= a and not b;
    layer0_outputs(4179) <= not b;
    layer0_outputs(4180) <= a and not b;
    layer0_outputs(4181) <= not (a or b);
    layer0_outputs(4182) <= a;
    layer0_outputs(4183) <= '0';
    layer0_outputs(4184) <= b;
    layer0_outputs(4185) <= a and not b;
    layer0_outputs(4186) <= a;
    layer0_outputs(4187) <= not (a and b);
    layer0_outputs(4188) <= a or b;
    layer0_outputs(4189) <= not b or a;
    layer0_outputs(4190) <= a;
    layer0_outputs(4191) <= not a or b;
    layer0_outputs(4192) <= a or b;
    layer0_outputs(4193) <= '1';
    layer0_outputs(4194) <= b;
    layer0_outputs(4195) <= not b or a;
    layer0_outputs(4196) <= not (a or b);
    layer0_outputs(4197) <= not (a xor b);
    layer0_outputs(4198) <= b;
    layer0_outputs(4199) <= a or b;
    layer0_outputs(4200) <= a;
    layer0_outputs(4201) <= a xor b;
    layer0_outputs(4202) <= not a;
    layer0_outputs(4203) <= not (a xor b);
    layer0_outputs(4204) <= '0';
    layer0_outputs(4205) <= a or b;
    layer0_outputs(4206) <= not b;
    layer0_outputs(4207) <= a xor b;
    layer0_outputs(4208) <= not (a or b);
    layer0_outputs(4209) <= a;
    layer0_outputs(4210) <= not a;
    layer0_outputs(4211) <= not (a and b);
    layer0_outputs(4212) <= not (a and b);
    layer0_outputs(4213) <= b and not a;
    layer0_outputs(4214) <= a xor b;
    layer0_outputs(4215) <= b;
    layer0_outputs(4216) <= a;
    layer0_outputs(4217) <= '0';
    layer0_outputs(4218) <= b and not a;
    layer0_outputs(4219) <= a xor b;
    layer0_outputs(4220) <= not (a or b);
    layer0_outputs(4221) <= a xor b;
    layer0_outputs(4222) <= a and not b;
    layer0_outputs(4223) <= b;
    layer0_outputs(4224) <= b and not a;
    layer0_outputs(4225) <= a;
    layer0_outputs(4226) <= not (a and b);
    layer0_outputs(4227) <= not b or a;
    layer0_outputs(4228) <= not a or b;
    layer0_outputs(4229) <= b and not a;
    layer0_outputs(4230) <= a;
    layer0_outputs(4231) <= a;
    layer0_outputs(4232) <= not (a xor b);
    layer0_outputs(4233) <= not b;
    layer0_outputs(4234) <= a and not b;
    layer0_outputs(4235) <= not b;
    layer0_outputs(4236) <= a and b;
    layer0_outputs(4237) <= not a or b;
    layer0_outputs(4238) <= not b;
    layer0_outputs(4239) <= not b;
    layer0_outputs(4240) <= not (a xor b);
    layer0_outputs(4241) <= a and b;
    layer0_outputs(4242) <= not b;
    layer0_outputs(4243) <= not (a or b);
    layer0_outputs(4244) <= b;
    layer0_outputs(4245) <= not b or a;
    layer0_outputs(4246) <= b;
    layer0_outputs(4247) <= a or b;
    layer0_outputs(4248) <= b and not a;
    layer0_outputs(4249) <= a or b;
    layer0_outputs(4250) <= not b or a;
    layer0_outputs(4251) <= not (a or b);
    layer0_outputs(4252) <= a and not b;
    layer0_outputs(4253) <= not a or b;
    layer0_outputs(4254) <= a and not b;
    layer0_outputs(4255) <= not b;
    layer0_outputs(4256) <= b and not a;
    layer0_outputs(4257) <= not a or b;
    layer0_outputs(4258) <= not (a or b);
    layer0_outputs(4259) <= b;
    layer0_outputs(4260) <= not a or b;
    layer0_outputs(4261) <= not b;
    layer0_outputs(4262) <= not a or b;
    layer0_outputs(4263) <= a;
    layer0_outputs(4264) <= not (a and b);
    layer0_outputs(4265) <= not b;
    layer0_outputs(4266) <= b and not a;
    layer0_outputs(4267) <= not a;
    layer0_outputs(4268) <= not a or b;
    layer0_outputs(4269) <= '1';
    layer0_outputs(4270) <= not (a xor b);
    layer0_outputs(4271) <= a and not b;
    layer0_outputs(4272) <= not (a or b);
    layer0_outputs(4273) <= b and not a;
    layer0_outputs(4274) <= '0';
    layer0_outputs(4275) <= b;
    layer0_outputs(4276) <= '0';
    layer0_outputs(4277) <= not b;
    layer0_outputs(4278) <= a or b;
    layer0_outputs(4279) <= a or b;
    layer0_outputs(4280) <= not b;
    layer0_outputs(4281) <= a xor b;
    layer0_outputs(4282) <= not (a xor b);
    layer0_outputs(4283) <= not (a xor b);
    layer0_outputs(4284) <= '0';
    layer0_outputs(4285) <= not (a or b);
    layer0_outputs(4286) <= not (a xor b);
    layer0_outputs(4287) <= a and b;
    layer0_outputs(4288) <= not (a xor b);
    layer0_outputs(4289) <= not a or b;
    layer0_outputs(4290) <= not a;
    layer0_outputs(4291) <= a and b;
    layer0_outputs(4292) <= not b or a;
    layer0_outputs(4293) <= not b;
    layer0_outputs(4294) <= not (a or b);
    layer0_outputs(4295) <= not b;
    layer0_outputs(4296) <= not (a or b);
    layer0_outputs(4297) <= a or b;
    layer0_outputs(4298) <= not (a and b);
    layer0_outputs(4299) <= a and b;
    layer0_outputs(4300) <= not (a xor b);
    layer0_outputs(4301) <= not (a or b);
    layer0_outputs(4302) <= a xor b;
    layer0_outputs(4303) <= '0';
    layer0_outputs(4304) <= '0';
    layer0_outputs(4305) <= '0';
    layer0_outputs(4306) <= not b or a;
    layer0_outputs(4307) <= not (a xor b);
    layer0_outputs(4308) <= not (a and b);
    layer0_outputs(4309) <= not a;
    layer0_outputs(4310) <= not b or a;
    layer0_outputs(4311) <= not a or b;
    layer0_outputs(4312) <= b;
    layer0_outputs(4313) <= not b or a;
    layer0_outputs(4314) <= a xor b;
    layer0_outputs(4315) <= not b or a;
    layer0_outputs(4316) <= not (a xor b);
    layer0_outputs(4317) <= not b;
    layer0_outputs(4318) <= b;
    layer0_outputs(4319) <= '0';
    layer0_outputs(4320) <= not (a or b);
    layer0_outputs(4321) <= not a;
    layer0_outputs(4322) <= not b;
    layer0_outputs(4323) <= '0';
    layer0_outputs(4324) <= not b or a;
    layer0_outputs(4325) <= not a;
    layer0_outputs(4326) <= b and not a;
    layer0_outputs(4327) <= not b;
    layer0_outputs(4328) <= '1';
    layer0_outputs(4329) <= b and not a;
    layer0_outputs(4330) <= not b;
    layer0_outputs(4331) <= a xor b;
    layer0_outputs(4332) <= a;
    layer0_outputs(4333) <= not b;
    layer0_outputs(4334) <= a and b;
    layer0_outputs(4335) <= a xor b;
    layer0_outputs(4336) <= a and not b;
    layer0_outputs(4337) <= a xor b;
    layer0_outputs(4338) <= not a or b;
    layer0_outputs(4339) <= a xor b;
    layer0_outputs(4340) <= '0';
    layer0_outputs(4341) <= a or b;
    layer0_outputs(4342) <= not (a xor b);
    layer0_outputs(4343) <= a xor b;
    layer0_outputs(4344) <= not b;
    layer0_outputs(4345) <= not (a and b);
    layer0_outputs(4346) <= not (a or b);
    layer0_outputs(4347) <= '1';
    layer0_outputs(4348) <= '1';
    layer0_outputs(4349) <= a or b;
    layer0_outputs(4350) <= a and not b;
    layer0_outputs(4351) <= a or b;
    layer0_outputs(4352) <= a or b;
    layer0_outputs(4353) <= not a;
    layer0_outputs(4354) <= '1';
    layer0_outputs(4355) <= not a;
    layer0_outputs(4356) <= not a;
    layer0_outputs(4357) <= a xor b;
    layer0_outputs(4358) <= not (a xor b);
    layer0_outputs(4359) <= not (a xor b);
    layer0_outputs(4360) <= b and not a;
    layer0_outputs(4361) <= not (a or b);
    layer0_outputs(4362) <= not (a xor b);
    layer0_outputs(4363) <= a;
    layer0_outputs(4364) <= not a;
    layer0_outputs(4365) <= b;
    layer0_outputs(4366) <= b;
    layer0_outputs(4367) <= not (a or b);
    layer0_outputs(4368) <= b;
    layer0_outputs(4369) <= not b or a;
    layer0_outputs(4370) <= a xor b;
    layer0_outputs(4371) <= a and not b;
    layer0_outputs(4372) <= not b or a;
    layer0_outputs(4373) <= not b;
    layer0_outputs(4374) <= not a or b;
    layer0_outputs(4375) <= not a;
    layer0_outputs(4376) <= a and not b;
    layer0_outputs(4377) <= not (a xor b);
    layer0_outputs(4378) <= not b or a;
    layer0_outputs(4379) <= not (a or b);
    layer0_outputs(4380) <= a and b;
    layer0_outputs(4381) <= b and not a;
    layer0_outputs(4382) <= a;
    layer0_outputs(4383) <= not b;
    layer0_outputs(4384) <= b;
    layer0_outputs(4385) <= a or b;
    layer0_outputs(4386) <= b and not a;
    layer0_outputs(4387) <= b and not a;
    layer0_outputs(4388) <= '0';
    layer0_outputs(4389) <= a and not b;
    layer0_outputs(4390) <= not (a and b);
    layer0_outputs(4391) <= '1';
    layer0_outputs(4392) <= not (a and b);
    layer0_outputs(4393) <= a;
    layer0_outputs(4394) <= a and b;
    layer0_outputs(4395) <= '0';
    layer0_outputs(4396) <= a and b;
    layer0_outputs(4397) <= '0';
    layer0_outputs(4398) <= b and not a;
    layer0_outputs(4399) <= '0';
    layer0_outputs(4400) <= a xor b;
    layer0_outputs(4401) <= '1';
    layer0_outputs(4402) <= not a;
    layer0_outputs(4403) <= a;
    layer0_outputs(4404) <= a and not b;
    layer0_outputs(4405) <= b;
    layer0_outputs(4406) <= '0';
    layer0_outputs(4407) <= not (a and b);
    layer0_outputs(4408) <= a or b;
    layer0_outputs(4409) <= b and not a;
    layer0_outputs(4410) <= a and b;
    layer0_outputs(4411) <= not (a or b);
    layer0_outputs(4412) <= b;
    layer0_outputs(4413) <= b and not a;
    layer0_outputs(4414) <= not (a xor b);
    layer0_outputs(4415) <= not (a and b);
    layer0_outputs(4416) <= not (a and b);
    layer0_outputs(4417) <= not b;
    layer0_outputs(4418) <= a xor b;
    layer0_outputs(4419) <= not b;
    layer0_outputs(4420) <= not a or b;
    layer0_outputs(4421) <= not b or a;
    layer0_outputs(4422) <= not b;
    layer0_outputs(4423) <= not a;
    layer0_outputs(4424) <= a xor b;
    layer0_outputs(4425) <= not (a xor b);
    layer0_outputs(4426) <= a xor b;
    layer0_outputs(4427) <= a or b;
    layer0_outputs(4428) <= not b;
    layer0_outputs(4429) <= a and not b;
    layer0_outputs(4430) <= not (a or b);
    layer0_outputs(4431) <= a;
    layer0_outputs(4432) <= a;
    layer0_outputs(4433) <= b and not a;
    layer0_outputs(4434) <= a or b;
    layer0_outputs(4435) <= a or b;
    layer0_outputs(4436) <= a xor b;
    layer0_outputs(4437) <= not (a and b);
    layer0_outputs(4438) <= a and b;
    layer0_outputs(4439) <= not (a or b);
    layer0_outputs(4440) <= not (a xor b);
    layer0_outputs(4441) <= a xor b;
    layer0_outputs(4442) <= a xor b;
    layer0_outputs(4443) <= a;
    layer0_outputs(4444) <= not (a and b);
    layer0_outputs(4445) <= not (a xor b);
    layer0_outputs(4446) <= '0';
    layer0_outputs(4447) <= a and not b;
    layer0_outputs(4448) <= not a;
    layer0_outputs(4449) <= a xor b;
    layer0_outputs(4450) <= not (a and b);
    layer0_outputs(4451) <= b and not a;
    layer0_outputs(4452) <= a or b;
    layer0_outputs(4453) <= '1';
    layer0_outputs(4454) <= a xor b;
    layer0_outputs(4455) <= a xor b;
    layer0_outputs(4456) <= '1';
    layer0_outputs(4457) <= a or b;
    layer0_outputs(4458) <= a or b;
    layer0_outputs(4459) <= not (a and b);
    layer0_outputs(4460) <= a;
    layer0_outputs(4461) <= not (a or b);
    layer0_outputs(4462) <= a and b;
    layer0_outputs(4463) <= not (a xor b);
    layer0_outputs(4464) <= b;
    layer0_outputs(4465) <= not (a or b);
    layer0_outputs(4466) <= not (a xor b);
    layer0_outputs(4467) <= not b;
    layer0_outputs(4468) <= '0';
    layer0_outputs(4469) <= not b;
    layer0_outputs(4470) <= a and b;
    layer0_outputs(4471) <= not a;
    layer0_outputs(4472) <= b and not a;
    layer0_outputs(4473) <= not (a and b);
    layer0_outputs(4474) <= not a or b;
    layer0_outputs(4475) <= not b;
    layer0_outputs(4476) <= not (a xor b);
    layer0_outputs(4477) <= not (a or b);
    layer0_outputs(4478) <= a and b;
    layer0_outputs(4479) <= a xor b;
    layer0_outputs(4480) <= a;
    layer0_outputs(4481) <= not (a xor b);
    layer0_outputs(4482) <= a or b;
    layer0_outputs(4483) <= '1';
    layer0_outputs(4484) <= not (a and b);
    layer0_outputs(4485) <= a or b;
    layer0_outputs(4486) <= a and b;
    layer0_outputs(4487) <= b and not a;
    layer0_outputs(4488) <= '1';
    layer0_outputs(4489) <= a;
    layer0_outputs(4490) <= a or b;
    layer0_outputs(4491) <= not a;
    layer0_outputs(4492) <= a or b;
    layer0_outputs(4493) <= a and not b;
    layer0_outputs(4494) <= a or b;
    layer0_outputs(4495) <= b and not a;
    layer0_outputs(4496) <= a and b;
    layer0_outputs(4497) <= not b;
    layer0_outputs(4498) <= a xor b;
    layer0_outputs(4499) <= a or b;
    layer0_outputs(4500) <= not (a and b);
    layer0_outputs(4501) <= not a or b;
    layer0_outputs(4502) <= '1';
    layer0_outputs(4503) <= not b or a;
    layer0_outputs(4504) <= b;
    layer0_outputs(4505) <= a or b;
    layer0_outputs(4506) <= a or b;
    layer0_outputs(4507) <= '1';
    layer0_outputs(4508) <= not b or a;
    layer0_outputs(4509) <= not a;
    layer0_outputs(4510) <= a and not b;
    layer0_outputs(4511) <= not b or a;
    layer0_outputs(4512) <= not (a or b);
    layer0_outputs(4513) <= a or b;
    layer0_outputs(4514) <= a or b;
    layer0_outputs(4515) <= b and not a;
    layer0_outputs(4516) <= not b or a;
    layer0_outputs(4517) <= not (a and b);
    layer0_outputs(4518) <= a or b;
    layer0_outputs(4519) <= not b or a;
    layer0_outputs(4520) <= b;
    layer0_outputs(4521) <= '1';
    layer0_outputs(4522) <= a and b;
    layer0_outputs(4523) <= not b;
    layer0_outputs(4524) <= not a;
    layer0_outputs(4525) <= a or b;
    layer0_outputs(4526) <= not (a xor b);
    layer0_outputs(4527) <= b;
    layer0_outputs(4528) <= not (a or b);
    layer0_outputs(4529) <= a xor b;
    layer0_outputs(4530) <= not (a or b);
    layer0_outputs(4531) <= not (a or b);
    layer0_outputs(4532) <= b and not a;
    layer0_outputs(4533) <= not b or a;
    layer0_outputs(4534) <= a;
    layer0_outputs(4535) <= not (a or b);
    layer0_outputs(4536) <= '0';
    layer0_outputs(4537) <= a or b;
    layer0_outputs(4538) <= not (a or b);
    layer0_outputs(4539) <= not (a and b);
    layer0_outputs(4540) <= not (a or b);
    layer0_outputs(4541) <= not (a or b);
    layer0_outputs(4542) <= not (a and b);
    layer0_outputs(4543) <= not a;
    layer0_outputs(4544) <= not (a or b);
    layer0_outputs(4545) <= not a;
    layer0_outputs(4546) <= not (a and b);
    layer0_outputs(4547) <= not (a or b);
    layer0_outputs(4548) <= a or b;
    layer0_outputs(4549) <= '1';
    layer0_outputs(4550) <= not (a xor b);
    layer0_outputs(4551) <= not b or a;
    layer0_outputs(4552) <= not (a xor b);
    layer0_outputs(4553) <= a and b;
    layer0_outputs(4554) <= not b;
    layer0_outputs(4555) <= b and not a;
    layer0_outputs(4556) <= not a;
    layer0_outputs(4557) <= not (a xor b);
    layer0_outputs(4558) <= b;
    layer0_outputs(4559) <= not a;
    layer0_outputs(4560) <= not a or b;
    layer0_outputs(4561) <= b;
    layer0_outputs(4562) <= not (a xor b);
    layer0_outputs(4563) <= a or b;
    layer0_outputs(4564) <= a or b;
    layer0_outputs(4565) <= not (a or b);
    layer0_outputs(4566) <= not a;
    layer0_outputs(4567) <= '1';
    layer0_outputs(4568) <= a and not b;
    layer0_outputs(4569) <= b;
    layer0_outputs(4570) <= a or b;
    layer0_outputs(4571) <= not b;
    layer0_outputs(4572) <= not a;
    layer0_outputs(4573) <= '1';
    layer0_outputs(4574) <= not a;
    layer0_outputs(4575) <= not (a xor b);
    layer0_outputs(4576) <= b;
    layer0_outputs(4577) <= a xor b;
    layer0_outputs(4578) <= a and not b;
    layer0_outputs(4579) <= '0';
    layer0_outputs(4580) <= a or b;
    layer0_outputs(4581) <= a xor b;
    layer0_outputs(4582) <= b;
    layer0_outputs(4583) <= a;
    layer0_outputs(4584) <= b and not a;
    layer0_outputs(4585) <= a xor b;
    layer0_outputs(4586) <= b;
    layer0_outputs(4587) <= a and b;
    layer0_outputs(4588) <= not (a or b);
    layer0_outputs(4589) <= not (a or b);
    layer0_outputs(4590) <= not a;
    layer0_outputs(4591) <= a;
    layer0_outputs(4592) <= b;
    layer0_outputs(4593) <= not (a or b);
    layer0_outputs(4594) <= '1';
    layer0_outputs(4595) <= b and not a;
    layer0_outputs(4596) <= '0';
    layer0_outputs(4597) <= not a;
    layer0_outputs(4598) <= not b;
    layer0_outputs(4599) <= not a;
    layer0_outputs(4600) <= not b;
    layer0_outputs(4601) <= a and not b;
    layer0_outputs(4602) <= b;
    layer0_outputs(4603) <= not a;
    layer0_outputs(4604) <= a;
    layer0_outputs(4605) <= b and not a;
    layer0_outputs(4606) <= not (a or b);
    layer0_outputs(4607) <= not b;
    layer0_outputs(4608) <= not (a or b);
    layer0_outputs(4609) <= not (a and b);
    layer0_outputs(4610) <= a and not b;
    layer0_outputs(4611) <= b;
    layer0_outputs(4612) <= b and not a;
    layer0_outputs(4613) <= b and not a;
    layer0_outputs(4614) <= not (a or b);
    layer0_outputs(4615) <= a;
    layer0_outputs(4616) <= b and not a;
    layer0_outputs(4617) <= a xor b;
    layer0_outputs(4618) <= not (a xor b);
    layer0_outputs(4619) <= a and b;
    layer0_outputs(4620) <= '1';
    layer0_outputs(4621) <= b;
    layer0_outputs(4622) <= a or b;
    layer0_outputs(4623) <= not (a and b);
    layer0_outputs(4624) <= a xor b;
    layer0_outputs(4625) <= a xor b;
    layer0_outputs(4626) <= a xor b;
    layer0_outputs(4627) <= not (a or b);
    layer0_outputs(4628) <= a or b;
    layer0_outputs(4629) <= not a or b;
    layer0_outputs(4630) <= not b or a;
    layer0_outputs(4631) <= not (a and b);
    layer0_outputs(4632) <= not b or a;
    layer0_outputs(4633) <= not a;
    layer0_outputs(4634) <= a or b;
    layer0_outputs(4635) <= b;
    layer0_outputs(4636) <= a or b;
    layer0_outputs(4637) <= not a or b;
    layer0_outputs(4638) <= not b or a;
    layer0_outputs(4639) <= a and b;
    layer0_outputs(4640) <= not b or a;
    layer0_outputs(4641) <= not b;
    layer0_outputs(4642) <= not b;
    layer0_outputs(4643) <= a and not b;
    layer0_outputs(4644) <= not a;
    layer0_outputs(4645) <= b;
    layer0_outputs(4646) <= b and not a;
    layer0_outputs(4647) <= not a;
    layer0_outputs(4648) <= a and not b;
    layer0_outputs(4649) <= not b or a;
    layer0_outputs(4650) <= a and b;
    layer0_outputs(4651) <= not a or b;
    layer0_outputs(4652) <= b;
    layer0_outputs(4653) <= not (a or b);
    layer0_outputs(4654) <= a;
    layer0_outputs(4655) <= a or b;
    layer0_outputs(4656) <= not b;
    layer0_outputs(4657) <= not (a or b);
    layer0_outputs(4658) <= b and not a;
    layer0_outputs(4659) <= not a;
    layer0_outputs(4660) <= '0';
    layer0_outputs(4661) <= '0';
    layer0_outputs(4662) <= not (a xor b);
    layer0_outputs(4663) <= a and not b;
    layer0_outputs(4664) <= a;
    layer0_outputs(4665) <= '1';
    layer0_outputs(4666) <= '1';
    layer0_outputs(4667) <= not b or a;
    layer0_outputs(4668) <= a;
    layer0_outputs(4669) <= a;
    layer0_outputs(4670) <= a;
    layer0_outputs(4671) <= a;
    layer0_outputs(4672) <= not (a or b);
    layer0_outputs(4673) <= not a or b;
    layer0_outputs(4674) <= not (a xor b);
    layer0_outputs(4675) <= not b or a;
    layer0_outputs(4676) <= a and not b;
    layer0_outputs(4677) <= not b;
    layer0_outputs(4678) <= not (a xor b);
    layer0_outputs(4679) <= a or b;
    layer0_outputs(4680) <= b and not a;
    layer0_outputs(4681) <= not (a xor b);
    layer0_outputs(4682) <= a;
    layer0_outputs(4683) <= a;
    layer0_outputs(4684) <= a and not b;
    layer0_outputs(4685) <= '0';
    layer0_outputs(4686) <= a and not b;
    layer0_outputs(4687) <= not a or b;
    layer0_outputs(4688) <= not (a xor b);
    layer0_outputs(4689) <= a;
    layer0_outputs(4690) <= not a;
    layer0_outputs(4691) <= '1';
    layer0_outputs(4692) <= b and not a;
    layer0_outputs(4693) <= not (a xor b);
    layer0_outputs(4694) <= a or b;
    layer0_outputs(4695) <= a and b;
    layer0_outputs(4696) <= a;
    layer0_outputs(4697) <= a or b;
    layer0_outputs(4698) <= not b or a;
    layer0_outputs(4699) <= not (a or b);
    layer0_outputs(4700) <= b;
    layer0_outputs(4701) <= not b;
    layer0_outputs(4702) <= not a or b;
    layer0_outputs(4703) <= a or b;
    layer0_outputs(4704) <= a and not b;
    layer0_outputs(4705) <= b and not a;
    layer0_outputs(4706) <= a and b;
    layer0_outputs(4707) <= '0';
    layer0_outputs(4708) <= '0';
    layer0_outputs(4709) <= a;
    layer0_outputs(4710) <= '0';
    layer0_outputs(4711) <= not a or b;
    layer0_outputs(4712) <= not b;
    layer0_outputs(4713) <= not (a or b);
    layer0_outputs(4714) <= not a;
    layer0_outputs(4715) <= a or b;
    layer0_outputs(4716) <= a;
    layer0_outputs(4717) <= b;
    layer0_outputs(4718) <= not (a and b);
    layer0_outputs(4719) <= not b or a;
    layer0_outputs(4720) <= not (a xor b);
    layer0_outputs(4721) <= '0';
    layer0_outputs(4722) <= '1';
    layer0_outputs(4723) <= a and not b;
    layer0_outputs(4724) <= not a or b;
    layer0_outputs(4725) <= not b or a;
    layer0_outputs(4726) <= b;
    layer0_outputs(4727) <= a and not b;
    layer0_outputs(4728) <= '0';
    layer0_outputs(4729) <= a;
    layer0_outputs(4730) <= a and b;
    layer0_outputs(4731) <= not b;
    layer0_outputs(4732) <= not (a or b);
    layer0_outputs(4733) <= b;
    layer0_outputs(4734) <= b;
    layer0_outputs(4735) <= a or b;
    layer0_outputs(4736) <= b;
    layer0_outputs(4737) <= not (a or b);
    layer0_outputs(4738) <= b and not a;
    layer0_outputs(4739) <= a xor b;
    layer0_outputs(4740) <= a or b;
    layer0_outputs(4741) <= not (a or b);
    layer0_outputs(4742) <= a and not b;
    layer0_outputs(4743) <= a and b;
    layer0_outputs(4744) <= not (a or b);
    layer0_outputs(4745) <= b and not a;
    layer0_outputs(4746) <= b;
    layer0_outputs(4747) <= '0';
    layer0_outputs(4748) <= not b;
    layer0_outputs(4749) <= a;
    layer0_outputs(4750) <= not a;
    layer0_outputs(4751) <= not (a xor b);
    layer0_outputs(4752) <= not (a or b);
    layer0_outputs(4753) <= '1';
    layer0_outputs(4754) <= not (a or b);
    layer0_outputs(4755) <= not a or b;
    layer0_outputs(4756) <= a or b;
    layer0_outputs(4757) <= a or b;
    layer0_outputs(4758) <= '0';
    layer0_outputs(4759) <= a xor b;
    layer0_outputs(4760) <= a and b;
    layer0_outputs(4761) <= a and b;
    layer0_outputs(4762) <= b and not a;
    layer0_outputs(4763) <= a or b;
    layer0_outputs(4764) <= b and not a;
    layer0_outputs(4765) <= not a or b;
    layer0_outputs(4766) <= a and b;
    layer0_outputs(4767) <= not a or b;
    layer0_outputs(4768) <= b and not a;
    layer0_outputs(4769) <= a;
    layer0_outputs(4770) <= b and not a;
    layer0_outputs(4771) <= not (a xor b);
    layer0_outputs(4772) <= a;
    layer0_outputs(4773) <= not a or b;
    layer0_outputs(4774) <= not a or b;
    layer0_outputs(4775) <= a or b;
    layer0_outputs(4776) <= a xor b;
    layer0_outputs(4777) <= not b;
    layer0_outputs(4778) <= not a;
    layer0_outputs(4779) <= not (a and b);
    layer0_outputs(4780) <= a xor b;
    layer0_outputs(4781) <= not b or a;
    layer0_outputs(4782) <= b;
    layer0_outputs(4783) <= not a;
    layer0_outputs(4784) <= not (a xor b);
    layer0_outputs(4785) <= not (a or b);
    layer0_outputs(4786) <= '0';
    layer0_outputs(4787) <= b and not a;
    layer0_outputs(4788) <= a xor b;
    layer0_outputs(4789) <= not b;
    layer0_outputs(4790) <= a and not b;
    layer0_outputs(4791) <= b and not a;
    layer0_outputs(4792) <= a xor b;
    layer0_outputs(4793) <= b and not a;
    layer0_outputs(4794) <= a and not b;
    layer0_outputs(4795) <= not a;
    layer0_outputs(4796) <= a or b;
    layer0_outputs(4797) <= a;
    layer0_outputs(4798) <= not b;
    layer0_outputs(4799) <= not a;
    layer0_outputs(4800) <= a;
    layer0_outputs(4801) <= not b or a;
    layer0_outputs(4802) <= b;
    layer0_outputs(4803) <= '0';
    layer0_outputs(4804) <= b;
    layer0_outputs(4805) <= not b or a;
    layer0_outputs(4806) <= a and b;
    layer0_outputs(4807) <= a;
    layer0_outputs(4808) <= a;
    layer0_outputs(4809) <= not (a and b);
    layer0_outputs(4810) <= not (a or b);
    layer0_outputs(4811) <= a xor b;
    layer0_outputs(4812) <= b;
    layer0_outputs(4813) <= '1';
    layer0_outputs(4814) <= a and not b;
    layer0_outputs(4815) <= a xor b;
    layer0_outputs(4816) <= not a or b;
    layer0_outputs(4817) <= not a;
    layer0_outputs(4818) <= a and b;
    layer0_outputs(4819) <= not (a or b);
    layer0_outputs(4820) <= not (a and b);
    layer0_outputs(4821) <= '0';
    layer0_outputs(4822) <= a and not b;
    layer0_outputs(4823) <= a xor b;
    layer0_outputs(4824) <= not b;
    layer0_outputs(4825) <= a xor b;
    layer0_outputs(4826) <= not b;
    layer0_outputs(4827) <= a and not b;
    layer0_outputs(4828) <= not b or a;
    layer0_outputs(4829) <= b;
    layer0_outputs(4830) <= not a or b;
    layer0_outputs(4831) <= '1';
    layer0_outputs(4832) <= b and not a;
    layer0_outputs(4833) <= not b;
    layer0_outputs(4834) <= not (a and b);
    layer0_outputs(4835) <= a xor b;
    layer0_outputs(4836) <= not a;
    layer0_outputs(4837) <= a or b;
    layer0_outputs(4838) <= not b;
    layer0_outputs(4839) <= '1';
    layer0_outputs(4840) <= a;
    layer0_outputs(4841) <= not (a or b);
    layer0_outputs(4842) <= '0';
    layer0_outputs(4843) <= a xor b;
    layer0_outputs(4844) <= a;
    layer0_outputs(4845) <= a xor b;
    layer0_outputs(4846) <= not a or b;
    layer0_outputs(4847) <= not (a xor b);
    layer0_outputs(4848) <= a and not b;
    layer0_outputs(4849) <= not (a or b);
    layer0_outputs(4850) <= b;
    layer0_outputs(4851) <= not (a or b);
    layer0_outputs(4852) <= '1';
    layer0_outputs(4853) <= a or b;
    layer0_outputs(4854) <= a and b;
    layer0_outputs(4855) <= a xor b;
    layer0_outputs(4856) <= not (a or b);
    layer0_outputs(4857) <= '1';
    layer0_outputs(4858) <= a;
    layer0_outputs(4859) <= a;
    layer0_outputs(4860) <= not b;
    layer0_outputs(4861) <= a xor b;
    layer0_outputs(4862) <= not a;
    layer0_outputs(4863) <= not (a xor b);
    layer0_outputs(4864) <= not a;
    layer0_outputs(4865) <= '0';
    layer0_outputs(4866) <= not a or b;
    layer0_outputs(4867) <= b and not a;
    layer0_outputs(4868) <= not (a xor b);
    layer0_outputs(4869) <= not (a xor b);
    layer0_outputs(4870) <= a;
    layer0_outputs(4871) <= a;
    layer0_outputs(4872) <= '1';
    layer0_outputs(4873) <= a or b;
    layer0_outputs(4874) <= a xor b;
    layer0_outputs(4875) <= a xor b;
    layer0_outputs(4876) <= b;
    layer0_outputs(4877) <= not (a or b);
    layer0_outputs(4878) <= not (a or b);
    layer0_outputs(4879) <= a or b;
    layer0_outputs(4880) <= not a or b;
    layer0_outputs(4881) <= not a;
    layer0_outputs(4882) <= a or b;
    layer0_outputs(4883) <= not (a xor b);
    layer0_outputs(4884) <= a and not b;
    layer0_outputs(4885) <= a or b;
    layer0_outputs(4886) <= a and not b;
    layer0_outputs(4887) <= '0';
    layer0_outputs(4888) <= a;
    layer0_outputs(4889) <= not b or a;
    layer0_outputs(4890) <= a;
    layer0_outputs(4891) <= a xor b;
    layer0_outputs(4892) <= not (a xor b);
    layer0_outputs(4893) <= a or b;
    layer0_outputs(4894) <= not (a or b);
    layer0_outputs(4895) <= not (a xor b);
    layer0_outputs(4896) <= a and not b;
    layer0_outputs(4897) <= not (a or b);
    layer0_outputs(4898) <= not a or b;
    layer0_outputs(4899) <= a or b;
    layer0_outputs(4900) <= not b or a;
    layer0_outputs(4901) <= a or b;
    layer0_outputs(4902) <= not a;
    layer0_outputs(4903) <= not a or b;
    layer0_outputs(4904) <= not a;
    layer0_outputs(4905) <= a;
    layer0_outputs(4906) <= not a or b;
    layer0_outputs(4907) <= not (a and b);
    layer0_outputs(4908) <= b and not a;
    layer0_outputs(4909) <= not (a xor b);
    layer0_outputs(4910) <= not (a and b);
    layer0_outputs(4911) <= not a or b;
    layer0_outputs(4912) <= a;
    layer0_outputs(4913) <= a xor b;
    layer0_outputs(4914) <= not b;
    layer0_outputs(4915) <= not b or a;
    layer0_outputs(4916) <= a;
    layer0_outputs(4917) <= not b;
    layer0_outputs(4918) <= b and not a;
    layer0_outputs(4919) <= not a;
    layer0_outputs(4920) <= not a;
    layer0_outputs(4921) <= not a or b;
    layer0_outputs(4922) <= not (a and b);
    layer0_outputs(4923) <= '0';
    layer0_outputs(4924) <= b and not a;
    layer0_outputs(4925) <= not a or b;
    layer0_outputs(4926) <= '0';
    layer0_outputs(4927) <= a;
    layer0_outputs(4928) <= a;
    layer0_outputs(4929) <= '1';
    layer0_outputs(4930) <= not (a and b);
    layer0_outputs(4931) <= b and not a;
    layer0_outputs(4932) <= a xor b;
    layer0_outputs(4933) <= a and b;
    layer0_outputs(4934) <= not a or b;
    layer0_outputs(4935) <= not b;
    layer0_outputs(4936) <= b;
    layer0_outputs(4937) <= a;
    layer0_outputs(4938) <= a and b;
    layer0_outputs(4939) <= not (a or b);
    layer0_outputs(4940) <= not b or a;
    layer0_outputs(4941) <= b;
    layer0_outputs(4942) <= a xor b;
    layer0_outputs(4943) <= '0';
    layer0_outputs(4944) <= not (a xor b);
    layer0_outputs(4945) <= not (a or b);
    layer0_outputs(4946) <= a or b;
    layer0_outputs(4947) <= not a or b;
    layer0_outputs(4948) <= not a or b;
    layer0_outputs(4949) <= a;
    layer0_outputs(4950) <= not b or a;
    layer0_outputs(4951) <= '1';
    layer0_outputs(4952) <= not a or b;
    layer0_outputs(4953) <= not a;
    layer0_outputs(4954) <= not a;
    layer0_outputs(4955) <= not (a or b);
    layer0_outputs(4956) <= a and b;
    layer0_outputs(4957) <= not a;
    layer0_outputs(4958) <= '0';
    layer0_outputs(4959) <= a or b;
    layer0_outputs(4960) <= '0';
    layer0_outputs(4961) <= not (a xor b);
    layer0_outputs(4962) <= b and not a;
    layer0_outputs(4963) <= a;
    layer0_outputs(4964) <= not (a or b);
    layer0_outputs(4965) <= b;
    layer0_outputs(4966) <= not a;
    layer0_outputs(4967) <= not (a and b);
    layer0_outputs(4968) <= not (a or b);
    layer0_outputs(4969) <= b;
    layer0_outputs(4970) <= not (a or b);
    layer0_outputs(4971) <= not (a and b);
    layer0_outputs(4972) <= not b;
    layer0_outputs(4973) <= not b or a;
    layer0_outputs(4974) <= b and not a;
    layer0_outputs(4975) <= a or b;
    layer0_outputs(4976) <= a and b;
    layer0_outputs(4977) <= not a;
    layer0_outputs(4978) <= not a;
    layer0_outputs(4979) <= b;
    layer0_outputs(4980) <= a and not b;
    layer0_outputs(4981) <= a or b;
    layer0_outputs(4982) <= a;
    layer0_outputs(4983) <= b;
    layer0_outputs(4984) <= not b;
    layer0_outputs(4985) <= b;
    layer0_outputs(4986) <= a or b;
    layer0_outputs(4987) <= a or b;
    layer0_outputs(4988) <= not a;
    layer0_outputs(4989) <= not b or a;
    layer0_outputs(4990) <= a or b;
    layer0_outputs(4991) <= a and not b;
    layer0_outputs(4992) <= '1';
    layer0_outputs(4993) <= '1';
    layer0_outputs(4994) <= not a;
    layer0_outputs(4995) <= a or b;
    layer0_outputs(4996) <= a or b;
    layer0_outputs(4997) <= not b;
    layer0_outputs(4998) <= b;
    layer0_outputs(4999) <= not (a and b);
    layer0_outputs(5000) <= not b;
    layer0_outputs(5001) <= '0';
    layer0_outputs(5002) <= not b;
    layer0_outputs(5003) <= a or b;
    layer0_outputs(5004) <= not a or b;
    layer0_outputs(5005) <= a or b;
    layer0_outputs(5006) <= not b;
    layer0_outputs(5007) <= a;
    layer0_outputs(5008) <= not (a or b);
    layer0_outputs(5009) <= not (a xor b);
    layer0_outputs(5010) <= a xor b;
    layer0_outputs(5011) <= not (a and b);
    layer0_outputs(5012) <= a xor b;
    layer0_outputs(5013) <= a xor b;
    layer0_outputs(5014) <= a;
    layer0_outputs(5015) <= not a;
    layer0_outputs(5016) <= not a or b;
    layer0_outputs(5017) <= not (a xor b);
    layer0_outputs(5018) <= a;
    layer0_outputs(5019) <= not a;
    layer0_outputs(5020) <= b and not a;
    layer0_outputs(5021) <= not a;
    layer0_outputs(5022) <= not (a and b);
    layer0_outputs(5023) <= not (a xor b);
    layer0_outputs(5024) <= a xor b;
    layer0_outputs(5025) <= a or b;
    layer0_outputs(5026) <= not b or a;
    layer0_outputs(5027) <= not a or b;
    layer0_outputs(5028) <= not (a xor b);
    layer0_outputs(5029) <= '1';
    layer0_outputs(5030) <= a or b;
    layer0_outputs(5031) <= not (a and b);
    layer0_outputs(5032) <= a;
    layer0_outputs(5033) <= not a or b;
    layer0_outputs(5034) <= not (a or b);
    layer0_outputs(5035) <= b;
    layer0_outputs(5036) <= not (a or b);
    layer0_outputs(5037) <= not a;
    layer0_outputs(5038) <= not b or a;
    layer0_outputs(5039) <= '0';
    layer0_outputs(5040) <= not (a and b);
    layer0_outputs(5041) <= not a or b;
    layer0_outputs(5042) <= b;
    layer0_outputs(5043) <= not (a xor b);
    layer0_outputs(5044) <= a xor b;
    layer0_outputs(5045) <= a xor b;
    layer0_outputs(5046) <= not (a and b);
    layer0_outputs(5047) <= '1';
    layer0_outputs(5048) <= a or b;
    layer0_outputs(5049) <= b;
    layer0_outputs(5050) <= b;
    layer0_outputs(5051) <= b and not a;
    layer0_outputs(5052) <= a or b;
    layer0_outputs(5053) <= not b;
    layer0_outputs(5054) <= a or b;
    layer0_outputs(5055) <= a xor b;
    layer0_outputs(5056) <= a;
    layer0_outputs(5057) <= not b;
    layer0_outputs(5058) <= not (a or b);
    layer0_outputs(5059) <= a;
    layer0_outputs(5060) <= not b;
    layer0_outputs(5061) <= a or b;
    layer0_outputs(5062) <= a and b;
    layer0_outputs(5063) <= not (a xor b);
    layer0_outputs(5064) <= not a or b;
    layer0_outputs(5065) <= not b or a;
    layer0_outputs(5066) <= not a;
    layer0_outputs(5067) <= a xor b;
    layer0_outputs(5068) <= not a;
    layer0_outputs(5069) <= not (a or b);
    layer0_outputs(5070) <= not (a or b);
    layer0_outputs(5071) <= b;
    layer0_outputs(5072) <= a;
    layer0_outputs(5073) <= a;
    layer0_outputs(5074) <= b;
    layer0_outputs(5075) <= a;
    layer0_outputs(5076) <= not a;
    layer0_outputs(5077) <= not a;
    layer0_outputs(5078) <= not a or b;
    layer0_outputs(5079) <= not b;
    layer0_outputs(5080) <= b;
    layer0_outputs(5081) <= not b;
    layer0_outputs(5082) <= '0';
    layer0_outputs(5083) <= '0';
    layer0_outputs(5084) <= a;
    layer0_outputs(5085) <= a and b;
    layer0_outputs(5086) <= not b or a;
    layer0_outputs(5087) <= a or b;
    layer0_outputs(5088) <= b and not a;
    layer0_outputs(5089) <= a and b;
    layer0_outputs(5090) <= '0';
    layer0_outputs(5091) <= a and b;
    layer0_outputs(5092) <= not a or b;
    layer0_outputs(5093) <= a;
    layer0_outputs(5094) <= not b or a;
    layer0_outputs(5095) <= not (a xor b);
    layer0_outputs(5096) <= not a;
    layer0_outputs(5097) <= not a or b;
    layer0_outputs(5098) <= not (a or b);
    layer0_outputs(5099) <= a or b;
    layer0_outputs(5100) <= not (a or b);
    layer0_outputs(5101) <= a xor b;
    layer0_outputs(5102) <= not (a xor b);
    layer0_outputs(5103) <= b and not a;
    layer0_outputs(5104) <= a;
    layer0_outputs(5105) <= b and not a;
    layer0_outputs(5106) <= a and not b;
    layer0_outputs(5107) <= not b or a;
    layer0_outputs(5108) <= b;
    layer0_outputs(5109) <= not a;
    layer0_outputs(5110) <= a and not b;
    layer0_outputs(5111) <= b;
    layer0_outputs(5112) <= a xor b;
    layer0_outputs(5113) <= not b or a;
    layer0_outputs(5114) <= not b or a;
    layer0_outputs(5115) <= b;
    layer0_outputs(5116) <= not a;
    layer0_outputs(5117) <= not (a and b);
    layer0_outputs(5118) <= not a or b;
    layer0_outputs(5119) <= a or b;
    layer0_outputs(5120) <= not a;
    layer0_outputs(5121) <= not b or a;
    layer0_outputs(5122) <= '1';
    layer0_outputs(5123) <= not (a or b);
    layer0_outputs(5124) <= not a or b;
    layer0_outputs(5125) <= a or b;
    layer0_outputs(5126) <= not (a and b);
    layer0_outputs(5127) <= a;
    layer0_outputs(5128) <= not a;
    layer0_outputs(5129) <= not (a or b);
    layer0_outputs(5130) <= a xor b;
    layer0_outputs(5131) <= a or b;
    layer0_outputs(5132) <= a;
    layer0_outputs(5133) <= a or b;
    layer0_outputs(5134) <= not a or b;
    layer0_outputs(5135) <= a;
    layer0_outputs(5136) <= not a;
    layer0_outputs(5137) <= a and b;
    layer0_outputs(5138) <= not (a or b);
    layer0_outputs(5139) <= a xor b;
    layer0_outputs(5140) <= not b or a;
    layer0_outputs(5141) <= a;
    layer0_outputs(5142) <= a xor b;
    layer0_outputs(5143) <= b and not a;
    layer0_outputs(5144) <= a and b;
    layer0_outputs(5145) <= b and not a;
    layer0_outputs(5146) <= not b;
    layer0_outputs(5147) <= not (a and b);
    layer0_outputs(5148) <= not (a xor b);
    layer0_outputs(5149) <= not a;
    layer0_outputs(5150) <= not b;
    layer0_outputs(5151) <= a or b;
    layer0_outputs(5152) <= not (a or b);
    layer0_outputs(5153) <= not (a xor b);
    layer0_outputs(5154) <= a xor b;
    layer0_outputs(5155) <= a xor b;
    layer0_outputs(5156) <= not (a xor b);
    layer0_outputs(5157) <= not a or b;
    layer0_outputs(5158) <= '1';
    layer0_outputs(5159) <= a xor b;
    layer0_outputs(5160) <= not (a and b);
    layer0_outputs(5161) <= b;
    layer0_outputs(5162) <= not (a xor b);
    layer0_outputs(5163) <= a and not b;
    layer0_outputs(5164) <= not b;
    layer0_outputs(5165) <= not (a or b);
    layer0_outputs(5166) <= a xor b;
    layer0_outputs(5167) <= not (a xor b);
    layer0_outputs(5168) <= a xor b;
    layer0_outputs(5169) <= a xor b;
    layer0_outputs(5170) <= not a;
    layer0_outputs(5171) <= not b;
    layer0_outputs(5172) <= a and b;
    layer0_outputs(5173) <= a xor b;
    layer0_outputs(5174) <= a;
    layer0_outputs(5175) <= a and not b;
    layer0_outputs(5176) <= '0';
    layer0_outputs(5177) <= not b or a;
    layer0_outputs(5178) <= b and not a;
    layer0_outputs(5179) <= b;
    layer0_outputs(5180) <= not (a and b);
    layer0_outputs(5181) <= a or b;
    layer0_outputs(5182) <= not a;
    layer0_outputs(5183) <= not (a or b);
    layer0_outputs(5184) <= not b;
    layer0_outputs(5185) <= '0';
    layer0_outputs(5186) <= not b or a;
    layer0_outputs(5187) <= not a;
    layer0_outputs(5188) <= a and b;
    layer0_outputs(5189) <= not (a xor b);
    layer0_outputs(5190) <= not b or a;
    layer0_outputs(5191) <= not (a and b);
    layer0_outputs(5192) <= a and not b;
    layer0_outputs(5193) <= not b or a;
    layer0_outputs(5194) <= a and b;
    layer0_outputs(5195) <= a and b;
    layer0_outputs(5196) <= a;
    layer0_outputs(5197) <= b and not a;
    layer0_outputs(5198) <= not (a or b);
    layer0_outputs(5199) <= a and not b;
    layer0_outputs(5200) <= not b;
    layer0_outputs(5201) <= not a;
    layer0_outputs(5202) <= not b or a;
    layer0_outputs(5203) <= b and not a;
    layer0_outputs(5204) <= a or b;
    layer0_outputs(5205) <= not a or b;
    layer0_outputs(5206) <= a and not b;
    layer0_outputs(5207) <= a and b;
    layer0_outputs(5208) <= not (a xor b);
    layer0_outputs(5209) <= b and not a;
    layer0_outputs(5210) <= not b;
    layer0_outputs(5211) <= not a;
    layer0_outputs(5212) <= a or b;
    layer0_outputs(5213) <= '0';
    layer0_outputs(5214) <= not b or a;
    layer0_outputs(5215) <= a and b;
    layer0_outputs(5216) <= not b;
    layer0_outputs(5217) <= a and not b;
    layer0_outputs(5218) <= not (a or b);
    layer0_outputs(5219) <= b and not a;
    layer0_outputs(5220) <= not b or a;
    layer0_outputs(5221) <= not (a or b);
    layer0_outputs(5222) <= not b;
    layer0_outputs(5223) <= not b;
    layer0_outputs(5224) <= not (a and b);
    layer0_outputs(5225) <= not (a and b);
    layer0_outputs(5226) <= not (a xor b);
    layer0_outputs(5227) <= a xor b;
    layer0_outputs(5228) <= a xor b;
    layer0_outputs(5229) <= a;
    layer0_outputs(5230) <= not b or a;
    layer0_outputs(5231) <= a;
    layer0_outputs(5232) <= b;
    layer0_outputs(5233) <= a xor b;
    layer0_outputs(5234) <= not b or a;
    layer0_outputs(5235) <= b;
    layer0_outputs(5236) <= not (a and b);
    layer0_outputs(5237) <= not a;
    layer0_outputs(5238) <= not a or b;
    layer0_outputs(5239) <= a and not b;
    layer0_outputs(5240) <= not b or a;
    layer0_outputs(5241) <= '1';
    layer0_outputs(5242) <= a;
    layer0_outputs(5243) <= not b or a;
    layer0_outputs(5244) <= not (a or b);
    layer0_outputs(5245) <= not (a and b);
    layer0_outputs(5246) <= a xor b;
    layer0_outputs(5247) <= not a;
    layer0_outputs(5248) <= not a;
    layer0_outputs(5249) <= not a or b;
    layer0_outputs(5250) <= not a;
    layer0_outputs(5251) <= b and not a;
    layer0_outputs(5252) <= not (a or b);
    layer0_outputs(5253) <= a or b;
    layer0_outputs(5254) <= b and not a;
    layer0_outputs(5255) <= a or b;
    layer0_outputs(5256) <= not b;
    layer0_outputs(5257) <= b;
    layer0_outputs(5258) <= not a;
    layer0_outputs(5259) <= b;
    layer0_outputs(5260) <= not a or b;
    layer0_outputs(5261) <= not (a and b);
    layer0_outputs(5262) <= not a;
    layer0_outputs(5263) <= not b;
    layer0_outputs(5264) <= a;
    layer0_outputs(5265) <= not (a and b);
    layer0_outputs(5266) <= not a;
    layer0_outputs(5267) <= b and not a;
    layer0_outputs(5268) <= a;
    layer0_outputs(5269) <= '1';
    layer0_outputs(5270) <= '0';
    layer0_outputs(5271) <= not (a or b);
    layer0_outputs(5272) <= b;
    layer0_outputs(5273) <= a and not b;
    layer0_outputs(5274) <= not a;
    layer0_outputs(5275) <= not b or a;
    layer0_outputs(5276) <= a and b;
    layer0_outputs(5277) <= not b or a;
    layer0_outputs(5278) <= a xor b;
    layer0_outputs(5279) <= a and b;
    layer0_outputs(5280) <= '0';
    layer0_outputs(5281) <= not b;
    layer0_outputs(5282) <= not a;
    layer0_outputs(5283) <= not b or a;
    layer0_outputs(5284) <= not a;
    layer0_outputs(5285) <= not (a or b);
    layer0_outputs(5286) <= a or b;
    layer0_outputs(5287) <= not (a xor b);
    layer0_outputs(5288) <= not b;
    layer0_outputs(5289) <= '0';
    layer0_outputs(5290) <= not b;
    layer0_outputs(5291) <= not (a or b);
    layer0_outputs(5292) <= a or b;
    layer0_outputs(5293) <= '0';
    layer0_outputs(5294) <= not a;
    layer0_outputs(5295) <= a;
    layer0_outputs(5296) <= b;
    layer0_outputs(5297) <= b;
    layer0_outputs(5298) <= not b;
    layer0_outputs(5299) <= a;
    layer0_outputs(5300) <= '1';
    layer0_outputs(5301) <= b;
    layer0_outputs(5302) <= not b;
    layer0_outputs(5303) <= a xor b;
    layer0_outputs(5304) <= b and not a;
    layer0_outputs(5305) <= b;
    layer0_outputs(5306) <= not b or a;
    layer0_outputs(5307) <= a xor b;
    layer0_outputs(5308) <= not (a and b);
    layer0_outputs(5309) <= '0';
    layer0_outputs(5310) <= not (a and b);
    layer0_outputs(5311) <= b and not a;
    layer0_outputs(5312) <= not a;
    layer0_outputs(5313) <= a xor b;
    layer0_outputs(5314) <= not b;
    layer0_outputs(5315) <= a;
    layer0_outputs(5316) <= b;
    layer0_outputs(5317) <= not b or a;
    layer0_outputs(5318) <= a xor b;
    layer0_outputs(5319) <= not (a xor b);
    layer0_outputs(5320) <= b and not a;
    layer0_outputs(5321) <= a and not b;
    layer0_outputs(5322) <= not a;
    layer0_outputs(5323) <= not (a or b);
    layer0_outputs(5324) <= a and not b;
    layer0_outputs(5325) <= b and not a;
    layer0_outputs(5326) <= a;
    layer0_outputs(5327) <= '1';
    layer0_outputs(5328) <= '0';
    layer0_outputs(5329) <= not b;
    layer0_outputs(5330) <= '0';
    layer0_outputs(5331) <= not b;
    layer0_outputs(5332) <= not a or b;
    layer0_outputs(5333) <= b and not a;
    layer0_outputs(5334) <= b;
    layer0_outputs(5335) <= a and not b;
    layer0_outputs(5336) <= not b;
    layer0_outputs(5337) <= not b;
    layer0_outputs(5338) <= a or b;
    layer0_outputs(5339) <= not a;
    layer0_outputs(5340) <= not b;
    layer0_outputs(5341) <= not a or b;
    layer0_outputs(5342) <= not (a or b);
    layer0_outputs(5343) <= not b;
    layer0_outputs(5344) <= '1';
    layer0_outputs(5345) <= a and b;
    layer0_outputs(5346) <= a xor b;
    layer0_outputs(5347) <= a and not b;
    layer0_outputs(5348) <= not b;
    layer0_outputs(5349) <= a and not b;
    layer0_outputs(5350) <= not (a xor b);
    layer0_outputs(5351) <= not (a and b);
    layer0_outputs(5352) <= b and not a;
    layer0_outputs(5353) <= b and not a;
    layer0_outputs(5354) <= a or b;
    layer0_outputs(5355) <= b and not a;
    layer0_outputs(5356) <= not (a and b);
    layer0_outputs(5357) <= b and not a;
    layer0_outputs(5358) <= not (a or b);
    layer0_outputs(5359) <= b;
    layer0_outputs(5360) <= a and b;
    layer0_outputs(5361) <= b;
    layer0_outputs(5362) <= '0';
    layer0_outputs(5363) <= a;
    layer0_outputs(5364) <= not b;
    layer0_outputs(5365) <= not b or a;
    layer0_outputs(5366) <= b;
    layer0_outputs(5367) <= a and not b;
    layer0_outputs(5368) <= '0';
    layer0_outputs(5369) <= b;
    layer0_outputs(5370) <= '1';
    layer0_outputs(5371) <= not (a xor b);
    layer0_outputs(5372) <= not b;
    layer0_outputs(5373) <= not (a and b);
    layer0_outputs(5374) <= b and not a;
    layer0_outputs(5375) <= not a;
    layer0_outputs(5376) <= not (a xor b);
    layer0_outputs(5377) <= '0';
    layer0_outputs(5378) <= not (a or b);
    layer0_outputs(5379) <= b and not a;
    layer0_outputs(5380) <= a and not b;
    layer0_outputs(5381) <= not b;
    layer0_outputs(5382) <= not (a and b);
    layer0_outputs(5383) <= a or b;
    layer0_outputs(5384) <= a and b;
    layer0_outputs(5385) <= b and not a;
    layer0_outputs(5386) <= '0';
    layer0_outputs(5387) <= a or b;
    layer0_outputs(5388) <= a and b;
    layer0_outputs(5389) <= not (a and b);
    layer0_outputs(5390) <= b and not a;
    layer0_outputs(5391) <= not a;
    layer0_outputs(5392) <= a or b;
    layer0_outputs(5393) <= not b;
    layer0_outputs(5394) <= not b or a;
    layer0_outputs(5395) <= not (a or b);
    layer0_outputs(5396) <= not (a or b);
    layer0_outputs(5397) <= b and not a;
    layer0_outputs(5398) <= a xor b;
    layer0_outputs(5399) <= a and b;
    layer0_outputs(5400) <= a xor b;
    layer0_outputs(5401) <= b;
    layer0_outputs(5402) <= not a;
    layer0_outputs(5403) <= a;
    layer0_outputs(5404) <= not (a xor b);
    layer0_outputs(5405) <= a or b;
    layer0_outputs(5406) <= a xor b;
    layer0_outputs(5407) <= a;
    layer0_outputs(5408) <= b;
    layer0_outputs(5409) <= b and not a;
    layer0_outputs(5410) <= not a or b;
    layer0_outputs(5411) <= b and not a;
    layer0_outputs(5412) <= a xor b;
    layer0_outputs(5413) <= a or b;
    layer0_outputs(5414) <= a or b;
    layer0_outputs(5415) <= a;
    layer0_outputs(5416) <= a;
    layer0_outputs(5417) <= not (a and b);
    layer0_outputs(5418) <= not (a xor b);
    layer0_outputs(5419) <= not b;
    layer0_outputs(5420) <= not a;
    layer0_outputs(5421) <= a or b;
    layer0_outputs(5422) <= a xor b;
    layer0_outputs(5423) <= not (a and b);
    layer0_outputs(5424) <= '0';
    layer0_outputs(5425) <= not b or a;
    layer0_outputs(5426) <= not (a or b);
    layer0_outputs(5427) <= not a or b;
    layer0_outputs(5428) <= '0';
    layer0_outputs(5429) <= not (a xor b);
    layer0_outputs(5430) <= not (a and b);
    layer0_outputs(5431) <= not b;
    layer0_outputs(5432) <= '0';
    layer0_outputs(5433) <= a or b;
    layer0_outputs(5434) <= a or b;
    layer0_outputs(5435) <= '1';
    layer0_outputs(5436) <= a and not b;
    layer0_outputs(5437) <= b;
    layer0_outputs(5438) <= a xor b;
    layer0_outputs(5439) <= not b or a;
    layer0_outputs(5440) <= not a;
    layer0_outputs(5441) <= not (a and b);
    layer0_outputs(5442) <= not a;
    layer0_outputs(5443) <= a;
    layer0_outputs(5444) <= a;
    layer0_outputs(5445) <= a;
    layer0_outputs(5446) <= not (a or b);
    layer0_outputs(5447) <= not (a or b);
    layer0_outputs(5448) <= not (a or b);
    layer0_outputs(5449) <= not b or a;
    layer0_outputs(5450) <= not b;
    layer0_outputs(5451) <= a;
    layer0_outputs(5452) <= b;
    layer0_outputs(5453) <= not (a xor b);
    layer0_outputs(5454) <= a or b;
    layer0_outputs(5455) <= '1';
    layer0_outputs(5456) <= not (a or b);
    layer0_outputs(5457) <= a and not b;
    layer0_outputs(5458) <= '0';
    layer0_outputs(5459) <= not b or a;
    layer0_outputs(5460) <= a and not b;
    layer0_outputs(5461) <= b and not a;
    layer0_outputs(5462) <= not a;
    layer0_outputs(5463) <= b and not a;
    layer0_outputs(5464) <= a xor b;
    layer0_outputs(5465) <= b and not a;
    layer0_outputs(5466) <= not (a and b);
    layer0_outputs(5467) <= a xor b;
    layer0_outputs(5468) <= b;
    layer0_outputs(5469) <= a xor b;
    layer0_outputs(5470) <= b;
    layer0_outputs(5471) <= not (a or b);
    layer0_outputs(5472) <= not a;
    layer0_outputs(5473) <= not b or a;
    layer0_outputs(5474) <= not (a xor b);
    layer0_outputs(5475) <= a xor b;
    layer0_outputs(5476) <= a and not b;
    layer0_outputs(5477) <= not b or a;
    layer0_outputs(5478) <= b and not a;
    layer0_outputs(5479) <= not b or a;
    layer0_outputs(5480) <= a and not b;
    layer0_outputs(5481) <= '1';
    layer0_outputs(5482) <= '1';
    layer0_outputs(5483) <= not a;
    layer0_outputs(5484) <= a and not b;
    layer0_outputs(5485) <= not a or b;
    layer0_outputs(5486) <= not (a and b);
    layer0_outputs(5487) <= not a;
    layer0_outputs(5488) <= not a or b;
    layer0_outputs(5489) <= not a;
    layer0_outputs(5490) <= not b or a;
    layer0_outputs(5491) <= b and not a;
    layer0_outputs(5492) <= '1';
    layer0_outputs(5493) <= not a;
    layer0_outputs(5494) <= a and not b;
    layer0_outputs(5495) <= not b;
    layer0_outputs(5496) <= not a or b;
    layer0_outputs(5497) <= a or b;
    layer0_outputs(5498) <= a or b;
    layer0_outputs(5499) <= a and not b;
    layer0_outputs(5500) <= a and not b;
    layer0_outputs(5501) <= a xor b;
    layer0_outputs(5502) <= b and not a;
    layer0_outputs(5503) <= '0';
    layer0_outputs(5504) <= not b or a;
    layer0_outputs(5505) <= a xor b;
    layer0_outputs(5506) <= not (a xor b);
    layer0_outputs(5507) <= a;
    layer0_outputs(5508) <= not b;
    layer0_outputs(5509) <= a and b;
    layer0_outputs(5510) <= not (a xor b);
    layer0_outputs(5511) <= not (a or b);
    layer0_outputs(5512) <= b;
    layer0_outputs(5513) <= not a or b;
    layer0_outputs(5514) <= not b or a;
    layer0_outputs(5515) <= not a or b;
    layer0_outputs(5516) <= a and not b;
    layer0_outputs(5517) <= b;
    layer0_outputs(5518) <= not b or a;
    layer0_outputs(5519) <= not (a or b);
    layer0_outputs(5520) <= not b;
    layer0_outputs(5521) <= not (a or b);
    layer0_outputs(5522) <= not b;
    layer0_outputs(5523) <= not (a and b);
    layer0_outputs(5524) <= a or b;
    layer0_outputs(5525) <= not (a or b);
    layer0_outputs(5526) <= not (a or b);
    layer0_outputs(5527) <= b and not a;
    layer0_outputs(5528) <= a;
    layer0_outputs(5529) <= a;
    layer0_outputs(5530) <= b and not a;
    layer0_outputs(5531) <= not (a xor b);
    layer0_outputs(5532) <= a and b;
    layer0_outputs(5533) <= a;
    layer0_outputs(5534) <= a and b;
    layer0_outputs(5535) <= not (a xor b);
    layer0_outputs(5536) <= not (a or b);
    layer0_outputs(5537) <= not b;
    layer0_outputs(5538) <= not b or a;
    layer0_outputs(5539) <= a or b;
    layer0_outputs(5540) <= not (a and b);
    layer0_outputs(5541) <= a or b;
    layer0_outputs(5542) <= '0';
    layer0_outputs(5543) <= a;
    layer0_outputs(5544) <= b and not a;
    layer0_outputs(5545) <= not a or b;
    layer0_outputs(5546) <= b and not a;
    layer0_outputs(5547) <= not b or a;
    layer0_outputs(5548) <= b and not a;
    layer0_outputs(5549) <= not a;
    layer0_outputs(5550) <= not b or a;
    layer0_outputs(5551) <= not a;
    layer0_outputs(5552) <= a and b;
    layer0_outputs(5553) <= a xor b;
    layer0_outputs(5554) <= not (a xor b);
    layer0_outputs(5555) <= not (a or b);
    layer0_outputs(5556) <= not b or a;
    layer0_outputs(5557) <= a;
    layer0_outputs(5558) <= not a;
    layer0_outputs(5559) <= not b or a;
    layer0_outputs(5560) <= not a or b;
    layer0_outputs(5561) <= not (a or b);
    layer0_outputs(5562) <= b;
    layer0_outputs(5563) <= b;
    layer0_outputs(5564) <= a xor b;
    layer0_outputs(5565) <= not b or a;
    layer0_outputs(5566) <= '0';
    layer0_outputs(5567) <= a and b;
    layer0_outputs(5568) <= a;
    layer0_outputs(5569) <= not a or b;
    layer0_outputs(5570) <= not a or b;
    layer0_outputs(5571) <= a xor b;
    layer0_outputs(5572) <= '1';
    layer0_outputs(5573) <= b;
    layer0_outputs(5574) <= not b;
    layer0_outputs(5575) <= b;
    layer0_outputs(5576) <= not (a or b);
    layer0_outputs(5577) <= '0';
    layer0_outputs(5578) <= a;
    layer0_outputs(5579) <= a and not b;
    layer0_outputs(5580) <= b and not a;
    layer0_outputs(5581) <= a;
    layer0_outputs(5582) <= not b or a;
    layer0_outputs(5583) <= not b or a;
    layer0_outputs(5584) <= a or b;
    layer0_outputs(5585) <= not (a and b);
    layer0_outputs(5586) <= not (a or b);
    layer0_outputs(5587) <= a or b;
    layer0_outputs(5588) <= a;
    layer0_outputs(5589) <= a;
    layer0_outputs(5590) <= not b or a;
    layer0_outputs(5591) <= '0';
    layer0_outputs(5592) <= not b;
    layer0_outputs(5593) <= b and not a;
    layer0_outputs(5594) <= a xor b;
    layer0_outputs(5595) <= a and not b;
    layer0_outputs(5596) <= not (a or b);
    layer0_outputs(5597) <= b and not a;
    layer0_outputs(5598) <= a xor b;
    layer0_outputs(5599) <= b and not a;
    layer0_outputs(5600) <= not b;
    layer0_outputs(5601) <= not a;
    layer0_outputs(5602) <= not (a or b);
    layer0_outputs(5603) <= a and b;
    layer0_outputs(5604) <= b and not a;
    layer0_outputs(5605) <= '1';
    layer0_outputs(5606) <= not (a xor b);
    layer0_outputs(5607) <= a;
    layer0_outputs(5608) <= '0';
    layer0_outputs(5609) <= a or b;
    layer0_outputs(5610) <= b;
    layer0_outputs(5611) <= not b;
    layer0_outputs(5612) <= a and not b;
    layer0_outputs(5613) <= a or b;
    layer0_outputs(5614) <= a or b;
    layer0_outputs(5615) <= not b or a;
    layer0_outputs(5616) <= b and not a;
    layer0_outputs(5617) <= b;
    layer0_outputs(5618) <= not a or b;
    layer0_outputs(5619) <= not a;
    layer0_outputs(5620) <= a;
    layer0_outputs(5621) <= a and not b;
    layer0_outputs(5622) <= a or b;
    layer0_outputs(5623) <= a xor b;
    layer0_outputs(5624) <= b and not a;
    layer0_outputs(5625) <= a;
    layer0_outputs(5626) <= not b or a;
    layer0_outputs(5627) <= b and not a;
    layer0_outputs(5628) <= a;
    layer0_outputs(5629) <= a or b;
    layer0_outputs(5630) <= '0';
    layer0_outputs(5631) <= not (a or b);
    layer0_outputs(5632) <= not b or a;
    layer0_outputs(5633) <= a or b;
    layer0_outputs(5634) <= a xor b;
    layer0_outputs(5635) <= not a;
    layer0_outputs(5636) <= not b or a;
    layer0_outputs(5637) <= a and not b;
    layer0_outputs(5638) <= not (a xor b);
    layer0_outputs(5639) <= b;
    layer0_outputs(5640) <= not (a and b);
    layer0_outputs(5641) <= '1';
    layer0_outputs(5642) <= a and b;
    layer0_outputs(5643) <= a xor b;
    layer0_outputs(5644) <= a or b;
    layer0_outputs(5645) <= a or b;
    layer0_outputs(5646) <= not (a or b);
    layer0_outputs(5647) <= b and not a;
    layer0_outputs(5648) <= not a;
    layer0_outputs(5649) <= not b or a;
    layer0_outputs(5650) <= b and not a;
    layer0_outputs(5651) <= not (a and b);
    layer0_outputs(5652) <= not b or a;
    layer0_outputs(5653) <= a and not b;
    layer0_outputs(5654) <= not (a or b);
    layer0_outputs(5655) <= '1';
    layer0_outputs(5656) <= a and not b;
    layer0_outputs(5657) <= a xor b;
    layer0_outputs(5658) <= '1';
    layer0_outputs(5659) <= a or b;
    layer0_outputs(5660) <= not a or b;
    layer0_outputs(5661) <= a and not b;
    layer0_outputs(5662) <= not (a and b);
    layer0_outputs(5663) <= a xor b;
    layer0_outputs(5664) <= not (a xor b);
    layer0_outputs(5665) <= not b or a;
    layer0_outputs(5666) <= not (a and b);
    layer0_outputs(5667) <= not a or b;
    layer0_outputs(5668) <= a or b;
    layer0_outputs(5669) <= not a;
    layer0_outputs(5670) <= not (a xor b);
    layer0_outputs(5671) <= a or b;
    layer0_outputs(5672) <= not b;
    layer0_outputs(5673) <= not a;
    layer0_outputs(5674) <= not a or b;
    layer0_outputs(5675) <= a xor b;
    layer0_outputs(5676) <= not b or a;
    layer0_outputs(5677) <= a;
    layer0_outputs(5678) <= not b or a;
    layer0_outputs(5679) <= a and not b;
    layer0_outputs(5680) <= not (a or b);
    layer0_outputs(5681) <= not (a or b);
    layer0_outputs(5682) <= not b;
    layer0_outputs(5683) <= a or b;
    layer0_outputs(5684) <= not (a and b);
    layer0_outputs(5685) <= a and not b;
    layer0_outputs(5686) <= not (a xor b);
    layer0_outputs(5687) <= b and not a;
    layer0_outputs(5688) <= not b;
    layer0_outputs(5689) <= a;
    layer0_outputs(5690) <= not a;
    layer0_outputs(5691) <= '1';
    layer0_outputs(5692) <= a xor b;
    layer0_outputs(5693) <= a;
    layer0_outputs(5694) <= a and b;
    layer0_outputs(5695) <= a xor b;
    layer0_outputs(5696) <= b;
    layer0_outputs(5697) <= a or b;
    layer0_outputs(5698) <= a and b;
    layer0_outputs(5699) <= a or b;
    layer0_outputs(5700) <= a or b;
    layer0_outputs(5701) <= '0';
    layer0_outputs(5702) <= not b or a;
    layer0_outputs(5703) <= a xor b;
    layer0_outputs(5704) <= a or b;
    layer0_outputs(5705) <= not (a or b);
    layer0_outputs(5706) <= not (a xor b);
    layer0_outputs(5707) <= not (a or b);
    layer0_outputs(5708) <= '1';
    layer0_outputs(5709) <= '1';
    layer0_outputs(5710) <= a xor b;
    layer0_outputs(5711) <= not (a xor b);
    layer0_outputs(5712) <= a or b;
    layer0_outputs(5713) <= not b or a;
    layer0_outputs(5714) <= not (a xor b);
    layer0_outputs(5715) <= not a;
    layer0_outputs(5716) <= '0';
    layer0_outputs(5717) <= a and not b;
    layer0_outputs(5718) <= not b;
    layer0_outputs(5719) <= a and b;
    layer0_outputs(5720) <= a;
    layer0_outputs(5721) <= '1';
    layer0_outputs(5722) <= a and not b;
    layer0_outputs(5723) <= '0';
    layer0_outputs(5724) <= not (a xor b);
    layer0_outputs(5725) <= not (a and b);
    layer0_outputs(5726) <= not (a or b);
    layer0_outputs(5727) <= not a or b;
    layer0_outputs(5728) <= not b;
    layer0_outputs(5729) <= a or b;
    layer0_outputs(5730) <= b and not a;
    layer0_outputs(5731) <= a xor b;
    layer0_outputs(5732) <= not a or b;
    layer0_outputs(5733) <= b and not a;
    layer0_outputs(5734) <= not (a or b);
    layer0_outputs(5735) <= not b or a;
    layer0_outputs(5736) <= a or b;
    layer0_outputs(5737) <= a and not b;
    layer0_outputs(5738) <= a and not b;
    layer0_outputs(5739) <= not (a xor b);
    layer0_outputs(5740) <= b;
    layer0_outputs(5741) <= not b or a;
    layer0_outputs(5742) <= a xor b;
    layer0_outputs(5743) <= not (a and b);
    layer0_outputs(5744) <= not (a or b);
    layer0_outputs(5745) <= a and not b;
    layer0_outputs(5746) <= b;
    layer0_outputs(5747) <= b and not a;
    layer0_outputs(5748) <= not b;
    layer0_outputs(5749) <= a and not b;
    layer0_outputs(5750) <= a and not b;
    layer0_outputs(5751) <= a xor b;
    layer0_outputs(5752) <= a xor b;
    layer0_outputs(5753) <= '0';
    layer0_outputs(5754) <= not b;
    layer0_outputs(5755) <= not b or a;
    layer0_outputs(5756) <= not (a or b);
    layer0_outputs(5757) <= a and not b;
    layer0_outputs(5758) <= a xor b;
    layer0_outputs(5759) <= not (a and b);
    layer0_outputs(5760) <= b and not a;
    layer0_outputs(5761) <= a;
    layer0_outputs(5762) <= a;
    layer0_outputs(5763) <= not b or a;
    layer0_outputs(5764) <= a or b;
    layer0_outputs(5765) <= a or b;
    layer0_outputs(5766) <= not (a or b);
    layer0_outputs(5767) <= b;
    layer0_outputs(5768) <= not (a or b);
    layer0_outputs(5769) <= not b or a;
    layer0_outputs(5770) <= '1';
    layer0_outputs(5771) <= not (a xor b);
    layer0_outputs(5772) <= a or b;
    layer0_outputs(5773) <= not (a or b);
    layer0_outputs(5774) <= not (a and b);
    layer0_outputs(5775) <= not b;
    layer0_outputs(5776) <= a and not b;
    layer0_outputs(5777) <= not (a xor b);
    layer0_outputs(5778) <= not a;
    layer0_outputs(5779) <= not (a or b);
    layer0_outputs(5780) <= a or b;
    layer0_outputs(5781) <= not (a or b);
    layer0_outputs(5782) <= a;
    layer0_outputs(5783) <= not b;
    layer0_outputs(5784) <= not a;
    layer0_outputs(5785) <= b;
    layer0_outputs(5786) <= not (a or b);
    layer0_outputs(5787) <= not b or a;
    layer0_outputs(5788) <= b and not a;
    layer0_outputs(5789) <= a or b;
    layer0_outputs(5790) <= a;
    layer0_outputs(5791) <= not b or a;
    layer0_outputs(5792) <= not a;
    layer0_outputs(5793) <= a;
    layer0_outputs(5794) <= a or b;
    layer0_outputs(5795) <= not (a xor b);
    layer0_outputs(5796) <= a or b;
    layer0_outputs(5797) <= a;
    layer0_outputs(5798) <= not a or b;
    layer0_outputs(5799) <= not b;
    layer0_outputs(5800) <= not (a and b);
    layer0_outputs(5801) <= b;
    layer0_outputs(5802) <= not (a or b);
    layer0_outputs(5803) <= b;
    layer0_outputs(5804) <= not (a or b);
    layer0_outputs(5805) <= not b or a;
    layer0_outputs(5806) <= a and not b;
    layer0_outputs(5807) <= '1';
    layer0_outputs(5808) <= not b;
    layer0_outputs(5809) <= a or b;
    layer0_outputs(5810) <= a or b;
    layer0_outputs(5811) <= a;
    layer0_outputs(5812) <= not b;
    layer0_outputs(5813) <= not b or a;
    layer0_outputs(5814) <= a or b;
    layer0_outputs(5815) <= a and not b;
    layer0_outputs(5816) <= b;
    layer0_outputs(5817) <= not a or b;
    layer0_outputs(5818) <= not a;
    layer0_outputs(5819) <= not (a and b);
    layer0_outputs(5820) <= a and b;
    layer0_outputs(5821) <= not (a and b);
    layer0_outputs(5822) <= a;
    layer0_outputs(5823) <= not b or a;
    layer0_outputs(5824) <= not (a or b);
    layer0_outputs(5825) <= not (a or b);
    layer0_outputs(5826) <= b;
    layer0_outputs(5827) <= a xor b;
    layer0_outputs(5828) <= not (a xor b);
    layer0_outputs(5829) <= '1';
    layer0_outputs(5830) <= a or b;
    layer0_outputs(5831) <= not (a or b);
    layer0_outputs(5832) <= b;
    layer0_outputs(5833) <= b;
    layer0_outputs(5834) <= b;
    layer0_outputs(5835) <= a and b;
    layer0_outputs(5836) <= '1';
    layer0_outputs(5837) <= not (a or b);
    layer0_outputs(5838) <= not a;
    layer0_outputs(5839) <= a;
    layer0_outputs(5840) <= b;
    layer0_outputs(5841) <= not a or b;
    layer0_outputs(5842) <= not b;
    layer0_outputs(5843) <= not (a and b);
    layer0_outputs(5844) <= '1';
    layer0_outputs(5845) <= not b or a;
    layer0_outputs(5846) <= '0';
    layer0_outputs(5847) <= a;
    layer0_outputs(5848) <= b;
    layer0_outputs(5849) <= a and b;
    layer0_outputs(5850) <= not b or a;
    layer0_outputs(5851) <= not (a or b);
    layer0_outputs(5852) <= a;
    layer0_outputs(5853) <= not a or b;
    layer0_outputs(5854) <= a;
    layer0_outputs(5855) <= not b;
    layer0_outputs(5856) <= not a;
    layer0_outputs(5857) <= a and not b;
    layer0_outputs(5858) <= not a;
    layer0_outputs(5859) <= '0';
    layer0_outputs(5860) <= not a;
    layer0_outputs(5861) <= not (a xor b);
    layer0_outputs(5862) <= b and not a;
    layer0_outputs(5863) <= b and not a;
    layer0_outputs(5864) <= not (a xor b);
    layer0_outputs(5865) <= not (a xor b);
    layer0_outputs(5866) <= a or b;
    layer0_outputs(5867) <= not (a or b);
    layer0_outputs(5868) <= a and not b;
    layer0_outputs(5869) <= not b;
    layer0_outputs(5870) <= b;
    layer0_outputs(5871) <= a or b;
    layer0_outputs(5872) <= a and not b;
    layer0_outputs(5873) <= a;
    layer0_outputs(5874) <= a xor b;
    layer0_outputs(5875) <= not b or a;
    layer0_outputs(5876) <= b;
    layer0_outputs(5877) <= a and not b;
    layer0_outputs(5878) <= a and not b;
    layer0_outputs(5879) <= not a or b;
    layer0_outputs(5880) <= not b;
    layer0_outputs(5881) <= a;
    layer0_outputs(5882) <= a or b;
    layer0_outputs(5883) <= not b;
    layer0_outputs(5884) <= a and b;
    layer0_outputs(5885) <= '0';
    layer0_outputs(5886) <= b and not a;
    layer0_outputs(5887) <= a;
    layer0_outputs(5888) <= not a;
    layer0_outputs(5889) <= b;
    layer0_outputs(5890) <= b and not a;
    layer0_outputs(5891) <= not (a or b);
    layer0_outputs(5892) <= not (a or b);
    layer0_outputs(5893) <= b;
    layer0_outputs(5894) <= not (a and b);
    layer0_outputs(5895) <= '0';
    layer0_outputs(5896) <= a;
    layer0_outputs(5897) <= not b;
    layer0_outputs(5898) <= not (a and b);
    layer0_outputs(5899) <= a;
    layer0_outputs(5900) <= not b or a;
    layer0_outputs(5901) <= '1';
    layer0_outputs(5902) <= a and not b;
    layer0_outputs(5903) <= b;
    layer0_outputs(5904) <= not b;
    layer0_outputs(5905) <= a and b;
    layer0_outputs(5906) <= '0';
    layer0_outputs(5907) <= a or b;
    layer0_outputs(5908) <= b;
    layer0_outputs(5909) <= not (a and b);
    layer0_outputs(5910) <= a or b;
    layer0_outputs(5911) <= a xor b;
    layer0_outputs(5912) <= a;
    layer0_outputs(5913) <= b;
    layer0_outputs(5914) <= a and b;
    layer0_outputs(5915) <= a xor b;
    layer0_outputs(5916) <= not (a and b);
    layer0_outputs(5917) <= a xor b;
    layer0_outputs(5918) <= not b;
    layer0_outputs(5919) <= a and not b;
    layer0_outputs(5920) <= not (a xor b);
    layer0_outputs(5921) <= a or b;
    layer0_outputs(5922) <= not (a or b);
    layer0_outputs(5923) <= not b or a;
    layer0_outputs(5924) <= not a;
    layer0_outputs(5925) <= not a;
    layer0_outputs(5926) <= a xor b;
    layer0_outputs(5927) <= not (a xor b);
    layer0_outputs(5928) <= not b;
    layer0_outputs(5929) <= not a or b;
    layer0_outputs(5930) <= b and not a;
    layer0_outputs(5931) <= not b or a;
    layer0_outputs(5932) <= a xor b;
    layer0_outputs(5933) <= '0';
    layer0_outputs(5934) <= not (a xor b);
    layer0_outputs(5935) <= not b;
    layer0_outputs(5936) <= a;
    layer0_outputs(5937) <= a;
    layer0_outputs(5938) <= not b;
    layer0_outputs(5939) <= not (a and b);
    layer0_outputs(5940) <= not (a and b);
    layer0_outputs(5941) <= not a;
    layer0_outputs(5942) <= '1';
    layer0_outputs(5943) <= b and not a;
    layer0_outputs(5944) <= a and not b;
    layer0_outputs(5945) <= a and not b;
    layer0_outputs(5946) <= a and not b;
    layer0_outputs(5947) <= a and b;
    layer0_outputs(5948) <= a or b;
    layer0_outputs(5949) <= not a;
    layer0_outputs(5950) <= a;
    layer0_outputs(5951) <= a and b;
    layer0_outputs(5952) <= not b;
    layer0_outputs(5953) <= a xor b;
    layer0_outputs(5954) <= not b;
    layer0_outputs(5955) <= not (a and b);
    layer0_outputs(5956) <= b and not a;
    layer0_outputs(5957) <= not b;
    layer0_outputs(5958) <= not b or a;
    layer0_outputs(5959) <= b and not a;
    layer0_outputs(5960) <= b and not a;
    layer0_outputs(5961) <= a and b;
    layer0_outputs(5962) <= not b or a;
    layer0_outputs(5963) <= a and b;
    layer0_outputs(5964) <= '1';
    layer0_outputs(5965) <= a xor b;
    layer0_outputs(5966) <= a and not b;
    layer0_outputs(5967) <= not (a or b);
    layer0_outputs(5968) <= a;
    layer0_outputs(5969) <= b;
    layer0_outputs(5970) <= a xor b;
    layer0_outputs(5971) <= not (a and b);
    layer0_outputs(5972) <= a xor b;
    layer0_outputs(5973) <= not a;
    layer0_outputs(5974) <= '1';
    layer0_outputs(5975) <= a xor b;
    layer0_outputs(5976) <= not a;
    layer0_outputs(5977) <= a;
    layer0_outputs(5978) <= not a or b;
    layer0_outputs(5979) <= b and not a;
    layer0_outputs(5980) <= not a or b;
    layer0_outputs(5981) <= b and not a;
    layer0_outputs(5982) <= not a;
    layer0_outputs(5983) <= a or b;
    layer0_outputs(5984) <= a and not b;
    layer0_outputs(5985) <= b and not a;
    layer0_outputs(5986) <= not (a or b);
    layer0_outputs(5987) <= not b or a;
    layer0_outputs(5988) <= '1';
    layer0_outputs(5989) <= a or b;
    layer0_outputs(5990) <= not b;
    layer0_outputs(5991) <= a;
    layer0_outputs(5992) <= not (a xor b);
    layer0_outputs(5993) <= '0';
    layer0_outputs(5994) <= a or b;
    layer0_outputs(5995) <= b;
    layer0_outputs(5996) <= a and b;
    layer0_outputs(5997) <= not a or b;
    layer0_outputs(5998) <= not b or a;
    layer0_outputs(5999) <= not (a xor b);
    layer0_outputs(6000) <= '1';
    layer0_outputs(6001) <= not (a xor b);
    layer0_outputs(6002) <= a or b;
    layer0_outputs(6003) <= not a or b;
    layer0_outputs(6004) <= b and not a;
    layer0_outputs(6005) <= b and not a;
    layer0_outputs(6006) <= a;
    layer0_outputs(6007) <= a or b;
    layer0_outputs(6008) <= not (a and b);
    layer0_outputs(6009) <= not a or b;
    layer0_outputs(6010) <= not b;
    layer0_outputs(6011) <= a and b;
    layer0_outputs(6012) <= a;
    layer0_outputs(6013) <= a xor b;
    layer0_outputs(6014) <= not b or a;
    layer0_outputs(6015) <= b and not a;
    layer0_outputs(6016) <= a and b;
    layer0_outputs(6017) <= a;
    layer0_outputs(6018) <= not (a or b);
    layer0_outputs(6019) <= a or b;
    layer0_outputs(6020) <= '0';
    layer0_outputs(6021) <= not b;
    layer0_outputs(6022) <= not b;
    layer0_outputs(6023) <= b;
    layer0_outputs(6024) <= not b or a;
    layer0_outputs(6025) <= a or b;
    layer0_outputs(6026) <= a or b;
    layer0_outputs(6027) <= a and b;
    layer0_outputs(6028) <= a and b;
    layer0_outputs(6029) <= '0';
    layer0_outputs(6030) <= not b;
    layer0_outputs(6031) <= a xor b;
    layer0_outputs(6032) <= not (a and b);
    layer0_outputs(6033) <= a or b;
    layer0_outputs(6034) <= a xor b;
    layer0_outputs(6035) <= not (a xor b);
    layer0_outputs(6036) <= not a or b;
    layer0_outputs(6037) <= a and b;
    layer0_outputs(6038) <= not (a xor b);
    layer0_outputs(6039) <= not b or a;
    layer0_outputs(6040) <= not a;
    layer0_outputs(6041) <= a or b;
    layer0_outputs(6042) <= a and b;
    layer0_outputs(6043) <= b and not a;
    layer0_outputs(6044) <= not b;
    layer0_outputs(6045) <= a and not b;
    layer0_outputs(6046) <= a and b;
    layer0_outputs(6047) <= not a or b;
    layer0_outputs(6048) <= not a;
    layer0_outputs(6049) <= a and not b;
    layer0_outputs(6050) <= not (a or b);
    layer0_outputs(6051) <= not a;
    layer0_outputs(6052) <= a;
    layer0_outputs(6053) <= a or b;
    layer0_outputs(6054) <= not a;
    layer0_outputs(6055) <= not a or b;
    layer0_outputs(6056) <= b;
    layer0_outputs(6057) <= a xor b;
    layer0_outputs(6058) <= a and not b;
    layer0_outputs(6059) <= not (a xor b);
    layer0_outputs(6060) <= a and not b;
    layer0_outputs(6061) <= '0';
    layer0_outputs(6062) <= not (a xor b);
    layer0_outputs(6063) <= a or b;
    layer0_outputs(6064) <= not (a or b);
    layer0_outputs(6065) <= a or b;
    layer0_outputs(6066) <= b;
    layer0_outputs(6067) <= a xor b;
    layer0_outputs(6068) <= a or b;
    layer0_outputs(6069) <= '0';
    layer0_outputs(6070) <= b;
    layer0_outputs(6071) <= not b or a;
    layer0_outputs(6072) <= a and b;
    layer0_outputs(6073) <= a and not b;
    layer0_outputs(6074) <= a xor b;
    layer0_outputs(6075) <= not (a and b);
    layer0_outputs(6076) <= not b or a;
    layer0_outputs(6077) <= a and b;
    layer0_outputs(6078) <= a or b;
    layer0_outputs(6079) <= not b;
    layer0_outputs(6080) <= '0';
    layer0_outputs(6081) <= not a or b;
    layer0_outputs(6082) <= a;
    layer0_outputs(6083) <= not (a xor b);
    layer0_outputs(6084) <= not (a or b);
    layer0_outputs(6085) <= not (a and b);
    layer0_outputs(6086) <= a;
    layer0_outputs(6087) <= not a or b;
    layer0_outputs(6088) <= not a;
    layer0_outputs(6089) <= not (a xor b);
    layer0_outputs(6090) <= not a or b;
    layer0_outputs(6091) <= a;
    layer0_outputs(6092) <= b;
    layer0_outputs(6093) <= '0';
    layer0_outputs(6094) <= not (a and b);
    layer0_outputs(6095) <= not (a or b);
    layer0_outputs(6096) <= a;
    layer0_outputs(6097) <= b and not a;
    layer0_outputs(6098) <= a xor b;
    layer0_outputs(6099) <= a xor b;
    layer0_outputs(6100) <= '1';
    layer0_outputs(6101) <= not (a xor b);
    layer0_outputs(6102) <= '1';
    layer0_outputs(6103) <= a or b;
    layer0_outputs(6104) <= not b or a;
    layer0_outputs(6105) <= not (a xor b);
    layer0_outputs(6106) <= a xor b;
    layer0_outputs(6107) <= '1';
    layer0_outputs(6108) <= not a or b;
    layer0_outputs(6109) <= a xor b;
    layer0_outputs(6110) <= a or b;
    layer0_outputs(6111) <= not a;
    layer0_outputs(6112) <= not (a or b);
    layer0_outputs(6113) <= not a;
    layer0_outputs(6114) <= not (a or b);
    layer0_outputs(6115) <= a xor b;
    layer0_outputs(6116) <= not (a and b);
    layer0_outputs(6117) <= a and not b;
    layer0_outputs(6118) <= a xor b;
    layer0_outputs(6119) <= b;
    layer0_outputs(6120) <= not (a xor b);
    layer0_outputs(6121) <= not (a or b);
    layer0_outputs(6122) <= not (a or b);
    layer0_outputs(6123) <= not (a or b);
    layer0_outputs(6124) <= a xor b;
    layer0_outputs(6125) <= a xor b;
    layer0_outputs(6126) <= not a;
    layer0_outputs(6127) <= not a or b;
    layer0_outputs(6128) <= not b;
    layer0_outputs(6129) <= a;
    layer0_outputs(6130) <= not a or b;
    layer0_outputs(6131) <= not a;
    layer0_outputs(6132) <= not (a or b);
    layer0_outputs(6133) <= a or b;
    layer0_outputs(6134) <= not (a or b);
    layer0_outputs(6135) <= a or b;
    layer0_outputs(6136) <= a and b;
    layer0_outputs(6137) <= not b;
    layer0_outputs(6138) <= not (a or b);
    layer0_outputs(6139) <= a;
    layer0_outputs(6140) <= a or b;
    layer0_outputs(6141) <= not b;
    layer0_outputs(6142) <= not b;
    layer0_outputs(6143) <= a xor b;
    layer0_outputs(6144) <= a;
    layer0_outputs(6145) <= a;
    layer0_outputs(6146) <= not a;
    layer0_outputs(6147) <= b;
    layer0_outputs(6148) <= not a or b;
    layer0_outputs(6149) <= not a or b;
    layer0_outputs(6150) <= '0';
    layer0_outputs(6151) <= a xor b;
    layer0_outputs(6152) <= not a;
    layer0_outputs(6153) <= not a or b;
    layer0_outputs(6154) <= a or b;
    layer0_outputs(6155) <= '0';
    layer0_outputs(6156) <= a and not b;
    layer0_outputs(6157) <= a xor b;
    layer0_outputs(6158) <= b;
    layer0_outputs(6159) <= a;
    layer0_outputs(6160) <= a and b;
    layer0_outputs(6161) <= b;
    layer0_outputs(6162) <= '1';
    layer0_outputs(6163) <= a xor b;
    layer0_outputs(6164) <= a xor b;
    layer0_outputs(6165) <= not (a or b);
    layer0_outputs(6166) <= a;
    layer0_outputs(6167) <= a;
    layer0_outputs(6168) <= not (a or b);
    layer0_outputs(6169) <= not (a or b);
    layer0_outputs(6170) <= a xor b;
    layer0_outputs(6171) <= not b or a;
    layer0_outputs(6172) <= not (a and b);
    layer0_outputs(6173) <= a;
    layer0_outputs(6174) <= not (a and b);
    layer0_outputs(6175) <= a or b;
    layer0_outputs(6176) <= a and not b;
    layer0_outputs(6177) <= not b;
    layer0_outputs(6178) <= '1';
    layer0_outputs(6179) <= '0';
    layer0_outputs(6180) <= not b or a;
    layer0_outputs(6181) <= a;
    layer0_outputs(6182) <= not (a and b);
    layer0_outputs(6183) <= not a;
    layer0_outputs(6184) <= not (a xor b);
    layer0_outputs(6185) <= b;
    layer0_outputs(6186) <= '1';
    layer0_outputs(6187) <= a and not b;
    layer0_outputs(6188) <= not (a and b);
    layer0_outputs(6189) <= a and not b;
    layer0_outputs(6190) <= a or b;
    layer0_outputs(6191) <= a;
    layer0_outputs(6192) <= a or b;
    layer0_outputs(6193) <= a xor b;
    layer0_outputs(6194) <= a;
    layer0_outputs(6195) <= b and not a;
    layer0_outputs(6196) <= a xor b;
    layer0_outputs(6197) <= b and not a;
    layer0_outputs(6198) <= a and b;
    layer0_outputs(6199) <= not b;
    layer0_outputs(6200) <= b;
    layer0_outputs(6201) <= not a;
    layer0_outputs(6202) <= not (a xor b);
    layer0_outputs(6203) <= not (a xor b);
    layer0_outputs(6204) <= '1';
    layer0_outputs(6205) <= not a or b;
    layer0_outputs(6206) <= a xor b;
    layer0_outputs(6207) <= '1';
    layer0_outputs(6208) <= not (a xor b);
    layer0_outputs(6209) <= a and not b;
    layer0_outputs(6210) <= not a or b;
    layer0_outputs(6211) <= a and b;
    layer0_outputs(6212) <= a and b;
    layer0_outputs(6213) <= a;
    layer0_outputs(6214) <= not b or a;
    layer0_outputs(6215) <= a and b;
    layer0_outputs(6216) <= '0';
    layer0_outputs(6217) <= a xor b;
    layer0_outputs(6218) <= not (a or b);
    layer0_outputs(6219) <= not b or a;
    layer0_outputs(6220) <= not a or b;
    layer0_outputs(6221) <= not (a and b);
    layer0_outputs(6222) <= a or b;
    layer0_outputs(6223) <= a;
    layer0_outputs(6224) <= not b or a;
    layer0_outputs(6225) <= a and not b;
    layer0_outputs(6226) <= a xor b;
    layer0_outputs(6227) <= a and b;
    layer0_outputs(6228) <= not a or b;
    layer0_outputs(6229) <= b;
    layer0_outputs(6230) <= not b or a;
    layer0_outputs(6231) <= '1';
    layer0_outputs(6232) <= a and not b;
    layer0_outputs(6233) <= not b or a;
    layer0_outputs(6234) <= b and not a;
    layer0_outputs(6235) <= not (a or b);
    layer0_outputs(6236) <= a;
    layer0_outputs(6237) <= '1';
    layer0_outputs(6238) <= a;
    layer0_outputs(6239) <= '0';
    layer0_outputs(6240) <= not (a xor b);
    layer0_outputs(6241) <= a and b;
    layer0_outputs(6242) <= a and b;
    layer0_outputs(6243) <= not b;
    layer0_outputs(6244) <= a or b;
    layer0_outputs(6245) <= b;
    layer0_outputs(6246) <= '1';
    layer0_outputs(6247) <= not (a xor b);
    layer0_outputs(6248) <= not (a or b);
    layer0_outputs(6249) <= b and not a;
    layer0_outputs(6250) <= a xor b;
    layer0_outputs(6251) <= b;
    layer0_outputs(6252) <= not a or b;
    layer0_outputs(6253) <= a;
    layer0_outputs(6254) <= a or b;
    layer0_outputs(6255) <= a and not b;
    layer0_outputs(6256) <= not a;
    layer0_outputs(6257) <= not a or b;
    layer0_outputs(6258) <= not (a and b);
    layer0_outputs(6259) <= a or b;
    layer0_outputs(6260) <= a and b;
    layer0_outputs(6261) <= a and b;
    layer0_outputs(6262) <= b;
    layer0_outputs(6263) <= b;
    layer0_outputs(6264) <= a or b;
    layer0_outputs(6265) <= not a;
    layer0_outputs(6266) <= not (a and b);
    layer0_outputs(6267) <= not a or b;
    layer0_outputs(6268) <= a and b;
    layer0_outputs(6269) <= b;
    layer0_outputs(6270) <= a;
    layer0_outputs(6271) <= b;
    layer0_outputs(6272) <= not (a or b);
    layer0_outputs(6273) <= a;
    layer0_outputs(6274) <= a and b;
    layer0_outputs(6275) <= a and b;
    layer0_outputs(6276) <= b and not a;
    layer0_outputs(6277) <= b and not a;
    layer0_outputs(6278) <= not (a xor b);
    layer0_outputs(6279) <= b and not a;
    layer0_outputs(6280) <= not (a or b);
    layer0_outputs(6281) <= not a;
    layer0_outputs(6282) <= not b;
    layer0_outputs(6283) <= not (a xor b);
    layer0_outputs(6284) <= not (a or b);
    layer0_outputs(6285) <= '1';
    layer0_outputs(6286) <= not a or b;
    layer0_outputs(6287) <= a;
    layer0_outputs(6288) <= a or b;
    layer0_outputs(6289) <= a;
    layer0_outputs(6290) <= b;
    layer0_outputs(6291) <= not b or a;
    layer0_outputs(6292) <= a and not b;
    layer0_outputs(6293) <= not (a or b);
    layer0_outputs(6294) <= a xor b;
    layer0_outputs(6295) <= b and not a;
    layer0_outputs(6296) <= a;
    layer0_outputs(6297) <= a or b;
    layer0_outputs(6298) <= not a or b;
    layer0_outputs(6299) <= a and not b;
    layer0_outputs(6300) <= a or b;
    layer0_outputs(6301) <= '0';
    layer0_outputs(6302) <= b and not a;
    layer0_outputs(6303) <= not (a xor b);
    layer0_outputs(6304) <= not (a or b);
    layer0_outputs(6305) <= not (a or b);
    layer0_outputs(6306) <= not (a and b);
    layer0_outputs(6307) <= not a;
    layer0_outputs(6308) <= not a;
    layer0_outputs(6309) <= not (a xor b);
    layer0_outputs(6310) <= a xor b;
    layer0_outputs(6311) <= not a or b;
    layer0_outputs(6312) <= a and b;
    layer0_outputs(6313) <= not (a or b);
    layer0_outputs(6314) <= not a or b;
    layer0_outputs(6315) <= not a or b;
    layer0_outputs(6316) <= not b;
    layer0_outputs(6317) <= not (a or b);
    layer0_outputs(6318) <= not (a or b);
    layer0_outputs(6319) <= a;
    layer0_outputs(6320) <= not b or a;
    layer0_outputs(6321) <= a xor b;
    layer0_outputs(6322) <= '1';
    layer0_outputs(6323) <= not (a xor b);
    layer0_outputs(6324) <= not a;
    layer0_outputs(6325) <= not (a and b);
    layer0_outputs(6326) <= a or b;
    layer0_outputs(6327) <= not b or a;
    layer0_outputs(6328) <= not (a and b);
    layer0_outputs(6329) <= not (a or b);
    layer0_outputs(6330) <= a;
    layer0_outputs(6331) <= a and not b;
    layer0_outputs(6332) <= not (a xor b);
    layer0_outputs(6333) <= a xor b;
    layer0_outputs(6334) <= not (a xor b);
    layer0_outputs(6335) <= a xor b;
    layer0_outputs(6336) <= not (a or b);
    layer0_outputs(6337) <= not a or b;
    layer0_outputs(6338) <= not b;
    layer0_outputs(6339) <= not b;
    layer0_outputs(6340) <= a xor b;
    layer0_outputs(6341) <= '1';
    layer0_outputs(6342) <= a;
    layer0_outputs(6343) <= a;
    layer0_outputs(6344) <= not a;
    layer0_outputs(6345) <= a xor b;
    layer0_outputs(6346) <= not b;
    layer0_outputs(6347) <= a;
    layer0_outputs(6348) <= b;
    layer0_outputs(6349) <= not a or b;
    layer0_outputs(6350) <= b;
    layer0_outputs(6351) <= a and not b;
    layer0_outputs(6352) <= b and not a;
    layer0_outputs(6353) <= not a;
    layer0_outputs(6354) <= b;
    layer0_outputs(6355) <= a and b;
    layer0_outputs(6356) <= not b;
    layer0_outputs(6357) <= a;
    layer0_outputs(6358) <= b and not a;
    layer0_outputs(6359) <= not a;
    layer0_outputs(6360) <= a and b;
    layer0_outputs(6361) <= not b or a;
    layer0_outputs(6362) <= a;
    layer0_outputs(6363) <= not a;
    layer0_outputs(6364) <= not (a xor b);
    layer0_outputs(6365) <= not (a or b);
    layer0_outputs(6366) <= a;
    layer0_outputs(6367) <= not b or a;
    layer0_outputs(6368) <= '1';
    layer0_outputs(6369) <= a;
    layer0_outputs(6370) <= not a;
    layer0_outputs(6371) <= not a;
    layer0_outputs(6372) <= b and not a;
    layer0_outputs(6373) <= a or b;
    layer0_outputs(6374) <= a xor b;
    layer0_outputs(6375) <= a xor b;
    layer0_outputs(6376) <= a and b;
    layer0_outputs(6377) <= not (a and b);
    layer0_outputs(6378) <= a xor b;
    layer0_outputs(6379) <= not (a or b);
    layer0_outputs(6380) <= not (a or b);
    layer0_outputs(6381) <= not a;
    layer0_outputs(6382) <= b and not a;
    layer0_outputs(6383) <= not (a or b);
    layer0_outputs(6384) <= not b;
    layer0_outputs(6385) <= not b or a;
    layer0_outputs(6386) <= not a;
    layer0_outputs(6387) <= a or b;
    layer0_outputs(6388) <= not (a and b);
    layer0_outputs(6389) <= not (a and b);
    layer0_outputs(6390) <= a;
    layer0_outputs(6391) <= not b;
    layer0_outputs(6392) <= '0';
    layer0_outputs(6393) <= not a;
    layer0_outputs(6394) <= not b;
    layer0_outputs(6395) <= b and not a;
    layer0_outputs(6396) <= '1';
    layer0_outputs(6397) <= not a or b;
    layer0_outputs(6398) <= not (a and b);
    layer0_outputs(6399) <= a xor b;
    layer0_outputs(6400) <= b and not a;
    layer0_outputs(6401) <= not (a or b);
    layer0_outputs(6402) <= not a;
    layer0_outputs(6403) <= a and not b;
    layer0_outputs(6404) <= a or b;
    layer0_outputs(6405) <= not a;
    layer0_outputs(6406) <= a or b;
    layer0_outputs(6407) <= '1';
    layer0_outputs(6408) <= not (a xor b);
    layer0_outputs(6409) <= b and not a;
    layer0_outputs(6410) <= a and b;
    layer0_outputs(6411) <= not b;
    layer0_outputs(6412) <= a or b;
    layer0_outputs(6413) <= b;
    layer0_outputs(6414) <= not (a and b);
    layer0_outputs(6415) <= b and not a;
    layer0_outputs(6416) <= not a;
    layer0_outputs(6417) <= '1';
    layer0_outputs(6418) <= b and not a;
    layer0_outputs(6419) <= a and b;
    layer0_outputs(6420) <= a;
    layer0_outputs(6421) <= not (a or b);
    layer0_outputs(6422) <= a and b;
    layer0_outputs(6423) <= not a or b;
    layer0_outputs(6424) <= not (a or b);
    layer0_outputs(6425) <= not b;
    layer0_outputs(6426) <= a;
    layer0_outputs(6427) <= not a;
    layer0_outputs(6428) <= '0';
    layer0_outputs(6429) <= a or b;
    layer0_outputs(6430) <= b and not a;
    layer0_outputs(6431) <= not (a and b);
    layer0_outputs(6432) <= not (a or b);
    layer0_outputs(6433) <= not a or b;
    layer0_outputs(6434) <= not b;
    layer0_outputs(6435) <= not (a or b);
    layer0_outputs(6436) <= a;
    layer0_outputs(6437) <= b and not a;
    layer0_outputs(6438) <= not a or b;
    layer0_outputs(6439) <= not a;
    layer0_outputs(6440) <= not b;
    layer0_outputs(6441) <= b and not a;
    layer0_outputs(6442) <= b and not a;
    layer0_outputs(6443) <= b;
    layer0_outputs(6444) <= '0';
    layer0_outputs(6445) <= not b;
    layer0_outputs(6446) <= not a;
    layer0_outputs(6447) <= a xor b;
    layer0_outputs(6448) <= not a or b;
    layer0_outputs(6449) <= not (a or b);
    layer0_outputs(6450) <= not b;
    layer0_outputs(6451) <= not (a xor b);
    layer0_outputs(6452) <= a;
    layer0_outputs(6453) <= '0';
    layer0_outputs(6454) <= not (a or b);
    layer0_outputs(6455) <= not b;
    layer0_outputs(6456) <= '0';
    layer0_outputs(6457) <= a and b;
    layer0_outputs(6458) <= not b or a;
    layer0_outputs(6459) <= a or b;
    layer0_outputs(6460) <= a and not b;
    layer0_outputs(6461) <= b;
    layer0_outputs(6462) <= '1';
    layer0_outputs(6463) <= a xor b;
    layer0_outputs(6464) <= not b;
    layer0_outputs(6465) <= a or b;
    layer0_outputs(6466) <= not a;
    layer0_outputs(6467) <= not (a xor b);
    layer0_outputs(6468) <= not (a or b);
    layer0_outputs(6469) <= not b or a;
    layer0_outputs(6470) <= b;
    layer0_outputs(6471) <= b;
    layer0_outputs(6472) <= a and not b;
    layer0_outputs(6473) <= a or b;
    layer0_outputs(6474) <= not b;
    layer0_outputs(6475) <= a or b;
    layer0_outputs(6476) <= not (a or b);
    layer0_outputs(6477) <= a and not b;
    layer0_outputs(6478) <= a and not b;
    layer0_outputs(6479) <= a;
    layer0_outputs(6480) <= b and not a;
    layer0_outputs(6481) <= not (a xor b);
    layer0_outputs(6482) <= not (a xor b);
    layer0_outputs(6483) <= b;
    layer0_outputs(6484) <= a and b;
    layer0_outputs(6485) <= '1';
    layer0_outputs(6486) <= not a or b;
    layer0_outputs(6487) <= b and not a;
    layer0_outputs(6488) <= not b;
    layer0_outputs(6489) <= not a;
    layer0_outputs(6490) <= '0';
    layer0_outputs(6491) <= not b or a;
    layer0_outputs(6492) <= not a;
    layer0_outputs(6493) <= not (a xor b);
    layer0_outputs(6494) <= b;
    layer0_outputs(6495) <= '1';
    layer0_outputs(6496) <= a;
    layer0_outputs(6497) <= not b;
    layer0_outputs(6498) <= a and not b;
    layer0_outputs(6499) <= b;
    layer0_outputs(6500) <= not b;
    layer0_outputs(6501) <= a or b;
    layer0_outputs(6502) <= b and not a;
    layer0_outputs(6503) <= a and not b;
    layer0_outputs(6504) <= not a;
    layer0_outputs(6505) <= not a or b;
    layer0_outputs(6506) <= not (a xor b);
    layer0_outputs(6507) <= a or b;
    layer0_outputs(6508) <= a or b;
    layer0_outputs(6509) <= not a or b;
    layer0_outputs(6510) <= not a;
    layer0_outputs(6511) <= not a;
    layer0_outputs(6512) <= a and b;
    layer0_outputs(6513) <= not a;
    layer0_outputs(6514) <= not b;
    layer0_outputs(6515) <= b and not a;
    layer0_outputs(6516) <= b and not a;
    layer0_outputs(6517) <= a and b;
    layer0_outputs(6518) <= a xor b;
    layer0_outputs(6519) <= not b;
    layer0_outputs(6520) <= b and not a;
    layer0_outputs(6521) <= not (a or b);
    layer0_outputs(6522) <= a and not b;
    layer0_outputs(6523) <= not a;
    layer0_outputs(6524) <= not (a xor b);
    layer0_outputs(6525) <= b and not a;
    layer0_outputs(6526) <= not a or b;
    layer0_outputs(6527) <= a and not b;
    layer0_outputs(6528) <= not b;
    layer0_outputs(6529) <= not a;
    layer0_outputs(6530) <= a xor b;
    layer0_outputs(6531) <= a;
    layer0_outputs(6532) <= a or b;
    layer0_outputs(6533) <= not a;
    layer0_outputs(6534) <= not a or b;
    layer0_outputs(6535) <= not (a and b);
    layer0_outputs(6536) <= '0';
    layer0_outputs(6537) <= a xor b;
    layer0_outputs(6538) <= '0';
    layer0_outputs(6539) <= b;
    layer0_outputs(6540) <= '0';
    layer0_outputs(6541) <= '0';
    layer0_outputs(6542) <= a and b;
    layer0_outputs(6543) <= '0';
    layer0_outputs(6544) <= b;
    layer0_outputs(6545) <= not a or b;
    layer0_outputs(6546) <= b;
    layer0_outputs(6547) <= '0';
    layer0_outputs(6548) <= a xor b;
    layer0_outputs(6549) <= a or b;
    layer0_outputs(6550) <= b;
    layer0_outputs(6551) <= not (a xor b);
    layer0_outputs(6552) <= not (a xor b);
    layer0_outputs(6553) <= not (a or b);
    layer0_outputs(6554) <= not b or a;
    layer0_outputs(6555) <= not b;
    layer0_outputs(6556) <= not (a xor b);
    layer0_outputs(6557) <= a and not b;
    layer0_outputs(6558) <= not (a or b);
    layer0_outputs(6559) <= not (a xor b);
    layer0_outputs(6560) <= not (a or b);
    layer0_outputs(6561) <= not (a and b);
    layer0_outputs(6562) <= not (a xor b);
    layer0_outputs(6563) <= '0';
    layer0_outputs(6564) <= not b or a;
    layer0_outputs(6565) <= b;
    layer0_outputs(6566) <= not (a and b);
    layer0_outputs(6567) <= b;
    layer0_outputs(6568) <= b;
    layer0_outputs(6569) <= '1';
    layer0_outputs(6570) <= b;
    layer0_outputs(6571) <= a;
    layer0_outputs(6572) <= a;
    layer0_outputs(6573) <= not a or b;
    layer0_outputs(6574) <= not (a xor b);
    layer0_outputs(6575) <= a xor b;
    layer0_outputs(6576) <= not (a xor b);
    layer0_outputs(6577) <= not (a or b);
    layer0_outputs(6578) <= a and not b;
    layer0_outputs(6579) <= not b;
    layer0_outputs(6580) <= a and b;
    layer0_outputs(6581) <= not a;
    layer0_outputs(6582) <= a;
    layer0_outputs(6583) <= '1';
    layer0_outputs(6584) <= b;
    layer0_outputs(6585) <= a;
    layer0_outputs(6586) <= not b or a;
    layer0_outputs(6587) <= not b or a;
    layer0_outputs(6588) <= a;
    layer0_outputs(6589) <= not (a or b);
    layer0_outputs(6590) <= a or b;
    layer0_outputs(6591) <= not a;
    layer0_outputs(6592) <= b;
    layer0_outputs(6593) <= '0';
    layer0_outputs(6594) <= not b;
    layer0_outputs(6595) <= a and not b;
    layer0_outputs(6596) <= '0';
    layer0_outputs(6597) <= a xor b;
    layer0_outputs(6598) <= not (a xor b);
    layer0_outputs(6599) <= not b;
    layer0_outputs(6600) <= not (a xor b);
    layer0_outputs(6601) <= a;
    layer0_outputs(6602) <= a xor b;
    layer0_outputs(6603) <= b and not a;
    layer0_outputs(6604) <= not b;
    layer0_outputs(6605) <= not a;
    layer0_outputs(6606) <= not (a and b);
    layer0_outputs(6607) <= b and not a;
    layer0_outputs(6608) <= a or b;
    layer0_outputs(6609) <= not (a xor b);
    layer0_outputs(6610) <= not (a or b);
    layer0_outputs(6611) <= a xor b;
    layer0_outputs(6612) <= not (a or b);
    layer0_outputs(6613) <= not a;
    layer0_outputs(6614) <= not a or b;
    layer0_outputs(6615) <= b and not a;
    layer0_outputs(6616) <= a and not b;
    layer0_outputs(6617) <= a and b;
    layer0_outputs(6618) <= a and not b;
    layer0_outputs(6619) <= not (a and b);
    layer0_outputs(6620) <= '0';
    layer0_outputs(6621) <= not b;
    layer0_outputs(6622) <= not (a or b);
    layer0_outputs(6623) <= not a;
    layer0_outputs(6624) <= not b or a;
    layer0_outputs(6625) <= '1';
    layer0_outputs(6626) <= not b or a;
    layer0_outputs(6627) <= not (a xor b);
    layer0_outputs(6628) <= a xor b;
    layer0_outputs(6629) <= a and b;
    layer0_outputs(6630) <= not (a or b);
    layer0_outputs(6631) <= b and not a;
    layer0_outputs(6632) <= '1';
    layer0_outputs(6633) <= not (a xor b);
    layer0_outputs(6634) <= not a or b;
    layer0_outputs(6635) <= b and not a;
    layer0_outputs(6636) <= '1';
    layer0_outputs(6637) <= not a;
    layer0_outputs(6638) <= b;
    layer0_outputs(6639) <= a and not b;
    layer0_outputs(6640) <= not a;
    layer0_outputs(6641) <= not a or b;
    layer0_outputs(6642) <= a and not b;
    layer0_outputs(6643) <= not a or b;
    layer0_outputs(6644) <= not (a xor b);
    layer0_outputs(6645) <= not (a or b);
    layer0_outputs(6646) <= not b or a;
    layer0_outputs(6647) <= a and not b;
    layer0_outputs(6648) <= '0';
    layer0_outputs(6649) <= a;
    layer0_outputs(6650) <= '1';
    layer0_outputs(6651) <= b and not a;
    layer0_outputs(6652) <= not a or b;
    layer0_outputs(6653) <= not (a and b);
    layer0_outputs(6654) <= a xor b;
    layer0_outputs(6655) <= not (a or b);
    layer0_outputs(6656) <= '0';
    layer0_outputs(6657) <= not a;
    layer0_outputs(6658) <= not (a xor b);
    layer0_outputs(6659) <= a or b;
    layer0_outputs(6660) <= a and b;
    layer0_outputs(6661) <= not b;
    layer0_outputs(6662) <= not b;
    layer0_outputs(6663) <= '0';
    layer0_outputs(6664) <= '1';
    layer0_outputs(6665) <= not (a or b);
    layer0_outputs(6666) <= b and not a;
    layer0_outputs(6667) <= a and not b;
    layer0_outputs(6668) <= '1';
    layer0_outputs(6669) <= a xor b;
    layer0_outputs(6670) <= not b or a;
    layer0_outputs(6671) <= '1';
    layer0_outputs(6672) <= a and b;
    layer0_outputs(6673) <= '1';
    layer0_outputs(6674) <= a;
    layer0_outputs(6675) <= a xor b;
    layer0_outputs(6676) <= not (a and b);
    layer0_outputs(6677) <= not (a and b);
    layer0_outputs(6678) <= not (a xor b);
    layer0_outputs(6679) <= a xor b;
    layer0_outputs(6680) <= not (a and b);
    layer0_outputs(6681) <= not (a or b);
    layer0_outputs(6682) <= '0';
    layer0_outputs(6683) <= not (a or b);
    layer0_outputs(6684) <= b and not a;
    layer0_outputs(6685) <= a or b;
    layer0_outputs(6686) <= '0';
    layer0_outputs(6687) <= a or b;
    layer0_outputs(6688) <= not (a xor b);
    layer0_outputs(6689) <= not (a or b);
    layer0_outputs(6690) <= a and not b;
    layer0_outputs(6691) <= a;
    layer0_outputs(6692) <= '0';
    layer0_outputs(6693) <= not a;
    layer0_outputs(6694) <= not a or b;
    layer0_outputs(6695) <= a and b;
    layer0_outputs(6696) <= a;
    layer0_outputs(6697) <= not a or b;
    layer0_outputs(6698) <= not a or b;
    layer0_outputs(6699) <= a or b;
    layer0_outputs(6700) <= '1';
    layer0_outputs(6701) <= a or b;
    layer0_outputs(6702) <= a and b;
    layer0_outputs(6703) <= a xor b;
    layer0_outputs(6704) <= '0';
    layer0_outputs(6705) <= not (a and b);
    layer0_outputs(6706) <= a or b;
    layer0_outputs(6707) <= '0';
    layer0_outputs(6708) <= a xor b;
    layer0_outputs(6709) <= not a;
    layer0_outputs(6710) <= b and not a;
    layer0_outputs(6711) <= not b;
    layer0_outputs(6712) <= b;
    layer0_outputs(6713) <= a xor b;
    layer0_outputs(6714) <= not a or b;
    layer0_outputs(6715) <= a xor b;
    layer0_outputs(6716) <= not a;
    layer0_outputs(6717) <= b;
    layer0_outputs(6718) <= not b or a;
    layer0_outputs(6719) <= not a;
    layer0_outputs(6720) <= not b or a;
    layer0_outputs(6721) <= not (a and b);
    layer0_outputs(6722) <= '0';
    layer0_outputs(6723) <= a and b;
    layer0_outputs(6724) <= b and not a;
    layer0_outputs(6725) <= '0';
    layer0_outputs(6726) <= not b;
    layer0_outputs(6727) <= not b;
    layer0_outputs(6728) <= a and b;
    layer0_outputs(6729) <= a and b;
    layer0_outputs(6730) <= '0';
    layer0_outputs(6731) <= not a or b;
    layer0_outputs(6732) <= not b;
    layer0_outputs(6733) <= not (a xor b);
    layer0_outputs(6734) <= '0';
    layer0_outputs(6735) <= not a;
    layer0_outputs(6736) <= not b or a;
    layer0_outputs(6737) <= not a;
    layer0_outputs(6738) <= b;
    layer0_outputs(6739) <= a or b;
    layer0_outputs(6740) <= not (a xor b);
    layer0_outputs(6741) <= a xor b;
    layer0_outputs(6742) <= a;
    layer0_outputs(6743) <= '1';
    layer0_outputs(6744) <= '1';
    layer0_outputs(6745) <= not a or b;
    layer0_outputs(6746) <= b;
    layer0_outputs(6747) <= not b or a;
    layer0_outputs(6748) <= not (a xor b);
    layer0_outputs(6749) <= '0';
    layer0_outputs(6750) <= a xor b;
    layer0_outputs(6751) <= a or b;
    layer0_outputs(6752) <= a or b;
    layer0_outputs(6753) <= a and not b;
    layer0_outputs(6754) <= a or b;
    layer0_outputs(6755) <= '0';
    layer0_outputs(6756) <= not b or a;
    layer0_outputs(6757) <= not (a or b);
    layer0_outputs(6758) <= a or b;
    layer0_outputs(6759) <= a and not b;
    layer0_outputs(6760) <= a xor b;
    layer0_outputs(6761) <= '1';
    layer0_outputs(6762) <= not b;
    layer0_outputs(6763) <= not (a or b);
    layer0_outputs(6764) <= b;
    layer0_outputs(6765) <= not (a xor b);
    layer0_outputs(6766) <= a and b;
    layer0_outputs(6767) <= a or b;
    layer0_outputs(6768) <= not a;
    layer0_outputs(6769) <= a or b;
    layer0_outputs(6770) <= b;
    layer0_outputs(6771) <= not (a and b);
    layer0_outputs(6772) <= not (a and b);
    layer0_outputs(6773) <= a xor b;
    layer0_outputs(6774) <= not b;
    layer0_outputs(6775) <= a or b;
    layer0_outputs(6776) <= '0';
    layer0_outputs(6777) <= not (a or b);
    layer0_outputs(6778) <= a and b;
    layer0_outputs(6779) <= a and not b;
    layer0_outputs(6780) <= a xor b;
    layer0_outputs(6781) <= not a;
    layer0_outputs(6782) <= not a;
    layer0_outputs(6783) <= not b;
    layer0_outputs(6784) <= a or b;
    layer0_outputs(6785) <= a;
    layer0_outputs(6786) <= a;
    layer0_outputs(6787) <= a or b;
    layer0_outputs(6788) <= b and not a;
    layer0_outputs(6789) <= a or b;
    layer0_outputs(6790) <= a xor b;
    layer0_outputs(6791) <= a xor b;
    layer0_outputs(6792) <= '1';
    layer0_outputs(6793) <= not (a xor b);
    layer0_outputs(6794) <= '1';
    layer0_outputs(6795) <= b and not a;
    layer0_outputs(6796) <= b and not a;
    layer0_outputs(6797) <= '1';
    layer0_outputs(6798) <= not a or b;
    layer0_outputs(6799) <= not b or a;
    layer0_outputs(6800) <= not a or b;
    layer0_outputs(6801) <= '0';
    layer0_outputs(6802) <= not (a or b);
    layer0_outputs(6803) <= b;
    layer0_outputs(6804) <= a;
    layer0_outputs(6805) <= a xor b;
    layer0_outputs(6806) <= not (a or b);
    layer0_outputs(6807) <= a and b;
    layer0_outputs(6808) <= '0';
    layer0_outputs(6809) <= a xor b;
    layer0_outputs(6810) <= not b;
    layer0_outputs(6811) <= b and not a;
    layer0_outputs(6812) <= a and not b;
    layer0_outputs(6813) <= not (a or b);
    layer0_outputs(6814) <= a and not b;
    layer0_outputs(6815) <= not (a or b);
    layer0_outputs(6816) <= not b;
    layer0_outputs(6817) <= a xor b;
    layer0_outputs(6818) <= a and b;
    layer0_outputs(6819) <= '0';
    layer0_outputs(6820) <= not a or b;
    layer0_outputs(6821) <= '1';
    layer0_outputs(6822) <= '0';
    layer0_outputs(6823) <= a and b;
    layer0_outputs(6824) <= '1';
    layer0_outputs(6825) <= b;
    layer0_outputs(6826) <= not (a or b);
    layer0_outputs(6827) <= not a;
    layer0_outputs(6828) <= a or b;
    layer0_outputs(6829) <= not a;
    layer0_outputs(6830) <= a or b;
    layer0_outputs(6831) <= not b;
    layer0_outputs(6832) <= not a;
    layer0_outputs(6833) <= not (a or b);
    layer0_outputs(6834) <= not a or b;
    layer0_outputs(6835) <= a xor b;
    layer0_outputs(6836) <= not (a and b);
    layer0_outputs(6837) <= not b or a;
    layer0_outputs(6838) <= b;
    layer0_outputs(6839) <= a;
    layer0_outputs(6840) <= not (a or b);
    layer0_outputs(6841) <= a;
    layer0_outputs(6842) <= not b;
    layer0_outputs(6843) <= not b or a;
    layer0_outputs(6844) <= a and b;
    layer0_outputs(6845) <= b;
    layer0_outputs(6846) <= b and not a;
    layer0_outputs(6847) <= b;
    layer0_outputs(6848) <= not b;
    layer0_outputs(6849) <= '0';
    layer0_outputs(6850) <= not b;
    layer0_outputs(6851) <= a xor b;
    layer0_outputs(6852) <= not a or b;
    layer0_outputs(6853) <= not b;
    layer0_outputs(6854) <= not b or a;
    layer0_outputs(6855) <= not b or a;
    layer0_outputs(6856) <= a and b;
    layer0_outputs(6857) <= a;
    layer0_outputs(6858) <= '1';
    layer0_outputs(6859) <= not b or a;
    layer0_outputs(6860) <= b and not a;
    layer0_outputs(6861) <= not (a or b);
    layer0_outputs(6862) <= b;
    layer0_outputs(6863) <= not b or a;
    layer0_outputs(6864) <= not a or b;
    layer0_outputs(6865) <= not (a and b);
    layer0_outputs(6866) <= not (a or b);
    layer0_outputs(6867) <= not b;
    layer0_outputs(6868) <= '0';
    layer0_outputs(6869) <= a or b;
    layer0_outputs(6870) <= a;
    layer0_outputs(6871) <= a and not b;
    layer0_outputs(6872) <= b and not a;
    layer0_outputs(6873) <= not b or a;
    layer0_outputs(6874) <= b and not a;
    layer0_outputs(6875) <= '0';
    layer0_outputs(6876) <= a;
    layer0_outputs(6877) <= not (a or b);
    layer0_outputs(6878) <= not (a or b);
    layer0_outputs(6879) <= not (a and b);
    layer0_outputs(6880) <= a;
    layer0_outputs(6881) <= '0';
    layer0_outputs(6882) <= a xor b;
    layer0_outputs(6883) <= not b or a;
    layer0_outputs(6884) <= a and b;
    layer0_outputs(6885) <= b and not a;
    layer0_outputs(6886) <= not a or b;
    layer0_outputs(6887) <= a or b;
    layer0_outputs(6888) <= not (a or b);
    layer0_outputs(6889) <= a xor b;
    layer0_outputs(6890) <= a xor b;
    layer0_outputs(6891) <= not (a xor b);
    layer0_outputs(6892) <= '1';
    layer0_outputs(6893) <= a or b;
    layer0_outputs(6894) <= not (a xor b);
    layer0_outputs(6895) <= b;
    layer0_outputs(6896) <= not (a or b);
    layer0_outputs(6897) <= not (a and b);
    layer0_outputs(6898) <= a and not b;
    layer0_outputs(6899) <= a and not b;
    layer0_outputs(6900) <= a or b;
    layer0_outputs(6901) <= not a;
    layer0_outputs(6902) <= not b or a;
    layer0_outputs(6903) <= b;
    layer0_outputs(6904) <= '1';
    layer0_outputs(6905) <= a xor b;
    layer0_outputs(6906) <= b and not a;
    layer0_outputs(6907) <= not a or b;
    layer0_outputs(6908) <= not b or a;
    layer0_outputs(6909) <= not a or b;
    layer0_outputs(6910) <= not b or a;
    layer0_outputs(6911) <= a and b;
    layer0_outputs(6912) <= a xor b;
    layer0_outputs(6913) <= not a;
    layer0_outputs(6914) <= a;
    layer0_outputs(6915) <= b;
    layer0_outputs(6916) <= a or b;
    layer0_outputs(6917) <= a;
    layer0_outputs(6918) <= not b;
    layer0_outputs(6919) <= not (a or b);
    layer0_outputs(6920) <= not a or b;
    layer0_outputs(6921) <= a xor b;
    layer0_outputs(6922) <= b and not a;
    layer0_outputs(6923) <= b and not a;
    layer0_outputs(6924) <= not b or a;
    layer0_outputs(6925) <= a and b;
    layer0_outputs(6926) <= not b;
    layer0_outputs(6927) <= not b or a;
    layer0_outputs(6928) <= a and b;
    layer0_outputs(6929) <= a and not b;
    layer0_outputs(6930) <= a xor b;
    layer0_outputs(6931) <= b and not a;
    layer0_outputs(6932) <= not (a xor b);
    layer0_outputs(6933) <= a and b;
    layer0_outputs(6934) <= a xor b;
    layer0_outputs(6935) <= a;
    layer0_outputs(6936) <= a or b;
    layer0_outputs(6937) <= '0';
    layer0_outputs(6938) <= b and not a;
    layer0_outputs(6939) <= b;
    layer0_outputs(6940) <= a or b;
    layer0_outputs(6941) <= a or b;
    layer0_outputs(6942) <= not b or a;
    layer0_outputs(6943) <= b;
    layer0_outputs(6944) <= b;
    layer0_outputs(6945) <= a;
    layer0_outputs(6946) <= not (a or b);
    layer0_outputs(6947) <= not a;
    layer0_outputs(6948) <= not b;
    layer0_outputs(6949) <= '0';
    layer0_outputs(6950) <= not (a xor b);
    layer0_outputs(6951) <= b and not a;
    layer0_outputs(6952) <= a xor b;
    layer0_outputs(6953) <= a xor b;
    layer0_outputs(6954) <= a and not b;
    layer0_outputs(6955) <= '0';
    layer0_outputs(6956) <= b and not a;
    layer0_outputs(6957) <= a and not b;
    layer0_outputs(6958) <= a or b;
    layer0_outputs(6959) <= not (a and b);
    layer0_outputs(6960) <= a;
    layer0_outputs(6961) <= b;
    layer0_outputs(6962) <= not (a or b);
    layer0_outputs(6963) <= not (a or b);
    layer0_outputs(6964) <= a;
    layer0_outputs(6965) <= b;
    layer0_outputs(6966) <= not a;
    layer0_outputs(6967) <= not (a xor b);
    layer0_outputs(6968) <= '0';
    layer0_outputs(6969) <= not b;
    layer0_outputs(6970) <= b and not a;
    layer0_outputs(6971) <= not (a or b);
    layer0_outputs(6972) <= a xor b;
    layer0_outputs(6973) <= not b;
    layer0_outputs(6974) <= '0';
    layer0_outputs(6975) <= '0';
    layer0_outputs(6976) <= not (a or b);
    layer0_outputs(6977) <= not b;
    layer0_outputs(6978) <= a and not b;
    layer0_outputs(6979) <= not (a or b);
    layer0_outputs(6980) <= not b;
    layer0_outputs(6981) <= not b or a;
    layer0_outputs(6982) <= a;
    layer0_outputs(6983) <= a or b;
    layer0_outputs(6984) <= a xor b;
    layer0_outputs(6985) <= a or b;
    layer0_outputs(6986) <= not b;
    layer0_outputs(6987) <= a and not b;
    layer0_outputs(6988) <= not b or a;
    layer0_outputs(6989) <= a and not b;
    layer0_outputs(6990) <= not b;
    layer0_outputs(6991) <= not (a or b);
    layer0_outputs(6992) <= '0';
    layer0_outputs(6993) <= not (a or b);
    layer0_outputs(6994) <= a;
    layer0_outputs(6995) <= a and not b;
    layer0_outputs(6996) <= a;
    layer0_outputs(6997) <= a xor b;
    layer0_outputs(6998) <= not a;
    layer0_outputs(6999) <= a and not b;
    layer0_outputs(7000) <= not (a and b);
    layer0_outputs(7001) <= not a or b;
    layer0_outputs(7002) <= '0';
    layer0_outputs(7003) <= not a or b;
    layer0_outputs(7004) <= not b or a;
    layer0_outputs(7005) <= not b;
    layer0_outputs(7006) <= not b or a;
    layer0_outputs(7007) <= not (a or b);
    layer0_outputs(7008) <= not b or a;
    layer0_outputs(7009) <= a and not b;
    layer0_outputs(7010) <= not (a and b);
    layer0_outputs(7011) <= b;
    layer0_outputs(7012) <= not (a or b);
    layer0_outputs(7013) <= a or b;
    layer0_outputs(7014) <= '0';
    layer0_outputs(7015) <= not b or a;
    layer0_outputs(7016) <= not (a and b);
    layer0_outputs(7017) <= a and not b;
    layer0_outputs(7018) <= b;
    layer0_outputs(7019) <= not (a or b);
    layer0_outputs(7020) <= a;
    layer0_outputs(7021) <= not (a or b);
    layer0_outputs(7022) <= not (a xor b);
    layer0_outputs(7023) <= a or b;
    layer0_outputs(7024) <= a;
    layer0_outputs(7025) <= not (a xor b);
    layer0_outputs(7026) <= not (a or b);
    layer0_outputs(7027) <= not b or a;
    layer0_outputs(7028) <= not b or a;
    layer0_outputs(7029) <= not a;
    layer0_outputs(7030) <= not (a and b);
    layer0_outputs(7031) <= b and not a;
    layer0_outputs(7032) <= '1';
    layer0_outputs(7033) <= not b or a;
    layer0_outputs(7034) <= a and not b;
    layer0_outputs(7035) <= b;
    layer0_outputs(7036) <= not a or b;
    layer0_outputs(7037) <= '0';
    layer0_outputs(7038) <= not (a xor b);
    layer0_outputs(7039) <= a and not b;
    layer0_outputs(7040) <= not (a and b);
    layer0_outputs(7041) <= not a;
    layer0_outputs(7042) <= not a;
    layer0_outputs(7043) <= a or b;
    layer0_outputs(7044) <= not (a and b);
    layer0_outputs(7045) <= not b;
    layer0_outputs(7046) <= b;
    layer0_outputs(7047) <= not (a and b);
    layer0_outputs(7048) <= not a;
    layer0_outputs(7049) <= b;
    layer0_outputs(7050) <= b and not a;
    layer0_outputs(7051) <= a;
    layer0_outputs(7052) <= a;
    layer0_outputs(7053) <= a and not b;
    layer0_outputs(7054) <= a or b;
    layer0_outputs(7055) <= b;
    layer0_outputs(7056) <= '1';
    layer0_outputs(7057) <= not (a xor b);
    layer0_outputs(7058) <= not b;
    layer0_outputs(7059) <= b;
    layer0_outputs(7060) <= a and not b;
    layer0_outputs(7061) <= not b;
    layer0_outputs(7062) <= a;
    layer0_outputs(7063) <= '1';
    layer0_outputs(7064) <= not b;
    layer0_outputs(7065) <= a and not b;
    layer0_outputs(7066) <= not b or a;
    layer0_outputs(7067) <= not (a and b);
    layer0_outputs(7068) <= a;
    layer0_outputs(7069) <= a;
    layer0_outputs(7070) <= b;
    layer0_outputs(7071) <= not a or b;
    layer0_outputs(7072) <= b and not a;
    layer0_outputs(7073) <= a xor b;
    layer0_outputs(7074) <= not a or b;
    layer0_outputs(7075) <= b;
    layer0_outputs(7076) <= a;
    layer0_outputs(7077) <= b;
    layer0_outputs(7078) <= not a;
    layer0_outputs(7079) <= not a or b;
    layer0_outputs(7080) <= not (a and b);
    layer0_outputs(7081) <= not (a and b);
    layer0_outputs(7082) <= a or b;
    layer0_outputs(7083) <= not (a and b);
    layer0_outputs(7084) <= b;
    layer0_outputs(7085) <= not (a xor b);
    layer0_outputs(7086) <= a xor b;
    layer0_outputs(7087) <= not (a and b);
    layer0_outputs(7088) <= a and b;
    layer0_outputs(7089) <= not (a or b);
    layer0_outputs(7090) <= a or b;
    layer0_outputs(7091) <= not b or a;
    layer0_outputs(7092) <= a or b;
    layer0_outputs(7093) <= not b;
    layer0_outputs(7094) <= a or b;
    layer0_outputs(7095) <= a or b;
    layer0_outputs(7096) <= '0';
    layer0_outputs(7097) <= not (a and b);
    layer0_outputs(7098) <= not b;
    layer0_outputs(7099) <= '0';
    layer0_outputs(7100) <= not b;
    layer0_outputs(7101) <= a xor b;
    layer0_outputs(7102) <= a and b;
    layer0_outputs(7103) <= a and not b;
    layer0_outputs(7104) <= a and not b;
    layer0_outputs(7105) <= a and b;
    layer0_outputs(7106) <= not b or a;
    layer0_outputs(7107) <= '1';
    layer0_outputs(7108) <= not (a and b);
    layer0_outputs(7109) <= not a;
    layer0_outputs(7110) <= a or b;
    layer0_outputs(7111) <= not (a or b);
    layer0_outputs(7112) <= not (a and b);
    layer0_outputs(7113) <= a;
    layer0_outputs(7114) <= b and not a;
    layer0_outputs(7115) <= not (a and b);
    layer0_outputs(7116) <= b;
    layer0_outputs(7117) <= not a or b;
    layer0_outputs(7118) <= a;
    layer0_outputs(7119) <= not b or a;
    layer0_outputs(7120) <= a and b;
    layer0_outputs(7121) <= a;
    layer0_outputs(7122) <= a and b;
    layer0_outputs(7123) <= not (a xor b);
    layer0_outputs(7124) <= a or b;
    layer0_outputs(7125) <= not b;
    layer0_outputs(7126) <= a or b;
    layer0_outputs(7127) <= a or b;
    layer0_outputs(7128) <= a xor b;
    layer0_outputs(7129) <= not (a xor b);
    layer0_outputs(7130) <= not a or b;
    layer0_outputs(7131) <= not (a or b);
    layer0_outputs(7132) <= b;
    layer0_outputs(7133) <= not b or a;
    layer0_outputs(7134) <= a xor b;
    layer0_outputs(7135) <= b and not a;
    layer0_outputs(7136) <= not (a or b);
    layer0_outputs(7137) <= a or b;
    layer0_outputs(7138) <= a xor b;
    layer0_outputs(7139) <= b and not a;
    layer0_outputs(7140) <= not a or b;
    layer0_outputs(7141) <= b;
    layer0_outputs(7142) <= b;
    layer0_outputs(7143) <= not (a xor b);
    layer0_outputs(7144) <= not (a or b);
    layer0_outputs(7145) <= not (a xor b);
    layer0_outputs(7146) <= b and not a;
    layer0_outputs(7147) <= a or b;
    layer0_outputs(7148) <= b and not a;
    layer0_outputs(7149) <= a and not b;
    layer0_outputs(7150) <= '1';
    layer0_outputs(7151) <= not (a or b);
    layer0_outputs(7152) <= not (a or b);
    layer0_outputs(7153) <= not a or b;
    layer0_outputs(7154) <= a xor b;
    layer0_outputs(7155) <= not (a or b);
    layer0_outputs(7156) <= a and not b;
    layer0_outputs(7157) <= not b;
    layer0_outputs(7158) <= not b;
    layer0_outputs(7159) <= b;
    layer0_outputs(7160) <= '0';
    layer0_outputs(7161) <= not (a or b);
    layer0_outputs(7162) <= '1';
    layer0_outputs(7163) <= a xor b;
    layer0_outputs(7164) <= not (a or b);
    layer0_outputs(7165) <= a and b;
    layer0_outputs(7166) <= not (a or b);
    layer0_outputs(7167) <= b;
    layer0_outputs(7168) <= '0';
    layer0_outputs(7169) <= a and b;
    layer0_outputs(7170) <= a or b;
    layer0_outputs(7171) <= not a or b;
    layer0_outputs(7172) <= a xor b;
    layer0_outputs(7173) <= a and not b;
    layer0_outputs(7174) <= not (a xor b);
    layer0_outputs(7175) <= '1';
    layer0_outputs(7176) <= not a or b;
    layer0_outputs(7177) <= not (a and b);
    layer0_outputs(7178) <= b;
    layer0_outputs(7179) <= b;
    layer0_outputs(7180) <= not (a or b);
    layer0_outputs(7181) <= not (a or b);
    layer0_outputs(7182) <= not a;
    layer0_outputs(7183) <= not a or b;
    layer0_outputs(7184) <= '0';
    layer0_outputs(7185) <= a and b;
    layer0_outputs(7186) <= not b;
    layer0_outputs(7187) <= '1';
    layer0_outputs(7188) <= '0';
    layer0_outputs(7189) <= a or b;
    layer0_outputs(7190) <= not a or b;
    layer0_outputs(7191) <= b;
    layer0_outputs(7192) <= a or b;
    layer0_outputs(7193) <= '0';
    layer0_outputs(7194) <= not a or b;
    layer0_outputs(7195) <= b and not a;
    layer0_outputs(7196) <= '1';
    layer0_outputs(7197) <= not a;
    layer0_outputs(7198) <= '1';
    layer0_outputs(7199) <= not b;
    layer0_outputs(7200) <= not a or b;
    layer0_outputs(7201) <= a xor b;
    layer0_outputs(7202) <= not (a or b);
    layer0_outputs(7203) <= not b or a;
    layer0_outputs(7204) <= not (a or b);
    layer0_outputs(7205) <= not b or a;
    layer0_outputs(7206) <= not (a and b);
    layer0_outputs(7207) <= not a or b;
    layer0_outputs(7208) <= not (a xor b);
    layer0_outputs(7209) <= b and not a;
    layer0_outputs(7210) <= not b or a;
    layer0_outputs(7211) <= a or b;
    layer0_outputs(7212) <= a or b;
    layer0_outputs(7213) <= '1';
    layer0_outputs(7214) <= not (a xor b);
    layer0_outputs(7215) <= not (a or b);
    layer0_outputs(7216) <= not b or a;
    layer0_outputs(7217) <= not a;
    layer0_outputs(7218) <= not b or a;
    layer0_outputs(7219) <= a and not b;
    layer0_outputs(7220) <= not a;
    layer0_outputs(7221) <= not (a and b);
    layer0_outputs(7222) <= not b or a;
    layer0_outputs(7223) <= a xor b;
    layer0_outputs(7224) <= b and not a;
    layer0_outputs(7225) <= a;
    layer0_outputs(7226) <= b;
    layer0_outputs(7227) <= b;
    layer0_outputs(7228) <= not (a or b);
    layer0_outputs(7229) <= a;
    layer0_outputs(7230) <= not b;
    layer0_outputs(7231) <= b and not a;
    layer0_outputs(7232) <= a;
    layer0_outputs(7233) <= not b or a;
    layer0_outputs(7234) <= not (a xor b);
    layer0_outputs(7235) <= a and not b;
    layer0_outputs(7236) <= a;
    layer0_outputs(7237) <= a and not b;
    layer0_outputs(7238) <= not (a and b);
    layer0_outputs(7239) <= a;
    layer0_outputs(7240) <= a xor b;
    layer0_outputs(7241) <= not (a or b);
    layer0_outputs(7242) <= a or b;
    layer0_outputs(7243) <= '0';
    layer0_outputs(7244) <= not b or a;
    layer0_outputs(7245) <= not b or a;
    layer0_outputs(7246) <= not b;
    layer0_outputs(7247) <= a or b;
    layer0_outputs(7248) <= a xor b;
    layer0_outputs(7249) <= not (a and b);
    layer0_outputs(7250) <= not (a xor b);
    layer0_outputs(7251) <= not (a xor b);
    layer0_outputs(7252) <= not b;
    layer0_outputs(7253) <= '1';
    layer0_outputs(7254) <= not (a and b);
    layer0_outputs(7255) <= b and not a;
    layer0_outputs(7256) <= not (a or b);
    layer0_outputs(7257) <= not (a xor b);
    layer0_outputs(7258) <= not (a xor b);
    layer0_outputs(7259) <= not (a xor b);
    layer0_outputs(7260) <= not (a xor b);
    layer0_outputs(7261) <= a and b;
    layer0_outputs(7262) <= a;
    layer0_outputs(7263) <= a or b;
    layer0_outputs(7264) <= not b;
    layer0_outputs(7265) <= b and not a;
    layer0_outputs(7266) <= a and b;
    layer0_outputs(7267) <= a;
    layer0_outputs(7268) <= not a;
    layer0_outputs(7269) <= a xor b;
    layer0_outputs(7270) <= not (a and b);
    layer0_outputs(7271) <= b;
    layer0_outputs(7272) <= not b or a;
    layer0_outputs(7273) <= '0';
    layer0_outputs(7274) <= '1';
    layer0_outputs(7275) <= b and not a;
    layer0_outputs(7276) <= '0';
    layer0_outputs(7277) <= a and not b;
    layer0_outputs(7278) <= not a;
    layer0_outputs(7279) <= not b;
    layer0_outputs(7280) <= not b;
    layer0_outputs(7281) <= b and not a;
    layer0_outputs(7282) <= b;
    layer0_outputs(7283) <= not (a xor b);
    layer0_outputs(7284) <= '0';
    layer0_outputs(7285) <= not a;
    layer0_outputs(7286) <= not a;
    layer0_outputs(7287) <= '0';
    layer0_outputs(7288) <= a or b;
    layer0_outputs(7289) <= b;
    layer0_outputs(7290) <= a and b;
    layer0_outputs(7291) <= '1';
    layer0_outputs(7292) <= not b or a;
    layer0_outputs(7293) <= b and not a;
    layer0_outputs(7294) <= '1';
    layer0_outputs(7295) <= a xor b;
    layer0_outputs(7296) <= a;
    layer0_outputs(7297) <= not a or b;
    layer0_outputs(7298) <= a or b;
    layer0_outputs(7299) <= '1';
    layer0_outputs(7300) <= a or b;
    layer0_outputs(7301) <= not (a and b);
    layer0_outputs(7302) <= not a or b;
    layer0_outputs(7303) <= b;
    layer0_outputs(7304) <= a and not b;
    layer0_outputs(7305) <= a xor b;
    layer0_outputs(7306) <= not (a or b);
    layer0_outputs(7307) <= b;
    layer0_outputs(7308) <= '1';
    layer0_outputs(7309) <= b;
    layer0_outputs(7310) <= not a or b;
    layer0_outputs(7311) <= not b;
    layer0_outputs(7312) <= b and not a;
    layer0_outputs(7313) <= '0';
    layer0_outputs(7314) <= a xor b;
    layer0_outputs(7315) <= not a;
    layer0_outputs(7316) <= a;
    layer0_outputs(7317) <= a or b;
    layer0_outputs(7318) <= not b;
    layer0_outputs(7319) <= not b or a;
    layer0_outputs(7320) <= not b;
    layer0_outputs(7321) <= not b;
    layer0_outputs(7322) <= a and not b;
    layer0_outputs(7323) <= not (a or b);
    layer0_outputs(7324) <= b and not a;
    layer0_outputs(7325) <= a xor b;
    layer0_outputs(7326) <= not a;
    layer0_outputs(7327) <= a and not b;
    layer0_outputs(7328) <= a;
    layer0_outputs(7329) <= not (a xor b);
    layer0_outputs(7330) <= not (a or b);
    layer0_outputs(7331) <= not (a or b);
    layer0_outputs(7332) <= not (a or b);
    layer0_outputs(7333) <= not a or b;
    layer0_outputs(7334) <= '0';
    layer0_outputs(7335) <= not b;
    layer0_outputs(7336) <= b;
    layer0_outputs(7337) <= not b or a;
    layer0_outputs(7338) <= not a or b;
    layer0_outputs(7339) <= b;
    layer0_outputs(7340) <= not b;
    layer0_outputs(7341) <= a and not b;
    layer0_outputs(7342) <= '0';
    layer0_outputs(7343) <= not b;
    layer0_outputs(7344) <= not b;
    layer0_outputs(7345) <= not a;
    layer0_outputs(7346) <= not a or b;
    layer0_outputs(7347) <= a or b;
    layer0_outputs(7348) <= a and not b;
    layer0_outputs(7349) <= not (a xor b);
    layer0_outputs(7350) <= a xor b;
    layer0_outputs(7351) <= not b;
    layer0_outputs(7352) <= a;
    layer0_outputs(7353) <= not b;
    layer0_outputs(7354) <= a or b;
    layer0_outputs(7355) <= not b or a;
    layer0_outputs(7356) <= not a;
    layer0_outputs(7357) <= not a;
    layer0_outputs(7358) <= not b;
    layer0_outputs(7359) <= not (a and b);
    layer0_outputs(7360) <= a and not b;
    layer0_outputs(7361) <= a;
    layer0_outputs(7362) <= not a or b;
    layer0_outputs(7363) <= not a;
    layer0_outputs(7364) <= b and not a;
    layer0_outputs(7365) <= not b;
    layer0_outputs(7366) <= '0';
    layer0_outputs(7367) <= not b;
    layer0_outputs(7368) <= '0';
    layer0_outputs(7369) <= not b;
    layer0_outputs(7370) <= a and not b;
    layer0_outputs(7371) <= '0';
    layer0_outputs(7372) <= '0';
    layer0_outputs(7373) <= a;
    layer0_outputs(7374) <= a and b;
    layer0_outputs(7375) <= a or b;
    layer0_outputs(7376) <= a xor b;
    layer0_outputs(7377) <= b and not a;
    layer0_outputs(7378) <= '0';
    layer0_outputs(7379) <= '1';
    layer0_outputs(7380) <= not b;
    layer0_outputs(7381) <= not a or b;
    layer0_outputs(7382) <= not (a or b);
    layer0_outputs(7383) <= not (a and b);
    layer0_outputs(7384) <= not b;
    layer0_outputs(7385) <= not b or a;
    layer0_outputs(7386) <= not (a or b);
    layer0_outputs(7387) <= a xor b;
    layer0_outputs(7388) <= a and b;
    layer0_outputs(7389) <= a and not b;
    layer0_outputs(7390) <= '1';
    layer0_outputs(7391) <= not (a or b);
    layer0_outputs(7392) <= a and b;
    layer0_outputs(7393) <= b;
    layer0_outputs(7394) <= b;
    layer0_outputs(7395) <= '0';
    layer0_outputs(7396) <= a and b;
    layer0_outputs(7397) <= not b;
    layer0_outputs(7398) <= a;
    layer0_outputs(7399) <= b;
    layer0_outputs(7400) <= b;
    layer0_outputs(7401) <= a and b;
    layer0_outputs(7402) <= not (a or b);
    layer0_outputs(7403) <= '0';
    layer0_outputs(7404) <= not (a xor b);
    layer0_outputs(7405) <= b and not a;
    layer0_outputs(7406) <= not (a or b);
    layer0_outputs(7407) <= '0';
    layer0_outputs(7408) <= b and not a;
    layer0_outputs(7409) <= a and not b;
    layer0_outputs(7410) <= '1';
    layer0_outputs(7411) <= '1';
    layer0_outputs(7412) <= not (a xor b);
    layer0_outputs(7413) <= not a or b;
    layer0_outputs(7414) <= not a or b;
    layer0_outputs(7415) <= not (a and b);
    layer0_outputs(7416) <= b and not a;
    layer0_outputs(7417) <= not b;
    layer0_outputs(7418) <= a and b;
    layer0_outputs(7419) <= not (a or b);
    layer0_outputs(7420) <= a;
    layer0_outputs(7421) <= '1';
    layer0_outputs(7422) <= not a or b;
    layer0_outputs(7423) <= a or b;
    layer0_outputs(7424) <= not b;
    layer0_outputs(7425) <= not b or a;
    layer0_outputs(7426) <= not a;
    layer0_outputs(7427) <= not (a xor b);
    layer0_outputs(7428) <= a and not b;
    layer0_outputs(7429) <= not (a and b);
    layer0_outputs(7430) <= a xor b;
    layer0_outputs(7431) <= a and not b;
    layer0_outputs(7432) <= a or b;
    layer0_outputs(7433) <= a or b;
    layer0_outputs(7434) <= not (a and b);
    layer0_outputs(7435) <= b;
    layer0_outputs(7436) <= not (a and b);
    layer0_outputs(7437) <= not b;
    layer0_outputs(7438) <= a and not b;
    layer0_outputs(7439) <= not (a xor b);
    layer0_outputs(7440) <= not (a xor b);
    layer0_outputs(7441) <= not (a xor b);
    layer0_outputs(7442) <= a xor b;
    layer0_outputs(7443) <= not (a or b);
    layer0_outputs(7444) <= b and not a;
    layer0_outputs(7445) <= a and b;
    layer0_outputs(7446) <= not b;
    layer0_outputs(7447) <= not a;
    layer0_outputs(7448) <= a;
    layer0_outputs(7449) <= not b;
    layer0_outputs(7450) <= '1';
    layer0_outputs(7451) <= a xor b;
    layer0_outputs(7452) <= a or b;
    layer0_outputs(7453) <= '1';
    layer0_outputs(7454) <= '1';
    layer0_outputs(7455) <= b and not a;
    layer0_outputs(7456) <= not (a xor b);
    layer0_outputs(7457) <= a or b;
    layer0_outputs(7458) <= a or b;
    layer0_outputs(7459) <= not b;
    layer0_outputs(7460) <= a or b;
    layer0_outputs(7461) <= not (a or b);
    layer0_outputs(7462) <= a or b;
    layer0_outputs(7463) <= a xor b;
    layer0_outputs(7464) <= b;
    layer0_outputs(7465) <= a and not b;
    layer0_outputs(7466) <= not a;
    layer0_outputs(7467) <= not (a or b);
    layer0_outputs(7468) <= b;
    layer0_outputs(7469) <= not b or a;
    layer0_outputs(7470) <= a and not b;
    layer0_outputs(7471) <= b;
    layer0_outputs(7472) <= not a or b;
    layer0_outputs(7473) <= not (a and b);
    layer0_outputs(7474) <= b;
    layer0_outputs(7475) <= not (a xor b);
    layer0_outputs(7476) <= a and b;
    layer0_outputs(7477) <= not b or a;
    layer0_outputs(7478) <= a or b;
    layer0_outputs(7479) <= not b;
    layer0_outputs(7480) <= '1';
    layer0_outputs(7481) <= not a;
    layer0_outputs(7482) <= not a;
    layer0_outputs(7483) <= a xor b;
    layer0_outputs(7484) <= '0';
    layer0_outputs(7485) <= a xor b;
    layer0_outputs(7486) <= not (a and b);
    layer0_outputs(7487) <= '1';
    layer0_outputs(7488) <= not b;
    layer0_outputs(7489) <= not a;
    layer0_outputs(7490) <= not (a or b);
    layer0_outputs(7491) <= not (a xor b);
    layer0_outputs(7492) <= not (a xor b);
    layer0_outputs(7493) <= a and b;
    layer0_outputs(7494) <= not (a xor b);
    layer0_outputs(7495) <= a;
    layer0_outputs(7496) <= not b;
    layer0_outputs(7497) <= not a or b;
    layer0_outputs(7498) <= '0';
    layer0_outputs(7499) <= not a;
    layer0_outputs(7500) <= not (a or b);
    layer0_outputs(7501) <= b;
    layer0_outputs(7502) <= a;
    layer0_outputs(7503) <= not (a or b);
    layer0_outputs(7504) <= a;
    layer0_outputs(7505) <= a and not b;
    layer0_outputs(7506) <= b and not a;
    layer0_outputs(7507) <= a;
    layer0_outputs(7508) <= not a;
    layer0_outputs(7509) <= a;
    layer0_outputs(7510) <= a;
    layer0_outputs(7511) <= a xor b;
    layer0_outputs(7512) <= b and not a;
    layer0_outputs(7513) <= b and not a;
    layer0_outputs(7514) <= a and b;
    layer0_outputs(7515) <= b;
    layer0_outputs(7516) <= not a or b;
    layer0_outputs(7517) <= a and not b;
    layer0_outputs(7518) <= not (a xor b);
    layer0_outputs(7519) <= not b;
    layer0_outputs(7520) <= a and not b;
    layer0_outputs(7521) <= a xor b;
    layer0_outputs(7522) <= a;
    layer0_outputs(7523) <= '1';
    layer0_outputs(7524) <= not a or b;
    layer0_outputs(7525) <= not (a xor b);
    layer0_outputs(7526) <= not (a or b);
    layer0_outputs(7527) <= '1';
    layer0_outputs(7528) <= '1';
    layer0_outputs(7529) <= a and b;
    layer0_outputs(7530) <= not b or a;
    layer0_outputs(7531) <= a or b;
    layer0_outputs(7532) <= a and not b;
    layer0_outputs(7533) <= a xor b;
    layer0_outputs(7534) <= a;
    layer0_outputs(7535) <= a xor b;
    layer0_outputs(7536) <= not a or b;
    layer0_outputs(7537) <= b;
    layer0_outputs(7538) <= not b;
    layer0_outputs(7539) <= not (a or b);
    layer0_outputs(7540) <= b;
    layer0_outputs(7541) <= not (a xor b);
    layer0_outputs(7542) <= not a or b;
    layer0_outputs(7543) <= not (a and b);
    layer0_outputs(7544) <= not (a xor b);
    layer0_outputs(7545) <= b;
    layer0_outputs(7546) <= not a;
    layer0_outputs(7547) <= not a;
    layer0_outputs(7548) <= not b;
    layer0_outputs(7549) <= a or b;
    layer0_outputs(7550) <= b and not a;
    layer0_outputs(7551) <= '1';
    layer0_outputs(7552) <= not (a or b);
    layer0_outputs(7553) <= not (a xor b);
    layer0_outputs(7554) <= not a or b;
    layer0_outputs(7555) <= a and b;
    layer0_outputs(7556) <= a and b;
    layer0_outputs(7557) <= b;
    layer0_outputs(7558) <= a or b;
    layer0_outputs(7559) <= not a;
    layer0_outputs(7560) <= b and not a;
    layer0_outputs(7561) <= not (a and b);
    layer0_outputs(7562) <= b;
    layer0_outputs(7563) <= '1';
    layer0_outputs(7564) <= a;
    layer0_outputs(7565) <= not a;
    layer0_outputs(7566) <= not a or b;
    layer0_outputs(7567) <= not (a xor b);
    layer0_outputs(7568) <= b and not a;
    layer0_outputs(7569) <= not a;
    layer0_outputs(7570) <= a and not b;
    layer0_outputs(7571) <= a and not b;
    layer0_outputs(7572) <= '0';
    layer0_outputs(7573) <= b and not a;
    layer0_outputs(7574) <= not (a or b);
    layer0_outputs(7575) <= b;
    layer0_outputs(7576) <= a;
    layer0_outputs(7577) <= a and not b;
    layer0_outputs(7578) <= b;
    layer0_outputs(7579) <= not a;
    layer0_outputs(7580) <= a;
    layer0_outputs(7581) <= a;
    layer0_outputs(7582) <= not a or b;
    layer0_outputs(7583) <= not (a and b);
    layer0_outputs(7584) <= not (a and b);
    layer0_outputs(7585) <= not (a or b);
    layer0_outputs(7586) <= a;
    layer0_outputs(7587) <= not a;
    layer0_outputs(7588) <= '1';
    layer0_outputs(7589) <= b and not a;
    layer0_outputs(7590) <= not (a or b);
    layer0_outputs(7591) <= not a;
    layer0_outputs(7592) <= b;
    layer0_outputs(7593) <= b and not a;
    layer0_outputs(7594) <= b;
    layer0_outputs(7595) <= b and not a;
    layer0_outputs(7596) <= a xor b;
    layer0_outputs(7597) <= not b or a;
    layer0_outputs(7598) <= not (a xor b);
    layer0_outputs(7599) <= not (a and b);
    layer0_outputs(7600) <= a or b;
    layer0_outputs(7601) <= b;
    layer0_outputs(7602) <= not (a or b);
    layer0_outputs(7603) <= '1';
    layer0_outputs(7604) <= a and not b;
    layer0_outputs(7605) <= not b or a;
    layer0_outputs(7606) <= not a;
    layer0_outputs(7607) <= a or b;
    layer0_outputs(7608) <= a;
    layer0_outputs(7609) <= '1';
    layer0_outputs(7610) <= not (a and b);
    layer0_outputs(7611) <= a;
    layer0_outputs(7612) <= '1';
    layer0_outputs(7613) <= a and not b;
    layer0_outputs(7614) <= not (a or b);
    layer0_outputs(7615) <= a xor b;
    layer0_outputs(7616) <= not a or b;
    layer0_outputs(7617) <= not (a or b);
    layer0_outputs(7618) <= b and not a;
    layer0_outputs(7619) <= b;
    layer0_outputs(7620) <= not b or a;
    layer0_outputs(7621) <= not b;
    layer0_outputs(7622) <= a and not b;
    layer0_outputs(7623) <= not a;
    layer0_outputs(7624) <= a xor b;
    layer0_outputs(7625) <= b;
    layer0_outputs(7626) <= a or b;
    layer0_outputs(7627) <= b and not a;
    layer0_outputs(7628) <= not (a xor b);
    layer0_outputs(7629) <= a or b;
    layer0_outputs(7630) <= not b;
    layer0_outputs(7631) <= not (a or b);
    layer0_outputs(7632) <= not (a or b);
    layer0_outputs(7633) <= not a or b;
    layer0_outputs(7634) <= not (a or b);
    layer0_outputs(7635) <= a and b;
    layer0_outputs(7636) <= '0';
    layer0_outputs(7637) <= b and not a;
    layer0_outputs(7638) <= b;
    layer0_outputs(7639) <= a xor b;
    layer0_outputs(7640) <= a xor b;
    layer0_outputs(7641) <= not a or b;
    layer0_outputs(7642) <= a xor b;
    layer0_outputs(7643) <= not a or b;
    layer0_outputs(7644) <= b and not a;
    layer0_outputs(7645) <= '0';
    layer0_outputs(7646) <= not b;
    layer0_outputs(7647) <= not (a xor b);
    layer0_outputs(7648) <= a xor b;
    layer0_outputs(7649) <= not (a or b);
    layer0_outputs(7650) <= not a or b;
    layer0_outputs(7651) <= not (a xor b);
    layer0_outputs(7652) <= a and not b;
    layer0_outputs(7653) <= not (a xor b);
    layer0_outputs(7654) <= not a or b;
    layer0_outputs(7655) <= not a;
    layer0_outputs(7656) <= b and not a;
    layer0_outputs(7657) <= a and b;
    layer0_outputs(7658) <= a and not b;
    layer0_outputs(7659) <= a;
    layer0_outputs(7660) <= not a;
    layer0_outputs(7661) <= not a;
    layer0_outputs(7662) <= a;
    layer0_outputs(7663) <= not (a or b);
    layer0_outputs(7664) <= not a;
    layer0_outputs(7665) <= b;
    layer0_outputs(7666) <= a xor b;
    layer0_outputs(7667) <= a and b;
    layer0_outputs(7668) <= a xor b;
    layer0_outputs(7669) <= not a or b;
    layer0_outputs(7670) <= not a;
    layer0_outputs(7671) <= not b;
    layer0_outputs(7672) <= a xor b;
    layer0_outputs(7673) <= a xor b;
    layer0_outputs(7674) <= a xor b;
    layer0_outputs(7675) <= a xor b;
    layer0_outputs(7676) <= a or b;
    layer0_outputs(7677) <= a;
    layer0_outputs(7678) <= a and b;
    layer0_outputs(7679) <= not (a xor b);
    layer0_outputs(7680) <= not (a or b);
    layer0_outputs(7681) <= a;
    layer0_outputs(7682) <= a;
    layer0_outputs(7683) <= a or b;
    layer0_outputs(7684) <= not b;
    layer0_outputs(7685) <= not b;
    layer0_outputs(7686) <= not a or b;
    layer0_outputs(7687) <= not (a and b);
    layer0_outputs(7688) <= not (a xor b);
    layer0_outputs(7689) <= '0';
    layer0_outputs(7690) <= not a or b;
    layer0_outputs(7691) <= not a;
    layer0_outputs(7692) <= not (a xor b);
    layer0_outputs(7693) <= '0';
    layer0_outputs(7694) <= not b or a;
    layer0_outputs(7695) <= a and b;
    layer0_outputs(7696) <= not (a xor b);
    layer0_outputs(7697) <= a and not b;
    layer0_outputs(7698) <= b;
    layer0_outputs(7699) <= b;
    layer0_outputs(7700) <= not (a and b);
    layer0_outputs(7701) <= '1';
    layer0_outputs(7702) <= '1';
    layer0_outputs(7703) <= not (a xor b);
    layer0_outputs(7704) <= not (a or b);
    layer0_outputs(7705) <= a;
    layer0_outputs(7706) <= a or b;
    layer0_outputs(7707) <= '0';
    layer0_outputs(7708) <= not a or b;
    layer0_outputs(7709) <= not (a xor b);
    layer0_outputs(7710) <= not a or b;
    layer0_outputs(7711) <= '1';
    layer0_outputs(7712) <= a and b;
    layer0_outputs(7713) <= b and not a;
    layer0_outputs(7714) <= b and not a;
    layer0_outputs(7715) <= '1';
    layer0_outputs(7716) <= a xor b;
    layer0_outputs(7717) <= a xor b;
    layer0_outputs(7718) <= b and not a;
    layer0_outputs(7719) <= not b or a;
    layer0_outputs(7720) <= b;
    layer0_outputs(7721) <= not a;
    layer0_outputs(7722) <= a and b;
    layer0_outputs(7723) <= b and not a;
    layer0_outputs(7724) <= a;
    layer0_outputs(7725) <= a xor b;
    layer0_outputs(7726) <= b and not a;
    layer0_outputs(7727) <= not (a xor b);
    layer0_outputs(7728) <= '1';
    layer0_outputs(7729) <= '0';
    layer0_outputs(7730) <= not (a xor b);
    layer0_outputs(7731) <= a;
    layer0_outputs(7732) <= not a or b;
    layer0_outputs(7733) <= a and not b;
    layer0_outputs(7734) <= a xor b;
    layer0_outputs(7735) <= not (a xor b);
    layer0_outputs(7736) <= not b;
    layer0_outputs(7737) <= a and not b;
    layer0_outputs(7738) <= not (a or b);
    layer0_outputs(7739) <= a and b;
    layer0_outputs(7740) <= a xor b;
    layer0_outputs(7741) <= not (a and b);
    layer0_outputs(7742) <= a or b;
    layer0_outputs(7743) <= a xor b;
    layer0_outputs(7744) <= not (a and b);
    layer0_outputs(7745) <= b and not a;
    layer0_outputs(7746) <= b and not a;
    layer0_outputs(7747) <= a or b;
    layer0_outputs(7748) <= b;
    layer0_outputs(7749) <= a xor b;
    layer0_outputs(7750) <= b;
    layer0_outputs(7751) <= not (a or b);
    layer0_outputs(7752) <= a or b;
    layer0_outputs(7753) <= not a or b;
    layer0_outputs(7754) <= not a;
    layer0_outputs(7755) <= not b or a;
    layer0_outputs(7756) <= b;
    layer0_outputs(7757) <= a and b;
    layer0_outputs(7758) <= a xor b;
    layer0_outputs(7759) <= not (a xor b);
    layer0_outputs(7760) <= a or b;
    layer0_outputs(7761) <= not a;
    layer0_outputs(7762) <= not a or b;
    layer0_outputs(7763) <= b;
    layer0_outputs(7764) <= b and not a;
    layer0_outputs(7765) <= not (a or b);
    layer0_outputs(7766) <= not a or b;
    layer0_outputs(7767) <= '1';
    layer0_outputs(7768) <= '1';
    layer0_outputs(7769) <= b and not a;
    layer0_outputs(7770) <= not b or a;
    layer0_outputs(7771) <= not a;
    layer0_outputs(7772) <= a xor b;
    layer0_outputs(7773) <= '1';
    layer0_outputs(7774) <= '0';
    layer0_outputs(7775) <= a xor b;
    layer0_outputs(7776) <= b and not a;
    layer0_outputs(7777) <= a xor b;
    layer0_outputs(7778) <= not b;
    layer0_outputs(7779) <= a;
    layer0_outputs(7780) <= a or b;
    layer0_outputs(7781) <= a and not b;
    layer0_outputs(7782) <= not (a or b);
    layer0_outputs(7783) <= not (a and b);
    layer0_outputs(7784) <= b;
    layer0_outputs(7785) <= '0';
    layer0_outputs(7786) <= not a;
    layer0_outputs(7787) <= not b;
    layer0_outputs(7788) <= not b or a;
    layer0_outputs(7789) <= not (a xor b);
    layer0_outputs(7790) <= '1';
    layer0_outputs(7791) <= a and b;
    layer0_outputs(7792) <= '0';
    layer0_outputs(7793) <= a and not b;
    layer0_outputs(7794) <= not (a and b);
    layer0_outputs(7795) <= not a;
    layer0_outputs(7796) <= not b;
    layer0_outputs(7797) <= not b;
    layer0_outputs(7798) <= not (a or b);
    layer0_outputs(7799) <= a xor b;
    layer0_outputs(7800) <= b and not a;
    layer0_outputs(7801) <= not (a or b);
    layer0_outputs(7802) <= a or b;
    layer0_outputs(7803) <= not (a xor b);
    layer0_outputs(7804) <= '1';
    layer0_outputs(7805) <= '0';
    layer0_outputs(7806) <= not (a or b);
    layer0_outputs(7807) <= a and b;
    layer0_outputs(7808) <= a xor b;
    layer0_outputs(7809) <= a;
    layer0_outputs(7810) <= '1';
    layer0_outputs(7811) <= a and b;
    layer0_outputs(7812) <= b and not a;
    layer0_outputs(7813) <= b and not a;
    layer0_outputs(7814) <= '0';
    layer0_outputs(7815) <= '0';
    layer0_outputs(7816) <= not (a or b);
    layer0_outputs(7817) <= a and not b;
    layer0_outputs(7818) <= a xor b;
    layer0_outputs(7819) <= not (a and b);
    layer0_outputs(7820) <= a and not b;
    layer0_outputs(7821) <= a xor b;
    layer0_outputs(7822) <= a;
    layer0_outputs(7823) <= a and b;
    layer0_outputs(7824) <= not (a and b);
    layer0_outputs(7825) <= not (a xor b);
    layer0_outputs(7826) <= b;
    layer0_outputs(7827) <= b;
    layer0_outputs(7828) <= not b;
    layer0_outputs(7829) <= not a;
    layer0_outputs(7830) <= not (a and b);
    layer0_outputs(7831) <= a;
    layer0_outputs(7832) <= not a or b;
    layer0_outputs(7833) <= not b or a;
    layer0_outputs(7834) <= not a;
    layer0_outputs(7835) <= b;
    layer0_outputs(7836) <= not (a xor b);
    layer0_outputs(7837) <= not b or a;
    layer0_outputs(7838) <= a and b;
    layer0_outputs(7839) <= not a;
    layer0_outputs(7840) <= not (a or b);
    layer0_outputs(7841) <= a;
    layer0_outputs(7842) <= not a or b;
    layer0_outputs(7843) <= a;
    layer0_outputs(7844) <= a and not b;
    layer0_outputs(7845) <= not a or b;
    layer0_outputs(7846) <= b;
    layer0_outputs(7847) <= '1';
    layer0_outputs(7848) <= not (a or b);
    layer0_outputs(7849) <= a;
    layer0_outputs(7850) <= b;
    layer0_outputs(7851) <= not b;
    layer0_outputs(7852) <= not b or a;
    layer0_outputs(7853) <= not b or a;
    layer0_outputs(7854) <= not a;
    layer0_outputs(7855) <= a;
    layer0_outputs(7856) <= '1';
    layer0_outputs(7857) <= b;
    layer0_outputs(7858) <= '1';
    layer0_outputs(7859) <= a and not b;
    layer0_outputs(7860) <= a or b;
    layer0_outputs(7861) <= not (a and b);
    layer0_outputs(7862) <= b and not a;
    layer0_outputs(7863) <= not a or b;
    layer0_outputs(7864) <= not (a or b);
    layer0_outputs(7865) <= a;
    layer0_outputs(7866) <= '1';
    layer0_outputs(7867) <= not (a or b);
    layer0_outputs(7868) <= not (a xor b);
    layer0_outputs(7869) <= not b;
    layer0_outputs(7870) <= a or b;
    layer0_outputs(7871) <= '1';
    layer0_outputs(7872) <= not (a or b);
    layer0_outputs(7873) <= not (a xor b);
    layer0_outputs(7874) <= b;
    layer0_outputs(7875) <= not (a or b);
    layer0_outputs(7876) <= not a or b;
    layer0_outputs(7877) <= a and b;
    layer0_outputs(7878) <= not a;
    layer0_outputs(7879) <= '0';
    layer0_outputs(7880) <= a and not b;
    layer0_outputs(7881) <= a and b;
    layer0_outputs(7882) <= not (a xor b);
    layer0_outputs(7883) <= a;
    layer0_outputs(7884) <= a or b;
    layer0_outputs(7885) <= a and b;
    layer0_outputs(7886) <= a or b;
    layer0_outputs(7887) <= a or b;
    layer0_outputs(7888) <= '1';
    layer0_outputs(7889) <= '1';
    layer0_outputs(7890) <= a;
    layer0_outputs(7891) <= not b;
    layer0_outputs(7892) <= a xor b;
    layer0_outputs(7893) <= b;
    layer0_outputs(7894) <= a;
    layer0_outputs(7895) <= a;
    layer0_outputs(7896) <= a;
    layer0_outputs(7897) <= not a or b;
    layer0_outputs(7898) <= not (a xor b);
    layer0_outputs(7899) <= a;
    layer0_outputs(7900) <= not a;
    layer0_outputs(7901) <= not (a or b);
    layer0_outputs(7902) <= a and not b;
    layer0_outputs(7903) <= not (a xor b);
    layer0_outputs(7904) <= '1';
    layer0_outputs(7905) <= b and not a;
    layer0_outputs(7906) <= a;
    layer0_outputs(7907) <= not (a or b);
    layer0_outputs(7908) <= not b;
    layer0_outputs(7909) <= b and not a;
    layer0_outputs(7910) <= a or b;
    layer0_outputs(7911) <= not (a or b);
    layer0_outputs(7912) <= '1';
    layer0_outputs(7913) <= a or b;
    layer0_outputs(7914) <= not a;
    layer0_outputs(7915) <= b and not a;
    layer0_outputs(7916) <= a or b;
    layer0_outputs(7917) <= b and not a;
    layer0_outputs(7918) <= a xor b;
    layer0_outputs(7919) <= not (a xor b);
    layer0_outputs(7920) <= b;
    layer0_outputs(7921) <= b;
    layer0_outputs(7922) <= not (a and b);
    layer0_outputs(7923) <= a and not b;
    layer0_outputs(7924) <= a or b;
    layer0_outputs(7925) <= a and not b;
    layer0_outputs(7926) <= '0';
    layer0_outputs(7927) <= not (a or b);
    layer0_outputs(7928) <= a or b;
    layer0_outputs(7929) <= a and b;
    layer0_outputs(7930) <= not (a and b);
    layer0_outputs(7931) <= a;
    layer0_outputs(7932) <= not (a or b);
    layer0_outputs(7933) <= a or b;
    layer0_outputs(7934) <= a and not b;
    layer0_outputs(7935) <= not a;
    layer0_outputs(7936) <= a or b;
    layer0_outputs(7937) <= a and not b;
    layer0_outputs(7938) <= not (a xor b);
    layer0_outputs(7939) <= not (a or b);
    layer0_outputs(7940) <= b and not a;
    layer0_outputs(7941) <= a and not b;
    layer0_outputs(7942) <= not a;
    layer0_outputs(7943) <= not (a and b);
    layer0_outputs(7944) <= a or b;
    layer0_outputs(7945) <= b;
    layer0_outputs(7946) <= not (a xor b);
    layer0_outputs(7947) <= not (a xor b);
    layer0_outputs(7948) <= a or b;
    layer0_outputs(7949) <= b and not a;
    layer0_outputs(7950) <= not (a or b);
    layer0_outputs(7951) <= a and b;
    layer0_outputs(7952) <= a;
    layer0_outputs(7953) <= not a or b;
    layer0_outputs(7954) <= not b;
    layer0_outputs(7955) <= not (a and b);
    layer0_outputs(7956) <= a xor b;
    layer0_outputs(7957) <= not a or b;
    layer0_outputs(7958) <= a and not b;
    layer0_outputs(7959) <= not (a xor b);
    layer0_outputs(7960) <= a;
    layer0_outputs(7961) <= not a;
    layer0_outputs(7962) <= not b;
    layer0_outputs(7963) <= a or b;
    layer0_outputs(7964) <= a xor b;
    layer0_outputs(7965) <= not (a or b);
    layer0_outputs(7966) <= a xor b;
    layer0_outputs(7967) <= '1';
    layer0_outputs(7968) <= a;
    layer0_outputs(7969) <= a xor b;
    layer0_outputs(7970) <= a and b;
    layer0_outputs(7971) <= a xor b;
    layer0_outputs(7972) <= a;
    layer0_outputs(7973) <= a or b;
    layer0_outputs(7974) <= not a or b;
    layer0_outputs(7975) <= not (a or b);
    layer0_outputs(7976) <= '1';
    layer0_outputs(7977) <= '1';
    layer0_outputs(7978) <= a xor b;
    layer0_outputs(7979) <= not a or b;
    layer0_outputs(7980) <= b;
    layer0_outputs(7981) <= '1';
    layer0_outputs(7982) <= a;
    layer0_outputs(7983) <= a;
    layer0_outputs(7984) <= not a;
    layer0_outputs(7985) <= not a;
    layer0_outputs(7986) <= not b or a;
    layer0_outputs(7987) <= '0';
    layer0_outputs(7988) <= a and not b;
    layer0_outputs(7989) <= not (a xor b);
    layer0_outputs(7990) <= not (a or b);
    layer0_outputs(7991) <= not (a xor b);
    layer0_outputs(7992) <= a xor b;
    layer0_outputs(7993) <= not (a xor b);
    layer0_outputs(7994) <= not a;
    layer0_outputs(7995) <= b;
    layer0_outputs(7996) <= not (a xor b);
    layer0_outputs(7997) <= a xor b;
    layer0_outputs(7998) <= b;
    layer0_outputs(7999) <= a or b;
    layer0_outputs(8000) <= not (a or b);
    layer0_outputs(8001) <= b and not a;
    layer0_outputs(8002) <= a;
    layer0_outputs(8003) <= b and not a;
    layer0_outputs(8004) <= a;
    layer0_outputs(8005) <= not b or a;
    layer0_outputs(8006) <= b;
    layer0_outputs(8007) <= a;
    layer0_outputs(8008) <= a xor b;
    layer0_outputs(8009) <= not (a xor b);
    layer0_outputs(8010) <= a or b;
    layer0_outputs(8011) <= not (a xor b);
    layer0_outputs(8012) <= not b or a;
    layer0_outputs(8013) <= a xor b;
    layer0_outputs(8014) <= not (a or b);
    layer0_outputs(8015) <= not a or b;
    layer0_outputs(8016) <= not (a xor b);
    layer0_outputs(8017) <= a;
    layer0_outputs(8018) <= not a or b;
    layer0_outputs(8019) <= not (a xor b);
    layer0_outputs(8020) <= not a;
    layer0_outputs(8021) <= b and not a;
    layer0_outputs(8022) <= not (a and b);
    layer0_outputs(8023) <= not (a or b);
    layer0_outputs(8024) <= not b or a;
    layer0_outputs(8025) <= '1';
    layer0_outputs(8026) <= a or b;
    layer0_outputs(8027) <= a;
    layer0_outputs(8028) <= a or b;
    layer0_outputs(8029) <= a;
    layer0_outputs(8030) <= a xor b;
    layer0_outputs(8031) <= not a;
    layer0_outputs(8032) <= not (a or b);
    layer0_outputs(8033) <= not a;
    layer0_outputs(8034) <= not a;
    layer0_outputs(8035) <= not a or b;
    layer0_outputs(8036) <= not (a xor b);
    layer0_outputs(8037) <= a and b;
    layer0_outputs(8038) <= not (a xor b);
    layer0_outputs(8039) <= not (a or b);
    layer0_outputs(8040) <= b;
    layer0_outputs(8041) <= not (a xor b);
    layer0_outputs(8042) <= not (a and b);
    layer0_outputs(8043) <= not (a xor b);
    layer0_outputs(8044) <= not (a or b);
    layer0_outputs(8045) <= not (a or b);
    layer0_outputs(8046) <= a;
    layer0_outputs(8047) <= a xor b;
    layer0_outputs(8048) <= a and not b;
    layer0_outputs(8049) <= b and not a;
    layer0_outputs(8050) <= not b;
    layer0_outputs(8051) <= a or b;
    layer0_outputs(8052) <= not (a or b);
    layer0_outputs(8053) <= '1';
    layer0_outputs(8054) <= not a;
    layer0_outputs(8055) <= a or b;
    layer0_outputs(8056) <= a xor b;
    layer0_outputs(8057) <= not (a and b);
    layer0_outputs(8058) <= not a;
    layer0_outputs(8059) <= b and not a;
    layer0_outputs(8060) <= not a;
    layer0_outputs(8061) <= not b;
    layer0_outputs(8062) <= a and not b;
    layer0_outputs(8063) <= not b or a;
    layer0_outputs(8064) <= not b;
    layer0_outputs(8065) <= not a;
    layer0_outputs(8066) <= a;
    layer0_outputs(8067) <= '1';
    layer0_outputs(8068) <= a and b;
    layer0_outputs(8069) <= not b or a;
    layer0_outputs(8070) <= not (a xor b);
    layer0_outputs(8071) <= not (a or b);
    layer0_outputs(8072) <= a or b;
    layer0_outputs(8073) <= not (a or b);
    layer0_outputs(8074) <= a and b;
    layer0_outputs(8075) <= a;
    layer0_outputs(8076) <= not (a and b);
    layer0_outputs(8077) <= a;
    layer0_outputs(8078) <= not b;
    layer0_outputs(8079) <= b;
    layer0_outputs(8080) <= not (a or b);
    layer0_outputs(8081) <= b and not a;
    layer0_outputs(8082) <= b;
    layer0_outputs(8083) <= a and b;
    layer0_outputs(8084) <= not (a xor b);
    layer0_outputs(8085) <= not (a and b);
    layer0_outputs(8086) <= a;
    layer0_outputs(8087) <= a or b;
    layer0_outputs(8088) <= not (a and b);
    layer0_outputs(8089) <= b and not a;
    layer0_outputs(8090) <= not a or b;
    layer0_outputs(8091) <= not (a or b);
    layer0_outputs(8092) <= b;
    layer0_outputs(8093) <= not (a xor b);
    layer0_outputs(8094) <= a or b;
    layer0_outputs(8095) <= a and not b;
    layer0_outputs(8096) <= not b;
    layer0_outputs(8097) <= not (a or b);
    layer0_outputs(8098) <= a or b;
    layer0_outputs(8099) <= a;
    layer0_outputs(8100) <= a or b;
    layer0_outputs(8101) <= b and not a;
    layer0_outputs(8102) <= not b;
    layer0_outputs(8103) <= not a;
    layer0_outputs(8104) <= b and not a;
    layer0_outputs(8105) <= not a or b;
    layer0_outputs(8106) <= not a;
    layer0_outputs(8107) <= not b;
    layer0_outputs(8108) <= a and not b;
    layer0_outputs(8109) <= not (a or b);
    layer0_outputs(8110) <= a and not b;
    layer0_outputs(8111) <= not (a or b);
    layer0_outputs(8112) <= not (a and b);
    layer0_outputs(8113) <= not (a or b);
    layer0_outputs(8114) <= not a;
    layer0_outputs(8115) <= not (a or b);
    layer0_outputs(8116) <= b;
    layer0_outputs(8117) <= a and b;
    layer0_outputs(8118) <= a xor b;
    layer0_outputs(8119) <= a;
    layer0_outputs(8120) <= not b;
    layer0_outputs(8121) <= not (a xor b);
    layer0_outputs(8122) <= not (a xor b);
    layer0_outputs(8123) <= not (a or b);
    layer0_outputs(8124) <= b;
    layer0_outputs(8125) <= not a or b;
    layer0_outputs(8126) <= not (a or b);
    layer0_outputs(8127) <= not a or b;
    layer0_outputs(8128) <= a and not b;
    layer0_outputs(8129) <= a;
    layer0_outputs(8130) <= a or b;
    layer0_outputs(8131) <= not b or a;
    layer0_outputs(8132) <= not (a xor b);
    layer0_outputs(8133) <= '1';
    layer0_outputs(8134) <= not (a and b);
    layer0_outputs(8135) <= not a;
    layer0_outputs(8136) <= b and not a;
    layer0_outputs(8137) <= b and not a;
    layer0_outputs(8138) <= a and not b;
    layer0_outputs(8139) <= a and b;
    layer0_outputs(8140) <= not a;
    layer0_outputs(8141) <= a and not b;
    layer0_outputs(8142) <= not b or a;
    layer0_outputs(8143) <= not (a or b);
    layer0_outputs(8144) <= not b;
    layer0_outputs(8145) <= not b or a;
    layer0_outputs(8146) <= not a;
    layer0_outputs(8147) <= a;
    layer0_outputs(8148) <= a and b;
    layer0_outputs(8149) <= '0';
    layer0_outputs(8150) <= '0';
    layer0_outputs(8151) <= a and not b;
    layer0_outputs(8152) <= '1';
    layer0_outputs(8153) <= b;
    layer0_outputs(8154) <= not a;
    layer0_outputs(8155) <= not a or b;
    layer0_outputs(8156) <= a and not b;
    layer0_outputs(8157) <= not b or a;
    layer0_outputs(8158) <= '0';
    layer0_outputs(8159) <= a;
    layer0_outputs(8160) <= b and not a;
    layer0_outputs(8161) <= a and b;
    layer0_outputs(8162) <= b and not a;
    layer0_outputs(8163) <= not (a or b);
    layer0_outputs(8164) <= not b;
    layer0_outputs(8165) <= b and not a;
    layer0_outputs(8166) <= not (a xor b);
    layer0_outputs(8167) <= not b or a;
    layer0_outputs(8168) <= a and b;
    layer0_outputs(8169) <= not a;
    layer0_outputs(8170) <= a and not b;
    layer0_outputs(8171) <= not (a xor b);
    layer0_outputs(8172) <= not b;
    layer0_outputs(8173) <= a or b;
    layer0_outputs(8174) <= not (a or b);
    layer0_outputs(8175) <= '0';
    layer0_outputs(8176) <= not a;
    layer0_outputs(8177) <= a;
    layer0_outputs(8178) <= not a;
    layer0_outputs(8179) <= not (a or b);
    layer0_outputs(8180) <= not (a or b);
    layer0_outputs(8181) <= not (a or b);
    layer0_outputs(8182) <= '1';
    layer0_outputs(8183) <= not a;
    layer0_outputs(8184) <= b;
    layer0_outputs(8185) <= '0';
    layer0_outputs(8186) <= a;
    layer0_outputs(8187) <= a;
    layer0_outputs(8188) <= a xor b;
    layer0_outputs(8189) <= not a;
    layer0_outputs(8190) <= not a;
    layer0_outputs(8191) <= not b;
    layer0_outputs(8192) <= '1';
    layer0_outputs(8193) <= b;
    layer0_outputs(8194) <= not b or a;
    layer0_outputs(8195) <= a or b;
    layer0_outputs(8196) <= not b or a;
    layer0_outputs(8197) <= b and not a;
    layer0_outputs(8198) <= not (a or b);
    layer0_outputs(8199) <= not a or b;
    layer0_outputs(8200) <= '0';
    layer0_outputs(8201) <= not (a or b);
    layer0_outputs(8202) <= '0';
    layer0_outputs(8203) <= not b;
    layer0_outputs(8204) <= not b or a;
    layer0_outputs(8205) <= not (a and b);
    layer0_outputs(8206) <= a xor b;
    layer0_outputs(8207) <= a xor b;
    layer0_outputs(8208) <= a or b;
    layer0_outputs(8209) <= not (a xor b);
    layer0_outputs(8210) <= not b or a;
    layer0_outputs(8211) <= '1';
    layer0_outputs(8212) <= '1';
    layer0_outputs(8213) <= not a;
    layer0_outputs(8214) <= b;
    layer0_outputs(8215) <= b;
    layer0_outputs(8216) <= a xor b;
    layer0_outputs(8217) <= a xor b;
    layer0_outputs(8218) <= a;
    layer0_outputs(8219) <= a or b;
    layer0_outputs(8220) <= a or b;
    layer0_outputs(8221) <= a or b;
    layer0_outputs(8222) <= not a;
    layer0_outputs(8223) <= a;
    layer0_outputs(8224) <= not b or a;
    layer0_outputs(8225) <= a and not b;
    layer0_outputs(8226) <= not (a xor b);
    layer0_outputs(8227) <= not (a or b);
    layer0_outputs(8228) <= not a;
    layer0_outputs(8229) <= not (a xor b);
    layer0_outputs(8230) <= b;
    layer0_outputs(8231) <= not a;
    layer0_outputs(8232) <= not b;
    layer0_outputs(8233) <= not (a or b);
    layer0_outputs(8234) <= not (a and b);
    layer0_outputs(8235) <= '0';
    layer0_outputs(8236) <= a and b;
    layer0_outputs(8237) <= not a;
    layer0_outputs(8238) <= b;
    layer0_outputs(8239) <= not a or b;
    layer0_outputs(8240) <= not b or a;
    layer0_outputs(8241) <= not (a and b);
    layer0_outputs(8242) <= not (a xor b);
    layer0_outputs(8243) <= not b or a;
    layer0_outputs(8244) <= a or b;
    layer0_outputs(8245) <= not a or b;
    layer0_outputs(8246) <= not (a or b);
    layer0_outputs(8247) <= not b or a;
    layer0_outputs(8248) <= not a;
    layer0_outputs(8249) <= b;
    layer0_outputs(8250) <= b;
    layer0_outputs(8251) <= a xor b;
    layer0_outputs(8252) <= a or b;
    layer0_outputs(8253) <= not a;
    layer0_outputs(8254) <= '1';
    layer0_outputs(8255) <= not a;
    layer0_outputs(8256) <= a or b;
    layer0_outputs(8257) <= not (a and b);
    layer0_outputs(8258) <= a xor b;
    layer0_outputs(8259) <= a and b;
    layer0_outputs(8260) <= b and not a;
    layer0_outputs(8261) <= a or b;
    layer0_outputs(8262) <= b and not a;
    layer0_outputs(8263) <= not a or b;
    layer0_outputs(8264) <= a or b;
    layer0_outputs(8265) <= not (a or b);
    layer0_outputs(8266) <= a xor b;
    layer0_outputs(8267) <= not a;
    layer0_outputs(8268) <= b and not a;
    layer0_outputs(8269) <= a and b;
    layer0_outputs(8270) <= not (a or b);
    layer0_outputs(8271) <= b and not a;
    layer0_outputs(8272) <= not (a and b);
    layer0_outputs(8273) <= not b or a;
    layer0_outputs(8274) <= a and not b;
    layer0_outputs(8275) <= not (a xor b);
    layer0_outputs(8276) <= a and b;
    layer0_outputs(8277) <= not (a or b);
    layer0_outputs(8278) <= a or b;
    layer0_outputs(8279) <= not a;
    layer0_outputs(8280) <= a xor b;
    layer0_outputs(8281) <= not b;
    layer0_outputs(8282) <= not a or b;
    layer0_outputs(8283) <= not b or a;
    layer0_outputs(8284) <= a and not b;
    layer0_outputs(8285) <= not (a or b);
    layer0_outputs(8286) <= not a;
    layer0_outputs(8287) <= not a;
    layer0_outputs(8288) <= a xor b;
    layer0_outputs(8289) <= a or b;
    layer0_outputs(8290) <= a and not b;
    layer0_outputs(8291) <= '0';
    layer0_outputs(8292) <= a and not b;
    layer0_outputs(8293) <= '1';
    layer0_outputs(8294) <= '1';
    layer0_outputs(8295) <= a xor b;
    layer0_outputs(8296) <= not a or b;
    layer0_outputs(8297) <= a and b;
    layer0_outputs(8298) <= a xor b;
    layer0_outputs(8299) <= a;
    layer0_outputs(8300) <= a and b;
    layer0_outputs(8301) <= b and not a;
    layer0_outputs(8302) <= a and not b;
    layer0_outputs(8303) <= not (a xor b);
    layer0_outputs(8304) <= a and not b;
    layer0_outputs(8305) <= a and b;
    layer0_outputs(8306) <= not a or b;
    layer0_outputs(8307) <= b;
    layer0_outputs(8308) <= not b;
    layer0_outputs(8309) <= not b or a;
    layer0_outputs(8310) <= not b;
    layer0_outputs(8311) <= not a or b;
    layer0_outputs(8312) <= '1';
    layer0_outputs(8313) <= b and not a;
    layer0_outputs(8314) <= b;
    layer0_outputs(8315) <= a and not b;
    layer0_outputs(8316) <= a and b;
    layer0_outputs(8317) <= not (a or b);
    layer0_outputs(8318) <= a and not b;
    layer0_outputs(8319) <= b and not a;
    layer0_outputs(8320) <= a and b;
    layer0_outputs(8321) <= not (a and b);
    layer0_outputs(8322) <= b and not a;
    layer0_outputs(8323) <= not b or a;
    layer0_outputs(8324) <= not a;
    layer0_outputs(8325) <= not a;
    layer0_outputs(8326) <= not b or a;
    layer0_outputs(8327) <= not b;
    layer0_outputs(8328) <= not a;
    layer0_outputs(8329) <= '0';
    layer0_outputs(8330) <= not a or b;
    layer0_outputs(8331) <= b;
    layer0_outputs(8332) <= a or b;
    layer0_outputs(8333) <= not a or b;
    layer0_outputs(8334) <= not a;
    layer0_outputs(8335) <= b;
    layer0_outputs(8336) <= a and not b;
    layer0_outputs(8337) <= a xor b;
    layer0_outputs(8338) <= not (a xor b);
    layer0_outputs(8339) <= not b or a;
    layer0_outputs(8340) <= not (a xor b);
    layer0_outputs(8341) <= not (a xor b);
    layer0_outputs(8342) <= a and b;
    layer0_outputs(8343) <= not (a xor b);
    layer0_outputs(8344) <= not (a xor b);
    layer0_outputs(8345) <= a or b;
    layer0_outputs(8346) <= not a or b;
    layer0_outputs(8347) <= not a or b;
    layer0_outputs(8348) <= b and not a;
    layer0_outputs(8349) <= not (a xor b);
    layer0_outputs(8350) <= a and not b;
    layer0_outputs(8351) <= not b;
    layer0_outputs(8352) <= b;
    layer0_outputs(8353) <= not b;
    layer0_outputs(8354) <= not (a or b);
    layer0_outputs(8355) <= not b;
    layer0_outputs(8356) <= b and not a;
    layer0_outputs(8357) <= a and not b;
    layer0_outputs(8358) <= a;
    layer0_outputs(8359) <= b;
    layer0_outputs(8360) <= a xor b;
    layer0_outputs(8361) <= a;
    layer0_outputs(8362) <= not (a or b);
    layer0_outputs(8363) <= not a or b;
    layer0_outputs(8364) <= '0';
    layer0_outputs(8365) <= '1';
    layer0_outputs(8366) <= a or b;
    layer0_outputs(8367) <= a;
    layer0_outputs(8368) <= '1';
    layer0_outputs(8369) <= not a or b;
    layer0_outputs(8370) <= not (a xor b);
    layer0_outputs(8371) <= not (a and b);
    layer0_outputs(8372) <= '0';
    layer0_outputs(8373) <= not (a and b);
    layer0_outputs(8374) <= a and b;
    layer0_outputs(8375) <= not (a xor b);
    layer0_outputs(8376) <= not a;
    layer0_outputs(8377) <= '0';
    layer0_outputs(8378) <= '1';
    layer0_outputs(8379) <= a xor b;
    layer0_outputs(8380) <= not (a or b);
    layer0_outputs(8381) <= b and not a;
    layer0_outputs(8382) <= '1';
    layer0_outputs(8383) <= not b or a;
    layer0_outputs(8384) <= b;
    layer0_outputs(8385) <= not b or a;
    layer0_outputs(8386) <= not a;
    layer0_outputs(8387) <= a and b;
    layer0_outputs(8388) <= a and not b;
    layer0_outputs(8389) <= '0';
    layer0_outputs(8390) <= a and b;
    layer0_outputs(8391) <= not b;
    layer0_outputs(8392) <= not (a and b);
    layer0_outputs(8393) <= not b;
    layer0_outputs(8394) <= '1';
    layer0_outputs(8395) <= a xor b;
    layer0_outputs(8396) <= '0';
    layer0_outputs(8397) <= '0';
    layer0_outputs(8398) <= b and not a;
    layer0_outputs(8399) <= not (a xor b);
    layer0_outputs(8400) <= not b;
    layer0_outputs(8401) <= not b;
    layer0_outputs(8402) <= not a or b;
    layer0_outputs(8403) <= a or b;
    layer0_outputs(8404) <= a and not b;
    layer0_outputs(8405) <= not b or a;
    layer0_outputs(8406) <= a and b;
    layer0_outputs(8407) <= not (a or b);
    layer0_outputs(8408) <= not (a or b);
    layer0_outputs(8409) <= not b;
    layer0_outputs(8410) <= not b or a;
    layer0_outputs(8411) <= a xor b;
    layer0_outputs(8412) <= b and not a;
    layer0_outputs(8413) <= a;
    layer0_outputs(8414) <= a;
    layer0_outputs(8415) <= a;
    layer0_outputs(8416) <= not b or a;
    layer0_outputs(8417) <= b;
    layer0_outputs(8418) <= b and not a;
    layer0_outputs(8419) <= a and b;
    layer0_outputs(8420) <= not a or b;
    layer0_outputs(8421) <= not a or b;
    layer0_outputs(8422) <= '0';
    layer0_outputs(8423) <= not a or b;
    layer0_outputs(8424) <= not b or a;
    layer0_outputs(8425) <= not (a and b);
    layer0_outputs(8426) <= a or b;
    layer0_outputs(8427) <= not a or b;
    layer0_outputs(8428) <= a and not b;
    layer0_outputs(8429) <= not a;
    layer0_outputs(8430) <= not (a xor b);
    layer0_outputs(8431) <= not b;
    layer0_outputs(8432) <= not a;
    layer0_outputs(8433) <= not a or b;
    layer0_outputs(8434) <= a and not b;
    layer0_outputs(8435) <= a;
    layer0_outputs(8436) <= not b;
    layer0_outputs(8437) <= a xor b;
    layer0_outputs(8438) <= a or b;
    layer0_outputs(8439) <= b;
    layer0_outputs(8440) <= not b;
    layer0_outputs(8441) <= b and not a;
    layer0_outputs(8442) <= a;
    layer0_outputs(8443) <= a or b;
    layer0_outputs(8444) <= a or b;
    layer0_outputs(8445) <= not (a or b);
    layer0_outputs(8446) <= not b or a;
    layer0_outputs(8447) <= a xor b;
    layer0_outputs(8448) <= not (a or b);
    layer0_outputs(8449) <= not (a or b);
    layer0_outputs(8450) <= not (a xor b);
    layer0_outputs(8451) <= '0';
    layer0_outputs(8452) <= b;
    layer0_outputs(8453) <= not (a or b);
    layer0_outputs(8454) <= not b;
    layer0_outputs(8455) <= a;
    layer0_outputs(8456) <= not a;
    layer0_outputs(8457) <= not a or b;
    layer0_outputs(8458) <= not b or a;
    layer0_outputs(8459) <= b;
    layer0_outputs(8460) <= b;
    layer0_outputs(8461) <= a and b;
    layer0_outputs(8462) <= a;
    layer0_outputs(8463) <= '0';
    layer0_outputs(8464) <= '0';
    layer0_outputs(8465) <= a xor b;
    layer0_outputs(8466) <= '0';
    layer0_outputs(8467) <= not (a xor b);
    layer0_outputs(8468) <= not a or b;
    layer0_outputs(8469) <= '1';
    layer0_outputs(8470) <= a;
    layer0_outputs(8471) <= not (a and b);
    layer0_outputs(8472) <= b and not a;
    layer0_outputs(8473) <= a or b;
    layer0_outputs(8474) <= not (a or b);
    layer0_outputs(8475) <= '1';
    layer0_outputs(8476) <= not a or b;
    layer0_outputs(8477) <= a or b;
    layer0_outputs(8478) <= not (a and b);
    layer0_outputs(8479) <= a xor b;
    layer0_outputs(8480) <= not b;
    layer0_outputs(8481) <= not (a xor b);
    layer0_outputs(8482) <= a;
    layer0_outputs(8483) <= not a or b;
    layer0_outputs(8484) <= not a or b;
    layer0_outputs(8485) <= not b;
    layer0_outputs(8486) <= a or b;
    layer0_outputs(8487) <= a;
    layer0_outputs(8488) <= b and not a;
    layer0_outputs(8489) <= '0';
    layer0_outputs(8490) <= a or b;
    layer0_outputs(8491) <= a or b;
    layer0_outputs(8492) <= a or b;
    layer0_outputs(8493) <= a;
    layer0_outputs(8494) <= not b or a;
    layer0_outputs(8495) <= not a;
    layer0_outputs(8496) <= a and b;
    layer0_outputs(8497) <= not b;
    layer0_outputs(8498) <= '1';
    layer0_outputs(8499) <= not a;
    layer0_outputs(8500) <= not (a or b);
    layer0_outputs(8501) <= a or b;
    layer0_outputs(8502) <= b;
    layer0_outputs(8503) <= not (a and b);
    layer0_outputs(8504) <= not b;
    layer0_outputs(8505) <= not (a or b);
    layer0_outputs(8506) <= not (a or b);
    layer0_outputs(8507) <= a or b;
    layer0_outputs(8508) <= not b;
    layer0_outputs(8509) <= a and not b;
    layer0_outputs(8510) <= b;
    layer0_outputs(8511) <= not a;
    layer0_outputs(8512) <= a;
    layer0_outputs(8513) <= a xor b;
    layer0_outputs(8514) <= a and b;
    layer0_outputs(8515) <= b and not a;
    layer0_outputs(8516) <= a and not b;
    layer0_outputs(8517) <= a;
    layer0_outputs(8518) <= '1';
    layer0_outputs(8519) <= not b or a;
    layer0_outputs(8520) <= b and not a;
    layer0_outputs(8521) <= not b or a;
    layer0_outputs(8522) <= not a or b;
    layer0_outputs(8523) <= a and b;
    layer0_outputs(8524) <= not (a xor b);
    layer0_outputs(8525) <= b;
    layer0_outputs(8526) <= b and not a;
    layer0_outputs(8527) <= a;
    layer0_outputs(8528) <= b;
    layer0_outputs(8529) <= b;
    layer0_outputs(8530) <= not (a or b);
    layer0_outputs(8531) <= not (a and b);
    layer0_outputs(8532) <= a;
    layer0_outputs(8533) <= not (a xor b);
    layer0_outputs(8534) <= b and not a;
    layer0_outputs(8535) <= a xor b;
    layer0_outputs(8536) <= a;
    layer0_outputs(8537) <= not (a and b);
    layer0_outputs(8538) <= b and not a;
    layer0_outputs(8539) <= not (a or b);
    layer0_outputs(8540) <= '0';
    layer0_outputs(8541) <= a xor b;
    layer0_outputs(8542) <= not (a and b);
    layer0_outputs(8543) <= not b;
    layer0_outputs(8544) <= a and b;
    layer0_outputs(8545) <= a and b;
    layer0_outputs(8546) <= not (a and b);
    layer0_outputs(8547) <= not a or b;
    layer0_outputs(8548) <= a xor b;
    layer0_outputs(8549) <= b and not a;
    layer0_outputs(8550) <= not (a or b);
    layer0_outputs(8551) <= b;
    layer0_outputs(8552) <= b;
    layer0_outputs(8553) <= a and b;
    layer0_outputs(8554) <= not (a xor b);
    layer0_outputs(8555) <= a xor b;
    layer0_outputs(8556) <= b;
    layer0_outputs(8557) <= '0';
    layer0_outputs(8558) <= a or b;
    layer0_outputs(8559) <= not b or a;
    layer0_outputs(8560) <= not b;
    layer0_outputs(8561) <= not (a or b);
    layer0_outputs(8562) <= a and not b;
    layer0_outputs(8563) <= a xor b;
    layer0_outputs(8564) <= '1';
    layer0_outputs(8565) <= not (a xor b);
    layer0_outputs(8566) <= not b or a;
    layer0_outputs(8567) <= not (a or b);
    layer0_outputs(8568) <= a;
    layer0_outputs(8569) <= not b;
    layer0_outputs(8570) <= not a or b;
    layer0_outputs(8571) <= not b or a;
    layer0_outputs(8572) <= not a;
    layer0_outputs(8573) <= not a;
    layer0_outputs(8574) <= a;
    layer0_outputs(8575) <= '1';
    layer0_outputs(8576) <= a xor b;
    layer0_outputs(8577) <= a xor b;
    layer0_outputs(8578) <= a xor b;
    layer0_outputs(8579) <= a or b;
    layer0_outputs(8580) <= '0';
    layer0_outputs(8581) <= a or b;
    layer0_outputs(8582) <= not a or b;
    layer0_outputs(8583) <= not (a or b);
    layer0_outputs(8584) <= '1';
    layer0_outputs(8585) <= not b;
    layer0_outputs(8586) <= a or b;
    layer0_outputs(8587) <= b;
    layer0_outputs(8588) <= a xor b;
    layer0_outputs(8589) <= a and b;
    layer0_outputs(8590) <= not (a or b);
    layer0_outputs(8591) <= a or b;
    layer0_outputs(8592) <= not (a and b);
    layer0_outputs(8593) <= not (a or b);
    layer0_outputs(8594) <= not (a and b);
    layer0_outputs(8595) <= '1';
    layer0_outputs(8596) <= not (a xor b);
    layer0_outputs(8597) <= not (a or b);
    layer0_outputs(8598) <= b and not a;
    layer0_outputs(8599) <= b;
    layer0_outputs(8600) <= '0';
    layer0_outputs(8601) <= a;
    layer0_outputs(8602) <= not a or b;
    layer0_outputs(8603) <= not b or a;
    layer0_outputs(8604) <= not a;
    layer0_outputs(8605) <= '0';
    layer0_outputs(8606) <= not a;
    layer0_outputs(8607) <= not (a or b);
    layer0_outputs(8608) <= a;
    layer0_outputs(8609) <= a xor b;
    layer0_outputs(8610) <= not b or a;
    layer0_outputs(8611) <= a or b;
    layer0_outputs(8612) <= not a;
    layer0_outputs(8613) <= not (a or b);
    layer0_outputs(8614) <= '0';
    layer0_outputs(8615) <= b;
    layer0_outputs(8616) <= a and b;
    layer0_outputs(8617) <= '0';
    layer0_outputs(8618) <= not (a or b);
    layer0_outputs(8619) <= '1';
    layer0_outputs(8620) <= '0';
    layer0_outputs(8621) <= a and b;
    layer0_outputs(8622) <= not a or b;
    layer0_outputs(8623) <= '0';
    layer0_outputs(8624) <= not b;
    layer0_outputs(8625) <= not a;
    layer0_outputs(8626) <= not (a or b);
    layer0_outputs(8627) <= a xor b;
    layer0_outputs(8628) <= not a or b;
    layer0_outputs(8629) <= not b or a;
    layer0_outputs(8630) <= a and b;
    layer0_outputs(8631) <= not a or b;
    layer0_outputs(8632) <= a and b;
    layer0_outputs(8633) <= a;
    layer0_outputs(8634) <= a xor b;
    layer0_outputs(8635) <= a or b;
    layer0_outputs(8636) <= b;
    layer0_outputs(8637) <= not b or a;
    layer0_outputs(8638) <= not (a xor b);
    layer0_outputs(8639) <= not (a or b);
    layer0_outputs(8640) <= not a or b;
    layer0_outputs(8641) <= not a;
    layer0_outputs(8642) <= not (a and b);
    layer0_outputs(8643) <= not b;
    layer0_outputs(8644) <= not (a and b);
    layer0_outputs(8645) <= not (a xor b);
    layer0_outputs(8646) <= not a or b;
    layer0_outputs(8647) <= not b;
    layer0_outputs(8648) <= '1';
    layer0_outputs(8649) <= not b;
    layer0_outputs(8650) <= not a or b;
    layer0_outputs(8651) <= b and not a;
    layer0_outputs(8652) <= b;
    layer0_outputs(8653) <= a;
    layer0_outputs(8654) <= '1';
    layer0_outputs(8655) <= not b or a;
    layer0_outputs(8656) <= a;
    layer0_outputs(8657) <= not a or b;
    layer0_outputs(8658) <= b;
    layer0_outputs(8659) <= b;
    layer0_outputs(8660) <= a;
    layer0_outputs(8661) <= a or b;
    layer0_outputs(8662) <= a or b;
    layer0_outputs(8663) <= '0';
    layer0_outputs(8664) <= not b or a;
    layer0_outputs(8665) <= '0';
    layer0_outputs(8666) <= '1';
    layer0_outputs(8667) <= not b;
    layer0_outputs(8668) <= not (a and b);
    layer0_outputs(8669) <= '0';
    layer0_outputs(8670) <= not b or a;
    layer0_outputs(8671) <= not (a xor b);
    layer0_outputs(8672) <= not (a or b);
    layer0_outputs(8673) <= a and b;
    layer0_outputs(8674) <= b;
    layer0_outputs(8675) <= not (a xor b);
    layer0_outputs(8676) <= a xor b;
    layer0_outputs(8677) <= not a;
    layer0_outputs(8678) <= not b or a;
    layer0_outputs(8679) <= '0';
    layer0_outputs(8680) <= a or b;
    layer0_outputs(8681) <= not a;
    layer0_outputs(8682) <= not (a and b);
    layer0_outputs(8683) <= not b or a;
    layer0_outputs(8684) <= a or b;
    layer0_outputs(8685) <= a or b;
    layer0_outputs(8686) <= a or b;
    layer0_outputs(8687) <= not (a and b);
    layer0_outputs(8688) <= not (a xor b);
    layer0_outputs(8689) <= a and not b;
    layer0_outputs(8690) <= not a;
    layer0_outputs(8691) <= not (a or b);
    layer0_outputs(8692) <= a or b;
    layer0_outputs(8693) <= a and not b;
    layer0_outputs(8694) <= '1';
    layer0_outputs(8695) <= a xor b;
    layer0_outputs(8696) <= b and not a;
    layer0_outputs(8697) <= a and not b;
    layer0_outputs(8698) <= '0';
    layer0_outputs(8699) <= not (a or b);
    layer0_outputs(8700) <= b and not a;
    layer0_outputs(8701) <= not (a or b);
    layer0_outputs(8702) <= not a or b;
    layer0_outputs(8703) <= a or b;
    layer0_outputs(8704) <= b and not a;
    layer0_outputs(8705) <= '0';
    layer0_outputs(8706) <= a and b;
    layer0_outputs(8707) <= not (a and b);
    layer0_outputs(8708) <= not a;
    layer0_outputs(8709) <= not b or a;
    layer0_outputs(8710) <= not a;
    layer0_outputs(8711) <= a and b;
    layer0_outputs(8712) <= b and not a;
    layer0_outputs(8713) <= not (a and b);
    layer0_outputs(8714) <= b and not a;
    layer0_outputs(8715) <= a;
    layer0_outputs(8716) <= not a;
    layer0_outputs(8717) <= not (a xor b);
    layer0_outputs(8718) <= not b;
    layer0_outputs(8719) <= a or b;
    layer0_outputs(8720) <= not b;
    layer0_outputs(8721) <= not (a xor b);
    layer0_outputs(8722) <= not (a or b);
    layer0_outputs(8723) <= b;
    layer0_outputs(8724) <= a or b;
    layer0_outputs(8725) <= a xor b;
    layer0_outputs(8726) <= not b or a;
    layer0_outputs(8727) <= not (a or b);
    layer0_outputs(8728) <= not b or a;
    layer0_outputs(8729) <= not b or a;
    layer0_outputs(8730) <= not b;
    layer0_outputs(8731) <= not a;
    layer0_outputs(8732) <= '0';
    layer0_outputs(8733) <= not (a or b);
    layer0_outputs(8734) <= a;
    layer0_outputs(8735) <= not (a or b);
    layer0_outputs(8736) <= not b;
    layer0_outputs(8737) <= not (a or b);
    layer0_outputs(8738) <= a and b;
    layer0_outputs(8739) <= not a;
    layer0_outputs(8740) <= '1';
    layer0_outputs(8741) <= not (a xor b);
    layer0_outputs(8742) <= '1';
    layer0_outputs(8743) <= a and not b;
    layer0_outputs(8744) <= not a;
    layer0_outputs(8745) <= not b;
    layer0_outputs(8746) <= a xor b;
    layer0_outputs(8747) <= not b or a;
    layer0_outputs(8748) <= not a or b;
    layer0_outputs(8749) <= not (a and b);
    layer0_outputs(8750) <= not b or a;
    layer0_outputs(8751) <= not (a or b);
    layer0_outputs(8752) <= not b;
    layer0_outputs(8753) <= a or b;
    layer0_outputs(8754) <= not (a or b);
    layer0_outputs(8755) <= '0';
    layer0_outputs(8756) <= a and b;
    layer0_outputs(8757) <= not a;
    layer0_outputs(8758) <= not (a or b);
    layer0_outputs(8759) <= a xor b;
    layer0_outputs(8760) <= not a;
    layer0_outputs(8761) <= not (a xor b);
    layer0_outputs(8762) <= not b;
    layer0_outputs(8763) <= b;
    layer0_outputs(8764) <= a and b;
    layer0_outputs(8765) <= a and not b;
    layer0_outputs(8766) <= not b;
    layer0_outputs(8767) <= not (a xor b);
    layer0_outputs(8768) <= not b;
    layer0_outputs(8769) <= not a or b;
    layer0_outputs(8770) <= a or b;
    layer0_outputs(8771) <= a;
    layer0_outputs(8772) <= not b;
    layer0_outputs(8773) <= not b;
    layer0_outputs(8774) <= a or b;
    layer0_outputs(8775) <= not a;
    layer0_outputs(8776) <= not a;
    layer0_outputs(8777) <= not a or b;
    layer0_outputs(8778) <= a;
    layer0_outputs(8779) <= not (a and b);
    layer0_outputs(8780) <= not b or a;
    layer0_outputs(8781) <= a;
    layer0_outputs(8782) <= not (a xor b);
    layer0_outputs(8783) <= '1';
    layer0_outputs(8784) <= not (a and b);
    layer0_outputs(8785) <= a or b;
    layer0_outputs(8786) <= not (a xor b);
    layer0_outputs(8787) <= not b or a;
    layer0_outputs(8788) <= a and not b;
    layer0_outputs(8789) <= a;
    layer0_outputs(8790) <= not a;
    layer0_outputs(8791) <= a;
    layer0_outputs(8792) <= b;
    layer0_outputs(8793) <= a;
    layer0_outputs(8794) <= not a or b;
    layer0_outputs(8795) <= not (a and b);
    layer0_outputs(8796) <= not (a and b);
    layer0_outputs(8797) <= a;
    layer0_outputs(8798) <= not (a or b);
    layer0_outputs(8799) <= b;
    layer0_outputs(8800) <= '1';
    layer0_outputs(8801) <= not a or b;
    layer0_outputs(8802) <= a xor b;
    layer0_outputs(8803) <= not (a or b);
    layer0_outputs(8804) <= not a;
    layer0_outputs(8805) <= a;
    layer0_outputs(8806) <= a and b;
    layer0_outputs(8807) <= not (a xor b);
    layer0_outputs(8808) <= b;
    layer0_outputs(8809) <= a or b;
    layer0_outputs(8810) <= not b or a;
    layer0_outputs(8811) <= not a or b;
    layer0_outputs(8812) <= a xor b;
    layer0_outputs(8813) <= not a;
    layer0_outputs(8814) <= not a;
    layer0_outputs(8815) <= a;
    layer0_outputs(8816) <= a or b;
    layer0_outputs(8817) <= b and not a;
    layer0_outputs(8818) <= a;
    layer0_outputs(8819) <= a and b;
    layer0_outputs(8820) <= not b or a;
    layer0_outputs(8821) <= a and not b;
    layer0_outputs(8822) <= a;
    layer0_outputs(8823) <= not (a or b);
    layer0_outputs(8824) <= a or b;
    layer0_outputs(8825) <= a or b;
    layer0_outputs(8826) <= a xor b;
    layer0_outputs(8827) <= '1';
    layer0_outputs(8828) <= '1';
    layer0_outputs(8829) <= not a or b;
    layer0_outputs(8830) <= not b;
    layer0_outputs(8831) <= '1';
    layer0_outputs(8832) <= not b;
    layer0_outputs(8833) <= b and not a;
    layer0_outputs(8834) <= b;
    layer0_outputs(8835) <= not (a xor b);
    layer0_outputs(8836) <= '1';
    layer0_outputs(8837) <= not (a xor b);
    layer0_outputs(8838) <= not a;
    layer0_outputs(8839) <= a or b;
    layer0_outputs(8840) <= not a;
    layer0_outputs(8841) <= not b;
    layer0_outputs(8842) <= '0';
    layer0_outputs(8843) <= not b;
    layer0_outputs(8844) <= not b or a;
    layer0_outputs(8845) <= not b;
    layer0_outputs(8846) <= a or b;
    layer0_outputs(8847) <= not b;
    layer0_outputs(8848) <= a xor b;
    layer0_outputs(8849) <= not b;
    layer0_outputs(8850) <= a xor b;
    layer0_outputs(8851) <= b and not a;
    layer0_outputs(8852) <= not (a xor b);
    layer0_outputs(8853) <= not (a or b);
    layer0_outputs(8854) <= not b;
    layer0_outputs(8855) <= not a;
    layer0_outputs(8856) <= a xor b;
    layer0_outputs(8857) <= a;
    layer0_outputs(8858) <= a;
    layer0_outputs(8859) <= a;
    layer0_outputs(8860) <= a or b;
    layer0_outputs(8861) <= b and not a;
    layer0_outputs(8862) <= not a;
    layer0_outputs(8863) <= not b;
    layer0_outputs(8864) <= b;
    layer0_outputs(8865) <= '0';
    layer0_outputs(8866) <= not (a and b);
    layer0_outputs(8867) <= not b;
    layer0_outputs(8868) <= not b;
    layer0_outputs(8869) <= not a or b;
    layer0_outputs(8870) <= not (a and b);
    layer0_outputs(8871) <= a and b;
    layer0_outputs(8872) <= '0';
    layer0_outputs(8873) <= a xor b;
    layer0_outputs(8874) <= '0';
    layer0_outputs(8875) <= not b;
    layer0_outputs(8876) <= not (a or b);
    layer0_outputs(8877) <= '0';
    layer0_outputs(8878) <= b;
    layer0_outputs(8879) <= not (a and b);
    layer0_outputs(8880) <= not a or b;
    layer0_outputs(8881) <= b and not a;
    layer0_outputs(8882) <= not b or a;
    layer0_outputs(8883) <= not (a or b);
    layer0_outputs(8884) <= a and not b;
    layer0_outputs(8885) <= a and not b;
    layer0_outputs(8886) <= a and b;
    layer0_outputs(8887) <= a or b;
    layer0_outputs(8888) <= not a;
    layer0_outputs(8889) <= not (a or b);
    layer0_outputs(8890) <= not b or a;
    layer0_outputs(8891) <= not (a xor b);
    layer0_outputs(8892) <= not b;
    layer0_outputs(8893) <= b;
    layer0_outputs(8894) <= b;
    layer0_outputs(8895) <= b;
    layer0_outputs(8896) <= not (a xor b);
    layer0_outputs(8897) <= a;
    layer0_outputs(8898) <= not (a xor b);
    layer0_outputs(8899) <= a or b;
    layer0_outputs(8900) <= '0';
    layer0_outputs(8901) <= b and not a;
    layer0_outputs(8902) <= a and not b;
    layer0_outputs(8903) <= not (a or b);
    layer0_outputs(8904) <= a xor b;
    layer0_outputs(8905) <= a and not b;
    layer0_outputs(8906) <= not (a xor b);
    layer0_outputs(8907) <= b;
    layer0_outputs(8908) <= not (a or b);
    layer0_outputs(8909) <= not b or a;
    layer0_outputs(8910) <= a xor b;
    layer0_outputs(8911) <= not a or b;
    layer0_outputs(8912) <= not (a and b);
    layer0_outputs(8913) <= not a or b;
    layer0_outputs(8914) <= '0';
    layer0_outputs(8915) <= a and b;
    layer0_outputs(8916) <= a or b;
    layer0_outputs(8917) <= not (a or b);
    layer0_outputs(8918) <= not b;
    layer0_outputs(8919) <= a xor b;
    layer0_outputs(8920) <= a;
    layer0_outputs(8921) <= not (a and b);
    layer0_outputs(8922) <= not b or a;
    layer0_outputs(8923) <= a and b;
    layer0_outputs(8924) <= b and not a;
    layer0_outputs(8925) <= not (a or b);
    layer0_outputs(8926) <= not (a or b);
    layer0_outputs(8927) <= not (a or b);
    layer0_outputs(8928) <= a and not b;
    layer0_outputs(8929) <= '0';
    layer0_outputs(8930) <= '1';
    layer0_outputs(8931) <= b and not a;
    layer0_outputs(8932) <= a and b;
    layer0_outputs(8933) <= '1';
    layer0_outputs(8934) <= not b;
    layer0_outputs(8935) <= not (a xor b);
    layer0_outputs(8936) <= a xor b;
    layer0_outputs(8937) <= a and b;
    layer0_outputs(8938) <= not (a xor b);
    layer0_outputs(8939) <= not a;
    layer0_outputs(8940) <= '0';
    layer0_outputs(8941) <= not a or b;
    layer0_outputs(8942) <= not b;
    layer0_outputs(8943) <= a or b;
    layer0_outputs(8944) <= '1';
    layer0_outputs(8945) <= '0';
    layer0_outputs(8946) <= a or b;
    layer0_outputs(8947) <= a;
    layer0_outputs(8948) <= not (a or b);
    layer0_outputs(8949) <= b;
    layer0_outputs(8950) <= b and not a;
    layer0_outputs(8951) <= b;
    layer0_outputs(8952) <= not (a or b);
    layer0_outputs(8953) <= b;
    layer0_outputs(8954) <= not (a xor b);
    layer0_outputs(8955) <= a;
    layer0_outputs(8956) <= a and not b;
    layer0_outputs(8957) <= not a;
    layer0_outputs(8958) <= not (a or b);
    layer0_outputs(8959) <= a;
    layer0_outputs(8960) <= not a or b;
    layer0_outputs(8961) <= not a;
    layer0_outputs(8962) <= a xor b;
    layer0_outputs(8963) <= not b or a;
    layer0_outputs(8964) <= a and not b;
    layer0_outputs(8965) <= not (a or b);
    layer0_outputs(8966) <= a and b;
    layer0_outputs(8967) <= a or b;
    layer0_outputs(8968) <= not (a and b);
    layer0_outputs(8969) <= a or b;
    layer0_outputs(8970) <= b and not a;
    layer0_outputs(8971) <= '0';
    layer0_outputs(8972) <= not (a or b);
    layer0_outputs(8973) <= a;
    layer0_outputs(8974) <= '1';
    layer0_outputs(8975) <= not (a xor b);
    layer0_outputs(8976) <= b;
    layer0_outputs(8977) <= not (a or b);
    layer0_outputs(8978) <= '0';
    layer0_outputs(8979) <= a and b;
    layer0_outputs(8980) <= a and not b;
    layer0_outputs(8981) <= a and not b;
    layer0_outputs(8982) <= not (a and b);
    layer0_outputs(8983) <= not (a and b);
    layer0_outputs(8984) <= a;
    layer0_outputs(8985) <= '0';
    layer0_outputs(8986) <= not a;
    layer0_outputs(8987) <= not a or b;
    layer0_outputs(8988) <= not a;
    layer0_outputs(8989) <= not (a or b);
    layer0_outputs(8990) <= not (a or b);
    layer0_outputs(8991) <= b;
    layer0_outputs(8992) <= not (a and b);
    layer0_outputs(8993) <= not (a or b);
    layer0_outputs(8994) <= '1';
    layer0_outputs(8995) <= b;
    layer0_outputs(8996) <= not (a and b);
    layer0_outputs(8997) <= a and not b;
    layer0_outputs(8998) <= b and not a;
    layer0_outputs(8999) <= not (a or b);
    layer0_outputs(9000) <= not b or a;
    layer0_outputs(9001) <= '0';
    layer0_outputs(9002) <= a or b;
    layer0_outputs(9003) <= a or b;
    layer0_outputs(9004) <= a or b;
    layer0_outputs(9005) <= b;
    layer0_outputs(9006) <= a xor b;
    layer0_outputs(9007) <= not (a and b);
    layer0_outputs(9008) <= not b;
    layer0_outputs(9009) <= not (a xor b);
    layer0_outputs(9010) <= a and b;
    layer0_outputs(9011) <= not a or b;
    layer0_outputs(9012) <= a or b;
    layer0_outputs(9013) <= not b or a;
    layer0_outputs(9014) <= not a or b;
    layer0_outputs(9015) <= a;
    layer0_outputs(9016) <= a or b;
    layer0_outputs(9017) <= b;
    layer0_outputs(9018) <= a and not b;
    layer0_outputs(9019) <= not a or b;
    layer0_outputs(9020) <= a and not b;
    layer0_outputs(9021) <= a;
    layer0_outputs(9022) <= not (a or b);
    layer0_outputs(9023) <= not (a or b);
    layer0_outputs(9024) <= '1';
    layer0_outputs(9025) <= a or b;
    layer0_outputs(9026) <= a xor b;
    layer0_outputs(9027) <= not b or a;
    layer0_outputs(9028) <= a or b;
    layer0_outputs(9029) <= not a;
    layer0_outputs(9030) <= not (a xor b);
    layer0_outputs(9031) <= not (a and b);
    layer0_outputs(9032) <= not a or b;
    layer0_outputs(9033) <= a or b;
    layer0_outputs(9034) <= not (a xor b);
    layer0_outputs(9035) <= a and not b;
    layer0_outputs(9036) <= '0';
    layer0_outputs(9037) <= not a or b;
    layer0_outputs(9038) <= '1';
    layer0_outputs(9039) <= not a;
    layer0_outputs(9040) <= '1';
    layer0_outputs(9041) <= a or b;
    layer0_outputs(9042) <= not a or b;
    layer0_outputs(9043) <= '1';
    layer0_outputs(9044) <= not (a and b);
    layer0_outputs(9045) <= '1';
    layer0_outputs(9046) <= not a;
    layer0_outputs(9047) <= '0';
    layer0_outputs(9048) <= '1';
    layer0_outputs(9049) <= '0';
    layer0_outputs(9050) <= a xor b;
    layer0_outputs(9051) <= a xor b;
    layer0_outputs(9052) <= a and not b;
    layer0_outputs(9053) <= not a;
    layer0_outputs(9054) <= not b;
    layer0_outputs(9055) <= a and not b;
    layer0_outputs(9056) <= '1';
    layer0_outputs(9057) <= b;
    layer0_outputs(9058) <= '1';
    layer0_outputs(9059) <= a or b;
    layer0_outputs(9060) <= not b or a;
    layer0_outputs(9061) <= not (a xor b);
    layer0_outputs(9062) <= a or b;
    layer0_outputs(9063) <= not (a or b);
    layer0_outputs(9064) <= not a or b;
    layer0_outputs(9065) <= not (a xor b);
    layer0_outputs(9066) <= a xor b;
    layer0_outputs(9067) <= b;
    layer0_outputs(9068) <= a xor b;
    layer0_outputs(9069) <= a xor b;
    layer0_outputs(9070) <= '0';
    layer0_outputs(9071) <= a or b;
    layer0_outputs(9072) <= not (a and b);
    layer0_outputs(9073) <= not (a and b);
    layer0_outputs(9074) <= a or b;
    layer0_outputs(9075) <= not (a and b);
    layer0_outputs(9076) <= not b or a;
    layer0_outputs(9077) <= b;
    layer0_outputs(9078) <= not a or b;
    layer0_outputs(9079) <= b;
    layer0_outputs(9080) <= '0';
    layer0_outputs(9081) <= a and not b;
    layer0_outputs(9082) <= not a or b;
    layer0_outputs(9083) <= '0';
    layer0_outputs(9084) <= not a;
    layer0_outputs(9085) <= not b;
    layer0_outputs(9086) <= a or b;
    layer0_outputs(9087) <= a xor b;
    layer0_outputs(9088) <= not b;
    layer0_outputs(9089) <= b;
    layer0_outputs(9090) <= a xor b;
    layer0_outputs(9091) <= '0';
    layer0_outputs(9092) <= a and b;
    layer0_outputs(9093) <= a and not b;
    layer0_outputs(9094) <= not (a xor b);
    layer0_outputs(9095) <= a or b;
    layer0_outputs(9096) <= b and not a;
    layer0_outputs(9097) <= a or b;
    layer0_outputs(9098) <= not (a xor b);
    layer0_outputs(9099) <= b and not a;
    layer0_outputs(9100) <= a and b;
    layer0_outputs(9101) <= b;
    layer0_outputs(9102) <= not b or a;
    layer0_outputs(9103) <= not (a or b);
    layer0_outputs(9104) <= a;
    layer0_outputs(9105) <= b;
    layer0_outputs(9106) <= b;
    layer0_outputs(9107) <= a and not b;
    layer0_outputs(9108) <= b;
    layer0_outputs(9109) <= not b or a;
    layer0_outputs(9110) <= not a or b;
    layer0_outputs(9111) <= a and b;
    layer0_outputs(9112) <= a and b;
    layer0_outputs(9113) <= a or b;
    layer0_outputs(9114) <= a xor b;
    layer0_outputs(9115) <= '0';
    layer0_outputs(9116) <= not (a or b);
    layer0_outputs(9117) <= not (a xor b);
    layer0_outputs(9118) <= a or b;
    layer0_outputs(9119) <= a and b;
    layer0_outputs(9120) <= a or b;
    layer0_outputs(9121) <= not (a and b);
    layer0_outputs(9122) <= not a or b;
    layer0_outputs(9123) <= not a or b;
    layer0_outputs(9124) <= not (a or b);
    layer0_outputs(9125) <= b;
    layer0_outputs(9126) <= '0';
    layer0_outputs(9127) <= not b or a;
    layer0_outputs(9128) <= not a or b;
    layer0_outputs(9129) <= b and not a;
    layer0_outputs(9130) <= a;
    layer0_outputs(9131) <= not b;
    layer0_outputs(9132) <= not b;
    layer0_outputs(9133) <= not a;
    layer0_outputs(9134) <= not (a and b);
    layer0_outputs(9135) <= b and not a;
    layer0_outputs(9136) <= not b or a;
    layer0_outputs(9137) <= not b;
    layer0_outputs(9138) <= a;
    layer0_outputs(9139) <= not (a and b);
    layer0_outputs(9140) <= a or b;
    layer0_outputs(9141) <= a or b;
    layer0_outputs(9142) <= not a or b;
    layer0_outputs(9143) <= not (a or b);
    layer0_outputs(9144) <= a or b;
    layer0_outputs(9145) <= not (a or b);
    layer0_outputs(9146) <= b;
    layer0_outputs(9147) <= a xor b;
    layer0_outputs(9148) <= a and not b;
    layer0_outputs(9149) <= a xor b;
    layer0_outputs(9150) <= not b;
    layer0_outputs(9151) <= b and not a;
    layer0_outputs(9152) <= '1';
    layer0_outputs(9153) <= a xor b;
    layer0_outputs(9154) <= a and not b;
    layer0_outputs(9155) <= a;
    layer0_outputs(9156) <= not b;
    layer0_outputs(9157) <= '1';
    layer0_outputs(9158) <= not a;
    layer0_outputs(9159) <= a xor b;
    layer0_outputs(9160) <= not (a or b);
    layer0_outputs(9161) <= b;
    layer0_outputs(9162) <= not a;
    layer0_outputs(9163) <= not (a xor b);
    layer0_outputs(9164) <= a or b;
    layer0_outputs(9165) <= a and b;
    layer0_outputs(9166) <= not (a xor b);
    layer0_outputs(9167) <= a or b;
    layer0_outputs(9168) <= not (a xor b);
    layer0_outputs(9169) <= not (a or b);
    layer0_outputs(9170) <= b and not a;
    layer0_outputs(9171) <= not (a and b);
    layer0_outputs(9172) <= not a;
    layer0_outputs(9173) <= not a or b;
    layer0_outputs(9174) <= not (a or b);
    layer0_outputs(9175) <= a;
    layer0_outputs(9176) <= a and b;
    layer0_outputs(9177) <= not (a or b);
    layer0_outputs(9178) <= not a or b;
    layer0_outputs(9179) <= a or b;
    layer0_outputs(9180) <= not (a xor b);
    layer0_outputs(9181) <= a;
    layer0_outputs(9182) <= a;
    layer0_outputs(9183) <= b and not a;
    layer0_outputs(9184) <= a and b;
    layer0_outputs(9185) <= not b;
    layer0_outputs(9186) <= b;
    layer0_outputs(9187) <= '0';
    layer0_outputs(9188) <= '1';
    layer0_outputs(9189) <= a or b;
    layer0_outputs(9190) <= a or b;
    layer0_outputs(9191) <= '1';
    layer0_outputs(9192) <= a or b;
    layer0_outputs(9193) <= not a;
    layer0_outputs(9194) <= not (a xor b);
    layer0_outputs(9195) <= not a or b;
    layer0_outputs(9196) <= not b;
    layer0_outputs(9197) <= a;
    layer0_outputs(9198) <= a;
    layer0_outputs(9199) <= b;
    layer0_outputs(9200) <= not b;
    layer0_outputs(9201) <= a xor b;
    layer0_outputs(9202) <= not (a or b);
    layer0_outputs(9203) <= not (a and b);
    layer0_outputs(9204) <= not (a and b);
    layer0_outputs(9205) <= not b or a;
    layer0_outputs(9206) <= '1';
    layer0_outputs(9207) <= a or b;
    layer0_outputs(9208) <= b and not a;
    layer0_outputs(9209) <= not a or b;
    layer0_outputs(9210) <= not a;
    layer0_outputs(9211) <= '0';
    layer0_outputs(9212) <= not a;
    layer0_outputs(9213) <= a or b;
    layer0_outputs(9214) <= a and not b;
    layer0_outputs(9215) <= b;
    layer0_outputs(9216) <= not (a and b);
    layer0_outputs(9217) <= not a or b;
    layer0_outputs(9218) <= a xor b;
    layer0_outputs(9219) <= a and b;
    layer0_outputs(9220) <= b;
    layer0_outputs(9221) <= not b;
    layer0_outputs(9222) <= a;
    layer0_outputs(9223) <= b;
    layer0_outputs(9224) <= a xor b;
    layer0_outputs(9225) <= b and not a;
    layer0_outputs(9226) <= not a or b;
    layer0_outputs(9227) <= b;
    layer0_outputs(9228) <= a and not b;
    layer0_outputs(9229) <= '0';
    layer0_outputs(9230) <= not a;
    layer0_outputs(9231) <= not (a or b);
    layer0_outputs(9232) <= not a or b;
    layer0_outputs(9233) <= not (a xor b);
    layer0_outputs(9234) <= not (a and b);
    layer0_outputs(9235) <= b and not a;
    layer0_outputs(9236) <= a;
    layer0_outputs(9237) <= not b;
    layer0_outputs(9238) <= not b or a;
    layer0_outputs(9239) <= not a;
    layer0_outputs(9240) <= a;
    layer0_outputs(9241) <= b;
    layer0_outputs(9242) <= not b or a;
    layer0_outputs(9243) <= b;
    layer0_outputs(9244) <= '1';
    layer0_outputs(9245) <= b;
    layer0_outputs(9246) <= a;
    layer0_outputs(9247) <= not a or b;
    layer0_outputs(9248) <= not (a or b);
    layer0_outputs(9249) <= b and not a;
    layer0_outputs(9250) <= a xor b;
    layer0_outputs(9251) <= not (a or b);
    layer0_outputs(9252) <= a and not b;
    layer0_outputs(9253) <= b and not a;
    layer0_outputs(9254) <= not a or b;
    layer0_outputs(9255) <= not a or b;
    layer0_outputs(9256) <= a or b;
    layer0_outputs(9257) <= not (a and b);
    layer0_outputs(9258) <= b;
    layer0_outputs(9259) <= not (a xor b);
    layer0_outputs(9260) <= '1';
    layer0_outputs(9261) <= not (a or b);
    layer0_outputs(9262) <= not (a and b);
    layer0_outputs(9263) <= '1';
    layer0_outputs(9264) <= not b;
    layer0_outputs(9265) <= a or b;
    layer0_outputs(9266) <= not (a or b);
    layer0_outputs(9267) <= not (a or b);
    layer0_outputs(9268) <= a or b;
    layer0_outputs(9269) <= not (a xor b);
    layer0_outputs(9270) <= a;
    layer0_outputs(9271) <= a;
    layer0_outputs(9272) <= not a;
    layer0_outputs(9273) <= b and not a;
    layer0_outputs(9274) <= not b;
    layer0_outputs(9275) <= a or b;
    layer0_outputs(9276) <= a xor b;
    layer0_outputs(9277) <= a xor b;
    layer0_outputs(9278) <= b;
    layer0_outputs(9279) <= b;
    layer0_outputs(9280) <= a xor b;
    layer0_outputs(9281) <= not a or b;
    layer0_outputs(9282) <= a and not b;
    layer0_outputs(9283) <= not a;
    layer0_outputs(9284) <= not (a or b);
    layer0_outputs(9285) <= b;
    layer0_outputs(9286) <= not a;
    layer0_outputs(9287) <= not (a or b);
    layer0_outputs(9288) <= not b;
    layer0_outputs(9289) <= not a;
    layer0_outputs(9290) <= a;
    layer0_outputs(9291) <= not a or b;
    layer0_outputs(9292) <= not b or a;
    layer0_outputs(9293) <= not (a xor b);
    layer0_outputs(9294) <= not (a xor b);
    layer0_outputs(9295) <= a;
    layer0_outputs(9296) <= a xor b;
    layer0_outputs(9297) <= a xor b;
    layer0_outputs(9298) <= a xor b;
    layer0_outputs(9299) <= a;
    layer0_outputs(9300) <= not b;
    layer0_outputs(9301) <= a and not b;
    layer0_outputs(9302) <= not b;
    layer0_outputs(9303) <= b and not a;
    layer0_outputs(9304) <= not (a xor b);
    layer0_outputs(9305) <= not (a or b);
    layer0_outputs(9306) <= a xor b;
    layer0_outputs(9307) <= b;
    layer0_outputs(9308) <= b and not a;
    layer0_outputs(9309) <= not a;
    layer0_outputs(9310) <= a and b;
    layer0_outputs(9311) <= a or b;
    layer0_outputs(9312) <= a;
    layer0_outputs(9313) <= b;
    layer0_outputs(9314) <= a or b;
    layer0_outputs(9315) <= not (a xor b);
    layer0_outputs(9316) <= a;
    layer0_outputs(9317) <= '1';
    layer0_outputs(9318) <= not (a or b);
    layer0_outputs(9319) <= b;
    layer0_outputs(9320) <= a and b;
    layer0_outputs(9321) <= b;
    layer0_outputs(9322) <= a and not b;
    layer0_outputs(9323) <= not b;
    layer0_outputs(9324) <= not a;
    layer0_outputs(9325) <= a;
    layer0_outputs(9326) <= a;
    layer0_outputs(9327) <= b and not a;
    layer0_outputs(9328) <= not a;
    layer0_outputs(9329) <= not a or b;
    layer0_outputs(9330) <= not (a and b);
    layer0_outputs(9331) <= a xor b;
    layer0_outputs(9332) <= not (a and b);
    layer0_outputs(9333) <= '1';
    layer0_outputs(9334) <= not b;
    layer0_outputs(9335) <= a or b;
    layer0_outputs(9336) <= not (a xor b);
    layer0_outputs(9337) <= not a;
    layer0_outputs(9338) <= not b;
    layer0_outputs(9339) <= b and not a;
    layer0_outputs(9340) <= b;
    layer0_outputs(9341) <= not (a xor b);
    layer0_outputs(9342) <= not a or b;
    layer0_outputs(9343) <= a xor b;
    layer0_outputs(9344) <= b and not a;
    layer0_outputs(9345) <= not (a and b);
    layer0_outputs(9346) <= not a;
    layer0_outputs(9347) <= not a;
    layer0_outputs(9348) <= '1';
    layer0_outputs(9349) <= a xor b;
    layer0_outputs(9350) <= a and b;
    layer0_outputs(9351) <= not a;
    layer0_outputs(9352) <= b;
    layer0_outputs(9353) <= not b;
    layer0_outputs(9354) <= not b;
    layer0_outputs(9355) <= a;
    layer0_outputs(9356) <= a;
    layer0_outputs(9357) <= a or b;
    layer0_outputs(9358) <= not a or b;
    layer0_outputs(9359) <= b;
    layer0_outputs(9360) <= b;
    layer0_outputs(9361) <= a xor b;
    layer0_outputs(9362) <= '1';
    layer0_outputs(9363) <= a;
    layer0_outputs(9364) <= not (a xor b);
    layer0_outputs(9365) <= not b;
    layer0_outputs(9366) <= not a or b;
    layer0_outputs(9367) <= '0';
    layer0_outputs(9368) <= a or b;
    layer0_outputs(9369) <= not (a or b);
    layer0_outputs(9370) <= not a or b;
    layer0_outputs(9371) <= a;
    layer0_outputs(9372) <= b and not a;
    layer0_outputs(9373) <= not (a or b);
    layer0_outputs(9374) <= not b;
    layer0_outputs(9375) <= '1';
    layer0_outputs(9376) <= not a;
    layer0_outputs(9377) <= not a or b;
    layer0_outputs(9378) <= a or b;
    layer0_outputs(9379) <= not (a xor b);
    layer0_outputs(9380) <= a xor b;
    layer0_outputs(9381) <= a or b;
    layer0_outputs(9382) <= a;
    layer0_outputs(9383) <= a xor b;
    layer0_outputs(9384) <= b;
    layer0_outputs(9385) <= not (a or b);
    layer0_outputs(9386) <= not a;
    layer0_outputs(9387) <= a or b;
    layer0_outputs(9388) <= a or b;
    layer0_outputs(9389) <= '0';
    layer0_outputs(9390) <= a and not b;
    layer0_outputs(9391) <= b;
    layer0_outputs(9392) <= not (a xor b);
    layer0_outputs(9393) <= not (a xor b);
    layer0_outputs(9394) <= not a or b;
    layer0_outputs(9395) <= not (a or b);
    layer0_outputs(9396) <= b and not a;
    layer0_outputs(9397) <= not (a or b);
    layer0_outputs(9398) <= not a;
    layer0_outputs(9399) <= '0';
    layer0_outputs(9400) <= a xor b;
    layer0_outputs(9401) <= '0';
    layer0_outputs(9402) <= '0';
    layer0_outputs(9403) <= a or b;
    layer0_outputs(9404) <= b and not a;
    layer0_outputs(9405) <= a and b;
    layer0_outputs(9406) <= not b or a;
    layer0_outputs(9407) <= b and not a;
    layer0_outputs(9408) <= b and not a;
    layer0_outputs(9409) <= a and b;
    layer0_outputs(9410) <= not (a xor b);
    layer0_outputs(9411) <= b;
    layer0_outputs(9412) <= not (a and b);
    layer0_outputs(9413) <= not (a and b);
    layer0_outputs(9414) <= a xor b;
    layer0_outputs(9415) <= a and not b;
    layer0_outputs(9416) <= not b or a;
    layer0_outputs(9417) <= b and not a;
    layer0_outputs(9418) <= not (a and b);
    layer0_outputs(9419) <= a or b;
    layer0_outputs(9420) <= b and not a;
    layer0_outputs(9421) <= not a;
    layer0_outputs(9422) <= not b;
    layer0_outputs(9423) <= not a;
    layer0_outputs(9424) <= '0';
    layer0_outputs(9425) <= '0';
    layer0_outputs(9426) <= '1';
    layer0_outputs(9427) <= a xor b;
    layer0_outputs(9428) <= a xor b;
    layer0_outputs(9429) <= not b;
    layer0_outputs(9430) <= b and not a;
    layer0_outputs(9431) <= not (a xor b);
    layer0_outputs(9432) <= '1';
    layer0_outputs(9433) <= not (a xor b);
    layer0_outputs(9434) <= not a;
    layer0_outputs(9435) <= not b or a;
    layer0_outputs(9436) <= a xor b;
    layer0_outputs(9437) <= a;
    layer0_outputs(9438) <= not b;
    layer0_outputs(9439) <= a;
    layer0_outputs(9440) <= '1';
    layer0_outputs(9441) <= b and not a;
    layer0_outputs(9442) <= not b or a;
    layer0_outputs(9443) <= a;
    layer0_outputs(9444) <= a and not b;
    layer0_outputs(9445) <= b and not a;
    layer0_outputs(9446) <= not (a or b);
    layer0_outputs(9447) <= not b;
    layer0_outputs(9448) <= not a or b;
    layer0_outputs(9449) <= not (a and b);
    layer0_outputs(9450) <= a;
    layer0_outputs(9451) <= a xor b;
    layer0_outputs(9452) <= '0';
    layer0_outputs(9453) <= not b or a;
    layer0_outputs(9454) <= not a;
    layer0_outputs(9455) <= not (a or b);
    layer0_outputs(9456) <= not a or b;
    layer0_outputs(9457) <= a and not b;
    layer0_outputs(9458) <= not b;
    layer0_outputs(9459) <= b;
    layer0_outputs(9460) <= not b or a;
    layer0_outputs(9461) <= a or b;
    layer0_outputs(9462) <= a and b;
    layer0_outputs(9463) <= a and b;
    layer0_outputs(9464) <= b and not a;
    layer0_outputs(9465) <= a or b;
    layer0_outputs(9466) <= b;
    layer0_outputs(9467) <= a and not b;
    layer0_outputs(9468) <= a;
    layer0_outputs(9469) <= '0';
    layer0_outputs(9470) <= a or b;
    layer0_outputs(9471) <= not (a and b);
    layer0_outputs(9472) <= b;
    layer0_outputs(9473) <= not (a and b);
    layer0_outputs(9474) <= not b or a;
    layer0_outputs(9475) <= a and not b;
    layer0_outputs(9476) <= not (a or b);
    layer0_outputs(9477) <= a;
    layer0_outputs(9478) <= not a or b;
    layer0_outputs(9479) <= '0';
    layer0_outputs(9480) <= a and b;
    layer0_outputs(9481) <= b and not a;
    layer0_outputs(9482) <= not b;
    layer0_outputs(9483) <= not b or a;
    layer0_outputs(9484) <= not (a or b);
    layer0_outputs(9485) <= a or b;
    layer0_outputs(9486) <= a or b;
    layer0_outputs(9487) <= not (a or b);
    layer0_outputs(9488) <= not b or a;
    layer0_outputs(9489) <= a;
    layer0_outputs(9490) <= not a or b;
    layer0_outputs(9491) <= not a;
    layer0_outputs(9492) <= a and not b;
    layer0_outputs(9493) <= not (a or b);
    layer0_outputs(9494) <= b and not a;
    layer0_outputs(9495) <= not (a xor b);
    layer0_outputs(9496) <= not (a or b);
    layer0_outputs(9497) <= a;
    layer0_outputs(9498) <= b;
    layer0_outputs(9499) <= a and not b;
    layer0_outputs(9500) <= a and not b;
    layer0_outputs(9501) <= a xor b;
    layer0_outputs(9502) <= a and b;
    layer0_outputs(9503) <= b;
    layer0_outputs(9504) <= not a or b;
    layer0_outputs(9505) <= a or b;
    layer0_outputs(9506) <= not b;
    layer0_outputs(9507) <= a or b;
    layer0_outputs(9508) <= not (a or b);
    layer0_outputs(9509) <= a and not b;
    layer0_outputs(9510) <= a and not b;
    layer0_outputs(9511) <= '1';
    layer0_outputs(9512) <= a xor b;
    layer0_outputs(9513) <= b and not a;
    layer0_outputs(9514) <= not a or b;
    layer0_outputs(9515) <= not a or b;
    layer0_outputs(9516) <= not (a xor b);
    layer0_outputs(9517) <= a and not b;
    layer0_outputs(9518) <= not (a and b);
    layer0_outputs(9519) <= a xor b;
    layer0_outputs(9520) <= not a;
    layer0_outputs(9521) <= a or b;
    layer0_outputs(9522) <= not b or a;
    layer0_outputs(9523) <= not b or a;
    layer0_outputs(9524) <= not (a or b);
    layer0_outputs(9525) <= a xor b;
    layer0_outputs(9526) <= b;
    layer0_outputs(9527) <= a xor b;
    layer0_outputs(9528) <= not b;
    layer0_outputs(9529) <= not (a xor b);
    layer0_outputs(9530) <= b;
    layer0_outputs(9531) <= a or b;
    layer0_outputs(9532) <= not (a xor b);
    layer0_outputs(9533) <= a and not b;
    layer0_outputs(9534) <= not a or b;
    layer0_outputs(9535) <= not a or b;
    layer0_outputs(9536) <= a or b;
    layer0_outputs(9537) <= not (a and b);
    layer0_outputs(9538) <= a xor b;
    layer0_outputs(9539) <= '1';
    layer0_outputs(9540) <= a xor b;
    layer0_outputs(9541) <= not b;
    layer0_outputs(9542) <= b and not a;
    layer0_outputs(9543) <= not a or b;
    layer0_outputs(9544) <= a or b;
    layer0_outputs(9545) <= not b;
    layer0_outputs(9546) <= not b or a;
    layer0_outputs(9547) <= b and not a;
    layer0_outputs(9548) <= b;
    layer0_outputs(9549) <= b and not a;
    layer0_outputs(9550) <= a xor b;
    layer0_outputs(9551) <= not b or a;
    layer0_outputs(9552) <= not b or a;
    layer0_outputs(9553) <= a and b;
    layer0_outputs(9554) <= not b;
    layer0_outputs(9555) <= b and not a;
    layer0_outputs(9556) <= a and not b;
    layer0_outputs(9557) <= b and not a;
    layer0_outputs(9558) <= b and not a;
    layer0_outputs(9559) <= '1';
    layer0_outputs(9560) <= a;
    layer0_outputs(9561) <= a and b;
    layer0_outputs(9562) <= not (a xor b);
    layer0_outputs(9563) <= a or b;
    layer0_outputs(9564) <= a and b;
    layer0_outputs(9565) <= not a;
    layer0_outputs(9566) <= not (a or b);
    layer0_outputs(9567) <= a xor b;
    layer0_outputs(9568) <= b;
    layer0_outputs(9569) <= a;
    layer0_outputs(9570) <= not a or b;
    layer0_outputs(9571) <= not b or a;
    layer0_outputs(9572) <= not a or b;
    layer0_outputs(9573) <= not (a and b);
    layer0_outputs(9574) <= not (a or b);
    layer0_outputs(9575) <= not (a and b);
    layer0_outputs(9576) <= a or b;
    layer0_outputs(9577) <= a;
    layer0_outputs(9578) <= a xor b;
    layer0_outputs(9579) <= a or b;
    layer0_outputs(9580) <= b;
    layer0_outputs(9581) <= b and not a;
    layer0_outputs(9582) <= b and not a;
    layer0_outputs(9583) <= a xor b;
    layer0_outputs(9584) <= a;
    layer0_outputs(9585) <= not a;
    layer0_outputs(9586) <= '1';
    layer0_outputs(9587) <= not (a and b);
    layer0_outputs(9588) <= not a;
    layer0_outputs(9589) <= '1';
    layer0_outputs(9590) <= a;
    layer0_outputs(9591) <= not b;
    layer0_outputs(9592) <= a and not b;
    layer0_outputs(9593) <= not (a or b);
    layer0_outputs(9594) <= '1';
    layer0_outputs(9595) <= a xor b;
    layer0_outputs(9596) <= a or b;
    layer0_outputs(9597) <= not b or a;
    layer0_outputs(9598) <= a and b;
    layer0_outputs(9599) <= not (a or b);
    layer0_outputs(9600) <= not b;
    layer0_outputs(9601) <= b and not a;
    layer0_outputs(9602) <= a xor b;
    layer0_outputs(9603) <= a and not b;
    layer0_outputs(9604) <= not a;
    layer0_outputs(9605) <= a or b;
    layer0_outputs(9606) <= b;
    layer0_outputs(9607) <= not b;
    layer0_outputs(9608) <= not (a or b);
    layer0_outputs(9609) <= not a or b;
    layer0_outputs(9610) <= b;
    layer0_outputs(9611) <= a or b;
    layer0_outputs(9612) <= not a or b;
    layer0_outputs(9613) <= not a or b;
    layer0_outputs(9614) <= '1';
    layer0_outputs(9615) <= a xor b;
    layer0_outputs(9616) <= not a;
    layer0_outputs(9617) <= '0';
    layer0_outputs(9618) <= not (a or b);
    layer0_outputs(9619) <= not (a xor b);
    layer0_outputs(9620) <= a xor b;
    layer0_outputs(9621) <= a xor b;
    layer0_outputs(9622) <= not b;
    layer0_outputs(9623) <= not (a xor b);
    layer0_outputs(9624) <= not a or b;
    layer0_outputs(9625) <= not (a or b);
    layer0_outputs(9626) <= '0';
    layer0_outputs(9627) <= not b;
    layer0_outputs(9628) <= not (a or b);
    layer0_outputs(9629) <= not (a xor b);
    layer0_outputs(9630) <= not (a xor b);
    layer0_outputs(9631) <= not (a xor b);
    layer0_outputs(9632) <= not b or a;
    layer0_outputs(9633) <= not b or a;
    layer0_outputs(9634) <= b;
    layer0_outputs(9635) <= not b;
    layer0_outputs(9636) <= a and b;
    layer0_outputs(9637) <= a or b;
    layer0_outputs(9638) <= not (a or b);
    layer0_outputs(9639) <= a and not b;
    layer0_outputs(9640) <= a and b;
    layer0_outputs(9641) <= not a;
    layer0_outputs(9642) <= '0';
    layer0_outputs(9643) <= '1';
    layer0_outputs(9644) <= b;
    layer0_outputs(9645) <= a;
    layer0_outputs(9646) <= '0';
    layer0_outputs(9647) <= a and b;
    layer0_outputs(9648) <= '0';
    layer0_outputs(9649) <= not a;
    layer0_outputs(9650) <= not a;
    layer0_outputs(9651) <= not a or b;
    layer0_outputs(9652) <= not (a or b);
    layer0_outputs(9653) <= '1';
    layer0_outputs(9654) <= not (a or b);
    layer0_outputs(9655) <= not a;
    layer0_outputs(9656) <= not a or b;
    layer0_outputs(9657) <= b;
    layer0_outputs(9658) <= a or b;
    layer0_outputs(9659) <= a;
    layer0_outputs(9660) <= not (a xor b);
    layer0_outputs(9661) <= not b;
    layer0_outputs(9662) <= not a or b;
    layer0_outputs(9663) <= a and not b;
    layer0_outputs(9664) <= not (a xor b);
    layer0_outputs(9665) <= '1';
    layer0_outputs(9666) <= '0';
    layer0_outputs(9667) <= '1';
    layer0_outputs(9668) <= '1';
    layer0_outputs(9669) <= not b;
    layer0_outputs(9670) <= a;
    layer0_outputs(9671) <= not b;
    layer0_outputs(9672) <= b and not a;
    layer0_outputs(9673) <= a xor b;
    layer0_outputs(9674) <= not (a or b);
    layer0_outputs(9675) <= not a or b;
    layer0_outputs(9676) <= '1';
    layer0_outputs(9677) <= not a or b;
    layer0_outputs(9678) <= a;
    layer0_outputs(9679) <= not b;
    layer0_outputs(9680) <= a xor b;
    layer0_outputs(9681) <= not b or a;
    layer0_outputs(9682) <= b and not a;
    layer0_outputs(9683) <= a;
    layer0_outputs(9684) <= '1';
    layer0_outputs(9685) <= a;
    layer0_outputs(9686) <= not (a or b);
    layer0_outputs(9687) <= b and not a;
    layer0_outputs(9688) <= not (a xor b);
    layer0_outputs(9689) <= b and not a;
    layer0_outputs(9690) <= not a or b;
    layer0_outputs(9691) <= not a or b;
    layer0_outputs(9692) <= a and b;
    layer0_outputs(9693) <= a;
    layer0_outputs(9694) <= a xor b;
    layer0_outputs(9695) <= not b or a;
    layer0_outputs(9696) <= a xor b;
    layer0_outputs(9697) <= a and b;
    layer0_outputs(9698) <= not (a xor b);
    layer0_outputs(9699) <= a and b;
    layer0_outputs(9700) <= not (a or b);
    layer0_outputs(9701) <= '0';
    layer0_outputs(9702) <= a;
    layer0_outputs(9703) <= not b;
    layer0_outputs(9704) <= not a;
    layer0_outputs(9705) <= not b;
    layer0_outputs(9706) <= b;
    layer0_outputs(9707) <= a;
    layer0_outputs(9708) <= a or b;
    layer0_outputs(9709) <= not a or b;
    layer0_outputs(9710) <= a;
    layer0_outputs(9711) <= a and b;
    layer0_outputs(9712) <= a or b;
    layer0_outputs(9713) <= not (a xor b);
    layer0_outputs(9714) <= not b or a;
    layer0_outputs(9715) <= not (a xor b);
    layer0_outputs(9716) <= not b;
    layer0_outputs(9717) <= not (a or b);
    layer0_outputs(9718) <= a and b;
    layer0_outputs(9719) <= not a;
    layer0_outputs(9720) <= a;
    layer0_outputs(9721) <= b;
    layer0_outputs(9722) <= '1';
    layer0_outputs(9723) <= '0';
    layer0_outputs(9724) <= not a;
    layer0_outputs(9725) <= a and not b;
    layer0_outputs(9726) <= a;
    layer0_outputs(9727) <= not b or a;
    layer0_outputs(9728) <= a and b;
    layer0_outputs(9729) <= '1';
    layer0_outputs(9730) <= not (a or b);
    layer0_outputs(9731) <= not a;
    layer0_outputs(9732) <= a or b;
    layer0_outputs(9733) <= not b or a;
    layer0_outputs(9734) <= a and not b;
    layer0_outputs(9735) <= not b;
    layer0_outputs(9736) <= not a or b;
    layer0_outputs(9737) <= b and not a;
    layer0_outputs(9738) <= not a;
    layer0_outputs(9739) <= not a or b;
    layer0_outputs(9740) <= not a;
    layer0_outputs(9741) <= not b;
    layer0_outputs(9742) <= not b;
    layer0_outputs(9743) <= a xor b;
    layer0_outputs(9744) <= not b;
    layer0_outputs(9745) <= not (a xor b);
    layer0_outputs(9746) <= b and not a;
    layer0_outputs(9747) <= not b;
    layer0_outputs(9748) <= a and b;
    layer0_outputs(9749) <= not (a or b);
    layer0_outputs(9750) <= not a or b;
    layer0_outputs(9751) <= not b;
    layer0_outputs(9752) <= a;
    layer0_outputs(9753) <= not (a xor b);
    layer0_outputs(9754) <= a;
    layer0_outputs(9755) <= a or b;
    layer0_outputs(9756) <= not b;
    layer0_outputs(9757) <= b and not a;
    layer0_outputs(9758) <= not a;
    layer0_outputs(9759) <= not b or a;
    layer0_outputs(9760) <= b;
    layer0_outputs(9761) <= a;
    layer0_outputs(9762) <= not (a and b);
    layer0_outputs(9763) <= not a;
    layer0_outputs(9764) <= not a;
    layer0_outputs(9765) <= '0';
    layer0_outputs(9766) <= a xor b;
    layer0_outputs(9767) <= b and not a;
    layer0_outputs(9768) <= b;
    layer0_outputs(9769) <= not a or b;
    layer0_outputs(9770) <= a xor b;
    layer0_outputs(9771) <= not a;
    layer0_outputs(9772) <= a xor b;
    layer0_outputs(9773) <= not a;
    layer0_outputs(9774) <= a;
    layer0_outputs(9775) <= not (a xor b);
    layer0_outputs(9776) <= '1';
    layer0_outputs(9777) <= a or b;
    layer0_outputs(9778) <= not (a or b);
    layer0_outputs(9779) <= not (a or b);
    layer0_outputs(9780) <= a xor b;
    layer0_outputs(9781) <= not (a xor b);
    layer0_outputs(9782) <= not (a xor b);
    layer0_outputs(9783) <= a or b;
    layer0_outputs(9784) <= not (a xor b);
    layer0_outputs(9785) <= not (a and b);
    layer0_outputs(9786) <= not b or a;
    layer0_outputs(9787) <= not b or a;
    layer0_outputs(9788) <= a or b;
    layer0_outputs(9789) <= '0';
    layer0_outputs(9790) <= '0';
    layer0_outputs(9791) <= not (a or b);
    layer0_outputs(9792) <= b and not a;
    layer0_outputs(9793) <= not (a and b);
    layer0_outputs(9794) <= a xor b;
    layer0_outputs(9795) <= a;
    layer0_outputs(9796) <= not (a and b);
    layer0_outputs(9797) <= a or b;
    layer0_outputs(9798) <= a;
    layer0_outputs(9799) <= not b;
    layer0_outputs(9800) <= not (a or b);
    layer0_outputs(9801) <= a and not b;
    layer0_outputs(9802) <= '1';
    layer0_outputs(9803) <= a;
    layer0_outputs(9804) <= a or b;
    layer0_outputs(9805) <= not a or b;
    layer0_outputs(9806) <= '1';
    layer0_outputs(9807) <= a xor b;
    layer0_outputs(9808) <= not b;
    layer0_outputs(9809) <= not (a or b);
    layer0_outputs(9810) <= not b;
    layer0_outputs(9811) <= b;
    layer0_outputs(9812) <= not (a xor b);
    layer0_outputs(9813) <= '1';
    layer0_outputs(9814) <= a xor b;
    layer0_outputs(9815) <= not a;
    layer0_outputs(9816) <= a xor b;
    layer0_outputs(9817) <= not (a or b);
    layer0_outputs(9818) <= not (a or b);
    layer0_outputs(9819) <= b;
    layer0_outputs(9820) <= not b or a;
    layer0_outputs(9821) <= a and b;
    layer0_outputs(9822) <= not (a and b);
    layer0_outputs(9823) <= b and not a;
    layer0_outputs(9824) <= a and b;
    layer0_outputs(9825) <= not b or a;
    layer0_outputs(9826) <= b;
    layer0_outputs(9827) <= '0';
    layer0_outputs(9828) <= a or b;
    layer0_outputs(9829) <= '1';
    layer0_outputs(9830) <= not (a or b);
    layer0_outputs(9831) <= not b or a;
    layer0_outputs(9832) <= not a;
    layer0_outputs(9833) <= not b;
    layer0_outputs(9834) <= a and not b;
    layer0_outputs(9835) <= not b or a;
    layer0_outputs(9836) <= not b;
    layer0_outputs(9837) <= b and not a;
    layer0_outputs(9838) <= not b or a;
    layer0_outputs(9839) <= not a;
    layer0_outputs(9840) <= b and not a;
    layer0_outputs(9841) <= not a;
    layer0_outputs(9842) <= a and not b;
    layer0_outputs(9843) <= not (a or b);
    layer0_outputs(9844) <= a and not b;
    layer0_outputs(9845) <= not (a xor b);
    layer0_outputs(9846) <= a xor b;
    layer0_outputs(9847) <= b;
    layer0_outputs(9848) <= a and b;
    layer0_outputs(9849) <= a xor b;
    layer0_outputs(9850) <= not (a or b);
    layer0_outputs(9851) <= a;
    layer0_outputs(9852) <= not a;
    layer0_outputs(9853) <= not (a or b);
    layer0_outputs(9854) <= a or b;
    layer0_outputs(9855) <= not (a xor b);
    layer0_outputs(9856) <= b;
    layer0_outputs(9857) <= '1';
    layer0_outputs(9858) <= '1';
    layer0_outputs(9859) <= not (a or b);
    layer0_outputs(9860) <= not (a or b);
    layer0_outputs(9861) <= a or b;
    layer0_outputs(9862) <= a;
    layer0_outputs(9863) <= not a;
    layer0_outputs(9864) <= not (a and b);
    layer0_outputs(9865) <= a or b;
    layer0_outputs(9866) <= a;
    layer0_outputs(9867) <= a and b;
    layer0_outputs(9868) <= a xor b;
    layer0_outputs(9869) <= not (a or b);
    layer0_outputs(9870) <= not (a xor b);
    layer0_outputs(9871) <= a and b;
    layer0_outputs(9872) <= not (a xor b);
    layer0_outputs(9873) <= a and not b;
    layer0_outputs(9874) <= a and not b;
    layer0_outputs(9875) <= a;
    layer0_outputs(9876) <= not (a and b);
    layer0_outputs(9877) <= a;
    layer0_outputs(9878) <= not (a or b);
    layer0_outputs(9879) <= b and not a;
    layer0_outputs(9880) <= not (a or b);
    layer0_outputs(9881) <= a;
    layer0_outputs(9882) <= not (a xor b);
    layer0_outputs(9883) <= not a;
    layer0_outputs(9884) <= a and not b;
    layer0_outputs(9885) <= not (a xor b);
    layer0_outputs(9886) <= b and not a;
    layer0_outputs(9887) <= a and b;
    layer0_outputs(9888) <= not b;
    layer0_outputs(9889) <= not (a xor b);
    layer0_outputs(9890) <= not b or a;
    layer0_outputs(9891) <= a;
    layer0_outputs(9892) <= not (a xor b);
    layer0_outputs(9893) <= not a;
    layer0_outputs(9894) <= b;
    layer0_outputs(9895) <= a xor b;
    layer0_outputs(9896) <= '0';
    layer0_outputs(9897) <= a and b;
    layer0_outputs(9898) <= not a or b;
    layer0_outputs(9899) <= '0';
    layer0_outputs(9900) <= not b;
    layer0_outputs(9901) <= a xor b;
    layer0_outputs(9902) <= not (a xor b);
    layer0_outputs(9903) <= b and not a;
    layer0_outputs(9904) <= a and not b;
    layer0_outputs(9905) <= not b;
    layer0_outputs(9906) <= not b;
    layer0_outputs(9907) <= not a;
    layer0_outputs(9908) <= a;
    layer0_outputs(9909) <= not a;
    layer0_outputs(9910) <= b;
    layer0_outputs(9911) <= not b or a;
    layer0_outputs(9912) <= not b;
    layer0_outputs(9913) <= a xor b;
    layer0_outputs(9914) <= '1';
    layer0_outputs(9915) <= '0';
    layer0_outputs(9916) <= a or b;
    layer0_outputs(9917) <= not (a or b);
    layer0_outputs(9918) <= not b;
    layer0_outputs(9919) <= b;
    layer0_outputs(9920) <= b and not a;
    layer0_outputs(9921) <= a and not b;
    layer0_outputs(9922) <= b;
    layer0_outputs(9923) <= not (a xor b);
    layer0_outputs(9924) <= not a or b;
    layer0_outputs(9925) <= not a;
    layer0_outputs(9926) <= '0';
    layer0_outputs(9927) <= a xor b;
    layer0_outputs(9928) <= not b;
    layer0_outputs(9929) <= not b;
    layer0_outputs(9930) <= b and not a;
    layer0_outputs(9931) <= not a or b;
    layer0_outputs(9932) <= not b;
    layer0_outputs(9933) <= a xor b;
    layer0_outputs(9934) <= a and not b;
    layer0_outputs(9935) <= not (a xor b);
    layer0_outputs(9936) <= b and not a;
    layer0_outputs(9937) <= '1';
    layer0_outputs(9938) <= a or b;
    layer0_outputs(9939) <= not (a xor b);
    layer0_outputs(9940) <= '1';
    layer0_outputs(9941) <= not (a xor b);
    layer0_outputs(9942) <= not a or b;
    layer0_outputs(9943) <= not (a and b);
    layer0_outputs(9944) <= b;
    layer0_outputs(9945) <= not b;
    layer0_outputs(9946) <= a xor b;
    layer0_outputs(9947) <= a;
    layer0_outputs(9948) <= not (a and b);
    layer0_outputs(9949) <= b and not a;
    layer0_outputs(9950) <= a and b;
    layer0_outputs(9951) <= b and not a;
    layer0_outputs(9952) <= a xor b;
    layer0_outputs(9953) <= not b;
    layer0_outputs(9954) <= b;
    layer0_outputs(9955) <= not a or b;
    layer0_outputs(9956) <= a and b;
    layer0_outputs(9957) <= not (a or b);
    layer0_outputs(9958) <= a xor b;
    layer0_outputs(9959) <= a and not b;
    layer0_outputs(9960) <= a xor b;
    layer0_outputs(9961) <= not (a xor b);
    layer0_outputs(9962) <= b;
    layer0_outputs(9963) <= not (a and b);
    layer0_outputs(9964) <= not b or a;
    layer0_outputs(9965) <= a or b;
    layer0_outputs(9966) <= not b or a;
    layer0_outputs(9967) <= not b or a;
    layer0_outputs(9968) <= not b;
    layer0_outputs(9969) <= '1';
    layer0_outputs(9970) <= not b;
    layer0_outputs(9971) <= a;
    layer0_outputs(9972) <= a xor b;
    layer0_outputs(9973) <= '0';
    layer0_outputs(9974) <= not b;
    layer0_outputs(9975) <= not b or a;
    layer0_outputs(9976) <= a or b;
    layer0_outputs(9977) <= not b;
    layer0_outputs(9978) <= not a or b;
    layer0_outputs(9979) <= b and not a;
    layer0_outputs(9980) <= '0';
    layer0_outputs(9981) <= a and b;
    layer0_outputs(9982) <= not a;
    layer0_outputs(9983) <= b;
    layer0_outputs(9984) <= a and b;
    layer0_outputs(9985) <= b and not a;
    layer0_outputs(9986) <= not b;
    layer0_outputs(9987) <= b and not a;
    layer0_outputs(9988) <= a or b;
    layer0_outputs(9989) <= a and not b;
    layer0_outputs(9990) <= not b;
    layer0_outputs(9991) <= not a;
    layer0_outputs(9992) <= not (a or b);
    layer0_outputs(9993) <= b;
    layer0_outputs(9994) <= b and not a;
    layer0_outputs(9995) <= a xor b;
    layer0_outputs(9996) <= not b or a;
    layer0_outputs(9997) <= a xor b;
    layer0_outputs(9998) <= not (a xor b);
    layer0_outputs(9999) <= a and not b;
    layer0_outputs(10000) <= b and not a;
    layer0_outputs(10001) <= not a or b;
    layer0_outputs(10002) <= not a;
    layer0_outputs(10003) <= not b;
    layer0_outputs(10004) <= not (a and b);
    layer0_outputs(10005) <= not (a and b);
    layer0_outputs(10006) <= a;
    layer0_outputs(10007) <= a or b;
    layer0_outputs(10008) <= not b or a;
    layer0_outputs(10009) <= a and not b;
    layer0_outputs(10010) <= not (a or b);
    layer0_outputs(10011) <= not b;
    layer0_outputs(10012) <= a;
    layer0_outputs(10013) <= a xor b;
    layer0_outputs(10014) <= b and not a;
    layer0_outputs(10015) <= b;
    layer0_outputs(10016) <= a xor b;
    layer0_outputs(10017) <= not (a or b);
    layer0_outputs(10018) <= not b;
    layer0_outputs(10019) <= a or b;
    layer0_outputs(10020) <= a xor b;
    layer0_outputs(10021) <= not b or a;
    layer0_outputs(10022) <= not a;
    layer0_outputs(10023) <= not b;
    layer0_outputs(10024) <= not a;
    layer0_outputs(10025) <= a and b;
    layer0_outputs(10026) <= b and not a;
    layer0_outputs(10027) <= b;
    layer0_outputs(10028) <= a and b;
    layer0_outputs(10029) <= not (a or b);
    layer0_outputs(10030) <= not a;
    layer0_outputs(10031) <= not b;
    layer0_outputs(10032) <= a;
    layer0_outputs(10033) <= a and b;
    layer0_outputs(10034) <= a or b;
    layer0_outputs(10035) <= not (a xor b);
    layer0_outputs(10036) <= not b or a;
    layer0_outputs(10037) <= not a;
    layer0_outputs(10038) <= not a;
    layer0_outputs(10039) <= '1';
    layer0_outputs(10040) <= b;
    layer0_outputs(10041) <= a or b;
    layer0_outputs(10042) <= a;
    layer0_outputs(10043) <= not (a and b);
    layer0_outputs(10044) <= not a;
    layer0_outputs(10045) <= not a;
    layer0_outputs(10046) <= a or b;
    layer0_outputs(10047) <= not a or b;
    layer0_outputs(10048) <= '0';
    layer0_outputs(10049) <= not (a xor b);
    layer0_outputs(10050) <= a or b;
    layer0_outputs(10051) <= '1';
    layer0_outputs(10052) <= not (a xor b);
    layer0_outputs(10053) <= not b;
    layer0_outputs(10054) <= not a;
    layer0_outputs(10055) <= a or b;
    layer0_outputs(10056) <= b;
    layer0_outputs(10057) <= b and not a;
    layer0_outputs(10058) <= a and not b;
    layer0_outputs(10059) <= a or b;
    layer0_outputs(10060) <= '0';
    layer0_outputs(10061) <= not (a or b);
    layer0_outputs(10062) <= a;
    layer0_outputs(10063) <= a or b;
    layer0_outputs(10064) <= not a or b;
    layer0_outputs(10065) <= a and not b;
    layer0_outputs(10066) <= a and not b;
    layer0_outputs(10067) <= '0';
    layer0_outputs(10068) <= not b;
    layer0_outputs(10069) <= not (a xor b);
    layer0_outputs(10070) <= not a or b;
    layer0_outputs(10071) <= not (a xor b);
    layer0_outputs(10072) <= '1';
    layer0_outputs(10073) <= not b;
    layer0_outputs(10074) <= a and not b;
    layer0_outputs(10075) <= not (a or b);
    layer0_outputs(10076) <= not (a and b);
    layer0_outputs(10077) <= not b;
    layer0_outputs(10078) <= a and not b;
    layer0_outputs(10079) <= not (a or b);
    layer0_outputs(10080) <= a and not b;
    layer0_outputs(10081) <= not b;
    layer0_outputs(10082) <= not b;
    layer0_outputs(10083) <= '0';
    layer0_outputs(10084) <= '0';
    layer0_outputs(10085) <= b;
    layer0_outputs(10086) <= not (a or b);
    layer0_outputs(10087) <= a;
    layer0_outputs(10088) <= not (a or b);
    layer0_outputs(10089) <= not a or b;
    layer0_outputs(10090) <= not b or a;
    layer0_outputs(10091) <= b and not a;
    layer0_outputs(10092) <= not (a and b);
    layer0_outputs(10093) <= a or b;
    layer0_outputs(10094) <= '1';
    layer0_outputs(10095) <= not b or a;
    layer0_outputs(10096) <= not (a or b);
    layer0_outputs(10097) <= a or b;
    layer0_outputs(10098) <= not (a or b);
    layer0_outputs(10099) <= not b or a;
    layer0_outputs(10100) <= not b or a;
    layer0_outputs(10101) <= '1';
    layer0_outputs(10102) <= b and not a;
    layer0_outputs(10103) <= not a or b;
    layer0_outputs(10104) <= not b;
    layer0_outputs(10105) <= not (a or b);
    layer0_outputs(10106) <= not (a and b);
    layer0_outputs(10107) <= not (a and b);
    layer0_outputs(10108) <= b;
    layer0_outputs(10109) <= not a;
    layer0_outputs(10110) <= '1';
    layer0_outputs(10111) <= '1';
    layer0_outputs(10112) <= b;
    layer0_outputs(10113) <= not (a xor b);
    layer0_outputs(10114) <= a;
    layer0_outputs(10115) <= not (a xor b);
    layer0_outputs(10116) <= not b or a;
    layer0_outputs(10117) <= not b;
    layer0_outputs(10118) <= not a or b;
    layer0_outputs(10119) <= not (a or b);
    layer0_outputs(10120) <= a;
    layer0_outputs(10121) <= a and b;
    layer0_outputs(10122) <= '0';
    layer0_outputs(10123) <= not a or b;
    layer0_outputs(10124) <= a and not b;
    layer0_outputs(10125) <= not (a xor b);
    layer0_outputs(10126) <= a and b;
    layer0_outputs(10127) <= a;
    layer0_outputs(10128) <= not a;
    layer0_outputs(10129) <= a;
    layer0_outputs(10130) <= a or b;
    layer0_outputs(10131) <= not a or b;
    layer0_outputs(10132) <= a or b;
    layer0_outputs(10133) <= a;
    layer0_outputs(10134) <= a and not b;
    layer0_outputs(10135) <= not b or a;
    layer0_outputs(10136) <= not (a or b);
    layer0_outputs(10137) <= not (a xor b);
    layer0_outputs(10138) <= b;
    layer0_outputs(10139) <= not b;
    layer0_outputs(10140) <= b and not a;
    layer0_outputs(10141) <= not a or b;
    layer0_outputs(10142) <= a or b;
    layer0_outputs(10143) <= a or b;
    layer0_outputs(10144) <= not b;
    layer0_outputs(10145) <= b;
    layer0_outputs(10146) <= b;
    layer0_outputs(10147) <= not b or a;
    layer0_outputs(10148) <= not (a or b);
    layer0_outputs(10149) <= a and b;
    layer0_outputs(10150) <= not (a or b);
    layer0_outputs(10151) <= not a or b;
    layer0_outputs(10152) <= b and not a;
    layer0_outputs(10153) <= not (a or b);
    layer0_outputs(10154) <= a;
    layer0_outputs(10155) <= not b;
    layer0_outputs(10156) <= a or b;
    layer0_outputs(10157) <= b and not a;
    layer0_outputs(10158) <= a xor b;
    layer0_outputs(10159) <= a xor b;
    layer0_outputs(10160) <= a xor b;
    layer0_outputs(10161) <= b and not a;
    layer0_outputs(10162) <= not a;
    layer0_outputs(10163) <= not a or b;
    layer0_outputs(10164) <= a;
    layer0_outputs(10165) <= a and b;
    layer0_outputs(10166) <= not (a or b);
    layer0_outputs(10167) <= not (a xor b);
    layer0_outputs(10168) <= not a or b;
    layer0_outputs(10169) <= not b;
    layer0_outputs(10170) <= a and b;
    layer0_outputs(10171) <= not b or a;
    layer0_outputs(10172) <= b;
    layer0_outputs(10173) <= not (a or b);
    layer0_outputs(10174) <= not (a xor b);
    layer0_outputs(10175) <= not b;
    layer0_outputs(10176) <= '0';
    layer0_outputs(10177) <= a and b;
    layer0_outputs(10178) <= a or b;
    layer0_outputs(10179) <= not (a or b);
    layer0_outputs(10180) <= a or b;
    layer0_outputs(10181) <= not b;
    layer0_outputs(10182) <= not a;
    layer0_outputs(10183) <= a or b;
    layer0_outputs(10184) <= b and not a;
    layer0_outputs(10185) <= '0';
    layer0_outputs(10186) <= not (a xor b);
    layer0_outputs(10187) <= not (a and b);
    layer0_outputs(10188) <= b;
    layer0_outputs(10189) <= a;
    layer0_outputs(10190) <= not b;
    layer0_outputs(10191) <= not b;
    layer0_outputs(10192) <= not b;
    layer0_outputs(10193) <= not b or a;
    layer0_outputs(10194) <= b and not a;
    layer0_outputs(10195) <= a and not b;
    layer0_outputs(10196) <= b;
    layer0_outputs(10197) <= not a or b;
    layer0_outputs(10198) <= not a;
    layer0_outputs(10199) <= not b or a;
    layer0_outputs(10200) <= b and not a;
    layer0_outputs(10201) <= not a or b;
    layer0_outputs(10202) <= a xor b;
    layer0_outputs(10203) <= not (a and b);
    layer0_outputs(10204) <= '1';
    layer0_outputs(10205) <= b;
    layer0_outputs(10206) <= not b;
    layer0_outputs(10207) <= b and not a;
    layer0_outputs(10208) <= not a;
    layer0_outputs(10209) <= not (a or b);
    layer0_outputs(10210) <= not b or a;
    layer0_outputs(10211) <= not b;
    layer0_outputs(10212) <= not a;
    layer0_outputs(10213) <= not a;
    layer0_outputs(10214) <= not b or a;
    layer0_outputs(10215) <= not (a or b);
    layer0_outputs(10216) <= not b;
    layer0_outputs(10217) <= '0';
    layer0_outputs(10218) <= not b;
    layer0_outputs(10219) <= a xor b;
    layer0_outputs(10220) <= not (a or b);
    layer0_outputs(10221) <= not (a or b);
    layer0_outputs(10222) <= a xor b;
    layer0_outputs(10223) <= '0';
    layer0_outputs(10224) <= a and b;
    layer0_outputs(10225) <= a or b;
    layer0_outputs(10226) <= not (a xor b);
    layer0_outputs(10227) <= a;
    layer0_outputs(10228) <= a or b;
    layer0_outputs(10229) <= a and b;
    layer0_outputs(10230) <= not (a or b);
    layer0_outputs(10231) <= a and not b;
    layer0_outputs(10232) <= not a;
    layer0_outputs(10233) <= a xor b;
    layer0_outputs(10234) <= not (a or b);
    layer0_outputs(10235) <= b;
    layer0_outputs(10236) <= a and b;
    layer0_outputs(10237) <= '1';
    layer0_outputs(10238) <= not (a xor b);
    layer0_outputs(10239) <= b;
    layer1_outputs(0) <= a;
    layer1_outputs(1) <= a and not b;
    layer1_outputs(2) <= a;
    layer1_outputs(3) <= a;
    layer1_outputs(4) <= not (a or b);
    layer1_outputs(5) <= a and not b;
    layer1_outputs(6) <= not (a or b);
    layer1_outputs(7) <= not b or a;
    layer1_outputs(8) <= b;
    layer1_outputs(9) <= a and b;
    layer1_outputs(10) <= not a or b;
    layer1_outputs(11) <= a;
    layer1_outputs(12) <= a and b;
    layer1_outputs(13) <= a and not b;
    layer1_outputs(14) <= '0';
    layer1_outputs(15) <= b;
    layer1_outputs(16) <= a or b;
    layer1_outputs(17) <= not b;
    layer1_outputs(18) <= a or b;
    layer1_outputs(19) <= '1';
    layer1_outputs(20) <= b;
    layer1_outputs(21) <= not b or a;
    layer1_outputs(22) <= not a;
    layer1_outputs(23) <= not (a and b);
    layer1_outputs(24) <= not (a or b);
    layer1_outputs(25) <= a xor b;
    layer1_outputs(26) <= b;
    layer1_outputs(27) <= not (a and b);
    layer1_outputs(28) <= a;
    layer1_outputs(29) <= not (a and b);
    layer1_outputs(30) <= not (a or b);
    layer1_outputs(31) <= b and not a;
    layer1_outputs(32) <= a or b;
    layer1_outputs(33) <= a and b;
    layer1_outputs(34) <= b;
    layer1_outputs(35) <= a xor b;
    layer1_outputs(36) <= '1';
    layer1_outputs(37) <= not a;
    layer1_outputs(38) <= b;
    layer1_outputs(39) <= b;
    layer1_outputs(40) <= not (a and b);
    layer1_outputs(41) <= not (a and b);
    layer1_outputs(42) <= not (a and b);
    layer1_outputs(43) <= not a;
    layer1_outputs(44) <= '0';
    layer1_outputs(45) <= a or b;
    layer1_outputs(46) <= a xor b;
    layer1_outputs(47) <= not a or b;
    layer1_outputs(48) <= not b;
    layer1_outputs(49) <= b;
    layer1_outputs(50) <= a and not b;
    layer1_outputs(51) <= a xor b;
    layer1_outputs(52) <= b and not a;
    layer1_outputs(53) <= not a;
    layer1_outputs(54) <= b;
    layer1_outputs(55) <= not b or a;
    layer1_outputs(56) <= '0';
    layer1_outputs(57) <= not b;
    layer1_outputs(58) <= a or b;
    layer1_outputs(59) <= a and b;
    layer1_outputs(60) <= b;
    layer1_outputs(61) <= not (a xor b);
    layer1_outputs(62) <= not a;
    layer1_outputs(63) <= a and b;
    layer1_outputs(64) <= b;
    layer1_outputs(65) <= not b or a;
    layer1_outputs(66) <= '0';
    layer1_outputs(67) <= not b or a;
    layer1_outputs(68) <= a and not b;
    layer1_outputs(69) <= a and not b;
    layer1_outputs(70) <= not a or b;
    layer1_outputs(71) <= '1';
    layer1_outputs(72) <= not a;
    layer1_outputs(73) <= not (a or b);
    layer1_outputs(74) <= a;
    layer1_outputs(75) <= not (a and b);
    layer1_outputs(76) <= a and not b;
    layer1_outputs(77) <= b;
    layer1_outputs(78) <= a or b;
    layer1_outputs(79) <= a and b;
    layer1_outputs(80) <= a and b;
    layer1_outputs(81) <= a;
    layer1_outputs(82) <= a;
    layer1_outputs(83) <= not (a or b);
    layer1_outputs(84) <= a and not b;
    layer1_outputs(85) <= b and not a;
    layer1_outputs(86) <= '0';
    layer1_outputs(87) <= not b;
    layer1_outputs(88) <= not b;
    layer1_outputs(89) <= not (a xor b);
    layer1_outputs(90) <= '0';
    layer1_outputs(91) <= b;
    layer1_outputs(92) <= a and b;
    layer1_outputs(93) <= not (a or b);
    layer1_outputs(94) <= not a or b;
    layer1_outputs(95) <= b and not a;
    layer1_outputs(96) <= not b;
    layer1_outputs(97) <= not a;
    layer1_outputs(98) <= b;
    layer1_outputs(99) <= not a;
    layer1_outputs(100) <= not a or b;
    layer1_outputs(101) <= '0';
    layer1_outputs(102) <= '1';
    layer1_outputs(103) <= a xor b;
    layer1_outputs(104) <= not b;
    layer1_outputs(105) <= b;
    layer1_outputs(106) <= not a;
    layer1_outputs(107) <= '1';
    layer1_outputs(108) <= a and b;
    layer1_outputs(109) <= not (a xor b);
    layer1_outputs(110) <= not (a or b);
    layer1_outputs(111) <= not (a and b);
    layer1_outputs(112) <= '0';
    layer1_outputs(113) <= b;
    layer1_outputs(114) <= b;
    layer1_outputs(115) <= a xor b;
    layer1_outputs(116) <= b and not a;
    layer1_outputs(117) <= a or b;
    layer1_outputs(118) <= a and b;
    layer1_outputs(119) <= not a;
    layer1_outputs(120) <= b and not a;
    layer1_outputs(121) <= a;
    layer1_outputs(122) <= '1';
    layer1_outputs(123) <= a and b;
    layer1_outputs(124) <= not (a or b);
    layer1_outputs(125) <= b;
    layer1_outputs(126) <= b;
    layer1_outputs(127) <= not a;
    layer1_outputs(128) <= '0';
    layer1_outputs(129) <= not a;
    layer1_outputs(130) <= b and not a;
    layer1_outputs(131) <= '1';
    layer1_outputs(132) <= a xor b;
    layer1_outputs(133) <= '0';
    layer1_outputs(134) <= b;
    layer1_outputs(135) <= '0';
    layer1_outputs(136) <= not (a or b);
    layer1_outputs(137) <= a and b;
    layer1_outputs(138) <= not b;
    layer1_outputs(139) <= b and not a;
    layer1_outputs(140) <= b and not a;
    layer1_outputs(141) <= not (a or b);
    layer1_outputs(142) <= not (a or b);
    layer1_outputs(143) <= a and not b;
    layer1_outputs(144) <= a and not b;
    layer1_outputs(145) <= a and b;
    layer1_outputs(146) <= b;
    layer1_outputs(147) <= a;
    layer1_outputs(148) <= a or b;
    layer1_outputs(149) <= not (a xor b);
    layer1_outputs(150) <= a and b;
    layer1_outputs(151) <= not (a and b);
    layer1_outputs(152) <= b;
    layer1_outputs(153) <= b;
    layer1_outputs(154) <= '0';
    layer1_outputs(155) <= a or b;
    layer1_outputs(156) <= a;
    layer1_outputs(157) <= not a or b;
    layer1_outputs(158) <= b;
    layer1_outputs(159) <= a or b;
    layer1_outputs(160) <= b and not a;
    layer1_outputs(161) <= b and not a;
    layer1_outputs(162) <= b and not a;
    layer1_outputs(163) <= not a;
    layer1_outputs(164) <= not a or b;
    layer1_outputs(165) <= not a;
    layer1_outputs(166) <= a and b;
    layer1_outputs(167) <= '0';
    layer1_outputs(168) <= not b or a;
    layer1_outputs(169) <= not (a and b);
    layer1_outputs(170) <= a and b;
    layer1_outputs(171) <= a and not b;
    layer1_outputs(172) <= b and not a;
    layer1_outputs(173) <= a xor b;
    layer1_outputs(174) <= b and not a;
    layer1_outputs(175) <= not a;
    layer1_outputs(176) <= a and b;
    layer1_outputs(177) <= b;
    layer1_outputs(178) <= a xor b;
    layer1_outputs(179) <= b;
    layer1_outputs(180) <= not (a or b);
    layer1_outputs(181) <= b;
    layer1_outputs(182) <= not b or a;
    layer1_outputs(183) <= a or b;
    layer1_outputs(184) <= not b or a;
    layer1_outputs(185) <= not b;
    layer1_outputs(186) <= a;
    layer1_outputs(187) <= a;
    layer1_outputs(188) <= not b;
    layer1_outputs(189) <= not b;
    layer1_outputs(190) <= not a;
    layer1_outputs(191) <= not (a xor b);
    layer1_outputs(192) <= a or b;
    layer1_outputs(193) <= a xor b;
    layer1_outputs(194) <= not a or b;
    layer1_outputs(195) <= '0';
    layer1_outputs(196) <= a and b;
    layer1_outputs(197) <= a and not b;
    layer1_outputs(198) <= not b;
    layer1_outputs(199) <= a and b;
    layer1_outputs(200) <= not (a xor b);
    layer1_outputs(201) <= not a;
    layer1_outputs(202) <= not b;
    layer1_outputs(203) <= a or b;
    layer1_outputs(204) <= a;
    layer1_outputs(205) <= not a or b;
    layer1_outputs(206) <= b;
    layer1_outputs(207) <= not (a and b);
    layer1_outputs(208) <= '1';
    layer1_outputs(209) <= not (a and b);
    layer1_outputs(210) <= a or b;
    layer1_outputs(211) <= not (a and b);
    layer1_outputs(212) <= b;
    layer1_outputs(213) <= not b or a;
    layer1_outputs(214) <= not a or b;
    layer1_outputs(215) <= not a;
    layer1_outputs(216) <= not a;
    layer1_outputs(217) <= a;
    layer1_outputs(218) <= b and not a;
    layer1_outputs(219) <= not b;
    layer1_outputs(220) <= a;
    layer1_outputs(221) <= a and b;
    layer1_outputs(222) <= not b;
    layer1_outputs(223) <= not b or a;
    layer1_outputs(224) <= b and not a;
    layer1_outputs(225) <= not a;
    layer1_outputs(226) <= a;
    layer1_outputs(227) <= a;
    layer1_outputs(228) <= a;
    layer1_outputs(229) <= not a;
    layer1_outputs(230) <= b;
    layer1_outputs(231) <= b and not a;
    layer1_outputs(232) <= not a;
    layer1_outputs(233) <= not a;
    layer1_outputs(234) <= a;
    layer1_outputs(235) <= not a;
    layer1_outputs(236) <= not b or a;
    layer1_outputs(237) <= a and not b;
    layer1_outputs(238) <= not b or a;
    layer1_outputs(239) <= '1';
    layer1_outputs(240) <= '0';
    layer1_outputs(241) <= b;
    layer1_outputs(242) <= a or b;
    layer1_outputs(243) <= a and not b;
    layer1_outputs(244) <= not a or b;
    layer1_outputs(245) <= a xor b;
    layer1_outputs(246) <= '1';
    layer1_outputs(247) <= not a;
    layer1_outputs(248) <= '1';
    layer1_outputs(249) <= a xor b;
    layer1_outputs(250) <= '0';
    layer1_outputs(251) <= not (a xor b);
    layer1_outputs(252) <= a xor b;
    layer1_outputs(253) <= not b;
    layer1_outputs(254) <= '0';
    layer1_outputs(255) <= a and not b;
    layer1_outputs(256) <= a or b;
    layer1_outputs(257) <= b;
    layer1_outputs(258) <= a or b;
    layer1_outputs(259) <= b and not a;
    layer1_outputs(260) <= '1';
    layer1_outputs(261) <= not a;
    layer1_outputs(262) <= not b or a;
    layer1_outputs(263) <= b and not a;
    layer1_outputs(264) <= a;
    layer1_outputs(265) <= a or b;
    layer1_outputs(266) <= b and not a;
    layer1_outputs(267) <= a;
    layer1_outputs(268) <= a and not b;
    layer1_outputs(269) <= not a or b;
    layer1_outputs(270) <= '0';
    layer1_outputs(271) <= not (a or b);
    layer1_outputs(272) <= b and not a;
    layer1_outputs(273) <= not b or a;
    layer1_outputs(274) <= '1';
    layer1_outputs(275) <= '1';
    layer1_outputs(276) <= a and not b;
    layer1_outputs(277) <= not (a or b);
    layer1_outputs(278) <= a and not b;
    layer1_outputs(279) <= a and not b;
    layer1_outputs(280) <= a and not b;
    layer1_outputs(281) <= a or b;
    layer1_outputs(282) <= a and b;
    layer1_outputs(283) <= not b;
    layer1_outputs(284) <= '0';
    layer1_outputs(285) <= not b;
    layer1_outputs(286) <= not a;
    layer1_outputs(287) <= b;
    layer1_outputs(288) <= not b;
    layer1_outputs(289) <= not (a or b);
    layer1_outputs(290) <= not (a xor b);
    layer1_outputs(291) <= a;
    layer1_outputs(292) <= not b or a;
    layer1_outputs(293) <= a or b;
    layer1_outputs(294) <= not a or b;
    layer1_outputs(295) <= b and not a;
    layer1_outputs(296) <= not (a or b);
    layer1_outputs(297) <= '1';
    layer1_outputs(298) <= not (a and b);
    layer1_outputs(299) <= b;
    layer1_outputs(300) <= not (a or b);
    layer1_outputs(301) <= '0';
    layer1_outputs(302) <= a and not b;
    layer1_outputs(303) <= not (a xor b);
    layer1_outputs(304) <= not (a or b);
    layer1_outputs(305) <= not a;
    layer1_outputs(306) <= b;
    layer1_outputs(307) <= not b or a;
    layer1_outputs(308) <= not b;
    layer1_outputs(309) <= not (a or b);
    layer1_outputs(310) <= not (a or b);
    layer1_outputs(311) <= not b or a;
    layer1_outputs(312) <= not b or a;
    layer1_outputs(313) <= b;
    layer1_outputs(314) <= not b;
    layer1_outputs(315) <= not b;
    layer1_outputs(316) <= not b;
    layer1_outputs(317) <= a and b;
    layer1_outputs(318) <= a and b;
    layer1_outputs(319) <= not a or b;
    layer1_outputs(320) <= not (a or b);
    layer1_outputs(321) <= not a or b;
    layer1_outputs(322) <= '0';
    layer1_outputs(323) <= not b;
    layer1_outputs(324) <= not a;
    layer1_outputs(325) <= a;
    layer1_outputs(326) <= b and not a;
    layer1_outputs(327) <= not a or b;
    layer1_outputs(328) <= a;
    layer1_outputs(329) <= not (a and b);
    layer1_outputs(330) <= b and not a;
    layer1_outputs(331) <= b;
    layer1_outputs(332) <= a;
    layer1_outputs(333) <= not b;
    layer1_outputs(334) <= b;
    layer1_outputs(335) <= b and not a;
    layer1_outputs(336) <= b;
    layer1_outputs(337) <= not b or a;
    layer1_outputs(338) <= not (a and b);
    layer1_outputs(339) <= '0';
    layer1_outputs(340) <= not b;
    layer1_outputs(341) <= a;
    layer1_outputs(342) <= not a;
    layer1_outputs(343) <= a and not b;
    layer1_outputs(344) <= b;
    layer1_outputs(345) <= b;
    layer1_outputs(346) <= a and b;
    layer1_outputs(347) <= not a;
    layer1_outputs(348) <= not b;
    layer1_outputs(349) <= not b;
    layer1_outputs(350) <= not (a or b);
    layer1_outputs(351) <= a and not b;
    layer1_outputs(352) <= a and not b;
    layer1_outputs(353) <= not (a or b);
    layer1_outputs(354) <= a or b;
    layer1_outputs(355) <= a or b;
    layer1_outputs(356) <= not a;
    layer1_outputs(357) <= a and not b;
    layer1_outputs(358) <= not (a xor b);
    layer1_outputs(359) <= b;
    layer1_outputs(360) <= not (a and b);
    layer1_outputs(361) <= not a;
    layer1_outputs(362) <= b;
    layer1_outputs(363) <= not a;
    layer1_outputs(364) <= a or b;
    layer1_outputs(365) <= not b or a;
    layer1_outputs(366) <= b and not a;
    layer1_outputs(367) <= not b or a;
    layer1_outputs(368) <= b;
    layer1_outputs(369) <= a xor b;
    layer1_outputs(370) <= not (a or b);
    layer1_outputs(371) <= a;
    layer1_outputs(372) <= not b or a;
    layer1_outputs(373) <= a;
    layer1_outputs(374) <= a or b;
    layer1_outputs(375) <= '1';
    layer1_outputs(376) <= '0';
    layer1_outputs(377) <= not a;
    layer1_outputs(378) <= not a;
    layer1_outputs(379) <= b and not a;
    layer1_outputs(380) <= a and b;
    layer1_outputs(381) <= not a;
    layer1_outputs(382) <= not (a or b);
    layer1_outputs(383) <= not b or a;
    layer1_outputs(384) <= not a or b;
    layer1_outputs(385) <= not (a and b);
    layer1_outputs(386) <= not (a or b);
    layer1_outputs(387) <= b and not a;
    layer1_outputs(388) <= '1';
    layer1_outputs(389) <= not a or b;
    layer1_outputs(390) <= not a or b;
    layer1_outputs(391) <= a or b;
    layer1_outputs(392) <= not b;
    layer1_outputs(393) <= a and not b;
    layer1_outputs(394) <= not b;
    layer1_outputs(395) <= b and not a;
    layer1_outputs(396) <= not b;
    layer1_outputs(397) <= not b or a;
    layer1_outputs(398) <= not (a or b);
    layer1_outputs(399) <= not (a xor b);
    layer1_outputs(400) <= not (a and b);
    layer1_outputs(401) <= not b or a;
    layer1_outputs(402) <= not a or b;
    layer1_outputs(403) <= not (a xor b);
    layer1_outputs(404) <= a or b;
    layer1_outputs(405) <= not (a or b);
    layer1_outputs(406) <= not a or b;
    layer1_outputs(407) <= not a or b;
    layer1_outputs(408) <= not b or a;
    layer1_outputs(409) <= a;
    layer1_outputs(410) <= b and not a;
    layer1_outputs(411) <= a;
    layer1_outputs(412) <= not a;
    layer1_outputs(413) <= not a;
    layer1_outputs(414) <= a and b;
    layer1_outputs(415) <= a and not b;
    layer1_outputs(416) <= a or b;
    layer1_outputs(417) <= b;
    layer1_outputs(418) <= not a;
    layer1_outputs(419) <= b and not a;
    layer1_outputs(420) <= a;
    layer1_outputs(421) <= a and b;
    layer1_outputs(422) <= a and b;
    layer1_outputs(423) <= not (a xor b);
    layer1_outputs(424) <= '1';
    layer1_outputs(425) <= a;
    layer1_outputs(426) <= a xor b;
    layer1_outputs(427) <= '1';
    layer1_outputs(428) <= a xor b;
    layer1_outputs(429) <= not a;
    layer1_outputs(430) <= not (a or b);
    layer1_outputs(431) <= not b;
    layer1_outputs(432) <= '0';
    layer1_outputs(433) <= b;
    layer1_outputs(434) <= not (a or b);
    layer1_outputs(435) <= b;
    layer1_outputs(436) <= not (a or b);
    layer1_outputs(437) <= not b or a;
    layer1_outputs(438) <= b and not a;
    layer1_outputs(439) <= not a or b;
    layer1_outputs(440) <= not b or a;
    layer1_outputs(441) <= not a;
    layer1_outputs(442) <= a or b;
    layer1_outputs(443) <= a;
    layer1_outputs(444) <= not a or b;
    layer1_outputs(445) <= a and b;
    layer1_outputs(446) <= b and not a;
    layer1_outputs(447) <= b and not a;
    layer1_outputs(448) <= not a or b;
    layer1_outputs(449) <= '0';
    layer1_outputs(450) <= a and not b;
    layer1_outputs(451) <= '0';
    layer1_outputs(452) <= '1';
    layer1_outputs(453) <= not (a xor b);
    layer1_outputs(454) <= '1';
    layer1_outputs(455) <= a or b;
    layer1_outputs(456) <= not a;
    layer1_outputs(457) <= b and not a;
    layer1_outputs(458) <= not a;
    layer1_outputs(459) <= not (a or b);
    layer1_outputs(460) <= b;
    layer1_outputs(461) <= '1';
    layer1_outputs(462) <= b and not a;
    layer1_outputs(463) <= a;
    layer1_outputs(464) <= a;
    layer1_outputs(465) <= not (a xor b);
    layer1_outputs(466) <= not b or a;
    layer1_outputs(467) <= b and not a;
    layer1_outputs(468) <= not (a xor b);
    layer1_outputs(469) <= not (a and b);
    layer1_outputs(470) <= b and not a;
    layer1_outputs(471) <= not a or b;
    layer1_outputs(472) <= not a;
    layer1_outputs(473) <= a and not b;
    layer1_outputs(474) <= '0';
    layer1_outputs(475) <= '1';
    layer1_outputs(476) <= not a;
    layer1_outputs(477) <= b;
    layer1_outputs(478) <= not a;
    layer1_outputs(479) <= not b;
    layer1_outputs(480) <= not (a or b);
    layer1_outputs(481) <= a and not b;
    layer1_outputs(482) <= not b;
    layer1_outputs(483) <= b;
    layer1_outputs(484) <= not (a and b);
    layer1_outputs(485) <= not (a and b);
    layer1_outputs(486) <= a and b;
    layer1_outputs(487) <= not b;
    layer1_outputs(488) <= '1';
    layer1_outputs(489) <= a;
    layer1_outputs(490) <= b and not a;
    layer1_outputs(491) <= b;
    layer1_outputs(492) <= a xor b;
    layer1_outputs(493) <= b;
    layer1_outputs(494) <= b and not a;
    layer1_outputs(495) <= not a or b;
    layer1_outputs(496) <= not (a and b);
    layer1_outputs(497) <= b;
    layer1_outputs(498) <= a;
    layer1_outputs(499) <= not (a and b);
    layer1_outputs(500) <= a and not b;
    layer1_outputs(501) <= a and not b;
    layer1_outputs(502) <= a xor b;
    layer1_outputs(503) <= not (a or b);
    layer1_outputs(504) <= not (a or b);
    layer1_outputs(505) <= a and not b;
    layer1_outputs(506) <= a or b;
    layer1_outputs(507) <= a and b;
    layer1_outputs(508) <= a;
    layer1_outputs(509) <= b;
    layer1_outputs(510) <= not a;
    layer1_outputs(511) <= a;
    layer1_outputs(512) <= a or b;
    layer1_outputs(513) <= not a;
    layer1_outputs(514) <= b;
    layer1_outputs(515) <= a xor b;
    layer1_outputs(516) <= not b or a;
    layer1_outputs(517) <= not b or a;
    layer1_outputs(518) <= a;
    layer1_outputs(519) <= not a or b;
    layer1_outputs(520) <= '0';
    layer1_outputs(521) <= not b;
    layer1_outputs(522) <= a;
    layer1_outputs(523) <= not a or b;
    layer1_outputs(524) <= '0';
    layer1_outputs(525) <= not (a and b);
    layer1_outputs(526) <= a;
    layer1_outputs(527) <= '0';
    layer1_outputs(528) <= a xor b;
    layer1_outputs(529) <= '0';
    layer1_outputs(530) <= '1';
    layer1_outputs(531) <= b;
    layer1_outputs(532) <= '0';
    layer1_outputs(533) <= not a;
    layer1_outputs(534) <= not a or b;
    layer1_outputs(535) <= not a;
    layer1_outputs(536) <= not b;
    layer1_outputs(537) <= a;
    layer1_outputs(538) <= not (a and b);
    layer1_outputs(539) <= a or b;
    layer1_outputs(540) <= not (a xor b);
    layer1_outputs(541) <= b and not a;
    layer1_outputs(542) <= not b;
    layer1_outputs(543) <= not (a xor b);
    layer1_outputs(544) <= b;
    layer1_outputs(545) <= not b or a;
    layer1_outputs(546) <= not a;
    layer1_outputs(547) <= a or b;
    layer1_outputs(548) <= a and not b;
    layer1_outputs(549) <= '0';
    layer1_outputs(550) <= '0';
    layer1_outputs(551) <= not (a and b);
    layer1_outputs(552) <= a or b;
    layer1_outputs(553) <= a or b;
    layer1_outputs(554) <= not a or b;
    layer1_outputs(555) <= '0';
    layer1_outputs(556) <= a;
    layer1_outputs(557) <= not (a or b);
    layer1_outputs(558) <= not b or a;
    layer1_outputs(559) <= not a or b;
    layer1_outputs(560) <= '0';
    layer1_outputs(561) <= '0';
    layer1_outputs(562) <= not a;
    layer1_outputs(563) <= not (a or b);
    layer1_outputs(564) <= not a;
    layer1_outputs(565) <= b and not a;
    layer1_outputs(566) <= not a or b;
    layer1_outputs(567) <= a and not b;
    layer1_outputs(568) <= not b;
    layer1_outputs(569) <= not b;
    layer1_outputs(570) <= not b or a;
    layer1_outputs(571) <= not (a or b);
    layer1_outputs(572) <= a or b;
    layer1_outputs(573) <= not b or a;
    layer1_outputs(574) <= a or b;
    layer1_outputs(575) <= a or b;
    layer1_outputs(576) <= not b or a;
    layer1_outputs(577) <= b;
    layer1_outputs(578) <= not b or a;
    layer1_outputs(579) <= not b;
    layer1_outputs(580) <= b and not a;
    layer1_outputs(581) <= a or b;
    layer1_outputs(582) <= not a or b;
    layer1_outputs(583) <= a;
    layer1_outputs(584) <= '1';
    layer1_outputs(585) <= not (a xor b);
    layer1_outputs(586) <= not b or a;
    layer1_outputs(587) <= not a;
    layer1_outputs(588) <= a or b;
    layer1_outputs(589) <= a or b;
    layer1_outputs(590) <= a and not b;
    layer1_outputs(591) <= not (a xor b);
    layer1_outputs(592) <= a or b;
    layer1_outputs(593) <= not a or b;
    layer1_outputs(594) <= '0';
    layer1_outputs(595) <= '0';
    layer1_outputs(596) <= a and not b;
    layer1_outputs(597) <= a;
    layer1_outputs(598) <= not a or b;
    layer1_outputs(599) <= b;
    layer1_outputs(600) <= '1';
    layer1_outputs(601) <= not b or a;
    layer1_outputs(602) <= b and not a;
    layer1_outputs(603) <= not (a or b);
    layer1_outputs(604) <= a;
    layer1_outputs(605) <= '0';
    layer1_outputs(606) <= b;
    layer1_outputs(607) <= a xor b;
    layer1_outputs(608) <= a and not b;
    layer1_outputs(609) <= not (a or b);
    layer1_outputs(610) <= not b;
    layer1_outputs(611) <= a and not b;
    layer1_outputs(612) <= a and not b;
    layer1_outputs(613) <= '0';
    layer1_outputs(614) <= a and not b;
    layer1_outputs(615) <= a;
    layer1_outputs(616) <= a or b;
    layer1_outputs(617) <= a and b;
    layer1_outputs(618) <= a and not b;
    layer1_outputs(619) <= a and b;
    layer1_outputs(620) <= not a;
    layer1_outputs(621) <= '1';
    layer1_outputs(622) <= a and not b;
    layer1_outputs(623) <= not b or a;
    layer1_outputs(624) <= not b or a;
    layer1_outputs(625) <= b;
    layer1_outputs(626) <= not (a and b);
    layer1_outputs(627) <= not b or a;
    layer1_outputs(628) <= a and not b;
    layer1_outputs(629) <= not b or a;
    layer1_outputs(630) <= b and not a;
    layer1_outputs(631) <= not b or a;
    layer1_outputs(632) <= not (a and b);
    layer1_outputs(633) <= a or b;
    layer1_outputs(634) <= not a;
    layer1_outputs(635) <= a and b;
    layer1_outputs(636) <= b and not a;
    layer1_outputs(637) <= not b or a;
    layer1_outputs(638) <= a;
    layer1_outputs(639) <= a xor b;
    layer1_outputs(640) <= not a;
    layer1_outputs(641) <= b;
    layer1_outputs(642) <= not a;
    layer1_outputs(643) <= a;
    layer1_outputs(644) <= a and b;
    layer1_outputs(645) <= a and not b;
    layer1_outputs(646) <= not (a and b);
    layer1_outputs(647) <= a and not b;
    layer1_outputs(648) <= not a or b;
    layer1_outputs(649) <= not (a or b);
    layer1_outputs(650) <= b;
    layer1_outputs(651) <= not (a xor b);
    layer1_outputs(652) <= b and not a;
    layer1_outputs(653) <= not (a and b);
    layer1_outputs(654) <= a xor b;
    layer1_outputs(655) <= a xor b;
    layer1_outputs(656) <= a and not b;
    layer1_outputs(657) <= b;
    layer1_outputs(658) <= b;
    layer1_outputs(659) <= not a or b;
    layer1_outputs(660) <= not (a xor b);
    layer1_outputs(661) <= not a;
    layer1_outputs(662) <= not b;
    layer1_outputs(663) <= a or b;
    layer1_outputs(664) <= b and not a;
    layer1_outputs(665) <= not b or a;
    layer1_outputs(666) <= b;
    layer1_outputs(667) <= '1';
    layer1_outputs(668) <= '0';
    layer1_outputs(669) <= not b;
    layer1_outputs(670) <= a and b;
    layer1_outputs(671) <= a and b;
    layer1_outputs(672) <= a and not b;
    layer1_outputs(673) <= b;
    layer1_outputs(674) <= a and b;
    layer1_outputs(675) <= a or b;
    layer1_outputs(676) <= b and not a;
    layer1_outputs(677) <= not a or b;
    layer1_outputs(678) <= '0';
    layer1_outputs(679) <= a;
    layer1_outputs(680) <= a and not b;
    layer1_outputs(681) <= a;
    layer1_outputs(682) <= a or b;
    layer1_outputs(683) <= not b or a;
    layer1_outputs(684) <= not a;
    layer1_outputs(685) <= not a;
    layer1_outputs(686) <= not a;
    layer1_outputs(687) <= b;
    layer1_outputs(688) <= not a;
    layer1_outputs(689) <= b and not a;
    layer1_outputs(690) <= a;
    layer1_outputs(691) <= not (a and b);
    layer1_outputs(692) <= b and not a;
    layer1_outputs(693) <= not b;
    layer1_outputs(694) <= b;
    layer1_outputs(695) <= not a or b;
    layer1_outputs(696) <= a;
    layer1_outputs(697) <= b;
    layer1_outputs(698) <= a;
    layer1_outputs(699) <= b;
    layer1_outputs(700) <= not a or b;
    layer1_outputs(701) <= a xor b;
    layer1_outputs(702) <= '0';
    layer1_outputs(703) <= not (a or b);
    layer1_outputs(704) <= b;
    layer1_outputs(705) <= a and not b;
    layer1_outputs(706) <= a;
    layer1_outputs(707) <= not a or b;
    layer1_outputs(708) <= not a;
    layer1_outputs(709) <= not (a and b);
    layer1_outputs(710) <= b;
    layer1_outputs(711) <= not b;
    layer1_outputs(712) <= not b;
    layer1_outputs(713) <= not b;
    layer1_outputs(714) <= not a;
    layer1_outputs(715) <= not (a or b);
    layer1_outputs(716) <= not (a xor b);
    layer1_outputs(717) <= '0';
    layer1_outputs(718) <= not b;
    layer1_outputs(719) <= a;
    layer1_outputs(720) <= a;
    layer1_outputs(721) <= a or b;
    layer1_outputs(722) <= a and b;
    layer1_outputs(723) <= '1';
    layer1_outputs(724) <= not (a or b);
    layer1_outputs(725) <= b;
    layer1_outputs(726) <= not b or a;
    layer1_outputs(727) <= '1';
    layer1_outputs(728) <= b;
    layer1_outputs(729) <= a xor b;
    layer1_outputs(730) <= not (a xor b);
    layer1_outputs(731) <= not (a xor b);
    layer1_outputs(732) <= a;
    layer1_outputs(733) <= not b;
    layer1_outputs(734) <= not (a or b);
    layer1_outputs(735) <= a and b;
    layer1_outputs(736) <= not a;
    layer1_outputs(737) <= not a;
    layer1_outputs(738) <= a or b;
    layer1_outputs(739) <= a and b;
    layer1_outputs(740) <= a and not b;
    layer1_outputs(741) <= a or b;
    layer1_outputs(742) <= a and not b;
    layer1_outputs(743) <= a and not b;
    layer1_outputs(744) <= not a;
    layer1_outputs(745) <= b and not a;
    layer1_outputs(746) <= not b or a;
    layer1_outputs(747) <= not (a and b);
    layer1_outputs(748) <= a or b;
    layer1_outputs(749) <= a and not b;
    layer1_outputs(750) <= not b;
    layer1_outputs(751) <= a or b;
    layer1_outputs(752) <= not a;
    layer1_outputs(753) <= b and not a;
    layer1_outputs(754) <= not b or a;
    layer1_outputs(755) <= not a;
    layer1_outputs(756) <= b;
    layer1_outputs(757) <= not a or b;
    layer1_outputs(758) <= a xor b;
    layer1_outputs(759) <= b and not a;
    layer1_outputs(760) <= b;
    layer1_outputs(761) <= not b;
    layer1_outputs(762) <= not a;
    layer1_outputs(763) <= a or b;
    layer1_outputs(764) <= a;
    layer1_outputs(765) <= a;
    layer1_outputs(766) <= a and not b;
    layer1_outputs(767) <= '1';
    layer1_outputs(768) <= a and not b;
    layer1_outputs(769) <= not b or a;
    layer1_outputs(770) <= b;
    layer1_outputs(771) <= '1';
    layer1_outputs(772) <= not (a and b);
    layer1_outputs(773) <= not b;
    layer1_outputs(774) <= '1';
    layer1_outputs(775) <= a or b;
    layer1_outputs(776) <= b and not a;
    layer1_outputs(777) <= b;
    layer1_outputs(778) <= a;
    layer1_outputs(779) <= a and b;
    layer1_outputs(780) <= a;
    layer1_outputs(781) <= a and b;
    layer1_outputs(782) <= not (a or b);
    layer1_outputs(783) <= not (a xor b);
    layer1_outputs(784) <= not (a and b);
    layer1_outputs(785) <= '0';
    layer1_outputs(786) <= not (a or b);
    layer1_outputs(787) <= not a;
    layer1_outputs(788) <= a or b;
    layer1_outputs(789) <= not a;
    layer1_outputs(790) <= a xor b;
    layer1_outputs(791) <= a and b;
    layer1_outputs(792) <= a xor b;
    layer1_outputs(793) <= not b or a;
    layer1_outputs(794) <= not b;
    layer1_outputs(795) <= not a;
    layer1_outputs(796) <= a and b;
    layer1_outputs(797) <= not b or a;
    layer1_outputs(798) <= a xor b;
    layer1_outputs(799) <= not b or a;
    layer1_outputs(800) <= a or b;
    layer1_outputs(801) <= '1';
    layer1_outputs(802) <= '0';
    layer1_outputs(803) <= b and not a;
    layer1_outputs(804) <= a or b;
    layer1_outputs(805) <= a xor b;
    layer1_outputs(806) <= not b or a;
    layer1_outputs(807) <= not a or b;
    layer1_outputs(808) <= not a or b;
    layer1_outputs(809) <= not (a and b);
    layer1_outputs(810) <= '1';
    layer1_outputs(811) <= not (a and b);
    layer1_outputs(812) <= not (a and b);
    layer1_outputs(813) <= a;
    layer1_outputs(814) <= not b or a;
    layer1_outputs(815) <= not (a or b);
    layer1_outputs(816) <= not a or b;
    layer1_outputs(817) <= not b or a;
    layer1_outputs(818) <= '0';
    layer1_outputs(819) <= a and b;
    layer1_outputs(820) <= a;
    layer1_outputs(821) <= b;
    layer1_outputs(822) <= not a;
    layer1_outputs(823) <= a and not b;
    layer1_outputs(824) <= '0';
    layer1_outputs(825) <= b;
    layer1_outputs(826) <= not b or a;
    layer1_outputs(827) <= not a or b;
    layer1_outputs(828) <= not a or b;
    layer1_outputs(829) <= a and b;
    layer1_outputs(830) <= not b;
    layer1_outputs(831) <= '0';
    layer1_outputs(832) <= not b or a;
    layer1_outputs(833) <= a;
    layer1_outputs(834) <= not b;
    layer1_outputs(835) <= '1';
    layer1_outputs(836) <= not b;
    layer1_outputs(837) <= not a;
    layer1_outputs(838) <= b;
    layer1_outputs(839) <= a or b;
    layer1_outputs(840) <= b;
    layer1_outputs(841) <= '0';
    layer1_outputs(842) <= a or b;
    layer1_outputs(843) <= not a;
    layer1_outputs(844) <= not (a and b);
    layer1_outputs(845) <= b;
    layer1_outputs(846) <= a xor b;
    layer1_outputs(847) <= not a or b;
    layer1_outputs(848) <= a and not b;
    layer1_outputs(849) <= not b;
    layer1_outputs(850) <= b;
    layer1_outputs(851) <= b;
    layer1_outputs(852) <= not (a and b);
    layer1_outputs(853) <= not b or a;
    layer1_outputs(854) <= b;
    layer1_outputs(855) <= b;
    layer1_outputs(856) <= not (a or b);
    layer1_outputs(857) <= not a or b;
    layer1_outputs(858) <= a and b;
    layer1_outputs(859) <= a or b;
    layer1_outputs(860) <= not b or a;
    layer1_outputs(861) <= not (a and b);
    layer1_outputs(862) <= a or b;
    layer1_outputs(863) <= a;
    layer1_outputs(864) <= not b or a;
    layer1_outputs(865) <= a;
    layer1_outputs(866) <= a and not b;
    layer1_outputs(867) <= b;
    layer1_outputs(868) <= b and not a;
    layer1_outputs(869) <= not b;
    layer1_outputs(870) <= b;
    layer1_outputs(871) <= '0';
    layer1_outputs(872) <= a or b;
    layer1_outputs(873) <= a;
    layer1_outputs(874) <= '1';
    layer1_outputs(875) <= not a or b;
    layer1_outputs(876) <= a and b;
    layer1_outputs(877) <= b and not a;
    layer1_outputs(878) <= not a or b;
    layer1_outputs(879) <= a and b;
    layer1_outputs(880) <= '0';
    layer1_outputs(881) <= b;
    layer1_outputs(882) <= a xor b;
    layer1_outputs(883) <= b;
    layer1_outputs(884) <= '1';
    layer1_outputs(885) <= a or b;
    layer1_outputs(886) <= not a or b;
    layer1_outputs(887) <= not a or b;
    layer1_outputs(888) <= not a or b;
    layer1_outputs(889) <= a and b;
    layer1_outputs(890) <= a and not b;
    layer1_outputs(891) <= not b;
    layer1_outputs(892) <= not (a and b);
    layer1_outputs(893) <= a xor b;
    layer1_outputs(894) <= not b;
    layer1_outputs(895) <= not (a or b);
    layer1_outputs(896) <= a and b;
    layer1_outputs(897) <= not a or b;
    layer1_outputs(898) <= b;
    layer1_outputs(899) <= '1';
    layer1_outputs(900) <= not (a and b);
    layer1_outputs(901) <= a xor b;
    layer1_outputs(902) <= a and b;
    layer1_outputs(903) <= b;
    layer1_outputs(904) <= not b;
    layer1_outputs(905) <= a;
    layer1_outputs(906) <= not a;
    layer1_outputs(907) <= not a or b;
    layer1_outputs(908) <= not (a or b);
    layer1_outputs(909) <= a;
    layer1_outputs(910) <= a xor b;
    layer1_outputs(911) <= not a;
    layer1_outputs(912) <= a and b;
    layer1_outputs(913) <= not b or a;
    layer1_outputs(914) <= a;
    layer1_outputs(915) <= not a or b;
    layer1_outputs(916) <= '1';
    layer1_outputs(917) <= '0';
    layer1_outputs(918) <= a;
    layer1_outputs(919) <= '1';
    layer1_outputs(920) <= a xor b;
    layer1_outputs(921) <= not (a or b);
    layer1_outputs(922) <= a and b;
    layer1_outputs(923) <= '0';
    layer1_outputs(924) <= not (a or b);
    layer1_outputs(925) <= '1';
    layer1_outputs(926) <= a;
    layer1_outputs(927) <= a;
    layer1_outputs(928) <= a and not b;
    layer1_outputs(929) <= a and not b;
    layer1_outputs(930) <= not a or b;
    layer1_outputs(931) <= b and not a;
    layer1_outputs(932) <= not (a or b);
    layer1_outputs(933) <= b;
    layer1_outputs(934) <= not b or a;
    layer1_outputs(935) <= a and not b;
    layer1_outputs(936) <= not a;
    layer1_outputs(937) <= not b;
    layer1_outputs(938) <= not b;
    layer1_outputs(939) <= b;
    layer1_outputs(940) <= b;
    layer1_outputs(941) <= a or b;
    layer1_outputs(942) <= a and b;
    layer1_outputs(943) <= not a;
    layer1_outputs(944) <= not a or b;
    layer1_outputs(945) <= a;
    layer1_outputs(946) <= not b;
    layer1_outputs(947) <= '1';
    layer1_outputs(948) <= not b or a;
    layer1_outputs(949) <= not (a or b);
    layer1_outputs(950) <= b;
    layer1_outputs(951) <= not (a or b);
    layer1_outputs(952) <= a;
    layer1_outputs(953) <= a xor b;
    layer1_outputs(954) <= a and not b;
    layer1_outputs(955) <= not (a and b);
    layer1_outputs(956) <= b;
    layer1_outputs(957) <= not b;
    layer1_outputs(958) <= '1';
    layer1_outputs(959) <= a;
    layer1_outputs(960) <= '0';
    layer1_outputs(961) <= not (a and b);
    layer1_outputs(962) <= not (a or b);
    layer1_outputs(963) <= not a;
    layer1_outputs(964) <= not a;
    layer1_outputs(965) <= '0';
    layer1_outputs(966) <= not b;
    layer1_outputs(967) <= not a;
    layer1_outputs(968) <= not (a or b);
    layer1_outputs(969) <= not a;
    layer1_outputs(970) <= not (a or b);
    layer1_outputs(971) <= not (a or b);
    layer1_outputs(972) <= b and not a;
    layer1_outputs(973) <= not a;
    layer1_outputs(974) <= not b;
    layer1_outputs(975) <= a or b;
    layer1_outputs(976) <= a or b;
    layer1_outputs(977) <= a and b;
    layer1_outputs(978) <= not b;
    layer1_outputs(979) <= a or b;
    layer1_outputs(980) <= not b;
    layer1_outputs(981) <= b and not a;
    layer1_outputs(982) <= '1';
    layer1_outputs(983) <= b and not a;
    layer1_outputs(984) <= not b or a;
    layer1_outputs(985) <= '1';
    layer1_outputs(986) <= a and b;
    layer1_outputs(987) <= b;
    layer1_outputs(988) <= b;
    layer1_outputs(989) <= '1';
    layer1_outputs(990) <= not b;
    layer1_outputs(991) <= a and not b;
    layer1_outputs(992) <= a and b;
    layer1_outputs(993) <= not (a and b);
    layer1_outputs(994) <= not (a and b);
    layer1_outputs(995) <= not b;
    layer1_outputs(996) <= a;
    layer1_outputs(997) <= not b;
    layer1_outputs(998) <= not a;
    layer1_outputs(999) <= not a or b;
    layer1_outputs(1000) <= '1';
    layer1_outputs(1001) <= a;
    layer1_outputs(1002) <= '0';
    layer1_outputs(1003) <= '1';
    layer1_outputs(1004) <= not a or b;
    layer1_outputs(1005) <= not a or b;
    layer1_outputs(1006) <= b;
    layer1_outputs(1007) <= b and not a;
    layer1_outputs(1008) <= '1';
    layer1_outputs(1009) <= not b or a;
    layer1_outputs(1010) <= not a;
    layer1_outputs(1011) <= not (a and b);
    layer1_outputs(1012) <= a or b;
    layer1_outputs(1013) <= a;
    layer1_outputs(1014) <= not a;
    layer1_outputs(1015) <= a;
    layer1_outputs(1016) <= not b or a;
    layer1_outputs(1017) <= a and b;
    layer1_outputs(1018) <= b;
    layer1_outputs(1019) <= not a;
    layer1_outputs(1020) <= not b;
    layer1_outputs(1021) <= not (a or b);
    layer1_outputs(1022) <= b and not a;
    layer1_outputs(1023) <= a and b;
    layer1_outputs(1024) <= a and b;
    layer1_outputs(1025) <= not (a xor b);
    layer1_outputs(1026) <= a or b;
    layer1_outputs(1027) <= a;
    layer1_outputs(1028) <= a or b;
    layer1_outputs(1029) <= '0';
    layer1_outputs(1030) <= '1';
    layer1_outputs(1031) <= b and not a;
    layer1_outputs(1032) <= not (a and b);
    layer1_outputs(1033) <= b;
    layer1_outputs(1034) <= a xor b;
    layer1_outputs(1035) <= not (a or b);
    layer1_outputs(1036) <= not b;
    layer1_outputs(1037) <= not (a or b);
    layer1_outputs(1038) <= a and b;
    layer1_outputs(1039) <= a and not b;
    layer1_outputs(1040) <= not b or a;
    layer1_outputs(1041) <= not b or a;
    layer1_outputs(1042) <= not (a and b);
    layer1_outputs(1043) <= not b;
    layer1_outputs(1044) <= not b;
    layer1_outputs(1045) <= a and not b;
    layer1_outputs(1046) <= not b or a;
    layer1_outputs(1047) <= not b;
    layer1_outputs(1048) <= a and not b;
    layer1_outputs(1049) <= not b;
    layer1_outputs(1050) <= b and not a;
    layer1_outputs(1051) <= b;
    layer1_outputs(1052) <= b and not a;
    layer1_outputs(1053) <= a or b;
    layer1_outputs(1054) <= not a;
    layer1_outputs(1055) <= '0';
    layer1_outputs(1056) <= not a or b;
    layer1_outputs(1057) <= not (a and b);
    layer1_outputs(1058) <= not b;
    layer1_outputs(1059) <= a and b;
    layer1_outputs(1060) <= a;
    layer1_outputs(1061) <= not b;
    layer1_outputs(1062) <= a;
    layer1_outputs(1063) <= a and b;
    layer1_outputs(1064) <= not (a and b);
    layer1_outputs(1065) <= '0';
    layer1_outputs(1066) <= b and not a;
    layer1_outputs(1067) <= a and b;
    layer1_outputs(1068) <= a;
    layer1_outputs(1069) <= not b or a;
    layer1_outputs(1070) <= '1';
    layer1_outputs(1071) <= not (a and b);
    layer1_outputs(1072) <= not b;
    layer1_outputs(1073) <= b and not a;
    layer1_outputs(1074) <= a;
    layer1_outputs(1075) <= a or b;
    layer1_outputs(1076) <= b and not a;
    layer1_outputs(1077) <= not (a or b);
    layer1_outputs(1078) <= not (a or b);
    layer1_outputs(1079) <= not b;
    layer1_outputs(1080) <= not (a or b);
    layer1_outputs(1081) <= not (a or b);
    layer1_outputs(1082) <= a or b;
    layer1_outputs(1083) <= a and b;
    layer1_outputs(1084) <= a or b;
    layer1_outputs(1085) <= b and not a;
    layer1_outputs(1086) <= a xor b;
    layer1_outputs(1087) <= a or b;
    layer1_outputs(1088) <= a and not b;
    layer1_outputs(1089) <= not (a and b);
    layer1_outputs(1090) <= not b or a;
    layer1_outputs(1091) <= a or b;
    layer1_outputs(1092) <= b;
    layer1_outputs(1093) <= a;
    layer1_outputs(1094) <= '1';
    layer1_outputs(1095) <= '1';
    layer1_outputs(1096) <= not (a xor b);
    layer1_outputs(1097) <= not a;
    layer1_outputs(1098) <= '0';
    layer1_outputs(1099) <= not (a or b);
    layer1_outputs(1100) <= not b;
    layer1_outputs(1101) <= not (a or b);
    layer1_outputs(1102) <= b;
    layer1_outputs(1103) <= b and not a;
    layer1_outputs(1104) <= a and not b;
    layer1_outputs(1105) <= a xor b;
    layer1_outputs(1106) <= b and not a;
    layer1_outputs(1107) <= not (a and b);
    layer1_outputs(1108) <= a and b;
    layer1_outputs(1109) <= not a or b;
    layer1_outputs(1110) <= a and b;
    layer1_outputs(1111) <= a or b;
    layer1_outputs(1112) <= a;
    layer1_outputs(1113) <= not (a and b);
    layer1_outputs(1114) <= not b;
    layer1_outputs(1115) <= not b;
    layer1_outputs(1116) <= a and b;
    layer1_outputs(1117) <= b;
    layer1_outputs(1118) <= b;
    layer1_outputs(1119) <= not (a xor b);
    layer1_outputs(1120) <= a xor b;
    layer1_outputs(1121) <= a;
    layer1_outputs(1122) <= a and b;
    layer1_outputs(1123) <= not (a or b);
    layer1_outputs(1124) <= a xor b;
    layer1_outputs(1125) <= a and not b;
    layer1_outputs(1126) <= not a;
    layer1_outputs(1127) <= not a or b;
    layer1_outputs(1128) <= not b or a;
    layer1_outputs(1129) <= a xor b;
    layer1_outputs(1130) <= a;
    layer1_outputs(1131) <= not a;
    layer1_outputs(1132) <= not (a and b);
    layer1_outputs(1133) <= a xor b;
    layer1_outputs(1134) <= b;
    layer1_outputs(1135) <= not (a and b);
    layer1_outputs(1136) <= not a;
    layer1_outputs(1137) <= not a or b;
    layer1_outputs(1138) <= a and not b;
    layer1_outputs(1139) <= a and b;
    layer1_outputs(1140) <= not b;
    layer1_outputs(1141) <= not (a or b);
    layer1_outputs(1142) <= not (a and b);
    layer1_outputs(1143) <= a xor b;
    layer1_outputs(1144) <= not a or b;
    layer1_outputs(1145) <= not b;
    layer1_outputs(1146) <= not (a or b);
    layer1_outputs(1147) <= b and not a;
    layer1_outputs(1148) <= b and not a;
    layer1_outputs(1149) <= a xor b;
    layer1_outputs(1150) <= '1';
    layer1_outputs(1151) <= not (a or b);
    layer1_outputs(1152) <= not a;
    layer1_outputs(1153) <= a xor b;
    layer1_outputs(1154) <= not b or a;
    layer1_outputs(1155) <= not (a or b);
    layer1_outputs(1156) <= '0';
    layer1_outputs(1157) <= not (a xor b);
    layer1_outputs(1158) <= a and b;
    layer1_outputs(1159) <= a or b;
    layer1_outputs(1160) <= a or b;
    layer1_outputs(1161) <= not a;
    layer1_outputs(1162) <= b;
    layer1_outputs(1163) <= a or b;
    layer1_outputs(1164) <= not a or b;
    layer1_outputs(1165) <= b and not a;
    layer1_outputs(1166) <= not (a xor b);
    layer1_outputs(1167) <= '0';
    layer1_outputs(1168) <= not (a xor b);
    layer1_outputs(1169) <= not a;
    layer1_outputs(1170) <= a;
    layer1_outputs(1171) <= '1';
    layer1_outputs(1172) <= b;
    layer1_outputs(1173) <= not b or a;
    layer1_outputs(1174) <= not b or a;
    layer1_outputs(1175) <= b;
    layer1_outputs(1176) <= a;
    layer1_outputs(1177) <= a and b;
    layer1_outputs(1178) <= b and not a;
    layer1_outputs(1179) <= not (a and b);
    layer1_outputs(1180) <= a and not b;
    layer1_outputs(1181) <= not a;
    layer1_outputs(1182) <= not b;
    layer1_outputs(1183) <= a xor b;
    layer1_outputs(1184) <= a;
    layer1_outputs(1185) <= b and not a;
    layer1_outputs(1186) <= b;
    layer1_outputs(1187) <= b;
    layer1_outputs(1188) <= a and not b;
    layer1_outputs(1189) <= not b;
    layer1_outputs(1190) <= not a or b;
    layer1_outputs(1191) <= a or b;
    layer1_outputs(1192) <= a or b;
    layer1_outputs(1193) <= a or b;
    layer1_outputs(1194) <= '1';
    layer1_outputs(1195) <= not (a and b);
    layer1_outputs(1196) <= a and not b;
    layer1_outputs(1197) <= a;
    layer1_outputs(1198) <= not b;
    layer1_outputs(1199) <= not b;
    layer1_outputs(1200) <= not (a or b);
    layer1_outputs(1201) <= not (a and b);
    layer1_outputs(1202) <= '0';
    layer1_outputs(1203) <= not a;
    layer1_outputs(1204) <= b and not a;
    layer1_outputs(1205) <= not b;
    layer1_outputs(1206) <= '0';
    layer1_outputs(1207) <= not a;
    layer1_outputs(1208) <= '0';
    layer1_outputs(1209) <= not (a and b);
    layer1_outputs(1210) <= a;
    layer1_outputs(1211) <= not a or b;
    layer1_outputs(1212) <= not a;
    layer1_outputs(1213) <= not (a or b);
    layer1_outputs(1214) <= a xor b;
    layer1_outputs(1215) <= a or b;
    layer1_outputs(1216) <= '1';
    layer1_outputs(1217) <= b and not a;
    layer1_outputs(1218) <= not (a or b);
    layer1_outputs(1219) <= not b;
    layer1_outputs(1220) <= not (a or b);
    layer1_outputs(1221) <= not b or a;
    layer1_outputs(1222) <= a;
    layer1_outputs(1223) <= not a;
    layer1_outputs(1224) <= a or b;
    layer1_outputs(1225) <= not b or a;
    layer1_outputs(1226) <= not (a or b);
    layer1_outputs(1227) <= not b or a;
    layer1_outputs(1228) <= a and b;
    layer1_outputs(1229) <= not a;
    layer1_outputs(1230) <= b and not a;
    layer1_outputs(1231) <= not b;
    layer1_outputs(1232) <= not (a xor b);
    layer1_outputs(1233) <= b and not a;
    layer1_outputs(1234) <= not a;
    layer1_outputs(1235) <= a or b;
    layer1_outputs(1236) <= '1';
    layer1_outputs(1237) <= '0';
    layer1_outputs(1238) <= a and b;
    layer1_outputs(1239) <= '1';
    layer1_outputs(1240) <= '1';
    layer1_outputs(1241) <= '0';
    layer1_outputs(1242) <= '1';
    layer1_outputs(1243) <= b;
    layer1_outputs(1244) <= not b or a;
    layer1_outputs(1245) <= not a or b;
    layer1_outputs(1246) <= not a;
    layer1_outputs(1247) <= b and not a;
    layer1_outputs(1248) <= b and not a;
    layer1_outputs(1249) <= a or b;
    layer1_outputs(1250) <= not b;
    layer1_outputs(1251) <= '1';
    layer1_outputs(1252) <= '1';
    layer1_outputs(1253) <= a xor b;
    layer1_outputs(1254) <= not (a and b);
    layer1_outputs(1255) <= a;
    layer1_outputs(1256) <= not (a and b);
    layer1_outputs(1257) <= not (a or b);
    layer1_outputs(1258) <= '0';
    layer1_outputs(1259) <= not b;
    layer1_outputs(1260) <= '1';
    layer1_outputs(1261) <= a and not b;
    layer1_outputs(1262) <= a and b;
    layer1_outputs(1263) <= not (a and b);
    layer1_outputs(1264) <= not b or a;
    layer1_outputs(1265) <= not a;
    layer1_outputs(1266) <= '1';
    layer1_outputs(1267) <= not (a xor b);
    layer1_outputs(1268) <= not a;
    layer1_outputs(1269) <= b and not a;
    layer1_outputs(1270) <= not b or a;
    layer1_outputs(1271) <= not (a xor b);
    layer1_outputs(1272) <= a and not b;
    layer1_outputs(1273) <= not (a and b);
    layer1_outputs(1274) <= '1';
    layer1_outputs(1275) <= not (a and b);
    layer1_outputs(1276) <= not (a and b);
    layer1_outputs(1277) <= not (a or b);
    layer1_outputs(1278) <= not b or a;
    layer1_outputs(1279) <= not a;
    layer1_outputs(1280) <= a or b;
    layer1_outputs(1281) <= not a;
    layer1_outputs(1282) <= not a or b;
    layer1_outputs(1283) <= a;
    layer1_outputs(1284) <= not b;
    layer1_outputs(1285) <= not b or a;
    layer1_outputs(1286) <= b;
    layer1_outputs(1287) <= b and not a;
    layer1_outputs(1288) <= a or b;
    layer1_outputs(1289) <= a;
    layer1_outputs(1290) <= a;
    layer1_outputs(1291) <= b and not a;
    layer1_outputs(1292) <= b and not a;
    layer1_outputs(1293) <= b;
    layer1_outputs(1294) <= '0';
    layer1_outputs(1295) <= '0';
    layer1_outputs(1296) <= '1';
    layer1_outputs(1297) <= a xor b;
    layer1_outputs(1298) <= a and not b;
    layer1_outputs(1299) <= not a;
    layer1_outputs(1300) <= '1';
    layer1_outputs(1301) <= '1';
    layer1_outputs(1302) <= a and not b;
    layer1_outputs(1303) <= not a;
    layer1_outputs(1304) <= '0';
    layer1_outputs(1305) <= a and b;
    layer1_outputs(1306) <= a;
    layer1_outputs(1307) <= a and not b;
    layer1_outputs(1308) <= not a or b;
    layer1_outputs(1309) <= not b or a;
    layer1_outputs(1310) <= not b;
    layer1_outputs(1311) <= not b;
    layer1_outputs(1312) <= not b;
    layer1_outputs(1313) <= not (a xor b);
    layer1_outputs(1314) <= a;
    layer1_outputs(1315) <= not (a or b);
    layer1_outputs(1316) <= '1';
    layer1_outputs(1317) <= not (a and b);
    layer1_outputs(1318) <= not a;
    layer1_outputs(1319) <= '0';
    layer1_outputs(1320) <= a and not b;
    layer1_outputs(1321) <= '0';
    layer1_outputs(1322) <= not b;
    layer1_outputs(1323) <= not a or b;
    layer1_outputs(1324) <= not (a xor b);
    layer1_outputs(1325) <= a or b;
    layer1_outputs(1326) <= not b;
    layer1_outputs(1327) <= not a;
    layer1_outputs(1328) <= b;
    layer1_outputs(1329) <= a or b;
    layer1_outputs(1330) <= '1';
    layer1_outputs(1331) <= not b or a;
    layer1_outputs(1332) <= not b;
    layer1_outputs(1333) <= '0';
    layer1_outputs(1334) <= not (a or b);
    layer1_outputs(1335) <= a and b;
    layer1_outputs(1336) <= b;
    layer1_outputs(1337) <= not b or a;
    layer1_outputs(1338) <= not a;
    layer1_outputs(1339) <= not b;
    layer1_outputs(1340) <= a and b;
    layer1_outputs(1341) <= not a;
    layer1_outputs(1342) <= not a;
    layer1_outputs(1343) <= not (a xor b);
    layer1_outputs(1344) <= '1';
    layer1_outputs(1345) <= not (a and b);
    layer1_outputs(1346) <= a or b;
    layer1_outputs(1347) <= a and b;
    layer1_outputs(1348) <= not a;
    layer1_outputs(1349) <= not (a and b);
    layer1_outputs(1350) <= not a;
    layer1_outputs(1351) <= a or b;
    layer1_outputs(1352) <= a;
    layer1_outputs(1353) <= a xor b;
    layer1_outputs(1354) <= '1';
    layer1_outputs(1355) <= a or b;
    layer1_outputs(1356) <= '0';
    layer1_outputs(1357) <= not a;
    layer1_outputs(1358) <= a xor b;
    layer1_outputs(1359) <= a and b;
    layer1_outputs(1360) <= b;
    layer1_outputs(1361) <= not b or a;
    layer1_outputs(1362) <= '0';
    layer1_outputs(1363) <= not a;
    layer1_outputs(1364) <= b and not a;
    layer1_outputs(1365) <= b and not a;
    layer1_outputs(1366) <= '1';
    layer1_outputs(1367) <= a or b;
    layer1_outputs(1368) <= b;
    layer1_outputs(1369) <= b;
    layer1_outputs(1370) <= a and not b;
    layer1_outputs(1371) <= a or b;
    layer1_outputs(1372) <= not a;
    layer1_outputs(1373) <= a and not b;
    layer1_outputs(1374) <= not (a and b);
    layer1_outputs(1375) <= '1';
    layer1_outputs(1376) <= not b or a;
    layer1_outputs(1377) <= '1';
    layer1_outputs(1378) <= b and not a;
    layer1_outputs(1379) <= not (a and b);
    layer1_outputs(1380) <= not (a or b);
    layer1_outputs(1381) <= '1';
    layer1_outputs(1382) <= a and not b;
    layer1_outputs(1383) <= a or b;
    layer1_outputs(1384) <= not b;
    layer1_outputs(1385) <= not a or b;
    layer1_outputs(1386) <= a xor b;
    layer1_outputs(1387) <= not (a xor b);
    layer1_outputs(1388) <= not b or a;
    layer1_outputs(1389) <= not a;
    layer1_outputs(1390) <= not (a or b);
    layer1_outputs(1391) <= not a or b;
    layer1_outputs(1392) <= a and b;
    layer1_outputs(1393) <= not a;
    layer1_outputs(1394) <= not a;
    layer1_outputs(1395) <= a and b;
    layer1_outputs(1396) <= not a or b;
    layer1_outputs(1397) <= not a;
    layer1_outputs(1398) <= not (a or b);
    layer1_outputs(1399) <= a;
    layer1_outputs(1400) <= not (a and b);
    layer1_outputs(1401) <= b and not a;
    layer1_outputs(1402) <= not a;
    layer1_outputs(1403) <= a and not b;
    layer1_outputs(1404) <= a and not b;
    layer1_outputs(1405) <= a;
    layer1_outputs(1406) <= not b or a;
    layer1_outputs(1407) <= b and not a;
    layer1_outputs(1408) <= a and b;
    layer1_outputs(1409) <= not b;
    layer1_outputs(1410) <= not b or a;
    layer1_outputs(1411) <= '0';
    layer1_outputs(1412) <= not a;
    layer1_outputs(1413) <= not a;
    layer1_outputs(1414) <= not (a xor b);
    layer1_outputs(1415) <= '0';
    layer1_outputs(1416) <= b;
    layer1_outputs(1417) <= not (a xor b);
    layer1_outputs(1418) <= not (a or b);
    layer1_outputs(1419) <= a or b;
    layer1_outputs(1420) <= not (a or b);
    layer1_outputs(1421) <= a and b;
    layer1_outputs(1422) <= not a or b;
    layer1_outputs(1423) <= a and not b;
    layer1_outputs(1424) <= not b or a;
    layer1_outputs(1425) <= a;
    layer1_outputs(1426) <= a and not b;
    layer1_outputs(1427) <= a and not b;
    layer1_outputs(1428) <= b;
    layer1_outputs(1429) <= not a or b;
    layer1_outputs(1430) <= '0';
    layer1_outputs(1431) <= not a or b;
    layer1_outputs(1432) <= not (a or b);
    layer1_outputs(1433) <= not a;
    layer1_outputs(1434) <= not (a or b);
    layer1_outputs(1435) <= not a;
    layer1_outputs(1436) <= not b or a;
    layer1_outputs(1437) <= '1';
    layer1_outputs(1438) <= a;
    layer1_outputs(1439) <= a and not b;
    layer1_outputs(1440) <= not (a or b);
    layer1_outputs(1441) <= a xor b;
    layer1_outputs(1442) <= not (a and b);
    layer1_outputs(1443) <= a and b;
    layer1_outputs(1444) <= not a;
    layer1_outputs(1445) <= '1';
    layer1_outputs(1446) <= a xor b;
    layer1_outputs(1447) <= not a;
    layer1_outputs(1448) <= a and not b;
    layer1_outputs(1449) <= a and not b;
    layer1_outputs(1450) <= not (a and b);
    layer1_outputs(1451) <= a and b;
    layer1_outputs(1452) <= a and b;
    layer1_outputs(1453) <= not (a and b);
    layer1_outputs(1454) <= not (a and b);
    layer1_outputs(1455) <= not a or b;
    layer1_outputs(1456) <= '1';
    layer1_outputs(1457) <= a or b;
    layer1_outputs(1458) <= not (a or b);
    layer1_outputs(1459) <= not b or a;
    layer1_outputs(1460) <= '0';
    layer1_outputs(1461) <= a and not b;
    layer1_outputs(1462) <= not b;
    layer1_outputs(1463) <= b and not a;
    layer1_outputs(1464) <= not (a and b);
    layer1_outputs(1465) <= not (a and b);
    layer1_outputs(1466) <= not b or a;
    layer1_outputs(1467) <= a or b;
    layer1_outputs(1468) <= not b or a;
    layer1_outputs(1469) <= not b;
    layer1_outputs(1470) <= '0';
    layer1_outputs(1471) <= not (a and b);
    layer1_outputs(1472) <= '1';
    layer1_outputs(1473) <= not a or b;
    layer1_outputs(1474) <= a and not b;
    layer1_outputs(1475) <= not a;
    layer1_outputs(1476) <= not (a and b);
    layer1_outputs(1477) <= not a;
    layer1_outputs(1478) <= not b or a;
    layer1_outputs(1479) <= a and b;
    layer1_outputs(1480) <= a;
    layer1_outputs(1481) <= not b;
    layer1_outputs(1482) <= b and not a;
    layer1_outputs(1483) <= not a or b;
    layer1_outputs(1484) <= b and not a;
    layer1_outputs(1485) <= '1';
    layer1_outputs(1486) <= not b;
    layer1_outputs(1487) <= not (a or b);
    layer1_outputs(1488) <= not b or a;
    layer1_outputs(1489) <= not b;
    layer1_outputs(1490) <= not b;
    layer1_outputs(1491) <= not a or b;
    layer1_outputs(1492) <= not b;
    layer1_outputs(1493) <= not (a or b);
    layer1_outputs(1494) <= not a or b;
    layer1_outputs(1495) <= not (a xor b);
    layer1_outputs(1496) <= not a or b;
    layer1_outputs(1497) <= a;
    layer1_outputs(1498) <= a or b;
    layer1_outputs(1499) <= a or b;
    layer1_outputs(1500) <= b;
    layer1_outputs(1501) <= not (a and b);
    layer1_outputs(1502) <= b;
    layer1_outputs(1503) <= not b;
    layer1_outputs(1504) <= a or b;
    layer1_outputs(1505) <= '0';
    layer1_outputs(1506) <= '1';
    layer1_outputs(1507) <= a and b;
    layer1_outputs(1508) <= not b or a;
    layer1_outputs(1509) <= a and b;
    layer1_outputs(1510) <= '1';
    layer1_outputs(1511) <= not b;
    layer1_outputs(1512) <= b and not a;
    layer1_outputs(1513) <= not (a xor b);
    layer1_outputs(1514) <= not a or b;
    layer1_outputs(1515) <= a;
    layer1_outputs(1516) <= a or b;
    layer1_outputs(1517) <= a or b;
    layer1_outputs(1518) <= not a or b;
    layer1_outputs(1519) <= not b;
    layer1_outputs(1520) <= '1';
    layer1_outputs(1521) <= b;
    layer1_outputs(1522) <= not (a and b);
    layer1_outputs(1523) <= '0';
    layer1_outputs(1524) <= '0';
    layer1_outputs(1525) <= not (a and b);
    layer1_outputs(1526) <= '1';
    layer1_outputs(1527) <= not b or a;
    layer1_outputs(1528) <= a;
    layer1_outputs(1529) <= a or b;
    layer1_outputs(1530) <= a;
    layer1_outputs(1531) <= a;
    layer1_outputs(1532) <= b and not a;
    layer1_outputs(1533) <= '1';
    layer1_outputs(1534) <= not (a and b);
    layer1_outputs(1535) <= '0';
    layer1_outputs(1536) <= '0';
    layer1_outputs(1537) <= not b;
    layer1_outputs(1538) <= not (a and b);
    layer1_outputs(1539) <= b and not a;
    layer1_outputs(1540) <= b;
    layer1_outputs(1541) <= '0';
    layer1_outputs(1542) <= b;
    layer1_outputs(1543) <= a and not b;
    layer1_outputs(1544) <= not a or b;
    layer1_outputs(1545) <= a;
    layer1_outputs(1546) <= not a;
    layer1_outputs(1547) <= not (a xor b);
    layer1_outputs(1548) <= a and b;
    layer1_outputs(1549) <= not (a or b);
    layer1_outputs(1550) <= not (a and b);
    layer1_outputs(1551) <= '0';
    layer1_outputs(1552) <= not a;
    layer1_outputs(1553) <= not (a xor b);
    layer1_outputs(1554) <= b;
    layer1_outputs(1555) <= b and not a;
    layer1_outputs(1556) <= a and b;
    layer1_outputs(1557) <= not b;
    layer1_outputs(1558) <= a;
    layer1_outputs(1559) <= b and not a;
    layer1_outputs(1560) <= not b or a;
    layer1_outputs(1561) <= a;
    layer1_outputs(1562) <= not b;
    layer1_outputs(1563) <= not a or b;
    layer1_outputs(1564) <= '1';
    layer1_outputs(1565) <= not b or a;
    layer1_outputs(1566) <= not a;
    layer1_outputs(1567) <= a and b;
    layer1_outputs(1568) <= a and b;
    layer1_outputs(1569) <= '1';
    layer1_outputs(1570) <= a;
    layer1_outputs(1571) <= '1';
    layer1_outputs(1572) <= b;
    layer1_outputs(1573) <= a and b;
    layer1_outputs(1574) <= '0';
    layer1_outputs(1575) <= '1';
    layer1_outputs(1576) <= not a or b;
    layer1_outputs(1577) <= b;
    layer1_outputs(1578) <= a;
    layer1_outputs(1579) <= b and not a;
    layer1_outputs(1580) <= not a or b;
    layer1_outputs(1581) <= not b or a;
    layer1_outputs(1582) <= a and b;
    layer1_outputs(1583) <= '0';
    layer1_outputs(1584) <= a or b;
    layer1_outputs(1585) <= a and not b;
    layer1_outputs(1586) <= not b or a;
    layer1_outputs(1587) <= not (a and b);
    layer1_outputs(1588) <= b and not a;
    layer1_outputs(1589) <= not b or a;
    layer1_outputs(1590) <= not b;
    layer1_outputs(1591) <= not b or a;
    layer1_outputs(1592) <= not (a or b);
    layer1_outputs(1593) <= b;
    layer1_outputs(1594) <= not (a or b);
    layer1_outputs(1595) <= not b or a;
    layer1_outputs(1596) <= not b;
    layer1_outputs(1597) <= not (a and b);
    layer1_outputs(1598) <= not (a xor b);
    layer1_outputs(1599) <= not (a or b);
    layer1_outputs(1600) <= b;
    layer1_outputs(1601) <= b and not a;
    layer1_outputs(1602) <= not a;
    layer1_outputs(1603) <= a xor b;
    layer1_outputs(1604) <= b;
    layer1_outputs(1605) <= b and not a;
    layer1_outputs(1606) <= not a or b;
    layer1_outputs(1607) <= not (a or b);
    layer1_outputs(1608) <= b;
    layer1_outputs(1609) <= '0';
    layer1_outputs(1610) <= a and b;
    layer1_outputs(1611) <= not (a or b);
    layer1_outputs(1612) <= b and not a;
    layer1_outputs(1613) <= b and not a;
    layer1_outputs(1614) <= b;
    layer1_outputs(1615) <= '0';
    layer1_outputs(1616) <= b;
    layer1_outputs(1617) <= '0';
    layer1_outputs(1618) <= a xor b;
    layer1_outputs(1619) <= '1';
    layer1_outputs(1620) <= not (a or b);
    layer1_outputs(1621) <= not (a or b);
    layer1_outputs(1622) <= not b;
    layer1_outputs(1623) <= not (a or b);
    layer1_outputs(1624) <= not b;
    layer1_outputs(1625) <= b;
    layer1_outputs(1626) <= not b or a;
    layer1_outputs(1627) <= a;
    layer1_outputs(1628) <= b;
    layer1_outputs(1629) <= a or b;
    layer1_outputs(1630) <= not b or a;
    layer1_outputs(1631) <= a and not b;
    layer1_outputs(1632) <= a;
    layer1_outputs(1633) <= '1';
    layer1_outputs(1634) <= a and not b;
    layer1_outputs(1635) <= b and not a;
    layer1_outputs(1636) <= a and b;
    layer1_outputs(1637) <= a;
    layer1_outputs(1638) <= '1';
    layer1_outputs(1639) <= not (a and b);
    layer1_outputs(1640) <= not a;
    layer1_outputs(1641) <= '1';
    layer1_outputs(1642) <= b;
    layer1_outputs(1643) <= not a;
    layer1_outputs(1644) <= '1';
    layer1_outputs(1645) <= b;
    layer1_outputs(1646) <= a and b;
    layer1_outputs(1647) <= not b or a;
    layer1_outputs(1648) <= a or b;
    layer1_outputs(1649) <= '0';
    layer1_outputs(1650) <= not b;
    layer1_outputs(1651) <= not b;
    layer1_outputs(1652) <= a and not b;
    layer1_outputs(1653) <= not b or a;
    layer1_outputs(1654) <= not (a or b);
    layer1_outputs(1655) <= a;
    layer1_outputs(1656) <= not a or b;
    layer1_outputs(1657) <= not (a or b);
    layer1_outputs(1658) <= not (a or b);
    layer1_outputs(1659) <= a or b;
    layer1_outputs(1660) <= a and b;
    layer1_outputs(1661) <= a and b;
    layer1_outputs(1662) <= a or b;
    layer1_outputs(1663) <= not b or a;
    layer1_outputs(1664) <= a and b;
    layer1_outputs(1665) <= not b or a;
    layer1_outputs(1666) <= '1';
    layer1_outputs(1667) <= not b;
    layer1_outputs(1668) <= not a or b;
    layer1_outputs(1669) <= not (a or b);
    layer1_outputs(1670) <= not b or a;
    layer1_outputs(1671) <= b;
    layer1_outputs(1672) <= a or b;
    layer1_outputs(1673) <= not a or b;
    layer1_outputs(1674) <= b;
    layer1_outputs(1675) <= not a or b;
    layer1_outputs(1676) <= a xor b;
    layer1_outputs(1677) <= not (a xor b);
    layer1_outputs(1678) <= not b or a;
    layer1_outputs(1679) <= b and not a;
    layer1_outputs(1680) <= not b;
    layer1_outputs(1681) <= a;
    layer1_outputs(1682) <= b;
    layer1_outputs(1683) <= not (a and b);
    layer1_outputs(1684) <= not (a and b);
    layer1_outputs(1685) <= b and not a;
    layer1_outputs(1686) <= b;
    layer1_outputs(1687) <= not b or a;
    layer1_outputs(1688) <= a xor b;
    layer1_outputs(1689) <= a and not b;
    layer1_outputs(1690) <= a and not b;
    layer1_outputs(1691) <= a xor b;
    layer1_outputs(1692) <= b and not a;
    layer1_outputs(1693) <= not a;
    layer1_outputs(1694) <= not b;
    layer1_outputs(1695) <= not a;
    layer1_outputs(1696) <= not b;
    layer1_outputs(1697) <= not (a and b);
    layer1_outputs(1698) <= not b or a;
    layer1_outputs(1699) <= not b;
    layer1_outputs(1700) <= a and b;
    layer1_outputs(1701) <= not a or b;
    layer1_outputs(1702) <= not a;
    layer1_outputs(1703) <= '1';
    layer1_outputs(1704) <= a xor b;
    layer1_outputs(1705) <= not b or a;
    layer1_outputs(1706) <= b and not a;
    layer1_outputs(1707) <= b and not a;
    layer1_outputs(1708) <= b;
    layer1_outputs(1709) <= '0';
    layer1_outputs(1710) <= not b;
    layer1_outputs(1711) <= not b or a;
    layer1_outputs(1712) <= not a or b;
    layer1_outputs(1713) <= not (a or b);
    layer1_outputs(1714) <= a and not b;
    layer1_outputs(1715) <= not b;
    layer1_outputs(1716) <= b and not a;
    layer1_outputs(1717) <= not b;
    layer1_outputs(1718) <= not b;
    layer1_outputs(1719) <= a and not b;
    layer1_outputs(1720) <= not b;
    layer1_outputs(1721) <= not b or a;
    layer1_outputs(1722) <= not b or a;
    layer1_outputs(1723) <= a xor b;
    layer1_outputs(1724) <= a and not b;
    layer1_outputs(1725) <= not b or a;
    layer1_outputs(1726) <= b and not a;
    layer1_outputs(1727) <= a xor b;
    layer1_outputs(1728) <= not a or b;
    layer1_outputs(1729) <= a and b;
    layer1_outputs(1730) <= not (a and b);
    layer1_outputs(1731) <= a or b;
    layer1_outputs(1732) <= not (a and b);
    layer1_outputs(1733) <= '0';
    layer1_outputs(1734) <= not b;
    layer1_outputs(1735) <= b and not a;
    layer1_outputs(1736) <= not b or a;
    layer1_outputs(1737) <= '0';
    layer1_outputs(1738) <= a and b;
    layer1_outputs(1739) <= '1';
    layer1_outputs(1740) <= not a;
    layer1_outputs(1741) <= not (a xor b);
    layer1_outputs(1742) <= b and not a;
    layer1_outputs(1743) <= not a or b;
    layer1_outputs(1744) <= b and not a;
    layer1_outputs(1745) <= a and not b;
    layer1_outputs(1746) <= not (a and b);
    layer1_outputs(1747) <= a and b;
    layer1_outputs(1748) <= a and b;
    layer1_outputs(1749) <= a or b;
    layer1_outputs(1750) <= not (a or b);
    layer1_outputs(1751) <= a or b;
    layer1_outputs(1752) <= '1';
    layer1_outputs(1753) <= a and b;
    layer1_outputs(1754) <= not a or b;
    layer1_outputs(1755) <= not b or a;
    layer1_outputs(1756) <= not (a and b);
    layer1_outputs(1757) <= not b;
    layer1_outputs(1758) <= not a or b;
    layer1_outputs(1759) <= a;
    layer1_outputs(1760) <= b;
    layer1_outputs(1761) <= b and not a;
    layer1_outputs(1762) <= a;
    layer1_outputs(1763) <= not (a or b);
    layer1_outputs(1764) <= a xor b;
    layer1_outputs(1765) <= a and not b;
    layer1_outputs(1766) <= a and b;
    layer1_outputs(1767) <= not a or b;
    layer1_outputs(1768) <= not (a or b);
    layer1_outputs(1769) <= not b;
    layer1_outputs(1770) <= a;
    layer1_outputs(1771) <= '0';
    layer1_outputs(1772) <= b;
    layer1_outputs(1773) <= not a or b;
    layer1_outputs(1774) <= a or b;
    layer1_outputs(1775) <= '0';
    layer1_outputs(1776) <= not b;
    layer1_outputs(1777) <= '1';
    layer1_outputs(1778) <= a;
    layer1_outputs(1779) <= not (a and b);
    layer1_outputs(1780) <= '0';
    layer1_outputs(1781) <= not a;
    layer1_outputs(1782) <= '1';
    layer1_outputs(1783) <= a and b;
    layer1_outputs(1784) <= b and not a;
    layer1_outputs(1785) <= not a;
    layer1_outputs(1786) <= not a;
    layer1_outputs(1787) <= not b;
    layer1_outputs(1788) <= a xor b;
    layer1_outputs(1789) <= not (a and b);
    layer1_outputs(1790) <= a and not b;
    layer1_outputs(1791) <= a or b;
    layer1_outputs(1792) <= a or b;
    layer1_outputs(1793) <= b and not a;
    layer1_outputs(1794) <= not a;
    layer1_outputs(1795) <= not b or a;
    layer1_outputs(1796) <= not (a or b);
    layer1_outputs(1797) <= a and not b;
    layer1_outputs(1798) <= b and not a;
    layer1_outputs(1799) <= '1';
    layer1_outputs(1800) <= not (a or b);
    layer1_outputs(1801) <= a xor b;
    layer1_outputs(1802) <= not b;
    layer1_outputs(1803) <= a xor b;
    layer1_outputs(1804) <= a;
    layer1_outputs(1805) <= a or b;
    layer1_outputs(1806) <= a or b;
    layer1_outputs(1807) <= b;
    layer1_outputs(1808) <= a or b;
    layer1_outputs(1809) <= not a;
    layer1_outputs(1810) <= a;
    layer1_outputs(1811) <= b;
    layer1_outputs(1812) <= '0';
    layer1_outputs(1813) <= not a;
    layer1_outputs(1814) <= a and not b;
    layer1_outputs(1815) <= a;
    layer1_outputs(1816) <= not a or b;
    layer1_outputs(1817) <= '1';
    layer1_outputs(1818) <= not (a xor b);
    layer1_outputs(1819) <= not (a xor b);
    layer1_outputs(1820) <= b and not a;
    layer1_outputs(1821) <= not a or b;
    layer1_outputs(1822) <= not a;
    layer1_outputs(1823) <= not a or b;
    layer1_outputs(1824) <= not a;
    layer1_outputs(1825) <= b and not a;
    layer1_outputs(1826) <= a and not b;
    layer1_outputs(1827) <= not (a or b);
    layer1_outputs(1828) <= not a or b;
    layer1_outputs(1829) <= '0';
    layer1_outputs(1830) <= not b;
    layer1_outputs(1831) <= not b;
    layer1_outputs(1832) <= not b;
    layer1_outputs(1833) <= b and not a;
    layer1_outputs(1834) <= not (a and b);
    layer1_outputs(1835) <= b;
    layer1_outputs(1836) <= b;
    layer1_outputs(1837) <= a and b;
    layer1_outputs(1838) <= b and not a;
    layer1_outputs(1839) <= a;
    layer1_outputs(1840) <= not (a and b);
    layer1_outputs(1841) <= not b or a;
    layer1_outputs(1842) <= a xor b;
    layer1_outputs(1843) <= not (a and b);
    layer1_outputs(1844) <= a;
    layer1_outputs(1845) <= not (a or b);
    layer1_outputs(1846) <= a or b;
    layer1_outputs(1847) <= b and not a;
    layer1_outputs(1848) <= a;
    layer1_outputs(1849) <= not (a or b);
    layer1_outputs(1850) <= '0';
    layer1_outputs(1851) <= not a or b;
    layer1_outputs(1852) <= b;
    layer1_outputs(1853) <= b and not a;
    layer1_outputs(1854) <= a;
    layer1_outputs(1855) <= a and b;
    layer1_outputs(1856) <= '1';
    layer1_outputs(1857) <= not (a and b);
    layer1_outputs(1858) <= not b or a;
    layer1_outputs(1859) <= a and b;
    layer1_outputs(1860) <= b;
    layer1_outputs(1861) <= not (a or b);
    layer1_outputs(1862) <= not (a and b);
    layer1_outputs(1863) <= b;
    layer1_outputs(1864) <= b and not a;
    layer1_outputs(1865) <= not (a and b);
    layer1_outputs(1866) <= '1';
    layer1_outputs(1867) <= b;
    layer1_outputs(1868) <= not (a or b);
    layer1_outputs(1869) <= b;
    layer1_outputs(1870) <= '0';
    layer1_outputs(1871) <= not (a and b);
    layer1_outputs(1872) <= b;
    layer1_outputs(1873) <= a;
    layer1_outputs(1874) <= not (a or b);
    layer1_outputs(1875) <= a and b;
    layer1_outputs(1876) <= not a;
    layer1_outputs(1877) <= a;
    layer1_outputs(1878) <= not b or a;
    layer1_outputs(1879) <= not b;
    layer1_outputs(1880) <= not b;
    layer1_outputs(1881) <= a or b;
    layer1_outputs(1882) <= not a or b;
    layer1_outputs(1883) <= b;
    layer1_outputs(1884) <= not (a and b);
    layer1_outputs(1885) <= not (a and b);
    layer1_outputs(1886) <= '0';
    layer1_outputs(1887) <= a and not b;
    layer1_outputs(1888) <= not b or a;
    layer1_outputs(1889) <= a;
    layer1_outputs(1890) <= not a;
    layer1_outputs(1891) <= not b or a;
    layer1_outputs(1892) <= a and not b;
    layer1_outputs(1893) <= not a or b;
    layer1_outputs(1894) <= a or b;
    layer1_outputs(1895) <= b and not a;
    layer1_outputs(1896) <= a;
    layer1_outputs(1897) <= not b or a;
    layer1_outputs(1898) <= '1';
    layer1_outputs(1899) <= '0';
    layer1_outputs(1900) <= a or b;
    layer1_outputs(1901) <= not b;
    layer1_outputs(1902) <= not b or a;
    layer1_outputs(1903) <= not (a or b);
    layer1_outputs(1904) <= '1';
    layer1_outputs(1905) <= not (a xor b);
    layer1_outputs(1906) <= not a;
    layer1_outputs(1907) <= a or b;
    layer1_outputs(1908) <= b;
    layer1_outputs(1909) <= not a;
    layer1_outputs(1910) <= '1';
    layer1_outputs(1911) <= not (a and b);
    layer1_outputs(1912) <= '0';
    layer1_outputs(1913) <= a;
    layer1_outputs(1914) <= b and not a;
    layer1_outputs(1915) <= not b or a;
    layer1_outputs(1916) <= a and not b;
    layer1_outputs(1917) <= not b or a;
    layer1_outputs(1918) <= not b or a;
    layer1_outputs(1919) <= a;
    layer1_outputs(1920) <= b;
    layer1_outputs(1921) <= not a or b;
    layer1_outputs(1922) <= not (a xor b);
    layer1_outputs(1923) <= not a;
    layer1_outputs(1924) <= b;
    layer1_outputs(1925) <= '0';
    layer1_outputs(1926) <= a;
    layer1_outputs(1927) <= not (a and b);
    layer1_outputs(1928) <= not a;
    layer1_outputs(1929) <= not a;
    layer1_outputs(1930) <= not b or a;
    layer1_outputs(1931) <= not (a xor b);
    layer1_outputs(1932) <= '0';
    layer1_outputs(1933) <= a;
    layer1_outputs(1934) <= not b or a;
    layer1_outputs(1935) <= not a;
    layer1_outputs(1936) <= a;
    layer1_outputs(1937) <= a xor b;
    layer1_outputs(1938) <= not b or a;
    layer1_outputs(1939) <= not a or b;
    layer1_outputs(1940) <= not a;
    layer1_outputs(1941) <= not (a xor b);
    layer1_outputs(1942) <= a;
    layer1_outputs(1943) <= not (a and b);
    layer1_outputs(1944) <= not b;
    layer1_outputs(1945) <= not (a or b);
    layer1_outputs(1946) <= a xor b;
    layer1_outputs(1947) <= not a;
    layer1_outputs(1948) <= a and not b;
    layer1_outputs(1949) <= '1';
    layer1_outputs(1950) <= not a;
    layer1_outputs(1951) <= not a;
    layer1_outputs(1952) <= not a or b;
    layer1_outputs(1953) <= not (a or b);
    layer1_outputs(1954) <= a or b;
    layer1_outputs(1955) <= a or b;
    layer1_outputs(1956) <= a and not b;
    layer1_outputs(1957) <= a and b;
    layer1_outputs(1958) <= b;
    layer1_outputs(1959) <= a and not b;
    layer1_outputs(1960) <= a and b;
    layer1_outputs(1961) <= not a;
    layer1_outputs(1962) <= not a or b;
    layer1_outputs(1963) <= '0';
    layer1_outputs(1964) <= not a;
    layer1_outputs(1965) <= not (a or b);
    layer1_outputs(1966) <= b;
    layer1_outputs(1967) <= not b;
    layer1_outputs(1968) <= a;
    layer1_outputs(1969) <= '0';
    layer1_outputs(1970) <= b and not a;
    layer1_outputs(1971) <= a and not b;
    layer1_outputs(1972) <= not a or b;
    layer1_outputs(1973) <= a and not b;
    layer1_outputs(1974) <= '1';
    layer1_outputs(1975) <= b;
    layer1_outputs(1976) <= b and not a;
    layer1_outputs(1977) <= not b or a;
    layer1_outputs(1978) <= not (a or b);
    layer1_outputs(1979) <= not (a and b);
    layer1_outputs(1980) <= not (a and b);
    layer1_outputs(1981) <= a;
    layer1_outputs(1982) <= a and not b;
    layer1_outputs(1983) <= not b or a;
    layer1_outputs(1984) <= '0';
    layer1_outputs(1985) <= b and not a;
    layer1_outputs(1986) <= not b;
    layer1_outputs(1987) <= not (a and b);
    layer1_outputs(1988) <= '0';
    layer1_outputs(1989) <= not b or a;
    layer1_outputs(1990) <= a and not b;
    layer1_outputs(1991) <= '0';
    layer1_outputs(1992) <= not b;
    layer1_outputs(1993) <= b and not a;
    layer1_outputs(1994) <= not b or a;
    layer1_outputs(1995) <= not a or b;
    layer1_outputs(1996) <= a;
    layer1_outputs(1997) <= a and not b;
    layer1_outputs(1998) <= a or b;
    layer1_outputs(1999) <= a xor b;
    layer1_outputs(2000) <= '1';
    layer1_outputs(2001) <= a or b;
    layer1_outputs(2002) <= not b or a;
    layer1_outputs(2003) <= not b;
    layer1_outputs(2004) <= not b;
    layer1_outputs(2005) <= not b;
    layer1_outputs(2006) <= not a;
    layer1_outputs(2007) <= not (a or b);
    layer1_outputs(2008) <= a and b;
    layer1_outputs(2009) <= b;
    layer1_outputs(2010) <= '1';
    layer1_outputs(2011) <= b;
    layer1_outputs(2012) <= not (a xor b);
    layer1_outputs(2013) <= '0';
    layer1_outputs(2014) <= '1';
    layer1_outputs(2015) <= not a or b;
    layer1_outputs(2016) <= '1';
    layer1_outputs(2017) <= a or b;
    layer1_outputs(2018) <= a xor b;
    layer1_outputs(2019) <= not a;
    layer1_outputs(2020) <= '0';
    layer1_outputs(2021) <= b;
    layer1_outputs(2022) <= not b or a;
    layer1_outputs(2023) <= '0';
    layer1_outputs(2024) <= b and not a;
    layer1_outputs(2025) <= a xor b;
    layer1_outputs(2026) <= not a or b;
    layer1_outputs(2027) <= a or b;
    layer1_outputs(2028) <= b;
    layer1_outputs(2029) <= not b or a;
    layer1_outputs(2030) <= not a or b;
    layer1_outputs(2031) <= a or b;
    layer1_outputs(2032) <= '1';
    layer1_outputs(2033) <= not (a or b);
    layer1_outputs(2034) <= not a or b;
    layer1_outputs(2035) <= not a;
    layer1_outputs(2036) <= '0';
    layer1_outputs(2037) <= not a;
    layer1_outputs(2038) <= a and not b;
    layer1_outputs(2039) <= not a;
    layer1_outputs(2040) <= not a;
    layer1_outputs(2041) <= not a;
    layer1_outputs(2042) <= not a;
    layer1_outputs(2043) <= '0';
    layer1_outputs(2044) <= '0';
    layer1_outputs(2045) <= a xor b;
    layer1_outputs(2046) <= not a;
    layer1_outputs(2047) <= '1';
    layer1_outputs(2048) <= not (a xor b);
    layer1_outputs(2049) <= not a;
    layer1_outputs(2050) <= not a;
    layer1_outputs(2051) <= a and b;
    layer1_outputs(2052) <= a;
    layer1_outputs(2053) <= not (a xor b);
    layer1_outputs(2054) <= not a or b;
    layer1_outputs(2055) <= '0';
    layer1_outputs(2056) <= not (a or b);
    layer1_outputs(2057) <= a and b;
    layer1_outputs(2058) <= not a or b;
    layer1_outputs(2059) <= a xor b;
    layer1_outputs(2060) <= b and not a;
    layer1_outputs(2061) <= '0';
    layer1_outputs(2062) <= not (a xor b);
    layer1_outputs(2063) <= not b;
    layer1_outputs(2064) <= b and not a;
    layer1_outputs(2065) <= not (a and b);
    layer1_outputs(2066) <= a and not b;
    layer1_outputs(2067) <= a or b;
    layer1_outputs(2068) <= not (a and b);
    layer1_outputs(2069) <= not b;
    layer1_outputs(2070) <= a;
    layer1_outputs(2071) <= a and not b;
    layer1_outputs(2072) <= '0';
    layer1_outputs(2073) <= a and not b;
    layer1_outputs(2074) <= b and not a;
    layer1_outputs(2075) <= not (a or b);
    layer1_outputs(2076) <= b and not a;
    layer1_outputs(2077) <= a and b;
    layer1_outputs(2078) <= a;
    layer1_outputs(2079) <= not b;
    layer1_outputs(2080) <= b and not a;
    layer1_outputs(2081) <= not a or b;
    layer1_outputs(2082) <= a;
    layer1_outputs(2083) <= '0';
    layer1_outputs(2084) <= not (a xor b);
    layer1_outputs(2085) <= not b or a;
    layer1_outputs(2086) <= not b or a;
    layer1_outputs(2087) <= not a or b;
    layer1_outputs(2088) <= b and not a;
    layer1_outputs(2089) <= a and b;
    layer1_outputs(2090) <= not b;
    layer1_outputs(2091) <= b and not a;
    layer1_outputs(2092) <= not (a or b);
    layer1_outputs(2093) <= a xor b;
    layer1_outputs(2094) <= not (a and b);
    layer1_outputs(2095) <= not b;
    layer1_outputs(2096) <= a and b;
    layer1_outputs(2097) <= a xor b;
    layer1_outputs(2098) <= a and not b;
    layer1_outputs(2099) <= a and not b;
    layer1_outputs(2100) <= not (a xor b);
    layer1_outputs(2101) <= not a;
    layer1_outputs(2102) <= '0';
    layer1_outputs(2103) <= b and not a;
    layer1_outputs(2104) <= not a or b;
    layer1_outputs(2105) <= not b;
    layer1_outputs(2106) <= a;
    layer1_outputs(2107) <= a xor b;
    layer1_outputs(2108) <= not a or b;
    layer1_outputs(2109) <= a and b;
    layer1_outputs(2110) <= a or b;
    layer1_outputs(2111) <= '1';
    layer1_outputs(2112) <= not a or b;
    layer1_outputs(2113) <= a and b;
    layer1_outputs(2114) <= a and not b;
    layer1_outputs(2115) <= b and not a;
    layer1_outputs(2116) <= not b or a;
    layer1_outputs(2117) <= not b;
    layer1_outputs(2118) <= a or b;
    layer1_outputs(2119) <= a and b;
    layer1_outputs(2120) <= a and b;
    layer1_outputs(2121) <= not b or a;
    layer1_outputs(2122) <= not b;
    layer1_outputs(2123) <= a xor b;
    layer1_outputs(2124) <= a;
    layer1_outputs(2125) <= b;
    layer1_outputs(2126) <= not (a and b);
    layer1_outputs(2127) <= a;
    layer1_outputs(2128) <= not a;
    layer1_outputs(2129) <= b and not a;
    layer1_outputs(2130) <= not b;
    layer1_outputs(2131) <= not a or b;
    layer1_outputs(2132) <= not a or b;
    layer1_outputs(2133) <= b and not a;
    layer1_outputs(2134) <= b and not a;
    layer1_outputs(2135) <= '0';
    layer1_outputs(2136) <= not b;
    layer1_outputs(2137) <= '1';
    layer1_outputs(2138) <= not b;
    layer1_outputs(2139) <= not a or b;
    layer1_outputs(2140) <= not (a and b);
    layer1_outputs(2141) <= b;
    layer1_outputs(2142) <= not a;
    layer1_outputs(2143) <= not b;
    layer1_outputs(2144) <= not (a or b);
    layer1_outputs(2145) <= b;
    layer1_outputs(2146) <= not b;
    layer1_outputs(2147) <= a and not b;
    layer1_outputs(2148) <= not a or b;
    layer1_outputs(2149) <= not b or a;
    layer1_outputs(2150) <= not a or b;
    layer1_outputs(2151) <= b;
    layer1_outputs(2152) <= not (a and b);
    layer1_outputs(2153) <= a or b;
    layer1_outputs(2154) <= a or b;
    layer1_outputs(2155) <= '1';
    layer1_outputs(2156) <= a xor b;
    layer1_outputs(2157) <= not b or a;
    layer1_outputs(2158) <= a;
    layer1_outputs(2159) <= not (a and b);
    layer1_outputs(2160) <= a and not b;
    layer1_outputs(2161) <= a xor b;
    layer1_outputs(2162) <= not (a or b);
    layer1_outputs(2163) <= a and b;
    layer1_outputs(2164) <= b and not a;
    layer1_outputs(2165) <= not a or b;
    layer1_outputs(2166) <= a xor b;
    layer1_outputs(2167) <= a or b;
    layer1_outputs(2168) <= not b or a;
    layer1_outputs(2169) <= a and b;
    layer1_outputs(2170) <= not b;
    layer1_outputs(2171) <= '1';
    layer1_outputs(2172) <= not a or b;
    layer1_outputs(2173) <= a and not b;
    layer1_outputs(2174) <= a and b;
    layer1_outputs(2175) <= not a;
    layer1_outputs(2176) <= a or b;
    layer1_outputs(2177) <= not (a or b);
    layer1_outputs(2178) <= not (a and b);
    layer1_outputs(2179) <= '0';
    layer1_outputs(2180) <= not b;
    layer1_outputs(2181) <= a and b;
    layer1_outputs(2182) <= '0';
    layer1_outputs(2183) <= '1';
    layer1_outputs(2184) <= a and not b;
    layer1_outputs(2185) <= not (a or b);
    layer1_outputs(2186) <= a or b;
    layer1_outputs(2187) <= a xor b;
    layer1_outputs(2188) <= b and not a;
    layer1_outputs(2189) <= a or b;
    layer1_outputs(2190) <= a or b;
    layer1_outputs(2191) <= not (a and b);
    layer1_outputs(2192) <= not b;
    layer1_outputs(2193) <= not (a and b);
    layer1_outputs(2194) <= not (a and b);
    layer1_outputs(2195) <= b and not a;
    layer1_outputs(2196) <= '1';
    layer1_outputs(2197) <= b;
    layer1_outputs(2198) <= b and not a;
    layer1_outputs(2199) <= '0';
    layer1_outputs(2200) <= b;
    layer1_outputs(2201) <= not a;
    layer1_outputs(2202) <= not a;
    layer1_outputs(2203) <= '0';
    layer1_outputs(2204) <= not (a or b);
    layer1_outputs(2205) <= b;
    layer1_outputs(2206) <= a and b;
    layer1_outputs(2207) <= a and b;
    layer1_outputs(2208) <= not (a and b);
    layer1_outputs(2209) <= not b;
    layer1_outputs(2210) <= a and not b;
    layer1_outputs(2211) <= not (a xor b);
    layer1_outputs(2212) <= not a or b;
    layer1_outputs(2213) <= b and not a;
    layer1_outputs(2214) <= not b or a;
    layer1_outputs(2215) <= a and b;
    layer1_outputs(2216) <= not a or b;
    layer1_outputs(2217) <= not a;
    layer1_outputs(2218) <= not b or a;
    layer1_outputs(2219) <= '0';
    layer1_outputs(2220) <= not a;
    layer1_outputs(2221) <= a and not b;
    layer1_outputs(2222) <= not b;
    layer1_outputs(2223) <= a or b;
    layer1_outputs(2224) <= not a;
    layer1_outputs(2225) <= not a;
    layer1_outputs(2226) <= a or b;
    layer1_outputs(2227) <= '1';
    layer1_outputs(2228) <= a;
    layer1_outputs(2229) <= '1';
    layer1_outputs(2230) <= b;
    layer1_outputs(2231) <= not a or b;
    layer1_outputs(2232) <= not (a and b);
    layer1_outputs(2233) <= a xor b;
    layer1_outputs(2234) <= a and b;
    layer1_outputs(2235) <= a and not b;
    layer1_outputs(2236) <= not b;
    layer1_outputs(2237) <= not a or b;
    layer1_outputs(2238) <= a;
    layer1_outputs(2239) <= a;
    layer1_outputs(2240) <= a and not b;
    layer1_outputs(2241) <= not (a and b);
    layer1_outputs(2242) <= '1';
    layer1_outputs(2243) <= not b or a;
    layer1_outputs(2244) <= '1';
    layer1_outputs(2245) <= not b or a;
    layer1_outputs(2246) <= not b;
    layer1_outputs(2247) <= not (a or b);
    layer1_outputs(2248) <= a or b;
    layer1_outputs(2249) <= not a;
    layer1_outputs(2250) <= not (a or b);
    layer1_outputs(2251) <= a and b;
    layer1_outputs(2252) <= '1';
    layer1_outputs(2253) <= b;
    layer1_outputs(2254) <= not b;
    layer1_outputs(2255) <= a or b;
    layer1_outputs(2256) <= not a;
    layer1_outputs(2257) <= not a or b;
    layer1_outputs(2258) <= not a or b;
    layer1_outputs(2259) <= not b;
    layer1_outputs(2260) <= '1';
    layer1_outputs(2261) <= a;
    layer1_outputs(2262) <= a and not b;
    layer1_outputs(2263) <= '1';
    layer1_outputs(2264) <= '1';
    layer1_outputs(2265) <= not (a and b);
    layer1_outputs(2266) <= not (a and b);
    layer1_outputs(2267) <= a;
    layer1_outputs(2268) <= not b;
    layer1_outputs(2269) <= not (a or b);
    layer1_outputs(2270) <= not b or a;
    layer1_outputs(2271) <= not a or b;
    layer1_outputs(2272) <= not (a xor b);
    layer1_outputs(2273) <= not (a xor b);
    layer1_outputs(2274) <= not (a and b);
    layer1_outputs(2275) <= b and not a;
    layer1_outputs(2276) <= a;
    layer1_outputs(2277) <= a or b;
    layer1_outputs(2278) <= b and not a;
    layer1_outputs(2279) <= b and not a;
    layer1_outputs(2280) <= not a;
    layer1_outputs(2281) <= not a;
    layer1_outputs(2282) <= not (a or b);
    layer1_outputs(2283) <= not a;
    layer1_outputs(2284) <= not (a or b);
    layer1_outputs(2285) <= '1';
    layer1_outputs(2286) <= a or b;
    layer1_outputs(2287) <= not b;
    layer1_outputs(2288) <= a and not b;
    layer1_outputs(2289) <= not b;
    layer1_outputs(2290) <= a or b;
    layer1_outputs(2291) <= '0';
    layer1_outputs(2292) <= '0';
    layer1_outputs(2293) <= not a or b;
    layer1_outputs(2294) <= not a;
    layer1_outputs(2295) <= not a;
    layer1_outputs(2296) <= not b;
    layer1_outputs(2297) <= not a;
    layer1_outputs(2298) <= b;
    layer1_outputs(2299) <= a or b;
    layer1_outputs(2300) <= b;
    layer1_outputs(2301) <= a xor b;
    layer1_outputs(2302) <= b and not a;
    layer1_outputs(2303) <= not (a and b);
    layer1_outputs(2304) <= b and not a;
    layer1_outputs(2305) <= not a or b;
    layer1_outputs(2306) <= '0';
    layer1_outputs(2307) <= b and not a;
    layer1_outputs(2308) <= '1';
    layer1_outputs(2309) <= a and b;
    layer1_outputs(2310) <= not (a or b);
    layer1_outputs(2311) <= b;
    layer1_outputs(2312) <= not (a and b);
    layer1_outputs(2313) <= '0';
    layer1_outputs(2314) <= '0';
    layer1_outputs(2315) <= not (a xor b);
    layer1_outputs(2316) <= not (a or b);
    layer1_outputs(2317) <= a or b;
    layer1_outputs(2318) <= not b;
    layer1_outputs(2319) <= '1';
    layer1_outputs(2320) <= not a or b;
    layer1_outputs(2321) <= not (a or b);
    layer1_outputs(2322) <= not b or a;
    layer1_outputs(2323) <= a and b;
    layer1_outputs(2324) <= a;
    layer1_outputs(2325) <= not a;
    layer1_outputs(2326) <= not (a and b);
    layer1_outputs(2327) <= a;
    layer1_outputs(2328) <= not a or b;
    layer1_outputs(2329) <= '1';
    layer1_outputs(2330) <= a and not b;
    layer1_outputs(2331) <= a and b;
    layer1_outputs(2332) <= not b;
    layer1_outputs(2333) <= b and not a;
    layer1_outputs(2334) <= not b or a;
    layer1_outputs(2335) <= not a;
    layer1_outputs(2336) <= not (a xor b);
    layer1_outputs(2337) <= a xor b;
    layer1_outputs(2338) <= a and b;
    layer1_outputs(2339) <= not (a and b);
    layer1_outputs(2340) <= a and b;
    layer1_outputs(2341) <= a xor b;
    layer1_outputs(2342) <= not a;
    layer1_outputs(2343) <= not a;
    layer1_outputs(2344) <= not a;
    layer1_outputs(2345) <= not a;
    layer1_outputs(2346) <= b;
    layer1_outputs(2347) <= a xor b;
    layer1_outputs(2348) <= not a;
    layer1_outputs(2349) <= not b;
    layer1_outputs(2350) <= '0';
    layer1_outputs(2351) <= not b;
    layer1_outputs(2352) <= b and not a;
    layer1_outputs(2353) <= not (a xor b);
    layer1_outputs(2354) <= a;
    layer1_outputs(2355) <= not a or b;
    layer1_outputs(2356) <= b;
    layer1_outputs(2357) <= not b;
    layer1_outputs(2358) <= '0';
    layer1_outputs(2359) <= not (a or b);
    layer1_outputs(2360) <= a and b;
    layer1_outputs(2361) <= '1';
    layer1_outputs(2362) <= not b or a;
    layer1_outputs(2363) <= not b or a;
    layer1_outputs(2364) <= not (a or b);
    layer1_outputs(2365) <= not (a or b);
    layer1_outputs(2366) <= b;
    layer1_outputs(2367) <= a;
    layer1_outputs(2368) <= '0';
    layer1_outputs(2369) <= not (a and b);
    layer1_outputs(2370) <= a and b;
    layer1_outputs(2371) <= a and not b;
    layer1_outputs(2372) <= '1';
    layer1_outputs(2373) <= b and not a;
    layer1_outputs(2374) <= not (a or b);
    layer1_outputs(2375) <= not b or a;
    layer1_outputs(2376) <= not (a and b);
    layer1_outputs(2377) <= not b or a;
    layer1_outputs(2378) <= not (a and b);
    layer1_outputs(2379) <= not b;
    layer1_outputs(2380) <= a xor b;
    layer1_outputs(2381) <= '0';
    layer1_outputs(2382) <= not b;
    layer1_outputs(2383) <= '1';
    layer1_outputs(2384) <= not b;
    layer1_outputs(2385) <= not (a or b);
    layer1_outputs(2386) <= not b;
    layer1_outputs(2387) <= not (a or b);
    layer1_outputs(2388) <= a;
    layer1_outputs(2389) <= a;
    layer1_outputs(2390) <= not b or a;
    layer1_outputs(2391) <= not b;
    layer1_outputs(2392) <= not (a or b);
    layer1_outputs(2393) <= not a;
    layer1_outputs(2394) <= a;
    layer1_outputs(2395) <= not b;
    layer1_outputs(2396) <= a and not b;
    layer1_outputs(2397) <= a and not b;
    layer1_outputs(2398) <= not (a or b);
    layer1_outputs(2399) <= not (a and b);
    layer1_outputs(2400) <= not (a or b);
    layer1_outputs(2401) <= b and not a;
    layer1_outputs(2402) <= not a;
    layer1_outputs(2403) <= a or b;
    layer1_outputs(2404) <= not (a or b);
    layer1_outputs(2405) <= not b;
    layer1_outputs(2406) <= a xor b;
    layer1_outputs(2407) <= not b or a;
    layer1_outputs(2408) <= a and b;
    layer1_outputs(2409) <= b;
    layer1_outputs(2410) <= not a;
    layer1_outputs(2411) <= not b;
    layer1_outputs(2412) <= not b;
    layer1_outputs(2413) <= not a;
    layer1_outputs(2414) <= b;
    layer1_outputs(2415) <= not (a and b);
    layer1_outputs(2416) <= '1';
    layer1_outputs(2417) <= b;
    layer1_outputs(2418) <= a and not b;
    layer1_outputs(2419) <= not (a and b);
    layer1_outputs(2420) <= not a;
    layer1_outputs(2421) <= '1';
    layer1_outputs(2422) <= not a;
    layer1_outputs(2423) <= a and not b;
    layer1_outputs(2424) <= a;
    layer1_outputs(2425) <= '0';
    layer1_outputs(2426) <= not b;
    layer1_outputs(2427) <= not a;
    layer1_outputs(2428) <= '1';
    layer1_outputs(2429) <= '1';
    layer1_outputs(2430) <= '1';
    layer1_outputs(2431) <= not (a or b);
    layer1_outputs(2432) <= a;
    layer1_outputs(2433) <= b;
    layer1_outputs(2434) <= b and not a;
    layer1_outputs(2435) <= '0';
    layer1_outputs(2436) <= a and not b;
    layer1_outputs(2437) <= not (a xor b);
    layer1_outputs(2438) <= not a;
    layer1_outputs(2439) <= a;
    layer1_outputs(2440) <= a and not b;
    layer1_outputs(2441) <= not b;
    layer1_outputs(2442) <= not b;
    layer1_outputs(2443) <= '0';
    layer1_outputs(2444) <= a;
    layer1_outputs(2445) <= not a;
    layer1_outputs(2446) <= not a or b;
    layer1_outputs(2447) <= not b;
    layer1_outputs(2448) <= not (a xor b);
    layer1_outputs(2449) <= a and not b;
    layer1_outputs(2450) <= not (a or b);
    layer1_outputs(2451) <= a and not b;
    layer1_outputs(2452) <= a;
    layer1_outputs(2453) <= '1';
    layer1_outputs(2454) <= not (a or b);
    layer1_outputs(2455) <= a;
    layer1_outputs(2456) <= not a or b;
    layer1_outputs(2457) <= a or b;
    layer1_outputs(2458) <= not b or a;
    layer1_outputs(2459) <= b and not a;
    layer1_outputs(2460) <= not b;
    layer1_outputs(2461) <= b and not a;
    layer1_outputs(2462) <= a and b;
    layer1_outputs(2463) <= b;
    layer1_outputs(2464) <= a;
    layer1_outputs(2465) <= not b;
    layer1_outputs(2466) <= a or b;
    layer1_outputs(2467) <= a;
    layer1_outputs(2468) <= b;
    layer1_outputs(2469) <= '0';
    layer1_outputs(2470) <= a;
    layer1_outputs(2471) <= a and not b;
    layer1_outputs(2472) <= not a;
    layer1_outputs(2473) <= b and not a;
    layer1_outputs(2474) <= '1';
    layer1_outputs(2475) <= not (a and b);
    layer1_outputs(2476) <= not a or b;
    layer1_outputs(2477) <= '0';
    layer1_outputs(2478) <= not a;
    layer1_outputs(2479) <= b;
    layer1_outputs(2480) <= a and not b;
    layer1_outputs(2481) <= a;
    layer1_outputs(2482) <= a;
    layer1_outputs(2483) <= '1';
    layer1_outputs(2484) <= a xor b;
    layer1_outputs(2485) <= a or b;
    layer1_outputs(2486) <= not (a and b);
    layer1_outputs(2487) <= not a;
    layer1_outputs(2488) <= not (a or b);
    layer1_outputs(2489) <= not (a or b);
    layer1_outputs(2490) <= not a or b;
    layer1_outputs(2491) <= not (a or b);
    layer1_outputs(2492) <= a xor b;
    layer1_outputs(2493) <= '0';
    layer1_outputs(2494) <= b;
    layer1_outputs(2495) <= '1';
    layer1_outputs(2496) <= b;
    layer1_outputs(2497) <= a and b;
    layer1_outputs(2498) <= b;
    layer1_outputs(2499) <= '1';
    layer1_outputs(2500) <= a or b;
    layer1_outputs(2501) <= not a or b;
    layer1_outputs(2502) <= b;
    layer1_outputs(2503) <= a and not b;
    layer1_outputs(2504) <= not b;
    layer1_outputs(2505) <= a or b;
    layer1_outputs(2506) <= b;
    layer1_outputs(2507) <= not b;
    layer1_outputs(2508) <= not (a or b);
    layer1_outputs(2509) <= a or b;
    layer1_outputs(2510) <= a or b;
    layer1_outputs(2511) <= b;
    layer1_outputs(2512) <= a or b;
    layer1_outputs(2513) <= '1';
    layer1_outputs(2514) <= b;
    layer1_outputs(2515) <= not b;
    layer1_outputs(2516) <= a or b;
    layer1_outputs(2517) <= not a or b;
    layer1_outputs(2518) <= '0';
    layer1_outputs(2519) <= a;
    layer1_outputs(2520) <= not b or a;
    layer1_outputs(2521) <= b;
    layer1_outputs(2522) <= a and not b;
    layer1_outputs(2523) <= not (a and b);
    layer1_outputs(2524) <= a;
    layer1_outputs(2525) <= not a or b;
    layer1_outputs(2526) <= a xor b;
    layer1_outputs(2527) <= not a;
    layer1_outputs(2528) <= not a or b;
    layer1_outputs(2529) <= a or b;
    layer1_outputs(2530) <= a and not b;
    layer1_outputs(2531) <= a and b;
    layer1_outputs(2532) <= a xor b;
    layer1_outputs(2533) <= not b;
    layer1_outputs(2534) <= '0';
    layer1_outputs(2535) <= b;
    layer1_outputs(2536) <= a or b;
    layer1_outputs(2537) <= not b;
    layer1_outputs(2538) <= not b;
    layer1_outputs(2539) <= b and not a;
    layer1_outputs(2540) <= not b or a;
    layer1_outputs(2541) <= not (a or b);
    layer1_outputs(2542) <= a or b;
    layer1_outputs(2543) <= not a;
    layer1_outputs(2544) <= a and not b;
    layer1_outputs(2545) <= a and b;
    layer1_outputs(2546) <= b and not a;
    layer1_outputs(2547) <= a and not b;
    layer1_outputs(2548) <= not (a and b);
    layer1_outputs(2549) <= b;
    layer1_outputs(2550) <= not b;
    layer1_outputs(2551) <= a or b;
    layer1_outputs(2552) <= a;
    layer1_outputs(2553) <= not b;
    layer1_outputs(2554) <= '0';
    layer1_outputs(2555) <= not a or b;
    layer1_outputs(2556) <= not a;
    layer1_outputs(2557) <= not b;
    layer1_outputs(2558) <= not b;
    layer1_outputs(2559) <= a or b;
    layer1_outputs(2560) <= not b or a;
    layer1_outputs(2561) <= a and b;
    layer1_outputs(2562) <= not b or a;
    layer1_outputs(2563) <= not b or a;
    layer1_outputs(2564) <= not b;
    layer1_outputs(2565) <= not a or b;
    layer1_outputs(2566) <= a or b;
    layer1_outputs(2567) <= a or b;
    layer1_outputs(2568) <= not b;
    layer1_outputs(2569) <= not a or b;
    layer1_outputs(2570) <= a and not b;
    layer1_outputs(2571) <= b;
    layer1_outputs(2572) <= b;
    layer1_outputs(2573) <= '1';
    layer1_outputs(2574) <= not (a xor b);
    layer1_outputs(2575) <= not a or b;
    layer1_outputs(2576) <= not b;
    layer1_outputs(2577) <= not (a or b);
    layer1_outputs(2578) <= not a;
    layer1_outputs(2579) <= not a or b;
    layer1_outputs(2580) <= a and b;
    layer1_outputs(2581) <= '0';
    layer1_outputs(2582) <= '0';
    layer1_outputs(2583) <= not a;
    layer1_outputs(2584) <= a or b;
    layer1_outputs(2585) <= not (a or b);
    layer1_outputs(2586) <= not (a and b);
    layer1_outputs(2587) <= b;
    layer1_outputs(2588) <= not b or a;
    layer1_outputs(2589) <= '1';
    layer1_outputs(2590) <= not (a xor b);
    layer1_outputs(2591) <= '1';
    layer1_outputs(2592) <= b;
    layer1_outputs(2593) <= not b;
    layer1_outputs(2594) <= not b or a;
    layer1_outputs(2595) <= not a or b;
    layer1_outputs(2596) <= not b or a;
    layer1_outputs(2597) <= a or b;
    layer1_outputs(2598) <= '1';
    layer1_outputs(2599) <= b and not a;
    layer1_outputs(2600) <= not (a and b);
    layer1_outputs(2601) <= not (a and b);
    layer1_outputs(2602) <= not b or a;
    layer1_outputs(2603) <= not a;
    layer1_outputs(2604) <= '1';
    layer1_outputs(2605) <= not b;
    layer1_outputs(2606) <= a and not b;
    layer1_outputs(2607) <= a;
    layer1_outputs(2608) <= a;
    layer1_outputs(2609) <= not (a xor b);
    layer1_outputs(2610) <= not b or a;
    layer1_outputs(2611) <= a and b;
    layer1_outputs(2612) <= a and b;
    layer1_outputs(2613) <= b and not a;
    layer1_outputs(2614) <= a and not b;
    layer1_outputs(2615) <= not (a and b);
    layer1_outputs(2616) <= not a or b;
    layer1_outputs(2617) <= a and b;
    layer1_outputs(2618) <= not a or b;
    layer1_outputs(2619) <= not (a or b);
    layer1_outputs(2620) <= b;
    layer1_outputs(2621) <= '0';
    layer1_outputs(2622) <= not (a or b);
    layer1_outputs(2623) <= not b or a;
    layer1_outputs(2624) <= a or b;
    layer1_outputs(2625) <= not b;
    layer1_outputs(2626) <= not a;
    layer1_outputs(2627) <= a;
    layer1_outputs(2628) <= a or b;
    layer1_outputs(2629) <= b;
    layer1_outputs(2630) <= not b or a;
    layer1_outputs(2631) <= a or b;
    layer1_outputs(2632) <= a and b;
    layer1_outputs(2633) <= not b;
    layer1_outputs(2634) <= not a or b;
    layer1_outputs(2635) <= not a;
    layer1_outputs(2636) <= not b;
    layer1_outputs(2637) <= a and b;
    layer1_outputs(2638) <= '1';
    layer1_outputs(2639) <= a or b;
    layer1_outputs(2640) <= not a;
    layer1_outputs(2641) <= not b;
    layer1_outputs(2642) <= b and not a;
    layer1_outputs(2643) <= not (a and b);
    layer1_outputs(2644) <= not b;
    layer1_outputs(2645) <= '0';
    layer1_outputs(2646) <= not (a or b);
    layer1_outputs(2647) <= not a;
    layer1_outputs(2648) <= not b or a;
    layer1_outputs(2649) <= a;
    layer1_outputs(2650) <= a or b;
    layer1_outputs(2651) <= a;
    layer1_outputs(2652) <= not (a or b);
    layer1_outputs(2653) <= not b;
    layer1_outputs(2654) <= not a or b;
    layer1_outputs(2655) <= not (a and b);
    layer1_outputs(2656) <= not (a and b);
    layer1_outputs(2657) <= not a;
    layer1_outputs(2658) <= not b or a;
    layer1_outputs(2659) <= not (a and b);
    layer1_outputs(2660) <= a;
    layer1_outputs(2661) <= a;
    layer1_outputs(2662) <= a;
    layer1_outputs(2663) <= b;
    layer1_outputs(2664) <= b and not a;
    layer1_outputs(2665) <= a and not b;
    layer1_outputs(2666) <= a;
    layer1_outputs(2667) <= b and not a;
    layer1_outputs(2668) <= a;
    layer1_outputs(2669) <= a and b;
    layer1_outputs(2670) <= not b or a;
    layer1_outputs(2671) <= a;
    layer1_outputs(2672) <= not (a and b);
    layer1_outputs(2673) <= not (a xor b);
    layer1_outputs(2674) <= not a or b;
    layer1_outputs(2675) <= b;
    layer1_outputs(2676) <= not a or b;
    layer1_outputs(2677) <= a;
    layer1_outputs(2678) <= a and not b;
    layer1_outputs(2679) <= b;
    layer1_outputs(2680) <= b;
    layer1_outputs(2681) <= '0';
    layer1_outputs(2682) <= not (a or b);
    layer1_outputs(2683) <= not b;
    layer1_outputs(2684) <= a;
    layer1_outputs(2685) <= not a or b;
    layer1_outputs(2686) <= '1';
    layer1_outputs(2687) <= not b;
    layer1_outputs(2688) <= a;
    layer1_outputs(2689) <= not b or a;
    layer1_outputs(2690) <= not (a or b);
    layer1_outputs(2691) <= a xor b;
    layer1_outputs(2692) <= a or b;
    layer1_outputs(2693) <= '0';
    layer1_outputs(2694) <= '1';
    layer1_outputs(2695) <= a or b;
    layer1_outputs(2696) <= a or b;
    layer1_outputs(2697) <= not (a and b);
    layer1_outputs(2698) <= not a or b;
    layer1_outputs(2699) <= not b or a;
    layer1_outputs(2700) <= a;
    layer1_outputs(2701) <= not (a or b);
    layer1_outputs(2702) <= b;
    layer1_outputs(2703) <= b and not a;
    layer1_outputs(2704) <= not (a xor b);
    layer1_outputs(2705) <= not (a or b);
    layer1_outputs(2706) <= '1';
    layer1_outputs(2707) <= not b or a;
    layer1_outputs(2708) <= a and not b;
    layer1_outputs(2709) <= '0';
    layer1_outputs(2710) <= b;
    layer1_outputs(2711) <= '1';
    layer1_outputs(2712) <= not (a and b);
    layer1_outputs(2713) <= a and not b;
    layer1_outputs(2714) <= not a;
    layer1_outputs(2715) <= not a or b;
    layer1_outputs(2716) <= not a;
    layer1_outputs(2717) <= '1';
    layer1_outputs(2718) <= b and not a;
    layer1_outputs(2719) <= not a;
    layer1_outputs(2720) <= b;
    layer1_outputs(2721) <= '1';
    layer1_outputs(2722) <= not (a xor b);
    layer1_outputs(2723) <= not (a xor b);
    layer1_outputs(2724) <= not b or a;
    layer1_outputs(2725) <= a and not b;
    layer1_outputs(2726) <= a;
    layer1_outputs(2727) <= not a;
    layer1_outputs(2728) <= a;
    layer1_outputs(2729) <= not a or b;
    layer1_outputs(2730) <= a;
    layer1_outputs(2731) <= not (a and b);
    layer1_outputs(2732) <= not a or b;
    layer1_outputs(2733) <= a and b;
    layer1_outputs(2734) <= a and not b;
    layer1_outputs(2735) <= a xor b;
    layer1_outputs(2736) <= a and not b;
    layer1_outputs(2737) <= a and b;
    layer1_outputs(2738) <= a and b;
    layer1_outputs(2739) <= '1';
    layer1_outputs(2740) <= a and b;
    layer1_outputs(2741) <= a;
    layer1_outputs(2742) <= not (a or b);
    layer1_outputs(2743) <= '1';
    layer1_outputs(2744) <= not (a or b);
    layer1_outputs(2745) <= a and b;
    layer1_outputs(2746) <= not a;
    layer1_outputs(2747) <= not a or b;
    layer1_outputs(2748) <= a or b;
    layer1_outputs(2749) <= a xor b;
    layer1_outputs(2750) <= '1';
    layer1_outputs(2751) <= not (a or b);
    layer1_outputs(2752) <= not (a and b);
    layer1_outputs(2753) <= a;
    layer1_outputs(2754) <= '1';
    layer1_outputs(2755) <= a;
    layer1_outputs(2756) <= not (a and b);
    layer1_outputs(2757) <= a;
    layer1_outputs(2758) <= a and not b;
    layer1_outputs(2759) <= b and not a;
    layer1_outputs(2760) <= a or b;
    layer1_outputs(2761) <= a or b;
    layer1_outputs(2762) <= '0';
    layer1_outputs(2763) <= b and not a;
    layer1_outputs(2764) <= b;
    layer1_outputs(2765) <= a and b;
    layer1_outputs(2766) <= a xor b;
    layer1_outputs(2767) <= not a;
    layer1_outputs(2768) <= not b;
    layer1_outputs(2769) <= '0';
    layer1_outputs(2770) <= not a or b;
    layer1_outputs(2771) <= b;
    layer1_outputs(2772) <= not (a xor b);
    layer1_outputs(2773) <= '0';
    layer1_outputs(2774) <= not (a and b);
    layer1_outputs(2775) <= '1';
    layer1_outputs(2776) <= b and not a;
    layer1_outputs(2777) <= not a or b;
    layer1_outputs(2778) <= '1';
    layer1_outputs(2779) <= not b;
    layer1_outputs(2780) <= '0';
    layer1_outputs(2781) <= b and not a;
    layer1_outputs(2782) <= not a;
    layer1_outputs(2783) <= not b or a;
    layer1_outputs(2784) <= not b or a;
    layer1_outputs(2785) <= b and not a;
    layer1_outputs(2786) <= not a;
    layer1_outputs(2787) <= not (a or b);
    layer1_outputs(2788) <= not b;
    layer1_outputs(2789) <= not b or a;
    layer1_outputs(2790) <= not b or a;
    layer1_outputs(2791) <= not (a or b);
    layer1_outputs(2792) <= a and not b;
    layer1_outputs(2793) <= not b or a;
    layer1_outputs(2794) <= a and b;
    layer1_outputs(2795) <= not (a and b);
    layer1_outputs(2796) <= not b;
    layer1_outputs(2797) <= a and b;
    layer1_outputs(2798) <= not (a xor b);
    layer1_outputs(2799) <= b;
    layer1_outputs(2800) <= a or b;
    layer1_outputs(2801) <= not b;
    layer1_outputs(2802) <= a;
    layer1_outputs(2803) <= b;
    layer1_outputs(2804) <= a;
    layer1_outputs(2805) <= a or b;
    layer1_outputs(2806) <= not a;
    layer1_outputs(2807) <= '1';
    layer1_outputs(2808) <= a or b;
    layer1_outputs(2809) <= not b;
    layer1_outputs(2810) <= not a;
    layer1_outputs(2811) <= not (a or b);
    layer1_outputs(2812) <= b and not a;
    layer1_outputs(2813) <= a or b;
    layer1_outputs(2814) <= a;
    layer1_outputs(2815) <= not b or a;
    layer1_outputs(2816) <= '1';
    layer1_outputs(2817) <= not (a xor b);
    layer1_outputs(2818) <= a or b;
    layer1_outputs(2819) <= not (a or b);
    layer1_outputs(2820) <= '0';
    layer1_outputs(2821) <= '1';
    layer1_outputs(2822) <= not a or b;
    layer1_outputs(2823) <= not (a xor b);
    layer1_outputs(2824) <= not a or b;
    layer1_outputs(2825) <= not (a or b);
    layer1_outputs(2826) <= b;
    layer1_outputs(2827) <= b and not a;
    layer1_outputs(2828) <= not b;
    layer1_outputs(2829) <= not b;
    layer1_outputs(2830) <= not b or a;
    layer1_outputs(2831) <= b and not a;
    layer1_outputs(2832) <= not b;
    layer1_outputs(2833) <= a xor b;
    layer1_outputs(2834) <= '0';
    layer1_outputs(2835) <= a;
    layer1_outputs(2836) <= a and b;
    layer1_outputs(2837) <= not a or b;
    layer1_outputs(2838) <= b;
    layer1_outputs(2839) <= '0';
    layer1_outputs(2840) <= a and b;
    layer1_outputs(2841) <= not a;
    layer1_outputs(2842) <= not a or b;
    layer1_outputs(2843) <= a;
    layer1_outputs(2844) <= not a or b;
    layer1_outputs(2845) <= not a;
    layer1_outputs(2846) <= '1';
    layer1_outputs(2847) <= not a;
    layer1_outputs(2848) <= a;
    layer1_outputs(2849) <= not b;
    layer1_outputs(2850) <= not b or a;
    layer1_outputs(2851) <= '1';
    layer1_outputs(2852) <= a and b;
    layer1_outputs(2853) <= a or b;
    layer1_outputs(2854) <= '1';
    layer1_outputs(2855) <= not a or b;
    layer1_outputs(2856) <= b and not a;
    layer1_outputs(2857) <= not (a and b);
    layer1_outputs(2858) <= a;
    layer1_outputs(2859) <= a or b;
    layer1_outputs(2860) <= not (a or b);
    layer1_outputs(2861) <= '0';
    layer1_outputs(2862) <= not a;
    layer1_outputs(2863) <= a or b;
    layer1_outputs(2864) <= b;
    layer1_outputs(2865) <= not a or b;
    layer1_outputs(2866) <= not b or a;
    layer1_outputs(2867) <= '1';
    layer1_outputs(2868) <= not (a and b);
    layer1_outputs(2869) <= a or b;
    layer1_outputs(2870) <= a xor b;
    layer1_outputs(2871) <= not a or b;
    layer1_outputs(2872) <= not (a or b);
    layer1_outputs(2873) <= not b;
    layer1_outputs(2874) <= '0';
    layer1_outputs(2875) <= b;
    layer1_outputs(2876) <= not b or a;
    layer1_outputs(2877) <= not a;
    layer1_outputs(2878) <= not a;
    layer1_outputs(2879) <= b and not a;
    layer1_outputs(2880) <= not a or b;
    layer1_outputs(2881) <= not (a and b);
    layer1_outputs(2882) <= '1';
    layer1_outputs(2883) <= b;
    layer1_outputs(2884) <= not b;
    layer1_outputs(2885) <= b;
    layer1_outputs(2886) <= a;
    layer1_outputs(2887) <= a and not b;
    layer1_outputs(2888) <= not (a and b);
    layer1_outputs(2889) <= a xor b;
    layer1_outputs(2890) <= not a;
    layer1_outputs(2891) <= not b;
    layer1_outputs(2892) <= not (a or b);
    layer1_outputs(2893) <= b and not a;
    layer1_outputs(2894) <= a;
    layer1_outputs(2895) <= not b or a;
    layer1_outputs(2896) <= not a;
    layer1_outputs(2897) <= not b;
    layer1_outputs(2898) <= not a or b;
    layer1_outputs(2899) <= b;
    layer1_outputs(2900) <= b;
    layer1_outputs(2901) <= b and not a;
    layer1_outputs(2902) <= not a;
    layer1_outputs(2903) <= '0';
    layer1_outputs(2904) <= not (a xor b);
    layer1_outputs(2905) <= not b;
    layer1_outputs(2906) <= '1';
    layer1_outputs(2907) <= not (a and b);
    layer1_outputs(2908) <= not b;
    layer1_outputs(2909) <= not (a and b);
    layer1_outputs(2910) <= not a or b;
    layer1_outputs(2911) <= b;
    layer1_outputs(2912) <= not b or a;
    layer1_outputs(2913) <= '0';
    layer1_outputs(2914) <= not (a and b);
    layer1_outputs(2915) <= not (a or b);
    layer1_outputs(2916) <= a and b;
    layer1_outputs(2917) <= a or b;
    layer1_outputs(2918) <= not a;
    layer1_outputs(2919) <= a or b;
    layer1_outputs(2920) <= not b or a;
    layer1_outputs(2921) <= a or b;
    layer1_outputs(2922) <= not a;
    layer1_outputs(2923) <= not (a xor b);
    layer1_outputs(2924) <= a;
    layer1_outputs(2925) <= '1';
    layer1_outputs(2926) <= not a or b;
    layer1_outputs(2927) <= b and not a;
    layer1_outputs(2928) <= a;
    layer1_outputs(2929) <= b;
    layer1_outputs(2930) <= not a;
    layer1_outputs(2931) <= not a or b;
    layer1_outputs(2932) <= not a;
    layer1_outputs(2933) <= a;
    layer1_outputs(2934) <= '0';
    layer1_outputs(2935) <= b and not a;
    layer1_outputs(2936) <= not (a or b);
    layer1_outputs(2937) <= not a or b;
    layer1_outputs(2938) <= '1';
    layer1_outputs(2939) <= a and b;
    layer1_outputs(2940) <= a xor b;
    layer1_outputs(2941) <= not a;
    layer1_outputs(2942) <= not a or b;
    layer1_outputs(2943) <= not (a or b);
    layer1_outputs(2944) <= not a;
    layer1_outputs(2945) <= not a;
    layer1_outputs(2946) <= not b or a;
    layer1_outputs(2947) <= '1';
    layer1_outputs(2948) <= a xor b;
    layer1_outputs(2949) <= a xor b;
    layer1_outputs(2950) <= b and not a;
    layer1_outputs(2951) <= '0';
    layer1_outputs(2952) <= b and not a;
    layer1_outputs(2953) <= not (a or b);
    layer1_outputs(2954) <= not a or b;
    layer1_outputs(2955) <= a and not b;
    layer1_outputs(2956) <= not (a and b);
    layer1_outputs(2957) <= '1';
    layer1_outputs(2958) <= not b;
    layer1_outputs(2959) <= not a or b;
    layer1_outputs(2960) <= a;
    layer1_outputs(2961) <= a or b;
    layer1_outputs(2962) <= b and not a;
    layer1_outputs(2963) <= '1';
    layer1_outputs(2964) <= a or b;
    layer1_outputs(2965) <= b and not a;
    layer1_outputs(2966) <= not b or a;
    layer1_outputs(2967) <= not (a xor b);
    layer1_outputs(2968) <= not (a or b);
    layer1_outputs(2969) <= not a or b;
    layer1_outputs(2970) <= not a;
    layer1_outputs(2971) <= a;
    layer1_outputs(2972) <= not (a and b);
    layer1_outputs(2973) <= not a;
    layer1_outputs(2974) <= a;
    layer1_outputs(2975) <= a xor b;
    layer1_outputs(2976) <= '0';
    layer1_outputs(2977) <= not b;
    layer1_outputs(2978) <= not b;
    layer1_outputs(2979) <= not a;
    layer1_outputs(2980) <= not a or b;
    layer1_outputs(2981) <= not b;
    layer1_outputs(2982) <= '0';
    layer1_outputs(2983) <= a and not b;
    layer1_outputs(2984) <= b;
    layer1_outputs(2985) <= b;
    layer1_outputs(2986) <= b and not a;
    layer1_outputs(2987) <= not a or b;
    layer1_outputs(2988) <= '1';
    layer1_outputs(2989) <= not b or a;
    layer1_outputs(2990) <= not a;
    layer1_outputs(2991) <= not a or b;
    layer1_outputs(2992) <= a and not b;
    layer1_outputs(2993) <= not (a or b);
    layer1_outputs(2994) <= a xor b;
    layer1_outputs(2995) <= '1';
    layer1_outputs(2996) <= '0';
    layer1_outputs(2997) <= a and not b;
    layer1_outputs(2998) <= a xor b;
    layer1_outputs(2999) <= not (a or b);
    layer1_outputs(3000) <= not (a xor b);
    layer1_outputs(3001) <= '1';
    layer1_outputs(3002) <= b and not a;
    layer1_outputs(3003) <= not a;
    layer1_outputs(3004) <= b and not a;
    layer1_outputs(3005) <= not b;
    layer1_outputs(3006) <= not a;
    layer1_outputs(3007) <= not b;
    layer1_outputs(3008) <= a and not b;
    layer1_outputs(3009) <= b and not a;
    layer1_outputs(3010) <= '0';
    layer1_outputs(3011) <= a and b;
    layer1_outputs(3012) <= b and not a;
    layer1_outputs(3013) <= a;
    layer1_outputs(3014) <= a;
    layer1_outputs(3015) <= a and b;
    layer1_outputs(3016) <= '1';
    layer1_outputs(3017) <= not a;
    layer1_outputs(3018) <= '1';
    layer1_outputs(3019) <= not (a or b);
    layer1_outputs(3020) <= '1';
    layer1_outputs(3021) <= a and b;
    layer1_outputs(3022) <= not (a and b);
    layer1_outputs(3023) <= a and not b;
    layer1_outputs(3024) <= '0';
    layer1_outputs(3025) <= a or b;
    layer1_outputs(3026) <= a;
    layer1_outputs(3027) <= a and not b;
    layer1_outputs(3028) <= not b;
    layer1_outputs(3029) <= not (a or b);
    layer1_outputs(3030) <= '1';
    layer1_outputs(3031) <= a;
    layer1_outputs(3032) <= a;
    layer1_outputs(3033) <= not (a and b);
    layer1_outputs(3034) <= a and not b;
    layer1_outputs(3035) <= '1';
    layer1_outputs(3036) <= a and not b;
    layer1_outputs(3037) <= not (a or b);
    layer1_outputs(3038) <= not (a and b);
    layer1_outputs(3039) <= a;
    layer1_outputs(3040) <= not a or b;
    layer1_outputs(3041) <= not b or a;
    layer1_outputs(3042) <= a;
    layer1_outputs(3043) <= a or b;
    layer1_outputs(3044) <= a or b;
    layer1_outputs(3045) <= not b;
    layer1_outputs(3046) <= b and not a;
    layer1_outputs(3047) <= b and not a;
    layer1_outputs(3048) <= a and b;
    layer1_outputs(3049) <= a and not b;
    layer1_outputs(3050) <= not b or a;
    layer1_outputs(3051) <= a and b;
    layer1_outputs(3052) <= b;
    layer1_outputs(3053) <= a or b;
    layer1_outputs(3054) <= not (a xor b);
    layer1_outputs(3055) <= '0';
    layer1_outputs(3056) <= a;
    layer1_outputs(3057) <= a and not b;
    layer1_outputs(3058) <= a or b;
    layer1_outputs(3059) <= not a;
    layer1_outputs(3060) <= not b or a;
    layer1_outputs(3061) <= '1';
    layer1_outputs(3062) <= not a or b;
    layer1_outputs(3063) <= not b;
    layer1_outputs(3064) <= '0';
    layer1_outputs(3065) <= not (a or b);
    layer1_outputs(3066) <= not b or a;
    layer1_outputs(3067) <= b;
    layer1_outputs(3068) <= a;
    layer1_outputs(3069) <= not (a xor b);
    layer1_outputs(3070) <= not (a or b);
    layer1_outputs(3071) <= '0';
    layer1_outputs(3072) <= a and not b;
    layer1_outputs(3073) <= not b;
    layer1_outputs(3074) <= a;
    layer1_outputs(3075) <= a;
    layer1_outputs(3076) <= not (a or b);
    layer1_outputs(3077) <= not a;
    layer1_outputs(3078) <= b;
    layer1_outputs(3079) <= not (a xor b);
    layer1_outputs(3080) <= a and b;
    layer1_outputs(3081) <= a or b;
    layer1_outputs(3082) <= not (a and b);
    layer1_outputs(3083) <= a and not b;
    layer1_outputs(3084) <= b;
    layer1_outputs(3085) <= not b;
    layer1_outputs(3086) <= a xor b;
    layer1_outputs(3087) <= '0';
    layer1_outputs(3088) <= not a or b;
    layer1_outputs(3089) <= not a;
    layer1_outputs(3090) <= not a;
    layer1_outputs(3091) <= not b;
    layer1_outputs(3092) <= not a or b;
    layer1_outputs(3093) <= not b or a;
    layer1_outputs(3094) <= not (a and b);
    layer1_outputs(3095) <= not a or b;
    layer1_outputs(3096) <= not b or a;
    layer1_outputs(3097) <= not (a or b);
    layer1_outputs(3098) <= '0';
    layer1_outputs(3099) <= not (a and b);
    layer1_outputs(3100) <= b;
    layer1_outputs(3101) <= not (a or b);
    layer1_outputs(3102) <= b;
    layer1_outputs(3103) <= not a;
    layer1_outputs(3104) <= not b or a;
    layer1_outputs(3105) <= '0';
    layer1_outputs(3106) <= a;
    layer1_outputs(3107) <= not (a and b);
    layer1_outputs(3108) <= not b;
    layer1_outputs(3109) <= not (a and b);
    layer1_outputs(3110) <= not (a and b);
    layer1_outputs(3111) <= not b or a;
    layer1_outputs(3112) <= a;
    layer1_outputs(3113) <= a or b;
    layer1_outputs(3114) <= a or b;
    layer1_outputs(3115) <= b;
    layer1_outputs(3116) <= not (a or b);
    layer1_outputs(3117) <= a;
    layer1_outputs(3118) <= not a or b;
    layer1_outputs(3119) <= not (a and b);
    layer1_outputs(3120) <= not (a and b);
    layer1_outputs(3121) <= b;
    layer1_outputs(3122) <= not a;
    layer1_outputs(3123) <= a or b;
    layer1_outputs(3124) <= not (a or b);
    layer1_outputs(3125) <= a and b;
    layer1_outputs(3126) <= not a or b;
    layer1_outputs(3127) <= not a;
    layer1_outputs(3128) <= '0';
    layer1_outputs(3129) <= a;
    layer1_outputs(3130) <= a or b;
    layer1_outputs(3131) <= not a or b;
    layer1_outputs(3132) <= b and not a;
    layer1_outputs(3133) <= '0';
    layer1_outputs(3134) <= '1';
    layer1_outputs(3135) <= a or b;
    layer1_outputs(3136) <= not (a or b);
    layer1_outputs(3137) <= a;
    layer1_outputs(3138) <= not (a xor b);
    layer1_outputs(3139) <= '0';
    layer1_outputs(3140) <= not a or b;
    layer1_outputs(3141) <= not a;
    layer1_outputs(3142) <= a;
    layer1_outputs(3143) <= a or b;
    layer1_outputs(3144) <= a and b;
    layer1_outputs(3145) <= b and not a;
    layer1_outputs(3146) <= not b;
    layer1_outputs(3147) <= not a or b;
    layer1_outputs(3148) <= '1';
    layer1_outputs(3149) <= not a or b;
    layer1_outputs(3150) <= a and b;
    layer1_outputs(3151) <= '1';
    layer1_outputs(3152) <= a;
    layer1_outputs(3153) <= a and not b;
    layer1_outputs(3154) <= not b;
    layer1_outputs(3155) <= b and not a;
    layer1_outputs(3156) <= not b;
    layer1_outputs(3157) <= not (a or b);
    layer1_outputs(3158) <= b and not a;
    layer1_outputs(3159) <= not a or b;
    layer1_outputs(3160) <= a xor b;
    layer1_outputs(3161) <= '1';
    layer1_outputs(3162) <= '1';
    layer1_outputs(3163) <= not a;
    layer1_outputs(3164) <= a;
    layer1_outputs(3165) <= '0';
    layer1_outputs(3166) <= not b;
    layer1_outputs(3167) <= '1';
    layer1_outputs(3168) <= '0';
    layer1_outputs(3169) <= a xor b;
    layer1_outputs(3170) <= not b or a;
    layer1_outputs(3171) <= a or b;
    layer1_outputs(3172) <= not a;
    layer1_outputs(3173) <= not b;
    layer1_outputs(3174) <= not b or a;
    layer1_outputs(3175) <= not (a and b);
    layer1_outputs(3176) <= '1';
    layer1_outputs(3177) <= a;
    layer1_outputs(3178) <= not (a or b);
    layer1_outputs(3179) <= '0';
    layer1_outputs(3180) <= not (a or b);
    layer1_outputs(3181) <= a and b;
    layer1_outputs(3182) <= not a;
    layer1_outputs(3183) <= a or b;
    layer1_outputs(3184) <= not (a and b);
    layer1_outputs(3185) <= b and not a;
    layer1_outputs(3186) <= not (a and b);
    layer1_outputs(3187) <= b and not a;
    layer1_outputs(3188) <= not (a and b);
    layer1_outputs(3189) <= not (a or b);
    layer1_outputs(3190) <= a;
    layer1_outputs(3191) <= a or b;
    layer1_outputs(3192) <= a and b;
    layer1_outputs(3193) <= not b or a;
    layer1_outputs(3194) <= b;
    layer1_outputs(3195) <= '1';
    layer1_outputs(3196) <= a or b;
    layer1_outputs(3197) <= not (a xor b);
    layer1_outputs(3198) <= b and not a;
    layer1_outputs(3199) <= '1';
    layer1_outputs(3200) <= a or b;
    layer1_outputs(3201) <= a;
    layer1_outputs(3202) <= a;
    layer1_outputs(3203) <= a and b;
    layer1_outputs(3204) <= b and not a;
    layer1_outputs(3205) <= a and b;
    layer1_outputs(3206) <= not b or a;
    layer1_outputs(3207) <= not (a and b);
    layer1_outputs(3208) <= '1';
    layer1_outputs(3209) <= not (a and b);
    layer1_outputs(3210) <= b;
    layer1_outputs(3211) <= b and not a;
    layer1_outputs(3212) <= '0';
    layer1_outputs(3213) <= not b or a;
    layer1_outputs(3214) <= not a;
    layer1_outputs(3215) <= '1';
    layer1_outputs(3216) <= b;
    layer1_outputs(3217) <= not b;
    layer1_outputs(3218) <= not (a and b);
    layer1_outputs(3219) <= not b;
    layer1_outputs(3220) <= not b;
    layer1_outputs(3221) <= not (a or b);
    layer1_outputs(3222) <= not (a xor b);
    layer1_outputs(3223) <= '0';
    layer1_outputs(3224) <= a;
    layer1_outputs(3225) <= a and not b;
    layer1_outputs(3226) <= not b or a;
    layer1_outputs(3227) <= not (a or b);
    layer1_outputs(3228) <= '0';
    layer1_outputs(3229) <= a;
    layer1_outputs(3230) <= '0';
    layer1_outputs(3231) <= '0';
    layer1_outputs(3232) <= a or b;
    layer1_outputs(3233) <= not a or b;
    layer1_outputs(3234) <= a xor b;
    layer1_outputs(3235) <= not a or b;
    layer1_outputs(3236) <= not (a or b);
    layer1_outputs(3237) <= not a or b;
    layer1_outputs(3238) <= not a;
    layer1_outputs(3239) <= '0';
    layer1_outputs(3240) <= not (a and b);
    layer1_outputs(3241) <= b and not a;
    layer1_outputs(3242) <= not (a and b);
    layer1_outputs(3243) <= not b;
    layer1_outputs(3244) <= not (a and b);
    layer1_outputs(3245) <= not (a or b);
    layer1_outputs(3246) <= not (a and b);
    layer1_outputs(3247) <= not b or a;
    layer1_outputs(3248) <= not b or a;
    layer1_outputs(3249) <= a;
    layer1_outputs(3250) <= not b or a;
    layer1_outputs(3251) <= not a;
    layer1_outputs(3252) <= a;
    layer1_outputs(3253) <= not a;
    layer1_outputs(3254) <= a;
    layer1_outputs(3255) <= '1';
    layer1_outputs(3256) <= a;
    layer1_outputs(3257) <= b;
    layer1_outputs(3258) <= b and not a;
    layer1_outputs(3259) <= a and not b;
    layer1_outputs(3260) <= a or b;
    layer1_outputs(3261) <= a and b;
    layer1_outputs(3262) <= not (a xor b);
    layer1_outputs(3263) <= not b;
    layer1_outputs(3264) <= not (a or b);
    layer1_outputs(3265) <= not a;
    layer1_outputs(3266) <= b;
    layer1_outputs(3267) <= b;
    layer1_outputs(3268) <= b and not a;
    layer1_outputs(3269) <= '0';
    layer1_outputs(3270) <= not b;
    layer1_outputs(3271) <= '1';
    layer1_outputs(3272) <= not b;
    layer1_outputs(3273) <= b;
    layer1_outputs(3274) <= '1';
    layer1_outputs(3275) <= not (a or b);
    layer1_outputs(3276) <= not a;
    layer1_outputs(3277) <= not (a and b);
    layer1_outputs(3278) <= b and not a;
    layer1_outputs(3279) <= a;
    layer1_outputs(3280) <= a and not b;
    layer1_outputs(3281) <= not (a or b);
    layer1_outputs(3282) <= not b or a;
    layer1_outputs(3283) <= '1';
    layer1_outputs(3284) <= not b;
    layer1_outputs(3285) <= not b;
    layer1_outputs(3286) <= not (a or b);
    layer1_outputs(3287) <= a and not b;
    layer1_outputs(3288) <= a;
    layer1_outputs(3289) <= '0';
    layer1_outputs(3290) <= a xor b;
    layer1_outputs(3291) <= a and b;
    layer1_outputs(3292) <= '0';
    layer1_outputs(3293) <= b and not a;
    layer1_outputs(3294) <= not a or b;
    layer1_outputs(3295) <= not (a or b);
    layer1_outputs(3296) <= not b or a;
    layer1_outputs(3297) <= b;
    layer1_outputs(3298) <= b and not a;
    layer1_outputs(3299) <= not (a and b);
    layer1_outputs(3300) <= not (a or b);
    layer1_outputs(3301) <= not (a xor b);
    layer1_outputs(3302) <= a or b;
    layer1_outputs(3303) <= not a or b;
    layer1_outputs(3304) <= '1';
    layer1_outputs(3305) <= a xor b;
    layer1_outputs(3306) <= a or b;
    layer1_outputs(3307) <= a xor b;
    layer1_outputs(3308) <= a and b;
    layer1_outputs(3309) <= not a or b;
    layer1_outputs(3310) <= not (a and b);
    layer1_outputs(3311) <= a and not b;
    layer1_outputs(3312) <= a or b;
    layer1_outputs(3313) <= not b or a;
    layer1_outputs(3314) <= b;
    layer1_outputs(3315) <= b and not a;
    layer1_outputs(3316) <= not b or a;
    layer1_outputs(3317) <= a or b;
    layer1_outputs(3318) <= not a;
    layer1_outputs(3319) <= not a or b;
    layer1_outputs(3320) <= not (a and b);
    layer1_outputs(3321) <= a and not b;
    layer1_outputs(3322) <= not (a and b);
    layer1_outputs(3323) <= not b or a;
    layer1_outputs(3324) <= not a or b;
    layer1_outputs(3325) <= b;
    layer1_outputs(3326) <= a and b;
    layer1_outputs(3327) <= not b or a;
    layer1_outputs(3328) <= not b or a;
    layer1_outputs(3329) <= b;
    layer1_outputs(3330) <= not a or b;
    layer1_outputs(3331) <= a;
    layer1_outputs(3332) <= not a or b;
    layer1_outputs(3333) <= not (a or b);
    layer1_outputs(3334) <= a or b;
    layer1_outputs(3335) <= a and not b;
    layer1_outputs(3336) <= b;
    layer1_outputs(3337) <= not b or a;
    layer1_outputs(3338) <= not b;
    layer1_outputs(3339) <= b and not a;
    layer1_outputs(3340) <= '0';
    layer1_outputs(3341) <= a and b;
    layer1_outputs(3342) <= a xor b;
    layer1_outputs(3343) <= a;
    layer1_outputs(3344) <= not a or b;
    layer1_outputs(3345) <= '0';
    layer1_outputs(3346) <= not a or b;
    layer1_outputs(3347) <= not (a and b);
    layer1_outputs(3348) <= b and not a;
    layer1_outputs(3349) <= not b or a;
    layer1_outputs(3350) <= not (a and b);
    layer1_outputs(3351) <= b;
    layer1_outputs(3352) <= '1';
    layer1_outputs(3353) <= '0';
    layer1_outputs(3354) <= not (a and b);
    layer1_outputs(3355) <= a or b;
    layer1_outputs(3356) <= not (a or b);
    layer1_outputs(3357) <= not a;
    layer1_outputs(3358) <= '1';
    layer1_outputs(3359) <= not b or a;
    layer1_outputs(3360) <= a xor b;
    layer1_outputs(3361) <= a xor b;
    layer1_outputs(3362) <= b and not a;
    layer1_outputs(3363) <= '0';
    layer1_outputs(3364) <= not a or b;
    layer1_outputs(3365) <= not (a or b);
    layer1_outputs(3366) <= a or b;
    layer1_outputs(3367) <= a and b;
    layer1_outputs(3368) <= a or b;
    layer1_outputs(3369) <= not a or b;
    layer1_outputs(3370) <= not b or a;
    layer1_outputs(3371) <= not (a and b);
    layer1_outputs(3372) <= a;
    layer1_outputs(3373) <= a;
    layer1_outputs(3374) <= not a;
    layer1_outputs(3375) <= b;
    layer1_outputs(3376) <= not a;
    layer1_outputs(3377) <= not a;
    layer1_outputs(3378) <= not b or a;
    layer1_outputs(3379) <= a or b;
    layer1_outputs(3380) <= not a or b;
    layer1_outputs(3381) <= b;
    layer1_outputs(3382) <= not (a or b);
    layer1_outputs(3383) <= not a or b;
    layer1_outputs(3384) <= b;
    layer1_outputs(3385) <= '0';
    layer1_outputs(3386) <= b and not a;
    layer1_outputs(3387) <= not b;
    layer1_outputs(3388) <= not (a xor b);
    layer1_outputs(3389) <= not (a or b);
    layer1_outputs(3390) <= '0';
    layer1_outputs(3391) <= not b;
    layer1_outputs(3392) <= '1';
    layer1_outputs(3393) <= a or b;
    layer1_outputs(3394) <= a and not b;
    layer1_outputs(3395) <= not (a or b);
    layer1_outputs(3396) <= not (a or b);
    layer1_outputs(3397) <= a xor b;
    layer1_outputs(3398) <= '1';
    layer1_outputs(3399) <= a;
    layer1_outputs(3400) <= a or b;
    layer1_outputs(3401) <= a and b;
    layer1_outputs(3402) <= a and b;
    layer1_outputs(3403) <= '1';
    layer1_outputs(3404) <= '0';
    layer1_outputs(3405) <= a and b;
    layer1_outputs(3406) <= not a;
    layer1_outputs(3407) <= not a or b;
    layer1_outputs(3408) <= not b or a;
    layer1_outputs(3409) <= a and b;
    layer1_outputs(3410) <= not (a or b);
    layer1_outputs(3411) <= a;
    layer1_outputs(3412) <= b;
    layer1_outputs(3413) <= not a or b;
    layer1_outputs(3414) <= not (a or b);
    layer1_outputs(3415) <= a;
    layer1_outputs(3416) <= not a;
    layer1_outputs(3417) <= b;
    layer1_outputs(3418) <= not a or b;
    layer1_outputs(3419) <= a;
    layer1_outputs(3420) <= b and not a;
    layer1_outputs(3421) <= not b;
    layer1_outputs(3422) <= not (a xor b);
    layer1_outputs(3423) <= not b;
    layer1_outputs(3424) <= not b;
    layer1_outputs(3425) <= not b or a;
    layer1_outputs(3426) <= not a or b;
    layer1_outputs(3427) <= not a or b;
    layer1_outputs(3428) <= not b or a;
    layer1_outputs(3429) <= a and not b;
    layer1_outputs(3430) <= a or b;
    layer1_outputs(3431) <= not (a or b);
    layer1_outputs(3432) <= not (a or b);
    layer1_outputs(3433) <= b;
    layer1_outputs(3434) <= a;
    layer1_outputs(3435) <= a;
    layer1_outputs(3436) <= a;
    layer1_outputs(3437) <= '0';
    layer1_outputs(3438) <= '1';
    layer1_outputs(3439) <= b and not a;
    layer1_outputs(3440) <= a and not b;
    layer1_outputs(3441) <= '1';
    layer1_outputs(3442) <= b;
    layer1_outputs(3443) <= a;
    layer1_outputs(3444) <= '1';
    layer1_outputs(3445) <= b and not a;
    layer1_outputs(3446) <= not b or a;
    layer1_outputs(3447) <= not (a xor b);
    layer1_outputs(3448) <= a or b;
    layer1_outputs(3449) <= not b;
    layer1_outputs(3450) <= not b;
    layer1_outputs(3451) <= not (a or b);
    layer1_outputs(3452) <= b;
    layer1_outputs(3453) <= not b;
    layer1_outputs(3454) <= not b or a;
    layer1_outputs(3455) <= b and not a;
    layer1_outputs(3456) <= not (a or b);
    layer1_outputs(3457) <= not b;
    layer1_outputs(3458) <= b and not a;
    layer1_outputs(3459) <= b;
    layer1_outputs(3460) <= a or b;
    layer1_outputs(3461) <= a;
    layer1_outputs(3462) <= a and not b;
    layer1_outputs(3463) <= b and not a;
    layer1_outputs(3464) <= '1';
    layer1_outputs(3465) <= a and b;
    layer1_outputs(3466) <= not (a xor b);
    layer1_outputs(3467) <= b;
    layer1_outputs(3468) <= '1';
    layer1_outputs(3469) <= b;
    layer1_outputs(3470) <= not a;
    layer1_outputs(3471) <= b and not a;
    layer1_outputs(3472) <= not b;
    layer1_outputs(3473) <= a or b;
    layer1_outputs(3474) <= b;
    layer1_outputs(3475) <= a and not b;
    layer1_outputs(3476) <= not a or b;
    layer1_outputs(3477) <= not b;
    layer1_outputs(3478) <= not (a or b);
    layer1_outputs(3479) <= not (a or b);
    layer1_outputs(3480) <= not (a and b);
    layer1_outputs(3481) <= b and not a;
    layer1_outputs(3482) <= b and not a;
    layer1_outputs(3483) <= a;
    layer1_outputs(3484) <= b;
    layer1_outputs(3485) <= not b;
    layer1_outputs(3486) <= not (a or b);
    layer1_outputs(3487) <= a xor b;
    layer1_outputs(3488) <= not (a or b);
    layer1_outputs(3489) <= a;
    layer1_outputs(3490) <= a and not b;
    layer1_outputs(3491) <= not (a xor b);
    layer1_outputs(3492) <= not a;
    layer1_outputs(3493) <= a or b;
    layer1_outputs(3494) <= a and not b;
    layer1_outputs(3495) <= a xor b;
    layer1_outputs(3496) <= '0';
    layer1_outputs(3497) <= a;
    layer1_outputs(3498) <= a and not b;
    layer1_outputs(3499) <= not (a xor b);
    layer1_outputs(3500) <= not b;
    layer1_outputs(3501) <= a;
    layer1_outputs(3502) <= not b or a;
    layer1_outputs(3503) <= not b or a;
    layer1_outputs(3504) <= a and not b;
    layer1_outputs(3505) <= not (a xor b);
    layer1_outputs(3506) <= not b or a;
    layer1_outputs(3507) <= not (a or b);
    layer1_outputs(3508) <= a and not b;
    layer1_outputs(3509) <= a;
    layer1_outputs(3510) <= '0';
    layer1_outputs(3511) <= a and not b;
    layer1_outputs(3512) <= b and not a;
    layer1_outputs(3513) <= '1';
    layer1_outputs(3514) <= not b or a;
    layer1_outputs(3515) <= a;
    layer1_outputs(3516) <= a or b;
    layer1_outputs(3517) <= a xor b;
    layer1_outputs(3518) <= not b;
    layer1_outputs(3519) <= '0';
    layer1_outputs(3520) <= b;
    layer1_outputs(3521) <= not a;
    layer1_outputs(3522) <= a or b;
    layer1_outputs(3523) <= b;
    layer1_outputs(3524) <= not b;
    layer1_outputs(3525) <= not (a or b);
    layer1_outputs(3526) <= a xor b;
    layer1_outputs(3527) <= a and b;
    layer1_outputs(3528) <= not a or b;
    layer1_outputs(3529) <= not a or b;
    layer1_outputs(3530) <= '0';
    layer1_outputs(3531) <= a xor b;
    layer1_outputs(3532) <= b;
    layer1_outputs(3533) <= b;
    layer1_outputs(3534) <= a xor b;
    layer1_outputs(3535) <= not (a and b);
    layer1_outputs(3536) <= not (a or b);
    layer1_outputs(3537) <= not b;
    layer1_outputs(3538) <= not b or a;
    layer1_outputs(3539) <= a and not b;
    layer1_outputs(3540) <= not (a or b);
    layer1_outputs(3541) <= a and b;
    layer1_outputs(3542) <= a;
    layer1_outputs(3543) <= '0';
    layer1_outputs(3544) <= a;
    layer1_outputs(3545) <= not b or a;
    layer1_outputs(3546) <= a;
    layer1_outputs(3547) <= a;
    layer1_outputs(3548) <= not (a or b);
    layer1_outputs(3549) <= not a;
    layer1_outputs(3550) <= not b;
    layer1_outputs(3551) <= a or b;
    layer1_outputs(3552) <= a xor b;
    layer1_outputs(3553) <= b;
    layer1_outputs(3554) <= b and not a;
    layer1_outputs(3555) <= a and b;
    layer1_outputs(3556) <= not (a and b);
    layer1_outputs(3557) <= a and b;
    layer1_outputs(3558) <= b;
    layer1_outputs(3559) <= a and b;
    layer1_outputs(3560) <= a;
    layer1_outputs(3561) <= not a or b;
    layer1_outputs(3562) <= a and b;
    layer1_outputs(3563) <= not (a xor b);
    layer1_outputs(3564) <= not (a and b);
    layer1_outputs(3565) <= b and not a;
    layer1_outputs(3566) <= '1';
    layer1_outputs(3567) <= a;
    layer1_outputs(3568) <= a or b;
    layer1_outputs(3569) <= not (a and b);
    layer1_outputs(3570) <= a or b;
    layer1_outputs(3571) <= '1';
    layer1_outputs(3572) <= a xor b;
    layer1_outputs(3573) <= not a or b;
    layer1_outputs(3574) <= a or b;
    layer1_outputs(3575) <= b;
    layer1_outputs(3576) <= not a;
    layer1_outputs(3577) <= a and not b;
    layer1_outputs(3578) <= '0';
    layer1_outputs(3579) <= not a;
    layer1_outputs(3580) <= not (a xor b);
    layer1_outputs(3581) <= b;
    layer1_outputs(3582) <= not b or a;
    layer1_outputs(3583) <= not a;
    layer1_outputs(3584) <= not (a or b);
    layer1_outputs(3585) <= a or b;
    layer1_outputs(3586) <= a or b;
    layer1_outputs(3587) <= not a or b;
    layer1_outputs(3588) <= a and not b;
    layer1_outputs(3589) <= not (a xor b);
    layer1_outputs(3590) <= not a;
    layer1_outputs(3591) <= a and b;
    layer1_outputs(3592) <= not (a or b);
    layer1_outputs(3593) <= not b;
    layer1_outputs(3594) <= not b;
    layer1_outputs(3595) <= b and not a;
    layer1_outputs(3596) <= a;
    layer1_outputs(3597) <= a and b;
    layer1_outputs(3598) <= not (a xor b);
    layer1_outputs(3599) <= not a;
    layer1_outputs(3600) <= not (a and b);
    layer1_outputs(3601) <= not b;
    layer1_outputs(3602) <= not (a xor b);
    layer1_outputs(3603) <= a or b;
    layer1_outputs(3604) <= b;
    layer1_outputs(3605) <= b and not a;
    layer1_outputs(3606) <= a;
    layer1_outputs(3607) <= not (a and b);
    layer1_outputs(3608) <= not a;
    layer1_outputs(3609) <= not b or a;
    layer1_outputs(3610) <= a and b;
    layer1_outputs(3611) <= a or b;
    layer1_outputs(3612) <= not b;
    layer1_outputs(3613) <= not a or b;
    layer1_outputs(3614) <= b and not a;
    layer1_outputs(3615) <= a and not b;
    layer1_outputs(3616) <= not a;
    layer1_outputs(3617) <= a or b;
    layer1_outputs(3618) <= a xor b;
    layer1_outputs(3619) <= a and not b;
    layer1_outputs(3620) <= not b or a;
    layer1_outputs(3621) <= '0';
    layer1_outputs(3622) <= b and not a;
    layer1_outputs(3623) <= b;
    layer1_outputs(3624) <= a or b;
    layer1_outputs(3625) <= not (a or b);
    layer1_outputs(3626) <= a xor b;
    layer1_outputs(3627) <= b;
    layer1_outputs(3628) <= b;
    layer1_outputs(3629) <= not (a and b);
    layer1_outputs(3630) <= a and not b;
    layer1_outputs(3631) <= '0';
    layer1_outputs(3632) <= not b or a;
    layer1_outputs(3633) <= not (a xor b);
    layer1_outputs(3634) <= a or b;
    layer1_outputs(3635) <= a xor b;
    layer1_outputs(3636) <= a or b;
    layer1_outputs(3637) <= not a;
    layer1_outputs(3638) <= not b;
    layer1_outputs(3639) <= not b or a;
    layer1_outputs(3640) <= not b or a;
    layer1_outputs(3641) <= not (a xor b);
    layer1_outputs(3642) <= '0';
    layer1_outputs(3643) <= a xor b;
    layer1_outputs(3644) <= not a or b;
    layer1_outputs(3645) <= not b or a;
    layer1_outputs(3646) <= b and not a;
    layer1_outputs(3647) <= '0';
    layer1_outputs(3648) <= a;
    layer1_outputs(3649) <= not (a xor b);
    layer1_outputs(3650) <= a;
    layer1_outputs(3651) <= a and not b;
    layer1_outputs(3652) <= b and not a;
    layer1_outputs(3653) <= not (a and b);
    layer1_outputs(3654) <= not a or b;
    layer1_outputs(3655) <= a and not b;
    layer1_outputs(3656) <= not (a and b);
    layer1_outputs(3657) <= not (a and b);
    layer1_outputs(3658) <= not b or a;
    layer1_outputs(3659) <= a;
    layer1_outputs(3660) <= a;
    layer1_outputs(3661) <= a;
    layer1_outputs(3662) <= b and not a;
    layer1_outputs(3663) <= '0';
    layer1_outputs(3664) <= not a;
    layer1_outputs(3665) <= not a;
    layer1_outputs(3666) <= '0';
    layer1_outputs(3667) <= b;
    layer1_outputs(3668) <= not (a or b);
    layer1_outputs(3669) <= b;
    layer1_outputs(3670) <= not b;
    layer1_outputs(3671) <= a and not b;
    layer1_outputs(3672) <= not a;
    layer1_outputs(3673) <= a;
    layer1_outputs(3674) <= a;
    layer1_outputs(3675) <= a;
    layer1_outputs(3676) <= a and not b;
    layer1_outputs(3677) <= '0';
    layer1_outputs(3678) <= a or b;
    layer1_outputs(3679) <= a;
    layer1_outputs(3680) <= b and not a;
    layer1_outputs(3681) <= not a or b;
    layer1_outputs(3682) <= not b or a;
    layer1_outputs(3683) <= not a;
    layer1_outputs(3684) <= '1';
    layer1_outputs(3685) <= not (a or b);
    layer1_outputs(3686) <= a xor b;
    layer1_outputs(3687) <= a or b;
    layer1_outputs(3688) <= a and not b;
    layer1_outputs(3689) <= not a;
    layer1_outputs(3690) <= a xor b;
    layer1_outputs(3691) <= '0';
    layer1_outputs(3692) <= not a;
    layer1_outputs(3693) <= b;
    layer1_outputs(3694) <= not a;
    layer1_outputs(3695) <= '1';
    layer1_outputs(3696) <= b and not a;
    layer1_outputs(3697) <= not (a and b);
    layer1_outputs(3698) <= not a;
    layer1_outputs(3699) <= a and not b;
    layer1_outputs(3700) <= a;
    layer1_outputs(3701) <= '1';
    layer1_outputs(3702) <= a and b;
    layer1_outputs(3703) <= not a;
    layer1_outputs(3704) <= '1';
    layer1_outputs(3705) <= b and not a;
    layer1_outputs(3706) <= not b or a;
    layer1_outputs(3707) <= a;
    layer1_outputs(3708) <= not (a xor b);
    layer1_outputs(3709) <= not a or b;
    layer1_outputs(3710) <= not b or a;
    layer1_outputs(3711) <= not a or b;
    layer1_outputs(3712) <= not b;
    layer1_outputs(3713) <= b;
    layer1_outputs(3714) <= not (a or b);
    layer1_outputs(3715) <= a and b;
    layer1_outputs(3716) <= b and not a;
    layer1_outputs(3717) <= not b or a;
    layer1_outputs(3718) <= a;
    layer1_outputs(3719) <= a or b;
    layer1_outputs(3720) <= '0';
    layer1_outputs(3721) <= not (a or b);
    layer1_outputs(3722) <= not a or b;
    layer1_outputs(3723) <= not (a and b);
    layer1_outputs(3724) <= b and not a;
    layer1_outputs(3725) <= '0';
    layer1_outputs(3726) <= a;
    layer1_outputs(3727) <= '1';
    layer1_outputs(3728) <= b;
    layer1_outputs(3729) <= '1';
    layer1_outputs(3730) <= not (a and b);
    layer1_outputs(3731) <= not (a and b);
    layer1_outputs(3732) <= b and not a;
    layer1_outputs(3733) <= a and not b;
    layer1_outputs(3734) <= a;
    layer1_outputs(3735) <= a or b;
    layer1_outputs(3736) <= a or b;
    layer1_outputs(3737) <= a and not b;
    layer1_outputs(3738) <= b;
    layer1_outputs(3739) <= a and not b;
    layer1_outputs(3740) <= a and not b;
    layer1_outputs(3741) <= '1';
    layer1_outputs(3742) <= b;
    layer1_outputs(3743) <= not a or b;
    layer1_outputs(3744) <= a or b;
    layer1_outputs(3745) <= b and not a;
    layer1_outputs(3746) <= a or b;
    layer1_outputs(3747) <= not a;
    layer1_outputs(3748) <= b and not a;
    layer1_outputs(3749) <= b;
    layer1_outputs(3750) <= b;
    layer1_outputs(3751) <= not (a xor b);
    layer1_outputs(3752) <= a or b;
    layer1_outputs(3753) <= a xor b;
    layer1_outputs(3754) <= not b;
    layer1_outputs(3755) <= a and b;
    layer1_outputs(3756) <= a and b;
    layer1_outputs(3757) <= not a or b;
    layer1_outputs(3758) <= not b;
    layer1_outputs(3759) <= b;
    layer1_outputs(3760) <= '0';
    layer1_outputs(3761) <= not (a xor b);
    layer1_outputs(3762) <= a xor b;
    layer1_outputs(3763) <= not (a and b);
    layer1_outputs(3764) <= b;
    layer1_outputs(3765) <= not (a and b);
    layer1_outputs(3766) <= a;
    layer1_outputs(3767) <= b;
    layer1_outputs(3768) <= a and b;
    layer1_outputs(3769) <= a and b;
    layer1_outputs(3770) <= a or b;
    layer1_outputs(3771) <= b;
    layer1_outputs(3772) <= a and b;
    layer1_outputs(3773) <= b;
    layer1_outputs(3774) <= not b or a;
    layer1_outputs(3775) <= '1';
    layer1_outputs(3776) <= a;
    layer1_outputs(3777) <= '0';
    layer1_outputs(3778) <= a and b;
    layer1_outputs(3779) <= not b or a;
    layer1_outputs(3780) <= a or b;
    layer1_outputs(3781) <= a or b;
    layer1_outputs(3782) <= not b;
    layer1_outputs(3783) <= not (a or b);
    layer1_outputs(3784) <= a or b;
    layer1_outputs(3785) <= not a;
    layer1_outputs(3786) <= b;
    layer1_outputs(3787) <= not a or b;
    layer1_outputs(3788) <= a and not b;
    layer1_outputs(3789) <= a xor b;
    layer1_outputs(3790) <= a xor b;
    layer1_outputs(3791) <= a or b;
    layer1_outputs(3792) <= not b;
    layer1_outputs(3793) <= not (a xor b);
    layer1_outputs(3794) <= a and not b;
    layer1_outputs(3795) <= '0';
    layer1_outputs(3796) <= b;
    layer1_outputs(3797) <= b and not a;
    layer1_outputs(3798) <= '0';
    layer1_outputs(3799) <= '0';
    layer1_outputs(3800) <= not a;
    layer1_outputs(3801) <= a;
    layer1_outputs(3802) <= not b or a;
    layer1_outputs(3803) <= '0';
    layer1_outputs(3804) <= b;
    layer1_outputs(3805) <= a or b;
    layer1_outputs(3806) <= a xor b;
    layer1_outputs(3807) <= a or b;
    layer1_outputs(3808) <= a or b;
    layer1_outputs(3809) <= not a;
    layer1_outputs(3810) <= not b or a;
    layer1_outputs(3811) <= not (a xor b);
    layer1_outputs(3812) <= a;
    layer1_outputs(3813) <= b and not a;
    layer1_outputs(3814) <= a or b;
    layer1_outputs(3815) <= a or b;
    layer1_outputs(3816) <= b and not a;
    layer1_outputs(3817) <= b;
    layer1_outputs(3818) <= '0';
    layer1_outputs(3819) <= '1';
    layer1_outputs(3820) <= a and not b;
    layer1_outputs(3821) <= b;
    layer1_outputs(3822) <= not (a or b);
    layer1_outputs(3823) <= a and not b;
    layer1_outputs(3824) <= not b;
    layer1_outputs(3825) <= a or b;
    layer1_outputs(3826) <= '0';
    layer1_outputs(3827) <= not (a and b);
    layer1_outputs(3828) <= not (a and b);
    layer1_outputs(3829) <= not (a or b);
    layer1_outputs(3830) <= a or b;
    layer1_outputs(3831) <= not (a xor b);
    layer1_outputs(3832) <= not b;
    layer1_outputs(3833) <= b;
    layer1_outputs(3834) <= a or b;
    layer1_outputs(3835) <= not b or a;
    layer1_outputs(3836) <= b and not a;
    layer1_outputs(3837) <= a xor b;
    layer1_outputs(3838) <= not (a and b);
    layer1_outputs(3839) <= a;
    layer1_outputs(3840) <= '1';
    layer1_outputs(3841) <= a and b;
    layer1_outputs(3842) <= not b or a;
    layer1_outputs(3843) <= '0';
    layer1_outputs(3844) <= a;
    layer1_outputs(3845) <= a;
    layer1_outputs(3846) <= not (a xor b);
    layer1_outputs(3847) <= a;
    layer1_outputs(3848) <= '0';
    layer1_outputs(3849) <= not (a and b);
    layer1_outputs(3850) <= not b or a;
    layer1_outputs(3851) <= a xor b;
    layer1_outputs(3852) <= '0';
    layer1_outputs(3853) <= not b;
    layer1_outputs(3854) <= not a;
    layer1_outputs(3855) <= '0';
    layer1_outputs(3856) <= a and b;
    layer1_outputs(3857) <= not (a and b);
    layer1_outputs(3858) <= not a;
    layer1_outputs(3859) <= b;
    layer1_outputs(3860) <= not a or b;
    layer1_outputs(3861) <= a and not b;
    layer1_outputs(3862) <= '1';
    layer1_outputs(3863) <= '1';
    layer1_outputs(3864) <= b;
    layer1_outputs(3865) <= a and not b;
    layer1_outputs(3866) <= not a;
    layer1_outputs(3867) <= a;
    layer1_outputs(3868) <= a or b;
    layer1_outputs(3869) <= not b;
    layer1_outputs(3870) <= a and b;
    layer1_outputs(3871) <= not b;
    layer1_outputs(3872) <= not (a or b);
    layer1_outputs(3873) <= a;
    layer1_outputs(3874) <= not a or b;
    layer1_outputs(3875) <= '0';
    layer1_outputs(3876) <= not a or b;
    layer1_outputs(3877) <= a;
    layer1_outputs(3878) <= not (a and b);
    layer1_outputs(3879) <= b;
    layer1_outputs(3880) <= not b or a;
    layer1_outputs(3881) <= b;
    layer1_outputs(3882) <= '1';
    layer1_outputs(3883) <= not (a or b);
    layer1_outputs(3884) <= not a or b;
    layer1_outputs(3885) <= a or b;
    layer1_outputs(3886) <= not (a or b);
    layer1_outputs(3887) <= not b or a;
    layer1_outputs(3888) <= not a;
    layer1_outputs(3889) <= not b or a;
    layer1_outputs(3890) <= b;
    layer1_outputs(3891) <= a;
    layer1_outputs(3892) <= a or b;
    layer1_outputs(3893) <= not a;
    layer1_outputs(3894) <= a and not b;
    layer1_outputs(3895) <= not (a or b);
    layer1_outputs(3896) <= a and b;
    layer1_outputs(3897) <= not (a or b);
    layer1_outputs(3898) <= '0';
    layer1_outputs(3899) <= '0';
    layer1_outputs(3900) <= b;
    layer1_outputs(3901) <= a and b;
    layer1_outputs(3902) <= not a;
    layer1_outputs(3903) <= a or b;
    layer1_outputs(3904) <= a;
    layer1_outputs(3905) <= not (a or b);
    layer1_outputs(3906) <= not b or a;
    layer1_outputs(3907) <= not a or b;
    layer1_outputs(3908) <= not (a xor b);
    layer1_outputs(3909) <= a or b;
    layer1_outputs(3910) <= a and not b;
    layer1_outputs(3911) <= not a;
    layer1_outputs(3912) <= not (a or b);
    layer1_outputs(3913) <= not b;
    layer1_outputs(3914) <= a and not b;
    layer1_outputs(3915) <= not (a or b);
    layer1_outputs(3916) <= '0';
    layer1_outputs(3917) <= not (a and b);
    layer1_outputs(3918) <= '0';
    layer1_outputs(3919) <= a and not b;
    layer1_outputs(3920) <= not a or b;
    layer1_outputs(3921) <= not a;
    layer1_outputs(3922) <= not a or b;
    layer1_outputs(3923) <= a or b;
    layer1_outputs(3924) <= a and b;
    layer1_outputs(3925) <= not b;
    layer1_outputs(3926) <= not b or a;
    layer1_outputs(3927) <= b and not a;
    layer1_outputs(3928) <= not b;
    layer1_outputs(3929) <= b;
    layer1_outputs(3930) <= '1';
    layer1_outputs(3931) <= b and not a;
    layer1_outputs(3932) <= a or b;
    layer1_outputs(3933) <= not a;
    layer1_outputs(3934) <= a;
    layer1_outputs(3935) <= a or b;
    layer1_outputs(3936) <= '0';
    layer1_outputs(3937) <= not (a xor b);
    layer1_outputs(3938) <= not (a and b);
    layer1_outputs(3939) <= b and not a;
    layer1_outputs(3940) <= not a;
    layer1_outputs(3941) <= not (a or b);
    layer1_outputs(3942) <= not b or a;
    layer1_outputs(3943) <= not b or a;
    layer1_outputs(3944) <= '0';
    layer1_outputs(3945) <= not a;
    layer1_outputs(3946) <= not b;
    layer1_outputs(3947) <= not b;
    layer1_outputs(3948) <= '0';
    layer1_outputs(3949) <= b;
    layer1_outputs(3950) <= not (a or b);
    layer1_outputs(3951) <= b;
    layer1_outputs(3952) <= not b;
    layer1_outputs(3953) <= not a;
    layer1_outputs(3954) <= '1';
    layer1_outputs(3955) <= b;
    layer1_outputs(3956) <= not (a or b);
    layer1_outputs(3957) <= b and not a;
    layer1_outputs(3958) <= '1';
    layer1_outputs(3959) <= a or b;
    layer1_outputs(3960) <= not b or a;
    layer1_outputs(3961) <= b and not a;
    layer1_outputs(3962) <= a and not b;
    layer1_outputs(3963) <= a;
    layer1_outputs(3964) <= not a or b;
    layer1_outputs(3965) <= a and b;
    layer1_outputs(3966) <= '0';
    layer1_outputs(3967) <= a and not b;
    layer1_outputs(3968) <= not (a or b);
    layer1_outputs(3969) <= a and not b;
    layer1_outputs(3970) <= a and b;
    layer1_outputs(3971) <= '1';
    layer1_outputs(3972) <= a and not b;
    layer1_outputs(3973) <= not b;
    layer1_outputs(3974) <= not (a or b);
    layer1_outputs(3975) <= b and not a;
    layer1_outputs(3976) <= not (a or b);
    layer1_outputs(3977) <= not b or a;
    layer1_outputs(3978) <= not (a or b);
    layer1_outputs(3979) <= a xor b;
    layer1_outputs(3980) <= '0';
    layer1_outputs(3981) <= a;
    layer1_outputs(3982) <= b;
    layer1_outputs(3983) <= a;
    layer1_outputs(3984) <= not b;
    layer1_outputs(3985) <= not b;
    layer1_outputs(3986) <= a;
    layer1_outputs(3987) <= a xor b;
    layer1_outputs(3988) <= not (a and b);
    layer1_outputs(3989) <= a and not b;
    layer1_outputs(3990) <= a or b;
    layer1_outputs(3991) <= a xor b;
    layer1_outputs(3992) <= not b;
    layer1_outputs(3993) <= not a;
    layer1_outputs(3994) <= a and not b;
    layer1_outputs(3995) <= a and b;
    layer1_outputs(3996) <= not a;
    layer1_outputs(3997) <= not b;
    layer1_outputs(3998) <= a;
    layer1_outputs(3999) <= a and not b;
    layer1_outputs(4000) <= not (a and b);
    layer1_outputs(4001) <= not (a xor b);
    layer1_outputs(4002) <= b and not a;
    layer1_outputs(4003) <= b;
    layer1_outputs(4004) <= a;
    layer1_outputs(4005) <= a or b;
    layer1_outputs(4006) <= '1';
    layer1_outputs(4007) <= not (a xor b);
    layer1_outputs(4008) <= not a;
    layer1_outputs(4009) <= not (a or b);
    layer1_outputs(4010) <= not b or a;
    layer1_outputs(4011) <= a and not b;
    layer1_outputs(4012) <= a;
    layer1_outputs(4013) <= a and not b;
    layer1_outputs(4014) <= b;
    layer1_outputs(4015) <= a and not b;
    layer1_outputs(4016) <= a;
    layer1_outputs(4017) <= a;
    layer1_outputs(4018) <= not b;
    layer1_outputs(4019) <= not b or a;
    layer1_outputs(4020) <= not (a and b);
    layer1_outputs(4021) <= not a;
    layer1_outputs(4022) <= not (a and b);
    layer1_outputs(4023) <= '0';
    layer1_outputs(4024) <= not a;
    layer1_outputs(4025) <= not (a and b);
    layer1_outputs(4026) <= a and not b;
    layer1_outputs(4027) <= a and not b;
    layer1_outputs(4028) <= a and not b;
    layer1_outputs(4029) <= not b;
    layer1_outputs(4030) <= a and not b;
    layer1_outputs(4031) <= not a;
    layer1_outputs(4032) <= a and b;
    layer1_outputs(4033) <= not a;
    layer1_outputs(4034) <= b;
    layer1_outputs(4035) <= b;
    layer1_outputs(4036) <= not b or a;
    layer1_outputs(4037) <= a or b;
    layer1_outputs(4038) <= b and not a;
    layer1_outputs(4039) <= not b or a;
    layer1_outputs(4040) <= a or b;
    layer1_outputs(4041) <= not b or a;
    layer1_outputs(4042) <= b;
    layer1_outputs(4043) <= a;
    layer1_outputs(4044) <= not b or a;
    layer1_outputs(4045) <= not (a and b);
    layer1_outputs(4046) <= not (a or b);
    layer1_outputs(4047) <= not a or b;
    layer1_outputs(4048) <= a or b;
    layer1_outputs(4049) <= not (a or b);
    layer1_outputs(4050) <= not (a and b);
    layer1_outputs(4051) <= not (a and b);
    layer1_outputs(4052) <= not b;
    layer1_outputs(4053) <= b and not a;
    layer1_outputs(4054) <= a and b;
    layer1_outputs(4055) <= a and b;
    layer1_outputs(4056) <= not (a or b);
    layer1_outputs(4057) <= a;
    layer1_outputs(4058) <= a;
    layer1_outputs(4059) <= not b or a;
    layer1_outputs(4060) <= not a;
    layer1_outputs(4061) <= a xor b;
    layer1_outputs(4062) <= not a or b;
    layer1_outputs(4063) <= b and not a;
    layer1_outputs(4064) <= not b;
    layer1_outputs(4065) <= not a or b;
    layer1_outputs(4066) <= not b or a;
    layer1_outputs(4067) <= a or b;
    layer1_outputs(4068) <= a and not b;
    layer1_outputs(4069) <= not b or a;
    layer1_outputs(4070) <= not a;
    layer1_outputs(4071) <= not (a or b);
    layer1_outputs(4072) <= not b or a;
    layer1_outputs(4073) <= not (a and b);
    layer1_outputs(4074) <= not (a and b);
    layer1_outputs(4075) <= '0';
    layer1_outputs(4076) <= a;
    layer1_outputs(4077) <= not (a or b);
    layer1_outputs(4078) <= '1';
    layer1_outputs(4079) <= a or b;
    layer1_outputs(4080) <= b;
    layer1_outputs(4081) <= a or b;
    layer1_outputs(4082) <= not b;
    layer1_outputs(4083) <= a xor b;
    layer1_outputs(4084) <= not (a or b);
    layer1_outputs(4085) <= a or b;
    layer1_outputs(4086) <= not (a or b);
    layer1_outputs(4087) <= '0';
    layer1_outputs(4088) <= not a;
    layer1_outputs(4089) <= b and not a;
    layer1_outputs(4090) <= not b;
    layer1_outputs(4091) <= '0';
    layer1_outputs(4092) <= not b or a;
    layer1_outputs(4093) <= not b;
    layer1_outputs(4094) <= '1';
    layer1_outputs(4095) <= b;
    layer1_outputs(4096) <= a;
    layer1_outputs(4097) <= a and not b;
    layer1_outputs(4098) <= not a;
    layer1_outputs(4099) <= not b;
    layer1_outputs(4100) <= a and not b;
    layer1_outputs(4101) <= '0';
    layer1_outputs(4102) <= a;
    layer1_outputs(4103) <= b;
    layer1_outputs(4104) <= a;
    layer1_outputs(4105) <= a and not b;
    layer1_outputs(4106) <= a and not b;
    layer1_outputs(4107) <= a and b;
    layer1_outputs(4108) <= not a;
    layer1_outputs(4109) <= b;
    layer1_outputs(4110) <= a and b;
    layer1_outputs(4111) <= not b;
    layer1_outputs(4112) <= a or b;
    layer1_outputs(4113) <= not a;
    layer1_outputs(4114) <= not (a and b);
    layer1_outputs(4115) <= a and b;
    layer1_outputs(4116) <= not a;
    layer1_outputs(4117) <= b and not a;
    layer1_outputs(4118) <= b;
    layer1_outputs(4119) <= b and not a;
    layer1_outputs(4120) <= '0';
    layer1_outputs(4121) <= a and b;
    layer1_outputs(4122) <= not b or a;
    layer1_outputs(4123) <= a and not b;
    layer1_outputs(4124) <= not a;
    layer1_outputs(4125) <= a;
    layer1_outputs(4126) <= not a;
    layer1_outputs(4127) <= a and not b;
    layer1_outputs(4128) <= b and not a;
    layer1_outputs(4129) <= not a;
    layer1_outputs(4130) <= '1';
    layer1_outputs(4131) <= b and not a;
    layer1_outputs(4132) <= a and not b;
    layer1_outputs(4133) <= not b;
    layer1_outputs(4134) <= not b or a;
    layer1_outputs(4135) <= b;
    layer1_outputs(4136) <= a xor b;
    layer1_outputs(4137) <= b and not a;
    layer1_outputs(4138) <= b and not a;
    layer1_outputs(4139) <= a;
    layer1_outputs(4140) <= '1';
    layer1_outputs(4141) <= a and not b;
    layer1_outputs(4142) <= not (a and b);
    layer1_outputs(4143) <= not (a xor b);
    layer1_outputs(4144) <= '1';
    layer1_outputs(4145) <= a and b;
    layer1_outputs(4146) <= not b;
    layer1_outputs(4147) <= '0';
    layer1_outputs(4148) <= not b or a;
    layer1_outputs(4149) <= '0';
    layer1_outputs(4150) <= a and not b;
    layer1_outputs(4151) <= a xor b;
    layer1_outputs(4152) <= not a or b;
    layer1_outputs(4153) <= b;
    layer1_outputs(4154) <= not b or a;
    layer1_outputs(4155) <= not a;
    layer1_outputs(4156) <= b and not a;
    layer1_outputs(4157) <= '1';
    layer1_outputs(4158) <= a;
    layer1_outputs(4159) <= not a or b;
    layer1_outputs(4160) <= '0';
    layer1_outputs(4161) <= not b;
    layer1_outputs(4162) <= a and not b;
    layer1_outputs(4163) <= not (a and b);
    layer1_outputs(4164) <= not b;
    layer1_outputs(4165) <= a and b;
    layer1_outputs(4166) <= not a or b;
    layer1_outputs(4167) <= a and b;
    layer1_outputs(4168) <= not b or a;
    layer1_outputs(4169) <= not a;
    layer1_outputs(4170) <= '1';
    layer1_outputs(4171) <= '1';
    layer1_outputs(4172) <= a or b;
    layer1_outputs(4173) <= '1';
    layer1_outputs(4174) <= a or b;
    layer1_outputs(4175) <= b;
    layer1_outputs(4176) <= not a;
    layer1_outputs(4177) <= not b;
    layer1_outputs(4178) <= b;
    layer1_outputs(4179) <= not a or b;
    layer1_outputs(4180) <= b;
    layer1_outputs(4181) <= not a;
    layer1_outputs(4182) <= a or b;
    layer1_outputs(4183) <= not (a xor b);
    layer1_outputs(4184) <= not a;
    layer1_outputs(4185) <= b;
    layer1_outputs(4186) <= not b or a;
    layer1_outputs(4187) <= not (a or b);
    layer1_outputs(4188) <= not b;
    layer1_outputs(4189) <= b;
    layer1_outputs(4190) <= b;
    layer1_outputs(4191) <= not (a and b);
    layer1_outputs(4192) <= not b;
    layer1_outputs(4193) <= b;
    layer1_outputs(4194) <= b;
    layer1_outputs(4195) <= a;
    layer1_outputs(4196) <= b;
    layer1_outputs(4197) <= not a;
    layer1_outputs(4198) <= not a;
    layer1_outputs(4199) <= not b or a;
    layer1_outputs(4200) <= not a;
    layer1_outputs(4201) <= a or b;
    layer1_outputs(4202) <= not b or a;
    layer1_outputs(4203) <= not a or b;
    layer1_outputs(4204) <= not b or a;
    layer1_outputs(4205) <= not a or b;
    layer1_outputs(4206) <= b and not a;
    layer1_outputs(4207) <= not b;
    layer1_outputs(4208) <= a and b;
    layer1_outputs(4209) <= a and b;
    layer1_outputs(4210) <= a and b;
    layer1_outputs(4211) <= b;
    layer1_outputs(4212) <= a;
    layer1_outputs(4213) <= not b;
    layer1_outputs(4214) <= a;
    layer1_outputs(4215) <= b;
    layer1_outputs(4216) <= '1';
    layer1_outputs(4217) <= a or b;
    layer1_outputs(4218) <= a;
    layer1_outputs(4219) <= a or b;
    layer1_outputs(4220) <= a and not b;
    layer1_outputs(4221) <= b;
    layer1_outputs(4222) <= a and not b;
    layer1_outputs(4223) <= a;
    layer1_outputs(4224) <= not (a and b);
    layer1_outputs(4225) <= '1';
    layer1_outputs(4226) <= not a;
    layer1_outputs(4227) <= a and b;
    layer1_outputs(4228) <= not b;
    layer1_outputs(4229) <= a and b;
    layer1_outputs(4230) <= a and b;
    layer1_outputs(4231) <= a;
    layer1_outputs(4232) <= a or b;
    layer1_outputs(4233) <= b;
    layer1_outputs(4234) <= not a;
    layer1_outputs(4235) <= a and not b;
    layer1_outputs(4236) <= '1';
    layer1_outputs(4237) <= not (a and b);
    layer1_outputs(4238) <= '0';
    layer1_outputs(4239) <= not a;
    layer1_outputs(4240) <= not b;
    layer1_outputs(4241) <= a and b;
    layer1_outputs(4242) <= b and not a;
    layer1_outputs(4243) <= not (a or b);
    layer1_outputs(4244) <= b;
    layer1_outputs(4245) <= a xor b;
    layer1_outputs(4246) <= not b;
    layer1_outputs(4247) <= not (a xor b);
    layer1_outputs(4248) <= a and not b;
    layer1_outputs(4249) <= not b or a;
    layer1_outputs(4250) <= not b;
    layer1_outputs(4251) <= not b;
    layer1_outputs(4252) <= b and not a;
    layer1_outputs(4253) <= a or b;
    layer1_outputs(4254) <= a;
    layer1_outputs(4255) <= not b;
    layer1_outputs(4256) <= a;
    layer1_outputs(4257) <= not b or a;
    layer1_outputs(4258) <= not (a and b);
    layer1_outputs(4259) <= a or b;
    layer1_outputs(4260) <= not (a or b);
    layer1_outputs(4261) <= '0';
    layer1_outputs(4262) <= a xor b;
    layer1_outputs(4263) <= b;
    layer1_outputs(4264) <= a;
    layer1_outputs(4265) <= '1';
    layer1_outputs(4266) <= '0';
    layer1_outputs(4267) <= not (a and b);
    layer1_outputs(4268) <= not a;
    layer1_outputs(4269) <= not b or a;
    layer1_outputs(4270) <= not (a and b);
    layer1_outputs(4271) <= '0';
    layer1_outputs(4272) <= b;
    layer1_outputs(4273) <= a or b;
    layer1_outputs(4274) <= not b;
    layer1_outputs(4275) <= a and b;
    layer1_outputs(4276) <= not b;
    layer1_outputs(4277) <= not (a and b);
    layer1_outputs(4278) <= a and b;
    layer1_outputs(4279) <= '1';
    layer1_outputs(4280) <= a;
    layer1_outputs(4281) <= not b;
    layer1_outputs(4282) <= not (a and b);
    layer1_outputs(4283) <= not a;
    layer1_outputs(4284) <= b;
    layer1_outputs(4285) <= '1';
    layer1_outputs(4286) <= not (a or b);
    layer1_outputs(4287) <= b and not a;
    layer1_outputs(4288) <= a and b;
    layer1_outputs(4289) <= a and b;
    layer1_outputs(4290) <= not (a or b);
    layer1_outputs(4291) <= a and not b;
    layer1_outputs(4292) <= not (a or b);
    layer1_outputs(4293) <= not a or b;
    layer1_outputs(4294) <= a and not b;
    layer1_outputs(4295) <= not b;
    layer1_outputs(4296) <= b and not a;
    layer1_outputs(4297) <= a or b;
    layer1_outputs(4298) <= not a;
    layer1_outputs(4299) <= not a or b;
    layer1_outputs(4300) <= b and not a;
    layer1_outputs(4301) <= '0';
    layer1_outputs(4302) <= not b or a;
    layer1_outputs(4303) <= not b;
    layer1_outputs(4304) <= b and not a;
    layer1_outputs(4305) <= b and not a;
    layer1_outputs(4306) <= a and b;
    layer1_outputs(4307) <= a or b;
    layer1_outputs(4308) <= a and b;
    layer1_outputs(4309) <= not b;
    layer1_outputs(4310) <= not (a and b);
    layer1_outputs(4311) <= not b or a;
    layer1_outputs(4312) <= a and b;
    layer1_outputs(4313) <= '1';
    layer1_outputs(4314) <= a or b;
    layer1_outputs(4315) <= not a;
    layer1_outputs(4316) <= b;
    layer1_outputs(4317) <= not b or a;
    layer1_outputs(4318) <= a or b;
    layer1_outputs(4319) <= a and b;
    layer1_outputs(4320) <= a;
    layer1_outputs(4321) <= not b or a;
    layer1_outputs(4322) <= '1';
    layer1_outputs(4323) <= b and not a;
    layer1_outputs(4324) <= not a or b;
    layer1_outputs(4325) <= not b or a;
    layer1_outputs(4326) <= a;
    layer1_outputs(4327) <= not (a and b);
    layer1_outputs(4328) <= not (a xor b);
    layer1_outputs(4329) <= not a or b;
    layer1_outputs(4330) <= a xor b;
    layer1_outputs(4331) <= a;
    layer1_outputs(4332) <= '1';
    layer1_outputs(4333) <= not b;
    layer1_outputs(4334) <= a and b;
    layer1_outputs(4335) <= b;
    layer1_outputs(4336) <= b;
    layer1_outputs(4337) <= not b;
    layer1_outputs(4338) <= a and not b;
    layer1_outputs(4339) <= not b or a;
    layer1_outputs(4340) <= b and not a;
    layer1_outputs(4341) <= not a or b;
    layer1_outputs(4342) <= not b;
    layer1_outputs(4343) <= a and not b;
    layer1_outputs(4344) <= a or b;
    layer1_outputs(4345) <= not a or b;
    layer1_outputs(4346) <= not a;
    layer1_outputs(4347) <= a or b;
    layer1_outputs(4348) <= '1';
    layer1_outputs(4349) <= not (a or b);
    layer1_outputs(4350) <= b and not a;
    layer1_outputs(4351) <= not a;
    layer1_outputs(4352) <= b;
    layer1_outputs(4353) <= b and not a;
    layer1_outputs(4354) <= not a;
    layer1_outputs(4355) <= not (a and b);
    layer1_outputs(4356) <= not a;
    layer1_outputs(4357) <= '1';
    layer1_outputs(4358) <= a and b;
    layer1_outputs(4359) <= a;
    layer1_outputs(4360) <= a;
    layer1_outputs(4361) <= '1';
    layer1_outputs(4362) <= not (a and b);
    layer1_outputs(4363) <= not a or b;
    layer1_outputs(4364) <= not a;
    layer1_outputs(4365) <= b;
    layer1_outputs(4366) <= not (a xor b);
    layer1_outputs(4367) <= not b;
    layer1_outputs(4368) <= b;
    layer1_outputs(4369) <= not b;
    layer1_outputs(4370) <= a;
    layer1_outputs(4371) <= a and not b;
    layer1_outputs(4372) <= a;
    layer1_outputs(4373) <= '1';
    layer1_outputs(4374) <= '1';
    layer1_outputs(4375) <= not b;
    layer1_outputs(4376) <= b and not a;
    layer1_outputs(4377) <= a;
    layer1_outputs(4378) <= a;
    layer1_outputs(4379) <= not b;
    layer1_outputs(4380) <= not (a and b);
    layer1_outputs(4381) <= not a or b;
    layer1_outputs(4382) <= not (a and b);
    layer1_outputs(4383) <= a or b;
    layer1_outputs(4384) <= not (a and b);
    layer1_outputs(4385) <= '1';
    layer1_outputs(4386) <= a and b;
    layer1_outputs(4387) <= a or b;
    layer1_outputs(4388) <= a xor b;
    layer1_outputs(4389) <= b and not a;
    layer1_outputs(4390) <= not (a and b);
    layer1_outputs(4391) <= not a;
    layer1_outputs(4392) <= a and not b;
    layer1_outputs(4393) <= a and b;
    layer1_outputs(4394) <= a and b;
    layer1_outputs(4395) <= not (a xor b);
    layer1_outputs(4396) <= not b or a;
    layer1_outputs(4397) <= not b or a;
    layer1_outputs(4398) <= '0';
    layer1_outputs(4399) <= a and b;
    layer1_outputs(4400) <= '1';
    layer1_outputs(4401) <= not (a or b);
    layer1_outputs(4402) <= a and not b;
    layer1_outputs(4403) <= not (a and b);
    layer1_outputs(4404) <= not (a or b);
    layer1_outputs(4405) <= not (a xor b);
    layer1_outputs(4406) <= not (a and b);
    layer1_outputs(4407) <= not a;
    layer1_outputs(4408) <= not (a or b);
    layer1_outputs(4409) <= not a;
    layer1_outputs(4410) <= not a;
    layer1_outputs(4411) <= a and not b;
    layer1_outputs(4412) <= not a;
    layer1_outputs(4413) <= a or b;
    layer1_outputs(4414) <= a xor b;
    layer1_outputs(4415) <= not (a or b);
    layer1_outputs(4416) <= a or b;
    layer1_outputs(4417) <= a;
    layer1_outputs(4418) <= not a or b;
    layer1_outputs(4419) <= not a;
    layer1_outputs(4420) <= b and not a;
    layer1_outputs(4421) <= not a or b;
    layer1_outputs(4422) <= not b;
    layer1_outputs(4423) <= not b or a;
    layer1_outputs(4424) <= a xor b;
    layer1_outputs(4425) <= not b or a;
    layer1_outputs(4426) <= not b;
    layer1_outputs(4427) <= a and b;
    layer1_outputs(4428) <= not a;
    layer1_outputs(4429) <= not (a and b);
    layer1_outputs(4430) <= not (a or b);
    layer1_outputs(4431) <= not b;
    layer1_outputs(4432) <= '1';
    layer1_outputs(4433) <= a;
    layer1_outputs(4434) <= a and not b;
    layer1_outputs(4435) <= a and not b;
    layer1_outputs(4436) <= not (a and b);
    layer1_outputs(4437) <= a;
    layer1_outputs(4438) <= '1';
    layer1_outputs(4439) <= b and not a;
    layer1_outputs(4440) <= '0';
    layer1_outputs(4441) <= '1';
    layer1_outputs(4442) <= '0';
    layer1_outputs(4443) <= not (a or b);
    layer1_outputs(4444) <= a and b;
    layer1_outputs(4445) <= a and not b;
    layer1_outputs(4446) <= '0';
    layer1_outputs(4447) <= a or b;
    layer1_outputs(4448) <= not (a and b);
    layer1_outputs(4449) <= not b;
    layer1_outputs(4450) <= a and not b;
    layer1_outputs(4451) <= b and not a;
    layer1_outputs(4452) <= not b or a;
    layer1_outputs(4453) <= not a or b;
    layer1_outputs(4454) <= a and b;
    layer1_outputs(4455) <= '0';
    layer1_outputs(4456) <= a and not b;
    layer1_outputs(4457) <= a and not b;
    layer1_outputs(4458) <= not a;
    layer1_outputs(4459) <= not a or b;
    layer1_outputs(4460) <= a;
    layer1_outputs(4461) <= a and not b;
    layer1_outputs(4462) <= a and not b;
    layer1_outputs(4463) <= '0';
    layer1_outputs(4464) <= b and not a;
    layer1_outputs(4465) <= not (a xor b);
    layer1_outputs(4466) <= a;
    layer1_outputs(4467) <= not b or a;
    layer1_outputs(4468) <= not a;
    layer1_outputs(4469) <= not a;
    layer1_outputs(4470) <= not (a and b);
    layer1_outputs(4471) <= a;
    layer1_outputs(4472) <= b and not a;
    layer1_outputs(4473) <= not a or b;
    layer1_outputs(4474) <= '1';
    layer1_outputs(4475) <= b and not a;
    layer1_outputs(4476) <= a or b;
    layer1_outputs(4477) <= a;
    layer1_outputs(4478) <= b and not a;
    layer1_outputs(4479) <= '1';
    layer1_outputs(4480) <= a;
    layer1_outputs(4481) <= not a;
    layer1_outputs(4482) <= not a or b;
    layer1_outputs(4483) <= not b;
    layer1_outputs(4484) <= not (a and b);
    layer1_outputs(4485) <= not (a or b);
    layer1_outputs(4486) <= not b or a;
    layer1_outputs(4487) <= not b or a;
    layer1_outputs(4488) <= a;
    layer1_outputs(4489) <= not a or b;
    layer1_outputs(4490) <= not a;
    layer1_outputs(4491) <= a;
    layer1_outputs(4492) <= a or b;
    layer1_outputs(4493) <= '1';
    layer1_outputs(4494) <= not a;
    layer1_outputs(4495) <= a;
    layer1_outputs(4496) <= b;
    layer1_outputs(4497) <= '0';
    layer1_outputs(4498) <= b and not a;
    layer1_outputs(4499) <= not (a or b);
    layer1_outputs(4500) <= not a;
    layer1_outputs(4501) <= a and b;
    layer1_outputs(4502) <= a and b;
    layer1_outputs(4503) <= '0';
    layer1_outputs(4504) <= a;
    layer1_outputs(4505) <= '0';
    layer1_outputs(4506) <= not (a and b);
    layer1_outputs(4507) <= not a or b;
    layer1_outputs(4508) <= b and not a;
    layer1_outputs(4509) <= '0';
    layer1_outputs(4510) <= not (a xor b);
    layer1_outputs(4511) <= not a or b;
    layer1_outputs(4512) <= not (a xor b);
    layer1_outputs(4513) <= a;
    layer1_outputs(4514) <= a or b;
    layer1_outputs(4515) <= not b;
    layer1_outputs(4516) <= not a;
    layer1_outputs(4517) <= a and not b;
    layer1_outputs(4518) <= '1';
    layer1_outputs(4519) <= a or b;
    layer1_outputs(4520) <= b;
    layer1_outputs(4521) <= a;
    layer1_outputs(4522) <= not a or b;
    layer1_outputs(4523) <= not b or a;
    layer1_outputs(4524) <= not a;
    layer1_outputs(4525) <= a or b;
    layer1_outputs(4526) <= '0';
    layer1_outputs(4527) <= not a or b;
    layer1_outputs(4528) <= a and b;
    layer1_outputs(4529) <= b;
    layer1_outputs(4530) <= not b;
    layer1_outputs(4531) <= not b or a;
    layer1_outputs(4532) <= not b;
    layer1_outputs(4533) <= b;
    layer1_outputs(4534) <= not a;
    layer1_outputs(4535) <= a and not b;
    layer1_outputs(4536) <= not a or b;
    layer1_outputs(4537) <= '0';
    layer1_outputs(4538) <= b;
    layer1_outputs(4539) <= a and b;
    layer1_outputs(4540) <= '0';
    layer1_outputs(4541) <= not a or b;
    layer1_outputs(4542) <= a and not b;
    layer1_outputs(4543) <= b;
    layer1_outputs(4544) <= not a;
    layer1_outputs(4545) <= a xor b;
    layer1_outputs(4546) <= not b or a;
    layer1_outputs(4547) <= not (a or b);
    layer1_outputs(4548) <= not a;
    layer1_outputs(4549) <= a and not b;
    layer1_outputs(4550) <= not a or b;
    layer1_outputs(4551) <= not b or a;
    layer1_outputs(4552) <= not a;
    layer1_outputs(4553) <= not a;
    layer1_outputs(4554) <= not b or a;
    layer1_outputs(4555) <= '1';
    layer1_outputs(4556) <= not b or a;
    layer1_outputs(4557) <= not (a and b);
    layer1_outputs(4558) <= a and not b;
    layer1_outputs(4559) <= '1';
    layer1_outputs(4560) <= not (a or b);
    layer1_outputs(4561) <= not a or b;
    layer1_outputs(4562) <= not a;
    layer1_outputs(4563) <= not b or a;
    layer1_outputs(4564) <= a and not b;
    layer1_outputs(4565) <= not (a or b);
    layer1_outputs(4566) <= a or b;
    layer1_outputs(4567) <= not a;
    layer1_outputs(4568) <= b;
    layer1_outputs(4569) <= a xor b;
    layer1_outputs(4570) <= b and not a;
    layer1_outputs(4571) <= not (a and b);
    layer1_outputs(4572) <= b and not a;
    layer1_outputs(4573) <= b;
    layer1_outputs(4574) <= not b or a;
    layer1_outputs(4575) <= not a;
    layer1_outputs(4576) <= not b;
    layer1_outputs(4577) <= a or b;
    layer1_outputs(4578) <= not b;
    layer1_outputs(4579) <= not b;
    layer1_outputs(4580) <= b;
    layer1_outputs(4581) <= not b;
    layer1_outputs(4582) <= not b;
    layer1_outputs(4583) <= not b;
    layer1_outputs(4584) <= b and not a;
    layer1_outputs(4585) <= not b;
    layer1_outputs(4586) <= a or b;
    layer1_outputs(4587) <= not (a xor b);
    layer1_outputs(4588) <= not b or a;
    layer1_outputs(4589) <= a and not b;
    layer1_outputs(4590) <= not (a xor b);
    layer1_outputs(4591) <= '1';
    layer1_outputs(4592) <= a;
    layer1_outputs(4593) <= b and not a;
    layer1_outputs(4594) <= a;
    layer1_outputs(4595) <= b;
    layer1_outputs(4596) <= '1';
    layer1_outputs(4597) <= a and not b;
    layer1_outputs(4598) <= not (a xor b);
    layer1_outputs(4599) <= a;
    layer1_outputs(4600) <= b and not a;
    layer1_outputs(4601) <= not a;
    layer1_outputs(4602) <= '0';
    layer1_outputs(4603) <= a or b;
    layer1_outputs(4604) <= not b or a;
    layer1_outputs(4605) <= '0';
    layer1_outputs(4606) <= not a;
    layer1_outputs(4607) <= not (a and b);
    layer1_outputs(4608) <= a;
    layer1_outputs(4609) <= not b;
    layer1_outputs(4610) <= not (a or b);
    layer1_outputs(4611) <= not b or a;
    layer1_outputs(4612) <= b;
    layer1_outputs(4613) <= '1';
    layer1_outputs(4614) <= b;
    layer1_outputs(4615) <= '1';
    layer1_outputs(4616) <= not (a or b);
    layer1_outputs(4617) <= not a;
    layer1_outputs(4618) <= not (a and b);
    layer1_outputs(4619) <= '1';
    layer1_outputs(4620) <= '0';
    layer1_outputs(4621) <= a or b;
    layer1_outputs(4622) <= a;
    layer1_outputs(4623) <= a or b;
    layer1_outputs(4624) <= not a or b;
    layer1_outputs(4625) <= a;
    layer1_outputs(4626) <= not (a and b);
    layer1_outputs(4627) <= b;
    layer1_outputs(4628) <= a;
    layer1_outputs(4629) <= not a or b;
    layer1_outputs(4630) <= '0';
    layer1_outputs(4631) <= not b or a;
    layer1_outputs(4632) <= a and b;
    layer1_outputs(4633) <= '1';
    layer1_outputs(4634) <= not b or a;
    layer1_outputs(4635) <= '0';
    layer1_outputs(4636) <= not (a or b);
    layer1_outputs(4637) <= '0';
    layer1_outputs(4638) <= '1';
    layer1_outputs(4639) <= b and not a;
    layer1_outputs(4640) <= b and not a;
    layer1_outputs(4641) <= a;
    layer1_outputs(4642) <= a or b;
    layer1_outputs(4643) <= not (a or b);
    layer1_outputs(4644) <= b and not a;
    layer1_outputs(4645) <= not (a xor b);
    layer1_outputs(4646) <= not (a xor b);
    layer1_outputs(4647) <= not (a and b);
    layer1_outputs(4648) <= not b or a;
    layer1_outputs(4649) <= a and not b;
    layer1_outputs(4650) <= '0';
    layer1_outputs(4651) <= b;
    layer1_outputs(4652) <= '1';
    layer1_outputs(4653) <= not b;
    layer1_outputs(4654) <= a and b;
    layer1_outputs(4655) <= not a;
    layer1_outputs(4656) <= not a;
    layer1_outputs(4657) <= a and not b;
    layer1_outputs(4658) <= a and not b;
    layer1_outputs(4659) <= not b or a;
    layer1_outputs(4660) <= not (a or b);
    layer1_outputs(4661) <= '0';
    layer1_outputs(4662) <= not b;
    layer1_outputs(4663) <= not (a or b);
    layer1_outputs(4664) <= not a;
    layer1_outputs(4665) <= not (a and b);
    layer1_outputs(4666) <= a and not b;
    layer1_outputs(4667) <= a xor b;
    layer1_outputs(4668) <= not a;
    layer1_outputs(4669) <= not (a or b);
    layer1_outputs(4670) <= '1';
    layer1_outputs(4671) <= not a or b;
    layer1_outputs(4672) <= not (a or b);
    layer1_outputs(4673) <= b;
    layer1_outputs(4674) <= a xor b;
    layer1_outputs(4675) <= a and b;
    layer1_outputs(4676) <= a and not b;
    layer1_outputs(4677) <= a or b;
    layer1_outputs(4678) <= '1';
    layer1_outputs(4679) <= not a;
    layer1_outputs(4680) <= not (a and b);
    layer1_outputs(4681) <= not (a and b);
    layer1_outputs(4682) <= not b or a;
    layer1_outputs(4683) <= '1';
    layer1_outputs(4684) <= not a or b;
    layer1_outputs(4685) <= a or b;
    layer1_outputs(4686) <= not a or b;
    layer1_outputs(4687) <= '0';
    layer1_outputs(4688) <= a and b;
    layer1_outputs(4689) <= a and b;
    layer1_outputs(4690) <= not a;
    layer1_outputs(4691) <= a or b;
    layer1_outputs(4692) <= b and not a;
    layer1_outputs(4693) <= not a or b;
    layer1_outputs(4694) <= a and b;
    layer1_outputs(4695) <= a;
    layer1_outputs(4696) <= not b or a;
    layer1_outputs(4697) <= a and b;
    layer1_outputs(4698) <= not (a and b);
    layer1_outputs(4699) <= '1';
    layer1_outputs(4700) <= b;
    layer1_outputs(4701) <= a or b;
    layer1_outputs(4702) <= '0';
    layer1_outputs(4703) <= a;
    layer1_outputs(4704) <= a and b;
    layer1_outputs(4705) <= a and b;
    layer1_outputs(4706) <= not a;
    layer1_outputs(4707) <= not b or a;
    layer1_outputs(4708) <= a and not b;
    layer1_outputs(4709) <= a and not b;
    layer1_outputs(4710) <= a and b;
    layer1_outputs(4711) <= not b or a;
    layer1_outputs(4712) <= not a;
    layer1_outputs(4713) <= not a;
    layer1_outputs(4714) <= not a;
    layer1_outputs(4715) <= a xor b;
    layer1_outputs(4716) <= not b;
    layer1_outputs(4717) <= b;
    layer1_outputs(4718) <= not (a xor b);
    layer1_outputs(4719) <= not (a xor b);
    layer1_outputs(4720) <= not a;
    layer1_outputs(4721) <= a or b;
    layer1_outputs(4722) <= not a;
    layer1_outputs(4723) <= '1';
    layer1_outputs(4724) <= a xor b;
    layer1_outputs(4725) <= '0';
    layer1_outputs(4726) <= b and not a;
    layer1_outputs(4727) <= not (a and b);
    layer1_outputs(4728) <= '1';
    layer1_outputs(4729) <= b and not a;
    layer1_outputs(4730) <= a or b;
    layer1_outputs(4731) <= a xor b;
    layer1_outputs(4732) <= not b or a;
    layer1_outputs(4733) <= b and not a;
    layer1_outputs(4734) <= a;
    layer1_outputs(4735) <= a and not b;
    layer1_outputs(4736) <= '0';
    layer1_outputs(4737) <= not a or b;
    layer1_outputs(4738) <= not (a and b);
    layer1_outputs(4739) <= not b or a;
    layer1_outputs(4740) <= not b or a;
    layer1_outputs(4741) <= not a;
    layer1_outputs(4742) <= a or b;
    layer1_outputs(4743) <= not b;
    layer1_outputs(4744) <= not (a and b);
    layer1_outputs(4745) <= a and not b;
    layer1_outputs(4746) <= b and not a;
    layer1_outputs(4747) <= b and not a;
    layer1_outputs(4748) <= not (a or b);
    layer1_outputs(4749) <= not (a and b);
    layer1_outputs(4750) <= b and not a;
    layer1_outputs(4751) <= not (a xor b);
    layer1_outputs(4752) <= a;
    layer1_outputs(4753) <= b;
    layer1_outputs(4754) <= a or b;
    layer1_outputs(4755) <= not (a or b);
    layer1_outputs(4756) <= a and b;
    layer1_outputs(4757) <= a and b;
    layer1_outputs(4758) <= a;
    layer1_outputs(4759) <= not (a or b);
    layer1_outputs(4760) <= a and not b;
    layer1_outputs(4761) <= '1';
    layer1_outputs(4762) <= not (a xor b);
    layer1_outputs(4763) <= not b;
    layer1_outputs(4764) <= '1';
    layer1_outputs(4765) <= a or b;
    layer1_outputs(4766) <= a;
    layer1_outputs(4767) <= a and b;
    layer1_outputs(4768) <= not (a and b);
    layer1_outputs(4769) <= a and b;
    layer1_outputs(4770) <= '0';
    layer1_outputs(4771) <= not b;
    layer1_outputs(4772) <= a;
    layer1_outputs(4773) <= not b;
    layer1_outputs(4774) <= a and b;
    layer1_outputs(4775) <= a xor b;
    layer1_outputs(4776) <= '0';
    layer1_outputs(4777) <= a;
    layer1_outputs(4778) <= a and b;
    layer1_outputs(4779) <= not (a or b);
    layer1_outputs(4780) <= not b or a;
    layer1_outputs(4781) <= a or b;
    layer1_outputs(4782) <= not a;
    layer1_outputs(4783) <= a xor b;
    layer1_outputs(4784) <= a;
    layer1_outputs(4785) <= not b;
    layer1_outputs(4786) <= a and not b;
    layer1_outputs(4787) <= a and not b;
    layer1_outputs(4788) <= a and not b;
    layer1_outputs(4789) <= not b;
    layer1_outputs(4790) <= not b or a;
    layer1_outputs(4791) <= not b;
    layer1_outputs(4792) <= b;
    layer1_outputs(4793) <= not b or a;
    layer1_outputs(4794) <= not (a and b);
    layer1_outputs(4795) <= '1';
    layer1_outputs(4796) <= not a;
    layer1_outputs(4797) <= not b;
    layer1_outputs(4798) <= not a;
    layer1_outputs(4799) <= not (a or b);
    layer1_outputs(4800) <= a;
    layer1_outputs(4801) <= '0';
    layer1_outputs(4802) <= a and not b;
    layer1_outputs(4803) <= not (a and b);
    layer1_outputs(4804) <= not (a and b);
    layer1_outputs(4805) <= b;
    layer1_outputs(4806) <= not b or a;
    layer1_outputs(4807) <= b and not a;
    layer1_outputs(4808) <= a or b;
    layer1_outputs(4809) <= not a;
    layer1_outputs(4810) <= a and b;
    layer1_outputs(4811) <= not a or b;
    layer1_outputs(4812) <= b and not a;
    layer1_outputs(4813) <= '0';
    layer1_outputs(4814) <= b;
    layer1_outputs(4815) <= not b or a;
    layer1_outputs(4816) <= not a;
    layer1_outputs(4817) <= '1';
    layer1_outputs(4818) <= not a or b;
    layer1_outputs(4819) <= a;
    layer1_outputs(4820) <= not b;
    layer1_outputs(4821) <= '0';
    layer1_outputs(4822) <= a and b;
    layer1_outputs(4823) <= '0';
    layer1_outputs(4824) <= a and not b;
    layer1_outputs(4825) <= b;
    layer1_outputs(4826) <= not b or a;
    layer1_outputs(4827) <= a or b;
    layer1_outputs(4828) <= not a;
    layer1_outputs(4829) <= a;
    layer1_outputs(4830) <= a or b;
    layer1_outputs(4831) <= not (a xor b);
    layer1_outputs(4832) <= not (a and b);
    layer1_outputs(4833) <= not a or b;
    layer1_outputs(4834) <= not b;
    layer1_outputs(4835) <= b and not a;
    layer1_outputs(4836) <= b and not a;
    layer1_outputs(4837) <= '1';
    layer1_outputs(4838) <= a;
    layer1_outputs(4839) <= b;
    layer1_outputs(4840) <= a and b;
    layer1_outputs(4841) <= a xor b;
    layer1_outputs(4842) <= a;
    layer1_outputs(4843) <= a and not b;
    layer1_outputs(4844) <= a and b;
    layer1_outputs(4845) <= b;
    layer1_outputs(4846) <= '0';
    layer1_outputs(4847) <= a xor b;
    layer1_outputs(4848) <= not (a and b);
    layer1_outputs(4849) <= a;
    layer1_outputs(4850) <= '0';
    layer1_outputs(4851) <= not (a or b);
    layer1_outputs(4852) <= a and b;
    layer1_outputs(4853) <= not (a or b);
    layer1_outputs(4854) <= '0';
    layer1_outputs(4855) <= not b;
    layer1_outputs(4856) <= not a;
    layer1_outputs(4857) <= b;
    layer1_outputs(4858) <= '0';
    layer1_outputs(4859) <= '0';
    layer1_outputs(4860) <= b and not a;
    layer1_outputs(4861) <= not b;
    layer1_outputs(4862) <= not b or a;
    layer1_outputs(4863) <= not (a or b);
    layer1_outputs(4864) <= a xor b;
    layer1_outputs(4865) <= not b;
    layer1_outputs(4866) <= not a or b;
    layer1_outputs(4867) <= a and not b;
    layer1_outputs(4868) <= a xor b;
    layer1_outputs(4869) <= not b;
    layer1_outputs(4870) <= not (a xor b);
    layer1_outputs(4871) <= not a;
    layer1_outputs(4872) <= a and not b;
    layer1_outputs(4873) <= not (a or b);
    layer1_outputs(4874) <= b and not a;
    layer1_outputs(4875) <= a;
    layer1_outputs(4876) <= not b or a;
    layer1_outputs(4877) <= not b or a;
    layer1_outputs(4878) <= not (a and b);
    layer1_outputs(4879) <= not b;
    layer1_outputs(4880) <= not b or a;
    layer1_outputs(4881) <= b;
    layer1_outputs(4882) <= not a or b;
    layer1_outputs(4883) <= not b or a;
    layer1_outputs(4884) <= a or b;
    layer1_outputs(4885) <= '1';
    layer1_outputs(4886) <= not a;
    layer1_outputs(4887) <= b;
    layer1_outputs(4888) <= a xor b;
    layer1_outputs(4889) <= not b;
    layer1_outputs(4890) <= not b or a;
    layer1_outputs(4891) <= '1';
    layer1_outputs(4892) <= not b or a;
    layer1_outputs(4893) <= a and b;
    layer1_outputs(4894) <= a;
    layer1_outputs(4895) <= a or b;
    layer1_outputs(4896) <= not (a or b);
    layer1_outputs(4897) <= a and not b;
    layer1_outputs(4898) <= a;
    layer1_outputs(4899) <= not a or b;
    layer1_outputs(4900) <= not b;
    layer1_outputs(4901) <= '1';
    layer1_outputs(4902) <= a;
    layer1_outputs(4903) <= not a;
    layer1_outputs(4904) <= b and not a;
    layer1_outputs(4905) <= not a;
    layer1_outputs(4906) <= a and not b;
    layer1_outputs(4907) <= not (a or b);
    layer1_outputs(4908) <= not b or a;
    layer1_outputs(4909) <= not a;
    layer1_outputs(4910) <= b;
    layer1_outputs(4911) <= a xor b;
    layer1_outputs(4912) <= '1';
    layer1_outputs(4913) <= not (a or b);
    layer1_outputs(4914) <= a and b;
    layer1_outputs(4915) <= '0';
    layer1_outputs(4916) <= not b or a;
    layer1_outputs(4917) <= a xor b;
    layer1_outputs(4918) <= b;
    layer1_outputs(4919) <= b;
    layer1_outputs(4920) <= not a or b;
    layer1_outputs(4921) <= not (a and b);
    layer1_outputs(4922) <= a;
    layer1_outputs(4923) <= '1';
    layer1_outputs(4924) <= not a;
    layer1_outputs(4925) <= not a or b;
    layer1_outputs(4926) <= '1';
    layer1_outputs(4927) <= b;
    layer1_outputs(4928) <= a or b;
    layer1_outputs(4929) <= not b;
    layer1_outputs(4930) <= b;
    layer1_outputs(4931) <= '0';
    layer1_outputs(4932) <= '0';
    layer1_outputs(4933) <= b;
    layer1_outputs(4934) <= a;
    layer1_outputs(4935) <= a and b;
    layer1_outputs(4936) <= not b or a;
    layer1_outputs(4937) <= not b;
    layer1_outputs(4938) <= not (a and b);
    layer1_outputs(4939) <= a and not b;
    layer1_outputs(4940) <= a xor b;
    layer1_outputs(4941) <= not (a and b);
    layer1_outputs(4942) <= not a;
    layer1_outputs(4943) <= a or b;
    layer1_outputs(4944) <= b and not a;
    layer1_outputs(4945) <= b and not a;
    layer1_outputs(4946) <= not (a xor b);
    layer1_outputs(4947) <= not a or b;
    layer1_outputs(4948) <= a;
    layer1_outputs(4949) <= '0';
    layer1_outputs(4950) <= b and not a;
    layer1_outputs(4951) <= a;
    layer1_outputs(4952) <= not a;
    layer1_outputs(4953) <= a and not b;
    layer1_outputs(4954) <= a and not b;
    layer1_outputs(4955) <= a xor b;
    layer1_outputs(4956) <= not a or b;
    layer1_outputs(4957) <= '1';
    layer1_outputs(4958) <= not (a or b);
    layer1_outputs(4959) <= a and not b;
    layer1_outputs(4960) <= not a or b;
    layer1_outputs(4961) <= '1';
    layer1_outputs(4962) <= b;
    layer1_outputs(4963) <= not a;
    layer1_outputs(4964) <= '1';
    layer1_outputs(4965) <= a xor b;
    layer1_outputs(4966) <= not a or b;
    layer1_outputs(4967) <= b;
    layer1_outputs(4968) <= a;
    layer1_outputs(4969) <= '1';
    layer1_outputs(4970) <= not a or b;
    layer1_outputs(4971) <= not b;
    layer1_outputs(4972) <= a;
    layer1_outputs(4973) <= not (a and b);
    layer1_outputs(4974) <= not (a or b);
    layer1_outputs(4975) <= not (a xor b);
    layer1_outputs(4976) <= b and not a;
    layer1_outputs(4977) <= a and not b;
    layer1_outputs(4978) <= not a or b;
    layer1_outputs(4979) <= a;
    layer1_outputs(4980) <= a xor b;
    layer1_outputs(4981) <= a and not b;
    layer1_outputs(4982) <= a;
    layer1_outputs(4983) <= a;
    layer1_outputs(4984) <= not (a and b);
    layer1_outputs(4985) <= '1';
    layer1_outputs(4986) <= not (a or b);
    layer1_outputs(4987) <= a and not b;
    layer1_outputs(4988) <= not a or b;
    layer1_outputs(4989) <= b and not a;
    layer1_outputs(4990) <= '0';
    layer1_outputs(4991) <= a and not b;
    layer1_outputs(4992) <= '0';
    layer1_outputs(4993) <= b;
    layer1_outputs(4994) <= not (a or b);
    layer1_outputs(4995) <= not b;
    layer1_outputs(4996) <= a and b;
    layer1_outputs(4997) <= not (a or b);
    layer1_outputs(4998) <= a or b;
    layer1_outputs(4999) <= a or b;
    layer1_outputs(5000) <= '0';
    layer1_outputs(5001) <= not b or a;
    layer1_outputs(5002) <= not a or b;
    layer1_outputs(5003) <= a and b;
    layer1_outputs(5004) <= not (a xor b);
    layer1_outputs(5005) <= a or b;
    layer1_outputs(5006) <= a and not b;
    layer1_outputs(5007) <= a or b;
    layer1_outputs(5008) <= b;
    layer1_outputs(5009) <= b;
    layer1_outputs(5010) <= not (a or b);
    layer1_outputs(5011) <= not a;
    layer1_outputs(5012) <= a;
    layer1_outputs(5013) <= not (a and b);
    layer1_outputs(5014) <= not a;
    layer1_outputs(5015) <= not (a or b);
    layer1_outputs(5016) <= b and not a;
    layer1_outputs(5017) <= a and not b;
    layer1_outputs(5018) <= a or b;
    layer1_outputs(5019) <= not (a and b);
    layer1_outputs(5020) <= not (a or b);
    layer1_outputs(5021) <= b;
    layer1_outputs(5022) <= not b;
    layer1_outputs(5023) <= b;
    layer1_outputs(5024) <= a;
    layer1_outputs(5025) <= not a;
    layer1_outputs(5026) <= b;
    layer1_outputs(5027) <= a;
    layer1_outputs(5028) <= a;
    layer1_outputs(5029) <= not (a and b);
    layer1_outputs(5030) <= a and b;
    layer1_outputs(5031) <= b;
    layer1_outputs(5032) <= not a;
    layer1_outputs(5033) <= not (a or b);
    layer1_outputs(5034) <= '1';
    layer1_outputs(5035) <= not (a xor b);
    layer1_outputs(5036) <= not (a and b);
    layer1_outputs(5037) <= b and not a;
    layer1_outputs(5038) <= not b;
    layer1_outputs(5039) <= not b or a;
    layer1_outputs(5040) <= not b;
    layer1_outputs(5041) <= not (a and b);
    layer1_outputs(5042) <= b;
    layer1_outputs(5043) <= not a;
    layer1_outputs(5044) <= a and not b;
    layer1_outputs(5045) <= a and b;
    layer1_outputs(5046) <= not a;
    layer1_outputs(5047) <= not a;
    layer1_outputs(5048) <= a xor b;
    layer1_outputs(5049) <= a and b;
    layer1_outputs(5050) <= not a;
    layer1_outputs(5051) <= not a or b;
    layer1_outputs(5052) <= not b;
    layer1_outputs(5053) <= not b;
    layer1_outputs(5054) <= a and b;
    layer1_outputs(5055) <= not a or b;
    layer1_outputs(5056) <= '0';
    layer1_outputs(5057) <= '0';
    layer1_outputs(5058) <= b and not a;
    layer1_outputs(5059) <= a;
    layer1_outputs(5060) <= '0';
    layer1_outputs(5061) <= not b or a;
    layer1_outputs(5062) <= not a;
    layer1_outputs(5063) <= b;
    layer1_outputs(5064) <= a and not b;
    layer1_outputs(5065) <= a;
    layer1_outputs(5066) <= not a or b;
    layer1_outputs(5067) <= not (a and b);
    layer1_outputs(5068) <= '0';
    layer1_outputs(5069) <= '1';
    layer1_outputs(5070) <= not (a and b);
    layer1_outputs(5071) <= b;
    layer1_outputs(5072) <= not b;
    layer1_outputs(5073) <= a and not b;
    layer1_outputs(5074) <= b;
    layer1_outputs(5075) <= not (a or b);
    layer1_outputs(5076) <= not b;
    layer1_outputs(5077) <= a or b;
    layer1_outputs(5078) <= not (a and b);
    layer1_outputs(5079) <= not b or a;
    layer1_outputs(5080) <= '1';
    layer1_outputs(5081) <= a or b;
    layer1_outputs(5082) <= '0';
    layer1_outputs(5083) <= '0';
    layer1_outputs(5084) <= not (a xor b);
    layer1_outputs(5085) <= not a or b;
    layer1_outputs(5086) <= b;
    layer1_outputs(5087) <= not (a and b);
    layer1_outputs(5088) <= not a;
    layer1_outputs(5089) <= not a;
    layer1_outputs(5090) <= a and b;
    layer1_outputs(5091) <= not a or b;
    layer1_outputs(5092) <= not b;
    layer1_outputs(5093) <= b;
    layer1_outputs(5094) <= a or b;
    layer1_outputs(5095) <= not a;
    layer1_outputs(5096) <= not a or b;
    layer1_outputs(5097) <= a xor b;
    layer1_outputs(5098) <= a or b;
    layer1_outputs(5099) <= '1';
    layer1_outputs(5100) <= not (a or b);
    layer1_outputs(5101) <= not (a or b);
    layer1_outputs(5102) <= not (a or b);
    layer1_outputs(5103) <= a or b;
    layer1_outputs(5104) <= not (a xor b);
    layer1_outputs(5105) <= not (a or b);
    layer1_outputs(5106) <= '0';
    layer1_outputs(5107) <= a and not b;
    layer1_outputs(5108) <= a and b;
    layer1_outputs(5109) <= b and not a;
    layer1_outputs(5110) <= a and b;
    layer1_outputs(5111) <= not a;
    layer1_outputs(5112) <= not (a or b);
    layer1_outputs(5113) <= a and b;
    layer1_outputs(5114) <= not a;
    layer1_outputs(5115) <= not (a and b);
    layer1_outputs(5116) <= not b or a;
    layer1_outputs(5117) <= not (a xor b);
    layer1_outputs(5118) <= not b;
    layer1_outputs(5119) <= a xor b;
    layer1_outputs(5120) <= not (a or b);
    layer1_outputs(5121) <= b and not a;
    layer1_outputs(5122) <= not (a and b);
    layer1_outputs(5123) <= a;
    layer1_outputs(5124) <= not (a or b);
    layer1_outputs(5125) <= b;
    layer1_outputs(5126) <= '1';
    layer1_outputs(5127) <= '0';
    layer1_outputs(5128) <= not b;
    layer1_outputs(5129) <= a or b;
    layer1_outputs(5130) <= a xor b;
    layer1_outputs(5131) <= a and b;
    layer1_outputs(5132) <= a and not b;
    layer1_outputs(5133) <= not (a or b);
    layer1_outputs(5134) <= not b or a;
    layer1_outputs(5135) <= not a;
    layer1_outputs(5136) <= not (a and b);
    layer1_outputs(5137) <= b;
    layer1_outputs(5138) <= not (a xor b);
    layer1_outputs(5139) <= a and b;
    layer1_outputs(5140) <= not (a or b);
    layer1_outputs(5141) <= not (a or b);
    layer1_outputs(5142) <= not b or a;
    layer1_outputs(5143) <= a and b;
    layer1_outputs(5144) <= not (a or b);
    layer1_outputs(5145) <= not a or b;
    layer1_outputs(5146) <= a or b;
    layer1_outputs(5147) <= not b;
    layer1_outputs(5148) <= b;
    layer1_outputs(5149) <= b;
    layer1_outputs(5150) <= not (a or b);
    layer1_outputs(5151) <= '1';
    layer1_outputs(5152) <= '1';
    layer1_outputs(5153) <= not (a and b);
    layer1_outputs(5154) <= b;
    layer1_outputs(5155) <= a and not b;
    layer1_outputs(5156) <= not b;
    layer1_outputs(5157) <= not a;
    layer1_outputs(5158) <= not b or a;
    layer1_outputs(5159) <= '1';
    layer1_outputs(5160) <= b and not a;
    layer1_outputs(5161) <= a xor b;
    layer1_outputs(5162) <= a xor b;
    layer1_outputs(5163) <= b and not a;
    layer1_outputs(5164) <= not a;
    layer1_outputs(5165) <= b and not a;
    layer1_outputs(5166) <= '0';
    layer1_outputs(5167) <= a or b;
    layer1_outputs(5168) <= b;
    layer1_outputs(5169) <= not (a or b);
    layer1_outputs(5170) <= a and not b;
    layer1_outputs(5171) <= not a;
    layer1_outputs(5172) <= '0';
    layer1_outputs(5173) <= b;
    layer1_outputs(5174) <= not b;
    layer1_outputs(5175) <= not b;
    layer1_outputs(5176) <= a;
    layer1_outputs(5177) <= b;
    layer1_outputs(5178) <= a and b;
    layer1_outputs(5179) <= b;
    layer1_outputs(5180) <= b and not a;
    layer1_outputs(5181) <= a;
    layer1_outputs(5182) <= not b;
    layer1_outputs(5183) <= not a;
    layer1_outputs(5184) <= not (a and b);
    layer1_outputs(5185) <= not (a and b);
    layer1_outputs(5186) <= b and not a;
    layer1_outputs(5187) <= a;
    layer1_outputs(5188) <= not a or b;
    layer1_outputs(5189) <= not a;
    layer1_outputs(5190) <= not a or b;
    layer1_outputs(5191) <= not (a and b);
    layer1_outputs(5192) <= not (a and b);
    layer1_outputs(5193) <= b and not a;
    layer1_outputs(5194) <= not (a or b);
    layer1_outputs(5195) <= not (a xor b);
    layer1_outputs(5196) <= not (a or b);
    layer1_outputs(5197) <= not b;
    layer1_outputs(5198) <= a;
    layer1_outputs(5199) <= not a;
    layer1_outputs(5200) <= not b or a;
    layer1_outputs(5201) <= not a;
    layer1_outputs(5202) <= a;
    layer1_outputs(5203) <= not (a or b);
    layer1_outputs(5204) <= '1';
    layer1_outputs(5205) <= not a or b;
    layer1_outputs(5206) <= not (a or b);
    layer1_outputs(5207) <= a and b;
    layer1_outputs(5208) <= b;
    layer1_outputs(5209) <= b and not a;
    layer1_outputs(5210) <= not a;
    layer1_outputs(5211) <= not b or a;
    layer1_outputs(5212) <= not a or b;
    layer1_outputs(5213) <= not a or b;
    layer1_outputs(5214) <= a and b;
    layer1_outputs(5215) <= not b or a;
    layer1_outputs(5216) <= not (a and b);
    layer1_outputs(5217) <= not a or b;
    layer1_outputs(5218) <= b;
    layer1_outputs(5219) <= b and not a;
    layer1_outputs(5220) <= not (a xor b);
    layer1_outputs(5221) <= not b;
    layer1_outputs(5222) <= not a;
    layer1_outputs(5223) <= not a or b;
    layer1_outputs(5224) <= b;
    layer1_outputs(5225) <= not b or a;
    layer1_outputs(5226) <= not (a or b);
    layer1_outputs(5227) <= not (a and b);
    layer1_outputs(5228) <= a and not b;
    layer1_outputs(5229) <= b and not a;
    layer1_outputs(5230) <= not a;
    layer1_outputs(5231) <= not a;
    layer1_outputs(5232) <= not b or a;
    layer1_outputs(5233) <= b;
    layer1_outputs(5234) <= not b;
    layer1_outputs(5235) <= a and b;
    layer1_outputs(5236) <= not (a xor b);
    layer1_outputs(5237) <= '0';
    layer1_outputs(5238) <= a or b;
    layer1_outputs(5239) <= not a or b;
    layer1_outputs(5240) <= b;
    layer1_outputs(5241) <= not (a or b);
    layer1_outputs(5242) <= not b or a;
    layer1_outputs(5243) <= a;
    layer1_outputs(5244) <= b;
    layer1_outputs(5245) <= not (a or b);
    layer1_outputs(5246) <= '0';
    layer1_outputs(5247) <= not (a and b);
    layer1_outputs(5248) <= not b;
    layer1_outputs(5249) <= a;
    layer1_outputs(5250) <= not (a or b);
    layer1_outputs(5251) <= not a;
    layer1_outputs(5252) <= not (a and b);
    layer1_outputs(5253) <= not (a and b);
    layer1_outputs(5254) <= not (a and b);
    layer1_outputs(5255) <= not b or a;
    layer1_outputs(5256) <= not b;
    layer1_outputs(5257) <= a or b;
    layer1_outputs(5258) <= b and not a;
    layer1_outputs(5259) <= a;
    layer1_outputs(5260) <= not b;
    layer1_outputs(5261) <= not (a and b);
    layer1_outputs(5262) <= not (a or b);
    layer1_outputs(5263) <= not a;
    layer1_outputs(5264) <= b and not a;
    layer1_outputs(5265) <= a or b;
    layer1_outputs(5266) <= a and not b;
    layer1_outputs(5267) <= a and b;
    layer1_outputs(5268) <= not (a and b);
    layer1_outputs(5269) <= a or b;
    layer1_outputs(5270) <= '0';
    layer1_outputs(5271) <= a or b;
    layer1_outputs(5272) <= not b;
    layer1_outputs(5273) <= a and b;
    layer1_outputs(5274) <= not (a or b);
    layer1_outputs(5275) <= a;
    layer1_outputs(5276) <= not a or b;
    layer1_outputs(5277) <= a and b;
    layer1_outputs(5278) <= not (a and b);
    layer1_outputs(5279) <= b;
    layer1_outputs(5280) <= not (a and b);
    layer1_outputs(5281) <= a or b;
    layer1_outputs(5282) <= not b;
    layer1_outputs(5283) <= not b;
    layer1_outputs(5284) <= not b or a;
    layer1_outputs(5285) <= b;
    layer1_outputs(5286) <= b;
    layer1_outputs(5287) <= a and b;
    layer1_outputs(5288) <= not a or b;
    layer1_outputs(5289) <= a xor b;
    layer1_outputs(5290) <= b;
    layer1_outputs(5291) <= b;
    layer1_outputs(5292) <= a and b;
    layer1_outputs(5293) <= '1';
    layer1_outputs(5294) <= not b;
    layer1_outputs(5295) <= b and not a;
    layer1_outputs(5296) <= '0';
    layer1_outputs(5297) <= '1';
    layer1_outputs(5298) <= '0';
    layer1_outputs(5299) <= a and not b;
    layer1_outputs(5300) <= b;
    layer1_outputs(5301) <= '0';
    layer1_outputs(5302) <= b;
    layer1_outputs(5303) <= b and not a;
    layer1_outputs(5304) <= '1';
    layer1_outputs(5305) <= '1';
    layer1_outputs(5306) <= b;
    layer1_outputs(5307) <= not (a xor b);
    layer1_outputs(5308) <= not a;
    layer1_outputs(5309) <= b and not a;
    layer1_outputs(5310) <= not b or a;
    layer1_outputs(5311) <= not b or a;
    layer1_outputs(5312) <= a and not b;
    layer1_outputs(5313) <= not b;
    layer1_outputs(5314) <= '1';
    layer1_outputs(5315) <= '1';
    layer1_outputs(5316) <= not a or b;
    layer1_outputs(5317) <= not a;
    layer1_outputs(5318) <= a and b;
    layer1_outputs(5319) <= b and not a;
    layer1_outputs(5320) <= not b;
    layer1_outputs(5321) <= not (a or b);
    layer1_outputs(5322) <= not b;
    layer1_outputs(5323) <= not (a or b);
    layer1_outputs(5324) <= '1';
    layer1_outputs(5325) <= not b;
    layer1_outputs(5326) <= not b;
    layer1_outputs(5327) <= not (a or b);
    layer1_outputs(5328) <= not b or a;
    layer1_outputs(5329) <= not b;
    layer1_outputs(5330) <= b;
    layer1_outputs(5331) <= not (a and b);
    layer1_outputs(5332) <= not (a or b);
    layer1_outputs(5333) <= not (a or b);
    layer1_outputs(5334) <= b and not a;
    layer1_outputs(5335) <= not b;
    layer1_outputs(5336) <= not (a and b);
    layer1_outputs(5337) <= b;
    layer1_outputs(5338) <= '0';
    layer1_outputs(5339) <= not (a or b);
    layer1_outputs(5340) <= a and b;
    layer1_outputs(5341) <= not b;
    layer1_outputs(5342) <= a;
    layer1_outputs(5343) <= '0';
    layer1_outputs(5344) <= b and not a;
    layer1_outputs(5345) <= not (a xor b);
    layer1_outputs(5346) <= a or b;
    layer1_outputs(5347) <= not b;
    layer1_outputs(5348) <= not a or b;
    layer1_outputs(5349) <= a and not b;
    layer1_outputs(5350) <= a and b;
    layer1_outputs(5351) <= a;
    layer1_outputs(5352) <= b and not a;
    layer1_outputs(5353) <= '0';
    layer1_outputs(5354) <= not a;
    layer1_outputs(5355) <= not b;
    layer1_outputs(5356) <= not b or a;
    layer1_outputs(5357) <= a and b;
    layer1_outputs(5358) <= a and b;
    layer1_outputs(5359) <= not a or b;
    layer1_outputs(5360) <= a and not b;
    layer1_outputs(5361) <= b;
    layer1_outputs(5362) <= '0';
    layer1_outputs(5363) <= not (a or b);
    layer1_outputs(5364) <= not (a xor b);
    layer1_outputs(5365) <= '1';
    layer1_outputs(5366) <= not b or a;
    layer1_outputs(5367) <= not a;
    layer1_outputs(5368) <= a;
    layer1_outputs(5369) <= not b or a;
    layer1_outputs(5370) <= not a or b;
    layer1_outputs(5371) <= not a or b;
    layer1_outputs(5372) <= not b or a;
    layer1_outputs(5373) <= b;
    layer1_outputs(5374) <= not b;
    layer1_outputs(5375) <= '0';
    layer1_outputs(5376) <= not (a or b);
    layer1_outputs(5377) <= not b or a;
    layer1_outputs(5378) <= a and b;
    layer1_outputs(5379) <= '0';
    layer1_outputs(5380) <= '0';
    layer1_outputs(5381) <= not a or b;
    layer1_outputs(5382) <= b and not a;
    layer1_outputs(5383) <= not b;
    layer1_outputs(5384) <= not (a and b);
    layer1_outputs(5385) <= not (a and b);
    layer1_outputs(5386) <= a or b;
    layer1_outputs(5387) <= not b or a;
    layer1_outputs(5388) <= not a;
    layer1_outputs(5389) <= not b or a;
    layer1_outputs(5390) <= not a;
    layer1_outputs(5391) <= not (a and b);
    layer1_outputs(5392) <= not a;
    layer1_outputs(5393) <= b;
    layer1_outputs(5394) <= not a or b;
    layer1_outputs(5395) <= a or b;
    layer1_outputs(5396) <= not (a xor b);
    layer1_outputs(5397) <= a or b;
    layer1_outputs(5398) <= '1';
    layer1_outputs(5399) <= not b or a;
    layer1_outputs(5400) <= not b;
    layer1_outputs(5401) <= b;
    layer1_outputs(5402) <= b;
    layer1_outputs(5403) <= a and b;
    layer1_outputs(5404) <= not (a and b);
    layer1_outputs(5405) <= b;
    layer1_outputs(5406) <= not (a or b);
    layer1_outputs(5407) <= '1';
    layer1_outputs(5408) <= not b or a;
    layer1_outputs(5409) <= not (a and b);
    layer1_outputs(5410) <= not b or a;
    layer1_outputs(5411) <= not (a or b);
    layer1_outputs(5412) <= a xor b;
    layer1_outputs(5413) <= a or b;
    layer1_outputs(5414) <= b and not a;
    layer1_outputs(5415) <= not (a and b);
    layer1_outputs(5416) <= not b;
    layer1_outputs(5417) <= '0';
    layer1_outputs(5418) <= a or b;
    layer1_outputs(5419) <= not b or a;
    layer1_outputs(5420) <= b;
    layer1_outputs(5421) <= not a;
    layer1_outputs(5422) <= a;
    layer1_outputs(5423) <= not (a or b);
    layer1_outputs(5424) <= a and b;
    layer1_outputs(5425) <= a;
    layer1_outputs(5426) <= not (a xor b);
    layer1_outputs(5427) <= '1';
    layer1_outputs(5428) <= a and b;
    layer1_outputs(5429) <= '1';
    layer1_outputs(5430) <= a or b;
    layer1_outputs(5431) <= not b or a;
    layer1_outputs(5432) <= b;
    layer1_outputs(5433) <= not b or a;
    layer1_outputs(5434) <= b;
    layer1_outputs(5435) <= a and not b;
    layer1_outputs(5436) <= b;
    layer1_outputs(5437) <= not a or b;
    layer1_outputs(5438) <= a;
    layer1_outputs(5439) <= not a;
    layer1_outputs(5440) <= b;
    layer1_outputs(5441) <= a;
    layer1_outputs(5442) <= '0';
    layer1_outputs(5443) <= a;
    layer1_outputs(5444) <= a and not b;
    layer1_outputs(5445) <= '0';
    layer1_outputs(5446) <= not b;
    layer1_outputs(5447) <= not (a and b);
    layer1_outputs(5448) <= a or b;
    layer1_outputs(5449) <= not a;
    layer1_outputs(5450) <= b and not a;
    layer1_outputs(5451) <= not (a and b);
    layer1_outputs(5452) <= not b;
    layer1_outputs(5453) <= a;
    layer1_outputs(5454) <= a;
    layer1_outputs(5455) <= not (a and b);
    layer1_outputs(5456) <= '0';
    layer1_outputs(5457) <= not b or a;
    layer1_outputs(5458) <= not b;
    layer1_outputs(5459) <= not b or a;
    layer1_outputs(5460) <= not (a or b);
    layer1_outputs(5461) <= a and not b;
    layer1_outputs(5462) <= a and b;
    layer1_outputs(5463) <= not (a and b);
    layer1_outputs(5464) <= not (a or b);
    layer1_outputs(5465) <= a or b;
    layer1_outputs(5466) <= a or b;
    layer1_outputs(5467) <= a and not b;
    layer1_outputs(5468) <= a xor b;
    layer1_outputs(5469) <= b;
    layer1_outputs(5470) <= not a;
    layer1_outputs(5471) <= not a or b;
    layer1_outputs(5472) <= not a or b;
    layer1_outputs(5473) <= not (a and b);
    layer1_outputs(5474) <= not a;
    layer1_outputs(5475) <= a and b;
    layer1_outputs(5476) <= not b;
    layer1_outputs(5477) <= a and b;
    layer1_outputs(5478) <= a xor b;
    layer1_outputs(5479) <= not (a and b);
    layer1_outputs(5480) <= not (a xor b);
    layer1_outputs(5481) <= b;
    layer1_outputs(5482) <= a and b;
    layer1_outputs(5483) <= b;
    layer1_outputs(5484) <= not a or b;
    layer1_outputs(5485) <= '0';
    layer1_outputs(5486) <= not b;
    layer1_outputs(5487) <= not b or a;
    layer1_outputs(5488) <= not (a and b);
    layer1_outputs(5489) <= a and b;
    layer1_outputs(5490) <= a and b;
    layer1_outputs(5491) <= not (a and b);
    layer1_outputs(5492) <= not (a and b);
    layer1_outputs(5493) <= not b;
    layer1_outputs(5494) <= not b;
    layer1_outputs(5495) <= not (a xor b);
    layer1_outputs(5496) <= a or b;
    layer1_outputs(5497) <= a;
    layer1_outputs(5498) <= b and not a;
    layer1_outputs(5499) <= not b or a;
    layer1_outputs(5500) <= not a or b;
    layer1_outputs(5501) <= '1';
    layer1_outputs(5502) <= b and not a;
    layer1_outputs(5503) <= a xor b;
    layer1_outputs(5504) <= a or b;
    layer1_outputs(5505) <= a or b;
    layer1_outputs(5506) <= a or b;
    layer1_outputs(5507) <= '1';
    layer1_outputs(5508) <= not b;
    layer1_outputs(5509) <= '1';
    layer1_outputs(5510) <= a;
    layer1_outputs(5511) <= b;
    layer1_outputs(5512) <= '1';
    layer1_outputs(5513) <= a;
    layer1_outputs(5514) <= not b;
    layer1_outputs(5515) <= not a;
    layer1_outputs(5516) <= b and not a;
    layer1_outputs(5517) <= not b or a;
    layer1_outputs(5518) <= '0';
    layer1_outputs(5519) <= '0';
    layer1_outputs(5520) <= a and b;
    layer1_outputs(5521) <= b and not a;
    layer1_outputs(5522) <= b;
    layer1_outputs(5523) <= a or b;
    layer1_outputs(5524) <= a;
    layer1_outputs(5525) <= a and not b;
    layer1_outputs(5526) <= '1';
    layer1_outputs(5527) <= a and not b;
    layer1_outputs(5528) <= not b;
    layer1_outputs(5529) <= a xor b;
    layer1_outputs(5530) <= not b;
    layer1_outputs(5531) <= not a or b;
    layer1_outputs(5532) <= not b;
    layer1_outputs(5533) <= b;
    layer1_outputs(5534) <= not a;
    layer1_outputs(5535) <= a xor b;
    layer1_outputs(5536) <= a or b;
    layer1_outputs(5537) <= not b or a;
    layer1_outputs(5538) <= not (a and b);
    layer1_outputs(5539) <= not b;
    layer1_outputs(5540) <= not (a or b);
    layer1_outputs(5541) <= a and not b;
    layer1_outputs(5542) <= a;
    layer1_outputs(5543) <= not b;
    layer1_outputs(5544) <= '1';
    layer1_outputs(5545) <= not (a or b);
    layer1_outputs(5546) <= not a;
    layer1_outputs(5547) <= '1';
    layer1_outputs(5548) <= b and not a;
    layer1_outputs(5549) <= not b or a;
    layer1_outputs(5550) <= not (a xor b);
    layer1_outputs(5551) <= not a or b;
    layer1_outputs(5552) <= '1';
    layer1_outputs(5553) <= b;
    layer1_outputs(5554) <= b and not a;
    layer1_outputs(5555) <= a or b;
    layer1_outputs(5556) <= not b or a;
    layer1_outputs(5557) <= a;
    layer1_outputs(5558) <= not (a and b);
    layer1_outputs(5559) <= not b or a;
    layer1_outputs(5560) <= b and not a;
    layer1_outputs(5561) <= not (a xor b);
    layer1_outputs(5562) <= b and not a;
    layer1_outputs(5563) <= a or b;
    layer1_outputs(5564) <= a;
    layer1_outputs(5565) <= a;
    layer1_outputs(5566) <= b;
    layer1_outputs(5567) <= not a;
    layer1_outputs(5568) <= b;
    layer1_outputs(5569) <= b and not a;
    layer1_outputs(5570) <= b and not a;
    layer1_outputs(5571) <= a xor b;
    layer1_outputs(5572) <= a;
    layer1_outputs(5573) <= a and b;
    layer1_outputs(5574) <= not a;
    layer1_outputs(5575) <= b;
    layer1_outputs(5576) <= b and not a;
    layer1_outputs(5577) <= '1';
    layer1_outputs(5578) <= a;
    layer1_outputs(5579) <= not b;
    layer1_outputs(5580) <= b;
    layer1_outputs(5581) <= not (a and b);
    layer1_outputs(5582) <= a;
    layer1_outputs(5583) <= not (a or b);
    layer1_outputs(5584) <= not a;
    layer1_outputs(5585) <= a and not b;
    layer1_outputs(5586) <= not (a xor b);
    layer1_outputs(5587) <= b;
    layer1_outputs(5588) <= not b;
    layer1_outputs(5589) <= a;
    layer1_outputs(5590) <= not b;
    layer1_outputs(5591) <= a and b;
    layer1_outputs(5592) <= a;
    layer1_outputs(5593) <= not (a or b);
    layer1_outputs(5594) <= not b;
    layer1_outputs(5595) <= '1';
    layer1_outputs(5596) <= not b;
    layer1_outputs(5597) <= b and not a;
    layer1_outputs(5598) <= a;
    layer1_outputs(5599) <= a and b;
    layer1_outputs(5600) <= not a or b;
    layer1_outputs(5601) <= not b;
    layer1_outputs(5602) <= not (a or b);
    layer1_outputs(5603) <= a and not b;
    layer1_outputs(5604) <= not (a or b);
    layer1_outputs(5605) <= a or b;
    layer1_outputs(5606) <= a or b;
    layer1_outputs(5607) <= not a;
    layer1_outputs(5608) <= a or b;
    layer1_outputs(5609) <= b;
    layer1_outputs(5610) <= a and not b;
    layer1_outputs(5611) <= b;
    layer1_outputs(5612) <= a or b;
    layer1_outputs(5613) <= not b or a;
    layer1_outputs(5614) <= not b;
    layer1_outputs(5615) <= b and not a;
    layer1_outputs(5616) <= a or b;
    layer1_outputs(5617) <= b;
    layer1_outputs(5618) <= not (a and b);
    layer1_outputs(5619) <= not (a xor b);
    layer1_outputs(5620) <= not a or b;
    layer1_outputs(5621) <= a and not b;
    layer1_outputs(5622) <= a;
    layer1_outputs(5623) <= '0';
    layer1_outputs(5624) <= b and not a;
    layer1_outputs(5625) <= not (a and b);
    layer1_outputs(5626) <= not a or b;
    layer1_outputs(5627) <= not b or a;
    layer1_outputs(5628) <= not (a or b);
    layer1_outputs(5629) <= a and not b;
    layer1_outputs(5630) <= b;
    layer1_outputs(5631) <= a and not b;
    layer1_outputs(5632) <= not b or a;
    layer1_outputs(5633) <= b and not a;
    layer1_outputs(5634) <= not a or b;
    layer1_outputs(5635) <= b and not a;
    layer1_outputs(5636) <= a and b;
    layer1_outputs(5637) <= not b or a;
    layer1_outputs(5638) <= b;
    layer1_outputs(5639) <= a or b;
    layer1_outputs(5640) <= a and not b;
    layer1_outputs(5641) <= a;
    layer1_outputs(5642) <= not b or a;
    layer1_outputs(5643) <= not (a xor b);
    layer1_outputs(5644) <= not b;
    layer1_outputs(5645) <= not (a xor b);
    layer1_outputs(5646) <= a;
    layer1_outputs(5647) <= not a;
    layer1_outputs(5648) <= '1';
    layer1_outputs(5649) <= not b;
    layer1_outputs(5650) <= not b or a;
    layer1_outputs(5651) <= a and not b;
    layer1_outputs(5652) <= a;
    layer1_outputs(5653) <= b;
    layer1_outputs(5654) <= '0';
    layer1_outputs(5655) <= not a or b;
    layer1_outputs(5656) <= a;
    layer1_outputs(5657) <= not (a or b);
    layer1_outputs(5658) <= b;
    layer1_outputs(5659) <= a;
    layer1_outputs(5660) <= '1';
    layer1_outputs(5661) <= b;
    layer1_outputs(5662) <= not (a xor b);
    layer1_outputs(5663) <= a and not b;
    layer1_outputs(5664) <= b;
    layer1_outputs(5665) <= not b or a;
    layer1_outputs(5666) <= not (a and b);
    layer1_outputs(5667) <= a xor b;
    layer1_outputs(5668) <= a;
    layer1_outputs(5669) <= a and not b;
    layer1_outputs(5670) <= not a or b;
    layer1_outputs(5671) <= not (a or b);
    layer1_outputs(5672) <= '1';
    layer1_outputs(5673) <= not (a and b);
    layer1_outputs(5674) <= b and not a;
    layer1_outputs(5675) <= a and b;
    layer1_outputs(5676) <= a;
    layer1_outputs(5677) <= a and not b;
    layer1_outputs(5678) <= a or b;
    layer1_outputs(5679) <= not a or b;
    layer1_outputs(5680) <= '1';
    layer1_outputs(5681) <= b;
    layer1_outputs(5682) <= not b;
    layer1_outputs(5683) <= not (a or b);
    layer1_outputs(5684) <= '1';
    layer1_outputs(5685) <= not a;
    layer1_outputs(5686) <= '1';
    layer1_outputs(5687) <= b;
    layer1_outputs(5688) <= b and not a;
    layer1_outputs(5689) <= a and not b;
    layer1_outputs(5690) <= not a or b;
    layer1_outputs(5691) <= a and b;
    layer1_outputs(5692) <= '1';
    layer1_outputs(5693) <= not (a or b);
    layer1_outputs(5694) <= b;
    layer1_outputs(5695) <= a and b;
    layer1_outputs(5696) <= a and b;
    layer1_outputs(5697) <= not (a or b);
    layer1_outputs(5698) <= not b;
    layer1_outputs(5699) <= '1';
    layer1_outputs(5700) <= not (a or b);
    layer1_outputs(5701) <= a or b;
    layer1_outputs(5702) <= '0';
    layer1_outputs(5703) <= a;
    layer1_outputs(5704) <= a and b;
    layer1_outputs(5705) <= a;
    layer1_outputs(5706) <= a or b;
    layer1_outputs(5707) <= '0';
    layer1_outputs(5708) <= '1';
    layer1_outputs(5709) <= not a or b;
    layer1_outputs(5710) <= a;
    layer1_outputs(5711) <= a or b;
    layer1_outputs(5712) <= not (a or b);
    layer1_outputs(5713) <= not b;
    layer1_outputs(5714) <= not (a and b);
    layer1_outputs(5715) <= not (a and b);
    layer1_outputs(5716) <= '0';
    layer1_outputs(5717) <= not b or a;
    layer1_outputs(5718) <= '0';
    layer1_outputs(5719) <= b;
    layer1_outputs(5720) <= not (a xor b);
    layer1_outputs(5721) <= not a;
    layer1_outputs(5722) <= a and not b;
    layer1_outputs(5723) <= '0';
    layer1_outputs(5724) <= a and not b;
    layer1_outputs(5725) <= not b;
    layer1_outputs(5726) <= not b or a;
    layer1_outputs(5727) <= '0';
    layer1_outputs(5728) <= not (a and b);
    layer1_outputs(5729) <= not a;
    layer1_outputs(5730) <= not b;
    layer1_outputs(5731) <= a and b;
    layer1_outputs(5732) <= b;
    layer1_outputs(5733) <= not (a and b);
    layer1_outputs(5734) <= not b;
    layer1_outputs(5735) <= not (a and b);
    layer1_outputs(5736) <= not (a and b);
    layer1_outputs(5737) <= a;
    layer1_outputs(5738) <= b;
    layer1_outputs(5739) <= a xor b;
    layer1_outputs(5740) <= '1';
    layer1_outputs(5741) <= a and b;
    layer1_outputs(5742) <= a or b;
    layer1_outputs(5743) <= b;
    layer1_outputs(5744) <= a and not b;
    layer1_outputs(5745) <= not b or a;
    layer1_outputs(5746) <= b;
    layer1_outputs(5747) <= not b;
    layer1_outputs(5748) <= not b;
    layer1_outputs(5749) <= b and not a;
    layer1_outputs(5750) <= a;
    layer1_outputs(5751) <= not a;
    layer1_outputs(5752) <= '1';
    layer1_outputs(5753) <= a xor b;
    layer1_outputs(5754) <= a and b;
    layer1_outputs(5755) <= not (a or b);
    layer1_outputs(5756) <= not a;
    layer1_outputs(5757) <= not (a and b);
    layer1_outputs(5758) <= b;
    layer1_outputs(5759) <= not b;
    layer1_outputs(5760) <= a and b;
    layer1_outputs(5761) <= b;
    layer1_outputs(5762) <= not a;
    layer1_outputs(5763) <= b and not a;
    layer1_outputs(5764) <= not a;
    layer1_outputs(5765) <= not b or a;
    layer1_outputs(5766) <= not b;
    layer1_outputs(5767) <= b;
    layer1_outputs(5768) <= a and not b;
    layer1_outputs(5769) <= b;
    layer1_outputs(5770) <= b;
    layer1_outputs(5771) <= not b or a;
    layer1_outputs(5772) <= a;
    layer1_outputs(5773) <= a and b;
    layer1_outputs(5774) <= not a or b;
    layer1_outputs(5775) <= not b;
    layer1_outputs(5776) <= b and not a;
    layer1_outputs(5777) <= a and b;
    layer1_outputs(5778) <= not b;
    layer1_outputs(5779) <= not b;
    layer1_outputs(5780) <= not b;
    layer1_outputs(5781) <= a and b;
    layer1_outputs(5782) <= not (a or b);
    layer1_outputs(5783) <= not a;
    layer1_outputs(5784) <= a and b;
    layer1_outputs(5785) <= not b or a;
    layer1_outputs(5786) <= not b;
    layer1_outputs(5787) <= not a;
    layer1_outputs(5788) <= not (a or b);
    layer1_outputs(5789) <= a or b;
    layer1_outputs(5790) <= a and b;
    layer1_outputs(5791) <= not (a or b);
    layer1_outputs(5792) <= not a;
    layer1_outputs(5793) <= not b or a;
    layer1_outputs(5794) <= not a or b;
    layer1_outputs(5795) <= '0';
    layer1_outputs(5796) <= not (a xor b);
    layer1_outputs(5797) <= a and b;
    layer1_outputs(5798) <= not b or a;
    layer1_outputs(5799) <= not b or a;
    layer1_outputs(5800) <= '0';
    layer1_outputs(5801) <= b;
    layer1_outputs(5802) <= '0';
    layer1_outputs(5803) <= not b;
    layer1_outputs(5804) <= not a;
    layer1_outputs(5805) <= not b or a;
    layer1_outputs(5806) <= not b or a;
    layer1_outputs(5807) <= not (a and b);
    layer1_outputs(5808) <= not (a xor b);
    layer1_outputs(5809) <= not (a or b);
    layer1_outputs(5810) <= b and not a;
    layer1_outputs(5811) <= not a;
    layer1_outputs(5812) <= not (a or b);
    layer1_outputs(5813) <= a or b;
    layer1_outputs(5814) <= b;
    layer1_outputs(5815) <= not (a and b);
    layer1_outputs(5816) <= not (a or b);
    layer1_outputs(5817) <= not a;
    layer1_outputs(5818) <= b;
    layer1_outputs(5819) <= b and not a;
    layer1_outputs(5820) <= b;
    layer1_outputs(5821) <= a;
    layer1_outputs(5822) <= not (a xor b);
    layer1_outputs(5823) <= not (a xor b);
    layer1_outputs(5824) <= b;
    layer1_outputs(5825) <= not b;
    layer1_outputs(5826) <= a xor b;
    layer1_outputs(5827) <= '0';
    layer1_outputs(5828) <= not a;
    layer1_outputs(5829) <= not (a and b);
    layer1_outputs(5830) <= b and not a;
    layer1_outputs(5831) <= a xor b;
    layer1_outputs(5832) <= not b or a;
    layer1_outputs(5833) <= a and not b;
    layer1_outputs(5834) <= a and b;
    layer1_outputs(5835) <= b;
    layer1_outputs(5836) <= a or b;
    layer1_outputs(5837) <= not (a or b);
    layer1_outputs(5838) <= not b;
    layer1_outputs(5839) <= b and not a;
    layer1_outputs(5840) <= not (a or b);
    layer1_outputs(5841) <= not b or a;
    layer1_outputs(5842) <= '1';
    layer1_outputs(5843) <= not (a or b);
    layer1_outputs(5844) <= a and not b;
    layer1_outputs(5845) <= not a or b;
    layer1_outputs(5846) <= not (a and b);
    layer1_outputs(5847) <= a and not b;
    layer1_outputs(5848) <= not b or a;
    layer1_outputs(5849) <= not a or b;
    layer1_outputs(5850) <= not a;
    layer1_outputs(5851) <= not b;
    layer1_outputs(5852) <= a or b;
    layer1_outputs(5853) <= '0';
    layer1_outputs(5854) <= not b or a;
    layer1_outputs(5855) <= not (a or b);
    layer1_outputs(5856) <= b and not a;
    layer1_outputs(5857) <= a;
    layer1_outputs(5858) <= a;
    layer1_outputs(5859) <= a and not b;
    layer1_outputs(5860) <= b and not a;
    layer1_outputs(5861) <= b;
    layer1_outputs(5862) <= a and b;
    layer1_outputs(5863) <= a or b;
    layer1_outputs(5864) <= b and not a;
    layer1_outputs(5865) <= not b;
    layer1_outputs(5866) <= not b;
    layer1_outputs(5867) <= b;
    layer1_outputs(5868) <= not a;
    layer1_outputs(5869) <= not b;
    layer1_outputs(5870) <= b;
    layer1_outputs(5871) <= a and not b;
    layer1_outputs(5872) <= a xor b;
    layer1_outputs(5873) <= not b;
    layer1_outputs(5874) <= not (a and b);
    layer1_outputs(5875) <= b and not a;
    layer1_outputs(5876) <= '1';
    layer1_outputs(5877) <= a;
    layer1_outputs(5878) <= a and b;
    layer1_outputs(5879) <= '1';
    layer1_outputs(5880) <= '1';
    layer1_outputs(5881) <= '1';
    layer1_outputs(5882) <= a or b;
    layer1_outputs(5883) <= not b;
    layer1_outputs(5884) <= '0';
    layer1_outputs(5885) <= not a or b;
    layer1_outputs(5886) <= '1';
    layer1_outputs(5887) <= '1';
    layer1_outputs(5888) <= a;
    layer1_outputs(5889) <= not (a and b);
    layer1_outputs(5890) <= a or b;
    layer1_outputs(5891) <= not b;
    layer1_outputs(5892) <= not (a or b);
    layer1_outputs(5893) <= not b or a;
    layer1_outputs(5894) <= not b;
    layer1_outputs(5895) <= not (a or b);
    layer1_outputs(5896) <= a and not b;
    layer1_outputs(5897) <= a or b;
    layer1_outputs(5898) <= not b;
    layer1_outputs(5899) <= '1';
    layer1_outputs(5900) <= not a;
    layer1_outputs(5901) <= not a or b;
    layer1_outputs(5902) <= '0';
    layer1_outputs(5903) <= a;
    layer1_outputs(5904) <= a and b;
    layer1_outputs(5905) <= a xor b;
    layer1_outputs(5906) <= a;
    layer1_outputs(5907) <= a;
    layer1_outputs(5908) <= not a;
    layer1_outputs(5909) <= a and b;
    layer1_outputs(5910) <= not b;
    layer1_outputs(5911) <= b and not a;
    layer1_outputs(5912) <= b;
    layer1_outputs(5913) <= '1';
    layer1_outputs(5914) <= b and not a;
    layer1_outputs(5915) <= a xor b;
    layer1_outputs(5916) <= not (a xor b);
    layer1_outputs(5917) <= not a or b;
    layer1_outputs(5918) <= not b;
    layer1_outputs(5919) <= b;
    layer1_outputs(5920) <= a and not b;
    layer1_outputs(5921) <= not b;
    layer1_outputs(5922) <= not b;
    layer1_outputs(5923) <= not a or b;
    layer1_outputs(5924) <= b;
    layer1_outputs(5925) <= a;
    layer1_outputs(5926) <= not b;
    layer1_outputs(5927) <= a and b;
    layer1_outputs(5928) <= '0';
    layer1_outputs(5929) <= a or b;
    layer1_outputs(5930) <= a and b;
    layer1_outputs(5931) <= a xor b;
    layer1_outputs(5932) <= not (a or b);
    layer1_outputs(5933) <= a and b;
    layer1_outputs(5934) <= a and b;
    layer1_outputs(5935) <= a or b;
    layer1_outputs(5936) <= not b;
    layer1_outputs(5937) <= not b or a;
    layer1_outputs(5938) <= not (a or b);
    layer1_outputs(5939) <= not (a and b);
    layer1_outputs(5940) <= not b or a;
    layer1_outputs(5941) <= b and not a;
    layer1_outputs(5942) <= b;
    layer1_outputs(5943) <= a xor b;
    layer1_outputs(5944) <= not (a or b);
    layer1_outputs(5945) <= not a;
    layer1_outputs(5946) <= a;
    layer1_outputs(5947) <= not b;
    layer1_outputs(5948) <= a and b;
    layer1_outputs(5949) <= a xor b;
    layer1_outputs(5950) <= not b;
    layer1_outputs(5951) <= not (a and b);
    layer1_outputs(5952) <= a;
    layer1_outputs(5953) <= a and not b;
    layer1_outputs(5954) <= not b;
    layer1_outputs(5955) <= not a;
    layer1_outputs(5956) <= not a;
    layer1_outputs(5957) <= not b;
    layer1_outputs(5958) <= '1';
    layer1_outputs(5959) <= b;
    layer1_outputs(5960) <= not a;
    layer1_outputs(5961) <= '1';
    layer1_outputs(5962) <= a;
    layer1_outputs(5963) <= not b;
    layer1_outputs(5964) <= b and not a;
    layer1_outputs(5965) <= a;
    layer1_outputs(5966) <= not (a and b);
    layer1_outputs(5967) <= not (a xor b);
    layer1_outputs(5968) <= not b or a;
    layer1_outputs(5969) <= b;
    layer1_outputs(5970) <= a or b;
    layer1_outputs(5971) <= '0';
    layer1_outputs(5972) <= not (a and b);
    layer1_outputs(5973) <= a xor b;
    layer1_outputs(5974) <= b and not a;
    layer1_outputs(5975) <= not b;
    layer1_outputs(5976) <= a xor b;
    layer1_outputs(5977) <= not (a and b);
    layer1_outputs(5978) <= not a;
    layer1_outputs(5979) <= b;
    layer1_outputs(5980) <= not (a or b);
    layer1_outputs(5981) <= '1';
    layer1_outputs(5982) <= a and b;
    layer1_outputs(5983) <= not b or a;
    layer1_outputs(5984) <= not a or b;
    layer1_outputs(5985) <= not b or a;
    layer1_outputs(5986) <= not (a and b);
    layer1_outputs(5987) <= not (a and b);
    layer1_outputs(5988) <= b and not a;
    layer1_outputs(5989) <= a and b;
    layer1_outputs(5990) <= not (a xor b);
    layer1_outputs(5991) <= not (a or b);
    layer1_outputs(5992) <= not a;
    layer1_outputs(5993) <= '1';
    layer1_outputs(5994) <= b and not a;
    layer1_outputs(5995) <= not a or b;
    layer1_outputs(5996) <= a xor b;
    layer1_outputs(5997) <= '1';
    layer1_outputs(5998) <= a and not b;
    layer1_outputs(5999) <= a;
    layer1_outputs(6000) <= a;
    layer1_outputs(6001) <= not a;
    layer1_outputs(6002) <= not b or a;
    layer1_outputs(6003) <= b;
    layer1_outputs(6004) <= not (a and b);
    layer1_outputs(6005) <= '1';
    layer1_outputs(6006) <= b and not a;
    layer1_outputs(6007) <= not a or b;
    layer1_outputs(6008) <= not a;
    layer1_outputs(6009) <= b;
    layer1_outputs(6010) <= not b;
    layer1_outputs(6011) <= b;
    layer1_outputs(6012) <= not (a and b);
    layer1_outputs(6013) <= not a or b;
    layer1_outputs(6014) <= a or b;
    layer1_outputs(6015) <= a or b;
    layer1_outputs(6016) <= not a or b;
    layer1_outputs(6017) <= '0';
    layer1_outputs(6018) <= a and b;
    layer1_outputs(6019) <= not (a or b);
    layer1_outputs(6020) <= a;
    layer1_outputs(6021) <= a;
    layer1_outputs(6022) <= b and not a;
    layer1_outputs(6023) <= b and not a;
    layer1_outputs(6024) <= a and b;
    layer1_outputs(6025) <= a and not b;
    layer1_outputs(6026) <= '1';
    layer1_outputs(6027) <= b;
    layer1_outputs(6028) <= b;
    layer1_outputs(6029) <= not (a or b);
    layer1_outputs(6030) <= not a or b;
    layer1_outputs(6031) <= '0';
    layer1_outputs(6032) <= a;
    layer1_outputs(6033) <= not (a and b);
    layer1_outputs(6034) <= a or b;
    layer1_outputs(6035) <= not (a or b);
    layer1_outputs(6036) <= a and b;
    layer1_outputs(6037) <= b;
    layer1_outputs(6038) <= a and b;
    layer1_outputs(6039) <= '1';
    layer1_outputs(6040) <= a;
    layer1_outputs(6041) <= a xor b;
    layer1_outputs(6042) <= not (a or b);
    layer1_outputs(6043) <= a or b;
    layer1_outputs(6044) <= not (a or b);
    layer1_outputs(6045) <= not a;
    layer1_outputs(6046) <= not b or a;
    layer1_outputs(6047) <= '1';
    layer1_outputs(6048) <= a and not b;
    layer1_outputs(6049) <= not b or a;
    layer1_outputs(6050) <= a and not b;
    layer1_outputs(6051) <= a and not b;
    layer1_outputs(6052) <= not (a xor b);
    layer1_outputs(6053) <= not b;
    layer1_outputs(6054) <= b;
    layer1_outputs(6055) <= not b or a;
    layer1_outputs(6056) <= b;
    layer1_outputs(6057) <= a xor b;
    layer1_outputs(6058) <= b;
    layer1_outputs(6059) <= b;
    layer1_outputs(6060) <= not a;
    layer1_outputs(6061) <= a and not b;
    layer1_outputs(6062) <= not b or a;
    layer1_outputs(6063) <= not b or a;
    layer1_outputs(6064) <= not (a and b);
    layer1_outputs(6065) <= a and not b;
    layer1_outputs(6066) <= b and not a;
    layer1_outputs(6067) <= a and not b;
    layer1_outputs(6068) <= a and b;
    layer1_outputs(6069) <= a or b;
    layer1_outputs(6070) <= not b or a;
    layer1_outputs(6071) <= a and not b;
    layer1_outputs(6072) <= not a;
    layer1_outputs(6073) <= '1';
    layer1_outputs(6074) <= not (a or b);
    layer1_outputs(6075) <= not a;
    layer1_outputs(6076) <= not b or a;
    layer1_outputs(6077) <= '1';
    layer1_outputs(6078) <= not b or a;
    layer1_outputs(6079) <= a;
    layer1_outputs(6080) <= '0';
    layer1_outputs(6081) <= '0';
    layer1_outputs(6082) <= a xor b;
    layer1_outputs(6083) <= not (a and b);
    layer1_outputs(6084) <= not a;
    layer1_outputs(6085) <= not (a or b);
    layer1_outputs(6086) <= not a or b;
    layer1_outputs(6087) <= a and not b;
    layer1_outputs(6088) <= not (a or b);
    layer1_outputs(6089) <= a and not b;
    layer1_outputs(6090) <= b;
    layer1_outputs(6091) <= not a or b;
    layer1_outputs(6092) <= not a;
    layer1_outputs(6093) <= not b;
    layer1_outputs(6094) <= not (a xor b);
    layer1_outputs(6095) <= not (a or b);
    layer1_outputs(6096) <= not b or a;
    layer1_outputs(6097) <= b;
    layer1_outputs(6098) <= b and not a;
    layer1_outputs(6099) <= a;
    layer1_outputs(6100) <= not a or b;
    layer1_outputs(6101) <= a or b;
    layer1_outputs(6102) <= not a;
    layer1_outputs(6103) <= b;
    layer1_outputs(6104) <= not b;
    layer1_outputs(6105) <= a or b;
    layer1_outputs(6106) <= not b;
    layer1_outputs(6107) <= not (a or b);
    layer1_outputs(6108) <= not a;
    layer1_outputs(6109) <= not a;
    layer1_outputs(6110) <= b;
    layer1_outputs(6111) <= '0';
    layer1_outputs(6112) <= a;
    layer1_outputs(6113) <= not b;
    layer1_outputs(6114) <= not (a or b);
    layer1_outputs(6115) <= a;
    layer1_outputs(6116) <= b;
    layer1_outputs(6117) <= not b;
    layer1_outputs(6118) <= b;
    layer1_outputs(6119) <= not (a or b);
    layer1_outputs(6120) <= not a;
    layer1_outputs(6121) <= a and b;
    layer1_outputs(6122) <= not (a and b);
    layer1_outputs(6123) <= not b or a;
    layer1_outputs(6124) <= a and b;
    layer1_outputs(6125) <= not b;
    layer1_outputs(6126) <= '1';
    layer1_outputs(6127) <= not (a or b);
    layer1_outputs(6128) <= not (a or b);
    layer1_outputs(6129) <= '1';
    layer1_outputs(6130) <= not (a or b);
    layer1_outputs(6131) <= not b or a;
    layer1_outputs(6132) <= b;
    layer1_outputs(6133) <= a and not b;
    layer1_outputs(6134) <= not b;
    layer1_outputs(6135) <= a xor b;
    layer1_outputs(6136) <= a and b;
    layer1_outputs(6137) <= a and b;
    layer1_outputs(6138) <= not a;
    layer1_outputs(6139) <= '0';
    layer1_outputs(6140) <= not (a or b);
    layer1_outputs(6141) <= a;
    layer1_outputs(6142) <= a;
    layer1_outputs(6143) <= a or b;
    layer1_outputs(6144) <= b and not a;
    layer1_outputs(6145) <= a xor b;
    layer1_outputs(6146) <= a;
    layer1_outputs(6147) <= not b;
    layer1_outputs(6148) <= not a;
    layer1_outputs(6149) <= a and b;
    layer1_outputs(6150) <= not b or a;
    layer1_outputs(6151) <= b;
    layer1_outputs(6152) <= a or b;
    layer1_outputs(6153) <= a;
    layer1_outputs(6154) <= a xor b;
    layer1_outputs(6155) <= a and not b;
    layer1_outputs(6156) <= b and not a;
    layer1_outputs(6157) <= b;
    layer1_outputs(6158) <= not b;
    layer1_outputs(6159) <= not b;
    layer1_outputs(6160) <= not a;
    layer1_outputs(6161) <= not b or a;
    layer1_outputs(6162) <= not a;
    layer1_outputs(6163) <= a and b;
    layer1_outputs(6164) <= not b;
    layer1_outputs(6165) <= not b or a;
    layer1_outputs(6166) <= b;
    layer1_outputs(6167) <= not a;
    layer1_outputs(6168) <= not (a or b);
    layer1_outputs(6169) <= a and b;
    layer1_outputs(6170) <= a;
    layer1_outputs(6171) <= not a;
    layer1_outputs(6172) <= a and not b;
    layer1_outputs(6173) <= b and not a;
    layer1_outputs(6174) <= not a;
    layer1_outputs(6175) <= b;
    layer1_outputs(6176) <= not b;
    layer1_outputs(6177) <= '0';
    layer1_outputs(6178) <= a and not b;
    layer1_outputs(6179) <= not b;
    layer1_outputs(6180) <= not b or a;
    layer1_outputs(6181) <= not b;
    layer1_outputs(6182) <= not b;
    layer1_outputs(6183) <= not b or a;
    layer1_outputs(6184) <= not (a or b);
    layer1_outputs(6185) <= not b or a;
    layer1_outputs(6186) <= not a;
    layer1_outputs(6187) <= a or b;
    layer1_outputs(6188) <= a and b;
    layer1_outputs(6189) <= a and b;
    layer1_outputs(6190) <= a;
    layer1_outputs(6191) <= not b;
    layer1_outputs(6192) <= a and not b;
    layer1_outputs(6193) <= b and not a;
    layer1_outputs(6194) <= not a;
    layer1_outputs(6195) <= not (a and b);
    layer1_outputs(6196) <= a;
    layer1_outputs(6197) <= not b or a;
    layer1_outputs(6198) <= '1';
    layer1_outputs(6199) <= not b;
    layer1_outputs(6200) <= a xor b;
    layer1_outputs(6201) <= a or b;
    layer1_outputs(6202) <= not a;
    layer1_outputs(6203) <= '0';
    layer1_outputs(6204) <= b;
    layer1_outputs(6205) <= a and not b;
    layer1_outputs(6206) <= b and not a;
    layer1_outputs(6207) <= a and b;
    layer1_outputs(6208) <= not (a or b);
    layer1_outputs(6209) <= not a or b;
    layer1_outputs(6210) <= not a;
    layer1_outputs(6211) <= b and not a;
    layer1_outputs(6212) <= not b or a;
    layer1_outputs(6213) <= a and not b;
    layer1_outputs(6214) <= not b or a;
    layer1_outputs(6215) <= b and not a;
    layer1_outputs(6216) <= not (a xor b);
    layer1_outputs(6217) <= not a;
    layer1_outputs(6218) <= b and not a;
    layer1_outputs(6219) <= a and not b;
    layer1_outputs(6220) <= a and not b;
    layer1_outputs(6221) <= not a;
    layer1_outputs(6222) <= a;
    layer1_outputs(6223) <= '0';
    layer1_outputs(6224) <= not b;
    layer1_outputs(6225) <= a and b;
    layer1_outputs(6226) <= a and b;
    layer1_outputs(6227) <= b;
    layer1_outputs(6228) <= '1';
    layer1_outputs(6229) <= a and not b;
    layer1_outputs(6230) <= not a;
    layer1_outputs(6231) <= not a;
    layer1_outputs(6232) <= b;
    layer1_outputs(6233) <= a or b;
    layer1_outputs(6234) <= not (a and b);
    layer1_outputs(6235) <= a and b;
    layer1_outputs(6236) <= a and b;
    layer1_outputs(6237) <= not (a or b);
    layer1_outputs(6238) <= '0';
    layer1_outputs(6239) <= a xor b;
    layer1_outputs(6240) <= not (a or b);
    layer1_outputs(6241) <= not a or b;
    layer1_outputs(6242) <= a or b;
    layer1_outputs(6243) <= b;
    layer1_outputs(6244) <= '0';
    layer1_outputs(6245) <= a and not b;
    layer1_outputs(6246) <= b and not a;
    layer1_outputs(6247) <= not a;
    layer1_outputs(6248) <= not b;
    layer1_outputs(6249) <= not (a and b);
    layer1_outputs(6250) <= not a or b;
    layer1_outputs(6251) <= a xor b;
    layer1_outputs(6252) <= not a or b;
    layer1_outputs(6253) <= a or b;
    layer1_outputs(6254) <= a and b;
    layer1_outputs(6255) <= not (a and b);
    layer1_outputs(6256) <= not a;
    layer1_outputs(6257) <= b;
    layer1_outputs(6258) <= '0';
    layer1_outputs(6259) <= '0';
    layer1_outputs(6260) <= not (a and b);
    layer1_outputs(6261) <= not a or b;
    layer1_outputs(6262) <= a or b;
    layer1_outputs(6263) <= not b or a;
    layer1_outputs(6264) <= a and b;
    layer1_outputs(6265) <= not b;
    layer1_outputs(6266) <= not a;
    layer1_outputs(6267) <= a or b;
    layer1_outputs(6268) <= not a or b;
    layer1_outputs(6269) <= not a;
    layer1_outputs(6270) <= '0';
    layer1_outputs(6271) <= '0';
    layer1_outputs(6272) <= not b or a;
    layer1_outputs(6273) <= a;
    layer1_outputs(6274) <= '1';
    layer1_outputs(6275) <= not (a or b);
    layer1_outputs(6276) <= a and not b;
    layer1_outputs(6277) <= a or b;
    layer1_outputs(6278) <= not (a xor b);
    layer1_outputs(6279) <= not (a or b);
    layer1_outputs(6280) <= not (a and b);
    layer1_outputs(6281) <= '0';
    layer1_outputs(6282) <= '1';
    layer1_outputs(6283) <= not a;
    layer1_outputs(6284) <= not b or a;
    layer1_outputs(6285) <= a or b;
    layer1_outputs(6286) <= a and not b;
    layer1_outputs(6287) <= not b;
    layer1_outputs(6288) <= not (a and b);
    layer1_outputs(6289) <= not a or b;
    layer1_outputs(6290) <= not (a or b);
    layer1_outputs(6291) <= a or b;
    layer1_outputs(6292) <= a or b;
    layer1_outputs(6293) <= not b or a;
    layer1_outputs(6294) <= a or b;
    layer1_outputs(6295) <= not b;
    layer1_outputs(6296) <= '0';
    layer1_outputs(6297) <= b;
    layer1_outputs(6298) <= a and b;
    layer1_outputs(6299) <= a and b;
    layer1_outputs(6300) <= not a;
    layer1_outputs(6301) <= not a;
    layer1_outputs(6302) <= not a;
    layer1_outputs(6303) <= not (a or b);
    layer1_outputs(6304) <= a;
    layer1_outputs(6305) <= not b;
    layer1_outputs(6306) <= a or b;
    layer1_outputs(6307) <= a and b;
    layer1_outputs(6308) <= not a or b;
    layer1_outputs(6309) <= not b or a;
    layer1_outputs(6310) <= b and not a;
    layer1_outputs(6311) <= not (a and b);
    layer1_outputs(6312) <= b and not a;
    layer1_outputs(6313) <= a;
    layer1_outputs(6314) <= not (a or b);
    layer1_outputs(6315) <= b and not a;
    layer1_outputs(6316) <= a and b;
    layer1_outputs(6317) <= not a;
    layer1_outputs(6318) <= '0';
    layer1_outputs(6319) <= b;
    layer1_outputs(6320) <= a or b;
    layer1_outputs(6321) <= '0';
    layer1_outputs(6322) <= a and b;
    layer1_outputs(6323) <= not a or b;
    layer1_outputs(6324) <= not (a and b);
    layer1_outputs(6325) <= not (a and b);
    layer1_outputs(6326) <= a;
    layer1_outputs(6327) <= b and not a;
    layer1_outputs(6328) <= a and not b;
    layer1_outputs(6329) <= not a;
    layer1_outputs(6330) <= not b;
    layer1_outputs(6331) <= '0';
    layer1_outputs(6332) <= not b or a;
    layer1_outputs(6333) <= a xor b;
    layer1_outputs(6334) <= a;
    layer1_outputs(6335) <= a and not b;
    layer1_outputs(6336) <= b;
    layer1_outputs(6337) <= not (a and b);
    layer1_outputs(6338) <= not b;
    layer1_outputs(6339) <= not (a or b);
    layer1_outputs(6340) <= a and not b;
    layer1_outputs(6341) <= a and not b;
    layer1_outputs(6342) <= not a or b;
    layer1_outputs(6343) <= b and not a;
    layer1_outputs(6344) <= '0';
    layer1_outputs(6345) <= a and not b;
    layer1_outputs(6346) <= not (a xor b);
    layer1_outputs(6347) <= a and not b;
    layer1_outputs(6348) <= '0';
    layer1_outputs(6349) <= a;
    layer1_outputs(6350) <= not (a or b);
    layer1_outputs(6351) <= b and not a;
    layer1_outputs(6352) <= b;
    layer1_outputs(6353) <= a or b;
    layer1_outputs(6354) <= not (a xor b);
    layer1_outputs(6355) <= a and b;
    layer1_outputs(6356) <= not a;
    layer1_outputs(6357) <= a and not b;
    layer1_outputs(6358) <= '1';
    layer1_outputs(6359) <= '0';
    layer1_outputs(6360) <= a;
    layer1_outputs(6361) <= a;
    layer1_outputs(6362) <= a or b;
    layer1_outputs(6363) <= a and b;
    layer1_outputs(6364) <= a and b;
    layer1_outputs(6365) <= a and b;
    layer1_outputs(6366) <= not b or a;
    layer1_outputs(6367) <= a and b;
    layer1_outputs(6368) <= not a;
    layer1_outputs(6369) <= not a or b;
    layer1_outputs(6370) <= b and not a;
    layer1_outputs(6371) <= not (a and b);
    layer1_outputs(6372) <= not (a and b);
    layer1_outputs(6373) <= a xor b;
    layer1_outputs(6374) <= not b;
    layer1_outputs(6375) <= '1';
    layer1_outputs(6376) <= b;
    layer1_outputs(6377) <= not (a or b);
    layer1_outputs(6378) <= not b;
    layer1_outputs(6379) <= not b;
    layer1_outputs(6380) <= a or b;
    layer1_outputs(6381) <= b;
    layer1_outputs(6382) <= '1';
    layer1_outputs(6383) <= a;
    layer1_outputs(6384) <= '0';
    layer1_outputs(6385) <= a;
    layer1_outputs(6386) <= a;
    layer1_outputs(6387) <= not b;
    layer1_outputs(6388) <= not b or a;
    layer1_outputs(6389) <= a or b;
    layer1_outputs(6390) <= not b or a;
    layer1_outputs(6391) <= '0';
    layer1_outputs(6392) <= b and not a;
    layer1_outputs(6393) <= '1';
    layer1_outputs(6394) <= not a or b;
    layer1_outputs(6395) <= not (a or b);
    layer1_outputs(6396) <= a or b;
    layer1_outputs(6397) <= not b or a;
    layer1_outputs(6398) <= '1';
    layer1_outputs(6399) <= not a;
    layer1_outputs(6400) <= b;
    layer1_outputs(6401) <= '0';
    layer1_outputs(6402) <= not a;
    layer1_outputs(6403) <= a xor b;
    layer1_outputs(6404) <= b and not a;
    layer1_outputs(6405) <= '1';
    layer1_outputs(6406) <= not b;
    layer1_outputs(6407) <= '1';
    layer1_outputs(6408) <= a or b;
    layer1_outputs(6409) <= a;
    layer1_outputs(6410) <= a;
    layer1_outputs(6411) <= not (a and b);
    layer1_outputs(6412) <= not (a or b);
    layer1_outputs(6413) <= a and b;
    layer1_outputs(6414) <= b;
    layer1_outputs(6415) <= not (a or b);
    layer1_outputs(6416) <= not (a and b);
    layer1_outputs(6417) <= not a;
    layer1_outputs(6418) <= not (a xor b);
    layer1_outputs(6419) <= a and b;
    layer1_outputs(6420) <= not a;
    layer1_outputs(6421) <= b and not a;
    layer1_outputs(6422) <= '0';
    layer1_outputs(6423) <= '0';
    layer1_outputs(6424) <= not a or b;
    layer1_outputs(6425) <= a or b;
    layer1_outputs(6426) <= not b;
    layer1_outputs(6427) <= a and b;
    layer1_outputs(6428) <= not b;
    layer1_outputs(6429) <= not (a or b);
    layer1_outputs(6430) <= not (a and b);
    layer1_outputs(6431) <= a;
    layer1_outputs(6432) <= a and not b;
    layer1_outputs(6433) <= not b;
    layer1_outputs(6434) <= '0';
    layer1_outputs(6435) <= b;
    layer1_outputs(6436) <= b;
    layer1_outputs(6437) <= not (a or b);
    layer1_outputs(6438) <= not (a or b);
    layer1_outputs(6439) <= not b or a;
    layer1_outputs(6440) <= b and not a;
    layer1_outputs(6441) <= a;
    layer1_outputs(6442) <= '1';
    layer1_outputs(6443) <= not (a and b);
    layer1_outputs(6444) <= not b or a;
    layer1_outputs(6445) <= a or b;
    layer1_outputs(6446) <= '0';
    layer1_outputs(6447) <= not b or a;
    layer1_outputs(6448) <= not (a or b);
    layer1_outputs(6449) <= not (a or b);
    layer1_outputs(6450) <= not b;
    layer1_outputs(6451) <= not a;
    layer1_outputs(6452) <= not (a xor b);
    layer1_outputs(6453) <= not (a and b);
    layer1_outputs(6454) <= not b or a;
    layer1_outputs(6455) <= '1';
    layer1_outputs(6456) <= '0';
    layer1_outputs(6457) <= a and b;
    layer1_outputs(6458) <= not (a xor b);
    layer1_outputs(6459) <= not b;
    layer1_outputs(6460) <= a and b;
    layer1_outputs(6461) <= b and not a;
    layer1_outputs(6462) <= not b or a;
    layer1_outputs(6463) <= a and b;
    layer1_outputs(6464) <= '1';
    layer1_outputs(6465) <= '0';
    layer1_outputs(6466) <= b;
    layer1_outputs(6467) <= not b;
    layer1_outputs(6468) <= not (a and b);
    layer1_outputs(6469) <= a xor b;
    layer1_outputs(6470) <= not (a and b);
    layer1_outputs(6471) <= b;
    layer1_outputs(6472) <= not a;
    layer1_outputs(6473) <= '0';
    layer1_outputs(6474) <= '0';
    layer1_outputs(6475) <= not a;
    layer1_outputs(6476) <= b and not a;
    layer1_outputs(6477) <= a or b;
    layer1_outputs(6478) <= a or b;
    layer1_outputs(6479) <= not a;
    layer1_outputs(6480) <= not (a xor b);
    layer1_outputs(6481) <= a and not b;
    layer1_outputs(6482) <= b;
    layer1_outputs(6483) <= not (a and b);
    layer1_outputs(6484) <= b and not a;
    layer1_outputs(6485) <= not (a or b);
    layer1_outputs(6486) <= a or b;
    layer1_outputs(6487) <= a;
    layer1_outputs(6488) <= not b;
    layer1_outputs(6489) <= a xor b;
    layer1_outputs(6490) <= a and not b;
    layer1_outputs(6491) <= a and not b;
    layer1_outputs(6492) <= a and not b;
    layer1_outputs(6493) <= not b or a;
    layer1_outputs(6494) <= b;
    layer1_outputs(6495) <= a and not b;
    layer1_outputs(6496) <= a xor b;
    layer1_outputs(6497) <= not a;
    layer1_outputs(6498) <= not a;
    layer1_outputs(6499) <= a and not b;
    layer1_outputs(6500) <= '1';
    layer1_outputs(6501) <= a and not b;
    layer1_outputs(6502) <= b;
    layer1_outputs(6503) <= not (a or b);
    layer1_outputs(6504) <= '0';
    layer1_outputs(6505) <= a;
    layer1_outputs(6506) <= not a;
    layer1_outputs(6507) <= not (a xor b);
    layer1_outputs(6508) <= not a or b;
    layer1_outputs(6509) <= b;
    layer1_outputs(6510) <= a and not b;
    layer1_outputs(6511) <= not (a or b);
    layer1_outputs(6512) <= '0';
    layer1_outputs(6513) <= not (a xor b);
    layer1_outputs(6514) <= a;
    layer1_outputs(6515) <= a or b;
    layer1_outputs(6516) <= a or b;
    layer1_outputs(6517) <= not (a xor b);
    layer1_outputs(6518) <= not a or b;
    layer1_outputs(6519) <= not a;
    layer1_outputs(6520) <= a and not b;
    layer1_outputs(6521) <= not a or b;
    layer1_outputs(6522) <= not b;
    layer1_outputs(6523) <= a xor b;
    layer1_outputs(6524) <= a or b;
    layer1_outputs(6525) <= a and not b;
    layer1_outputs(6526) <= a;
    layer1_outputs(6527) <= not a or b;
    layer1_outputs(6528) <= b;
    layer1_outputs(6529) <= not b or a;
    layer1_outputs(6530) <= a or b;
    layer1_outputs(6531) <= '0';
    layer1_outputs(6532) <= b;
    layer1_outputs(6533) <= a;
    layer1_outputs(6534) <= '1';
    layer1_outputs(6535) <= a and b;
    layer1_outputs(6536) <= '0';
    layer1_outputs(6537) <= a and not b;
    layer1_outputs(6538) <= not (a xor b);
    layer1_outputs(6539) <= a;
    layer1_outputs(6540) <= a or b;
    layer1_outputs(6541) <= b;
    layer1_outputs(6542) <= not a;
    layer1_outputs(6543) <= a and b;
    layer1_outputs(6544) <= a;
    layer1_outputs(6545) <= not (a or b);
    layer1_outputs(6546) <= b;
    layer1_outputs(6547) <= b and not a;
    layer1_outputs(6548) <= a;
    layer1_outputs(6549) <= a and not b;
    layer1_outputs(6550) <= not b or a;
    layer1_outputs(6551) <= not b or a;
    layer1_outputs(6552) <= not (a and b);
    layer1_outputs(6553) <= not b;
    layer1_outputs(6554) <= not (a and b);
    layer1_outputs(6555) <= not a or b;
    layer1_outputs(6556) <= '1';
    layer1_outputs(6557) <= '0';
    layer1_outputs(6558) <= not a or b;
    layer1_outputs(6559) <= b;
    layer1_outputs(6560) <= not b or a;
    layer1_outputs(6561) <= '1';
    layer1_outputs(6562) <= a;
    layer1_outputs(6563) <= a;
    layer1_outputs(6564) <= '1';
    layer1_outputs(6565) <= not b or a;
    layer1_outputs(6566) <= a or b;
    layer1_outputs(6567) <= a and b;
    layer1_outputs(6568) <= b and not a;
    layer1_outputs(6569) <= a xor b;
    layer1_outputs(6570) <= not a;
    layer1_outputs(6571) <= a and not b;
    layer1_outputs(6572) <= not b or a;
    layer1_outputs(6573) <= not a or b;
    layer1_outputs(6574) <= b;
    layer1_outputs(6575) <= not (a and b);
    layer1_outputs(6576) <= not a;
    layer1_outputs(6577) <= '0';
    layer1_outputs(6578) <= a and b;
    layer1_outputs(6579) <= not (a and b);
    layer1_outputs(6580) <= a and not b;
    layer1_outputs(6581) <= b and not a;
    layer1_outputs(6582) <= not (a xor b);
    layer1_outputs(6583) <= a and b;
    layer1_outputs(6584) <= not (a and b);
    layer1_outputs(6585) <= '1';
    layer1_outputs(6586) <= b and not a;
    layer1_outputs(6587) <= not (a and b);
    layer1_outputs(6588) <= not (a and b);
    layer1_outputs(6589) <= a and not b;
    layer1_outputs(6590) <= a and not b;
    layer1_outputs(6591) <= a or b;
    layer1_outputs(6592) <= '0';
    layer1_outputs(6593) <= '1';
    layer1_outputs(6594) <= not (a and b);
    layer1_outputs(6595) <= not a;
    layer1_outputs(6596) <= not (a and b);
    layer1_outputs(6597) <= not b;
    layer1_outputs(6598) <= not (a or b);
    layer1_outputs(6599) <= b and not a;
    layer1_outputs(6600) <= a and not b;
    layer1_outputs(6601) <= a;
    layer1_outputs(6602) <= not a or b;
    layer1_outputs(6603) <= not (a and b);
    layer1_outputs(6604) <= b;
    layer1_outputs(6605) <= a and not b;
    layer1_outputs(6606) <= b;
    layer1_outputs(6607) <= '1';
    layer1_outputs(6608) <= not b;
    layer1_outputs(6609) <= a and b;
    layer1_outputs(6610) <= not b;
    layer1_outputs(6611) <= not (a or b);
    layer1_outputs(6612) <= a xor b;
    layer1_outputs(6613) <= '0';
    layer1_outputs(6614) <= not a;
    layer1_outputs(6615) <= not (a xor b);
    layer1_outputs(6616) <= a;
    layer1_outputs(6617) <= not (a and b);
    layer1_outputs(6618) <= not (a or b);
    layer1_outputs(6619) <= not b;
    layer1_outputs(6620) <= '1';
    layer1_outputs(6621) <= b;
    layer1_outputs(6622) <= not a or b;
    layer1_outputs(6623) <= a or b;
    layer1_outputs(6624) <= not (a xor b);
    layer1_outputs(6625) <= a or b;
    layer1_outputs(6626) <= not a;
    layer1_outputs(6627) <= not b or a;
    layer1_outputs(6628) <= a and not b;
    layer1_outputs(6629) <= not a;
    layer1_outputs(6630) <= not a or b;
    layer1_outputs(6631) <= not (a and b);
    layer1_outputs(6632) <= not (a xor b);
    layer1_outputs(6633) <= a and b;
    layer1_outputs(6634) <= a xor b;
    layer1_outputs(6635) <= a or b;
    layer1_outputs(6636) <= not b or a;
    layer1_outputs(6637) <= a or b;
    layer1_outputs(6638) <= b;
    layer1_outputs(6639) <= not (a and b);
    layer1_outputs(6640) <= '1';
    layer1_outputs(6641) <= not b or a;
    layer1_outputs(6642) <= a or b;
    layer1_outputs(6643) <= a and not b;
    layer1_outputs(6644) <= '0';
    layer1_outputs(6645) <= a;
    layer1_outputs(6646) <= not (a and b);
    layer1_outputs(6647) <= '1';
    layer1_outputs(6648) <= '1';
    layer1_outputs(6649) <= not b or a;
    layer1_outputs(6650) <= not b or a;
    layer1_outputs(6651) <= not a;
    layer1_outputs(6652) <= '0';
    layer1_outputs(6653) <= not (a or b);
    layer1_outputs(6654) <= a and b;
    layer1_outputs(6655) <= not a;
    layer1_outputs(6656) <= b;
    layer1_outputs(6657) <= not a or b;
    layer1_outputs(6658) <= b and not a;
    layer1_outputs(6659) <= not b;
    layer1_outputs(6660) <= '1';
    layer1_outputs(6661) <= '1';
    layer1_outputs(6662) <= not a or b;
    layer1_outputs(6663) <= b and not a;
    layer1_outputs(6664) <= '0';
    layer1_outputs(6665) <= a xor b;
    layer1_outputs(6666) <= not a or b;
    layer1_outputs(6667) <= not b;
    layer1_outputs(6668) <= b;
    layer1_outputs(6669) <= b;
    layer1_outputs(6670) <= b;
    layer1_outputs(6671) <= a;
    layer1_outputs(6672) <= a and not b;
    layer1_outputs(6673) <= b;
    layer1_outputs(6674) <= a and not b;
    layer1_outputs(6675) <= not b;
    layer1_outputs(6676) <= not (a xor b);
    layer1_outputs(6677) <= a or b;
    layer1_outputs(6678) <= b;
    layer1_outputs(6679) <= not (a and b);
    layer1_outputs(6680) <= a or b;
    layer1_outputs(6681) <= not (a and b);
    layer1_outputs(6682) <= '0';
    layer1_outputs(6683) <= not b;
    layer1_outputs(6684) <= a xor b;
    layer1_outputs(6685) <= b;
    layer1_outputs(6686) <= not b or a;
    layer1_outputs(6687) <= not a or b;
    layer1_outputs(6688) <= b;
    layer1_outputs(6689) <= not (a or b);
    layer1_outputs(6690) <= '1';
    layer1_outputs(6691) <= not b or a;
    layer1_outputs(6692) <= not (a and b);
    layer1_outputs(6693) <= a xor b;
    layer1_outputs(6694) <= not b or a;
    layer1_outputs(6695) <= not a;
    layer1_outputs(6696) <= a xor b;
    layer1_outputs(6697) <= a or b;
    layer1_outputs(6698) <= not b;
    layer1_outputs(6699) <= a;
    layer1_outputs(6700) <= a xor b;
    layer1_outputs(6701) <= not (a xor b);
    layer1_outputs(6702) <= not (a xor b);
    layer1_outputs(6703) <= a;
    layer1_outputs(6704) <= a;
    layer1_outputs(6705) <= a and b;
    layer1_outputs(6706) <= not (a and b);
    layer1_outputs(6707) <= a and not b;
    layer1_outputs(6708) <= a or b;
    layer1_outputs(6709) <= not a;
    layer1_outputs(6710) <= not a;
    layer1_outputs(6711) <= a and not b;
    layer1_outputs(6712) <= not a or b;
    layer1_outputs(6713) <= b;
    layer1_outputs(6714) <= a;
    layer1_outputs(6715) <= a or b;
    layer1_outputs(6716) <= not a;
    layer1_outputs(6717) <= not b;
    layer1_outputs(6718) <= '1';
    layer1_outputs(6719) <= b and not a;
    layer1_outputs(6720) <= a;
    layer1_outputs(6721) <= a or b;
    layer1_outputs(6722) <= not b;
    layer1_outputs(6723) <= not b;
    layer1_outputs(6724) <= not (a or b);
    layer1_outputs(6725) <= not b;
    layer1_outputs(6726) <= '0';
    layer1_outputs(6727) <= b and not a;
    layer1_outputs(6728) <= not a;
    layer1_outputs(6729) <= not a;
    layer1_outputs(6730) <= not (a xor b);
    layer1_outputs(6731) <= not (a and b);
    layer1_outputs(6732) <= not (a or b);
    layer1_outputs(6733) <= not (a and b);
    layer1_outputs(6734) <= not a;
    layer1_outputs(6735) <= b and not a;
    layer1_outputs(6736) <= not b;
    layer1_outputs(6737) <= '1';
    layer1_outputs(6738) <= a;
    layer1_outputs(6739) <= not b;
    layer1_outputs(6740) <= not b;
    layer1_outputs(6741) <= not b;
    layer1_outputs(6742) <= not a;
    layer1_outputs(6743) <= not b or a;
    layer1_outputs(6744) <= not a;
    layer1_outputs(6745) <= '0';
    layer1_outputs(6746) <= a and b;
    layer1_outputs(6747) <= b and not a;
    layer1_outputs(6748) <= b;
    layer1_outputs(6749) <= not a;
    layer1_outputs(6750) <= not a;
    layer1_outputs(6751) <= b;
    layer1_outputs(6752) <= not a or b;
    layer1_outputs(6753) <= '1';
    layer1_outputs(6754) <= not a or b;
    layer1_outputs(6755) <= not b or a;
    layer1_outputs(6756) <= '1';
    layer1_outputs(6757) <= '0';
    layer1_outputs(6758) <= not b;
    layer1_outputs(6759) <= '1';
    layer1_outputs(6760) <= not b or a;
    layer1_outputs(6761) <= not (a and b);
    layer1_outputs(6762) <= '1';
    layer1_outputs(6763) <= not b;
    layer1_outputs(6764) <= '0';
    layer1_outputs(6765) <= a;
    layer1_outputs(6766) <= a;
    layer1_outputs(6767) <= not b or a;
    layer1_outputs(6768) <= a and not b;
    layer1_outputs(6769) <= not b;
    layer1_outputs(6770) <= not b;
    layer1_outputs(6771) <= '0';
    layer1_outputs(6772) <= '1';
    layer1_outputs(6773) <= a and b;
    layer1_outputs(6774) <= a or b;
    layer1_outputs(6775) <= b and not a;
    layer1_outputs(6776) <= not a;
    layer1_outputs(6777) <= b;
    layer1_outputs(6778) <= a and not b;
    layer1_outputs(6779) <= not (a and b);
    layer1_outputs(6780) <= b;
    layer1_outputs(6781) <= not (a xor b);
    layer1_outputs(6782) <= a and not b;
    layer1_outputs(6783) <= not a;
    layer1_outputs(6784) <= not (a and b);
    layer1_outputs(6785) <= not (a or b);
    layer1_outputs(6786) <= a and b;
    layer1_outputs(6787) <= not a;
    layer1_outputs(6788) <= '1';
    layer1_outputs(6789) <= a and not b;
    layer1_outputs(6790) <= not b;
    layer1_outputs(6791) <= not (a and b);
    layer1_outputs(6792) <= not (a or b);
    layer1_outputs(6793) <= a;
    layer1_outputs(6794) <= not b or a;
    layer1_outputs(6795) <= not (a xor b);
    layer1_outputs(6796) <= a xor b;
    layer1_outputs(6797) <= not b;
    layer1_outputs(6798) <= b;
    layer1_outputs(6799) <= a or b;
    layer1_outputs(6800) <= not b;
    layer1_outputs(6801) <= not (a and b);
    layer1_outputs(6802) <= not b;
    layer1_outputs(6803) <= a xor b;
    layer1_outputs(6804) <= not a;
    layer1_outputs(6805) <= a and b;
    layer1_outputs(6806) <= a or b;
    layer1_outputs(6807) <= not b;
    layer1_outputs(6808) <= not (a and b);
    layer1_outputs(6809) <= b and not a;
    layer1_outputs(6810) <= b;
    layer1_outputs(6811) <= a and b;
    layer1_outputs(6812) <= not a;
    layer1_outputs(6813) <= not (a and b);
    layer1_outputs(6814) <= not b;
    layer1_outputs(6815) <= a xor b;
    layer1_outputs(6816) <= a and not b;
    layer1_outputs(6817) <= a xor b;
    layer1_outputs(6818) <= a or b;
    layer1_outputs(6819) <= not (a and b);
    layer1_outputs(6820) <= a;
    layer1_outputs(6821) <= not a or b;
    layer1_outputs(6822) <= not b;
    layer1_outputs(6823) <= '1';
    layer1_outputs(6824) <= not b or a;
    layer1_outputs(6825) <= not b;
    layer1_outputs(6826) <= b;
    layer1_outputs(6827) <= not a;
    layer1_outputs(6828) <= not a;
    layer1_outputs(6829) <= b;
    layer1_outputs(6830) <= b;
    layer1_outputs(6831) <= b and not a;
    layer1_outputs(6832) <= not a;
    layer1_outputs(6833) <= a;
    layer1_outputs(6834) <= a and b;
    layer1_outputs(6835) <= b;
    layer1_outputs(6836) <= b;
    layer1_outputs(6837) <= b;
    layer1_outputs(6838) <= not b;
    layer1_outputs(6839) <= b and not a;
    layer1_outputs(6840) <= a;
    layer1_outputs(6841) <= not (a and b);
    layer1_outputs(6842) <= b and not a;
    layer1_outputs(6843) <= a or b;
    layer1_outputs(6844) <= not b or a;
    layer1_outputs(6845) <= a xor b;
    layer1_outputs(6846) <= not b;
    layer1_outputs(6847) <= not a;
    layer1_outputs(6848) <= not b;
    layer1_outputs(6849) <= not a or b;
    layer1_outputs(6850) <= not b;
    layer1_outputs(6851) <= a or b;
    layer1_outputs(6852) <= not (a and b);
    layer1_outputs(6853) <= '0';
    layer1_outputs(6854) <= not (a xor b);
    layer1_outputs(6855) <= a;
    layer1_outputs(6856) <= not a;
    layer1_outputs(6857) <= not b;
    layer1_outputs(6858) <= not b or a;
    layer1_outputs(6859) <= not b;
    layer1_outputs(6860) <= a and b;
    layer1_outputs(6861) <= a;
    layer1_outputs(6862) <= not a;
    layer1_outputs(6863) <= '0';
    layer1_outputs(6864) <= not (a xor b);
    layer1_outputs(6865) <= not a;
    layer1_outputs(6866) <= not b or a;
    layer1_outputs(6867) <= not b;
    layer1_outputs(6868) <= a and not b;
    layer1_outputs(6869) <= not (a and b);
    layer1_outputs(6870) <= not a;
    layer1_outputs(6871) <= not (a xor b);
    layer1_outputs(6872) <= not b or a;
    layer1_outputs(6873) <= a and not b;
    layer1_outputs(6874) <= not (a xor b);
    layer1_outputs(6875) <= a and not b;
    layer1_outputs(6876) <= not a;
    layer1_outputs(6877) <= not (a and b);
    layer1_outputs(6878) <= b;
    layer1_outputs(6879) <= not a;
    layer1_outputs(6880) <= not a;
    layer1_outputs(6881) <= not (a and b);
    layer1_outputs(6882) <= a;
    layer1_outputs(6883) <= not a or b;
    layer1_outputs(6884) <= '1';
    layer1_outputs(6885) <= not (a and b);
    layer1_outputs(6886) <= b;
    layer1_outputs(6887) <= '1';
    layer1_outputs(6888) <= not a or b;
    layer1_outputs(6889) <= '1';
    layer1_outputs(6890) <= not b;
    layer1_outputs(6891) <= not b;
    layer1_outputs(6892) <= b;
    layer1_outputs(6893) <= not a or b;
    layer1_outputs(6894) <= a;
    layer1_outputs(6895) <= '1';
    layer1_outputs(6896) <= a or b;
    layer1_outputs(6897) <= not b;
    layer1_outputs(6898) <= not (a xor b);
    layer1_outputs(6899) <= not a;
    layer1_outputs(6900) <= not a or b;
    layer1_outputs(6901) <= not (a or b);
    layer1_outputs(6902) <= not (a and b);
    layer1_outputs(6903) <= '0';
    layer1_outputs(6904) <= a and b;
    layer1_outputs(6905) <= not (a xor b);
    layer1_outputs(6906) <= b and not a;
    layer1_outputs(6907) <= a or b;
    layer1_outputs(6908) <= a or b;
    layer1_outputs(6909) <= a;
    layer1_outputs(6910) <= not (a or b);
    layer1_outputs(6911) <= a or b;
    layer1_outputs(6912) <= not a;
    layer1_outputs(6913) <= not (a or b);
    layer1_outputs(6914) <= a or b;
    layer1_outputs(6915) <= not b or a;
    layer1_outputs(6916) <= '1';
    layer1_outputs(6917) <= not (a xor b);
    layer1_outputs(6918) <= b and not a;
    layer1_outputs(6919) <= b and not a;
    layer1_outputs(6920) <= not (a or b);
    layer1_outputs(6921) <= not (a or b);
    layer1_outputs(6922) <= a;
    layer1_outputs(6923) <= not b;
    layer1_outputs(6924) <= '1';
    layer1_outputs(6925) <= b;
    layer1_outputs(6926) <= '0';
    layer1_outputs(6927) <= '0';
    layer1_outputs(6928) <= not a;
    layer1_outputs(6929) <= a or b;
    layer1_outputs(6930) <= a and not b;
    layer1_outputs(6931) <= not (a or b);
    layer1_outputs(6932) <= not (a or b);
    layer1_outputs(6933) <= b and not a;
    layer1_outputs(6934) <= b;
    layer1_outputs(6935) <= not (a or b);
    layer1_outputs(6936) <= a and b;
    layer1_outputs(6937) <= b;
    layer1_outputs(6938) <= not a;
    layer1_outputs(6939) <= '1';
    layer1_outputs(6940) <= not b;
    layer1_outputs(6941) <= not a;
    layer1_outputs(6942) <= not a;
    layer1_outputs(6943) <= not a or b;
    layer1_outputs(6944) <= not a or b;
    layer1_outputs(6945) <= not b or a;
    layer1_outputs(6946) <= not (a or b);
    layer1_outputs(6947) <= a and b;
    layer1_outputs(6948) <= a;
    layer1_outputs(6949) <= not b;
    layer1_outputs(6950) <= '0';
    layer1_outputs(6951) <= a and not b;
    layer1_outputs(6952) <= '1';
    layer1_outputs(6953) <= not b or a;
    layer1_outputs(6954) <= not (a and b);
    layer1_outputs(6955) <= '1';
    layer1_outputs(6956) <= '0';
    layer1_outputs(6957) <= a and not b;
    layer1_outputs(6958) <= b and not a;
    layer1_outputs(6959) <= not a;
    layer1_outputs(6960) <= a;
    layer1_outputs(6961) <= not b;
    layer1_outputs(6962) <= not (a or b);
    layer1_outputs(6963) <= not a;
    layer1_outputs(6964) <= '1';
    layer1_outputs(6965) <= b;
    layer1_outputs(6966) <= not a;
    layer1_outputs(6967) <= not b or a;
    layer1_outputs(6968) <= a or b;
    layer1_outputs(6969) <= not a;
    layer1_outputs(6970) <= not a;
    layer1_outputs(6971) <= a and not b;
    layer1_outputs(6972) <= not a or b;
    layer1_outputs(6973) <= not b or a;
    layer1_outputs(6974) <= b;
    layer1_outputs(6975) <= '1';
    layer1_outputs(6976) <= a xor b;
    layer1_outputs(6977) <= a;
    layer1_outputs(6978) <= a xor b;
    layer1_outputs(6979) <= '1';
    layer1_outputs(6980) <= not b;
    layer1_outputs(6981) <= '1';
    layer1_outputs(6982) <= a and b;
    layer1_outputs(6983) <= not (a and b);
    layer1_outputs(6984) <= a;
    layer1_outputs(6985) <= not (a or b);
    layer1_outputs(6986) <= a;
    layer1_outputs(6987) <= b;
    layer1_outputs(6988) <= not b;
    layer1_outputs(6989) <= not b;
    layer1_outputs(6990) <= a or b;
    layer1_outputs(6991) <= a xor b;
    layer1_outputs(6992) <= not a or b;
    layer1_outputs(6993) <= a;
    layer1_outputs(6994) <= '0';
    layer1_outputs(6995) <= b and not a;
    layer1_outputs(6996) <= a;
    layer1_outputs(6997) <= not b;
    layer1_outputs(6998) <= not (a or b);
    layer1_outputs(6999) <= a and b;
    layer1_outputs(7000) <= b;
    layer1_outputs(7001) <= a and not b;
    layer1_outputs(7002) <= not a or b;
    layer1_outputs(7003) <= not a or b;
    layer1_outputs(7004) <= not a;
    layer1_outputs(7005) <= b and not a;
    layer1_outputs(7006) <= not a;
    layer1_outputs(7007) <= not a or b;
    layer1_outputs(7008) <= not b or a;
    layer1_outputs(7009) <= a or b;
    layer1_outputs(7010) <= a or b;
    layer1_outputs(7011) <= not a or b;
    layer1_outputs(7012) <= a xor b;
    layer1_outputs(7013) <= a and b;
    layer1_outputs(7014) <= '1';
    layer1_outputs(7015) <= not b;
    layer1_outputs(7016) <= a xor b;
    layer1_outputs(7017) <= not (a and b);
    layer1_outputs(7018) <= not (a or b);
    layer1_outputs(7019) <= '1';
    layer1_outputs(7020) <= not b or a;
    layer1_outputs(7021) <= '1';
    layer1_outputs(7022) <= '1';
    layer1_outputs(7023) <= not (a or b);
    layer1_outputs(7024) <= not b;
    layer1_outputs(7025) <= a and b;
    layer1_outputs(7026) <= a;
    layer1_outputs(7027) <= b;
    layer1_outputs(7028) <= not b;
    layer1_outputs(7029) <= not (a and b);
    layer1_outputs(7030) <= not (a or b);
    layer1_outputs(7031) <= not a;
    layer1_outputs(7032) <= not a or b;
    layer1_outputs(7033) <= '1';
    layer1_outputs(7034) <= '1';
    layer1_outputs(7035) <= not (a and b);
    layer1_outputs(7036) <= a;
    layer1_outputs(7037) <= a or b;
    layer1_outputs(7038) <= a and b;
    layer1_outputs(7039) <= not (a or b);
    layer1_outputs(7040) <= b;
    layer1_outputs(7041) <= a or b;
    layer1_outputs(7042) <= not a;
    layer1_outputs(7043) <= b;
    layer1_outputs(7044) <= a or b;
    layer1_outputs(7045) <= a and b;
    layer1_outputs(7046) <= a and not b;
    layer1_outputs(7047) <= not b or a;
    layer1_outputs(7048) <= a or b;
    layer1_outputs(7049) <= not (a and b);
    layer1_outputs(7050) <= not a or b;
    layer1_outputs(7051) <= '0';
    layer1_outputs(7052) <= not a;
    layer1_outputs(7053) <= not (a and b);
    layer1_outputs(7054) <= '1';
    layer1_outputs(7055) <= not (a or b);
    layer1_outputs(7056) <= not (a xor b);
    layer1_outputs(7057) <= not a;
    layer1_outputs(7058) <= b;
    layer1_outputs(7059) <= '0';
    layer1_outputs(7060) <= not a;
    layer1_outputs(7061) <= not (a or b);
    layer1_outputs(7062) <= not b;
    layer1_outputs(7063) <= not b;
    layer1_outputs(7064) <= b;
    layer1_outputs(7065) <= a or b;
    layer1_outputs(7066) <= not b or a;
    layer1_outputs(7067) <= not b;
    layer1_outputs(7068) <= not b or a;
    layer1_outputs(7069) <= a or b;
    layer1_outputs(7070) <= '0';
    layer1_outputs(7071) <= a and b;
    layer1_outputs(7072) <= a;
    layer1_outputs(7073) <= '1';
    layer1_outputs(7074) <= a or b;
    layer1_outputs(7075) <= a and b;
    layer1_outputs(7076) <= a or b;
    layer1_outputs(7077) <= not a or b;
    layer1_outputs(7078) <= not a;
    layer1_outputs(7079) <= '1';
    layer1_outputs(7080) <= not a or b;
    layer1_outputs(7081) <= a;
    layer1_outputs(7082) <= not a or b;
    layer1_outputs(7083) <= not b;
    layer1_outputs(7084) <= not a;
    layer1_outputs(7085) <= not b or a;
    layer1_outputs(7086) <= '0';
    layer1_outputs(7087) <= not a or b;
    layer1_outputs(7088) <= a or b;
    layer1_outputs(7089) <= a;
    layer1_outputs(7090) <= a;
    layer1_outputs(7091) <= b;
    layer1_outputs(7092) <= not b;
    layer1_outputs(7093) <= a xor b;
    layer1_outputs(7094) <= a and not b;
    layer1_outputs(7095) <= not (a or b);
    layer1_outputs(7096) <= b;
    layer1_outputs(7097) <= b;
    layer1_outputs(7098) <= b;
    layer1_outputs(7099) <= a;
    layer1_outputs(7100) <= a or b;
    layer1_outputs(7101) <= not a or b;
    layer1_outputs(7102) <= a;
    layer1_outputs(7103) <= not (a or b);
    layer1_outputs(7104) <= b and not a;
    layer1_outputs(7105) <= a;
    layer1_outputs(7106) <= not b or a;
    layer1_outputs(7107) <= a xor b;
    layer1_outputs(7108) <= a xor b;
    layer1_outputs(7109) <= not (a xor b);
    layer1_outputs(7110) <= not b or a;
    layer1_outputs(7111) <= not (a and b);
    layer1_outputs(7112) <= '1';
    layer1_outputs(7113) <= '1';
    layer1_outputs(7114) <= not (a and b);
    layer1_outputs(7115) <= b;
    layer1_outputs(7116) <= not b;
    layer1_outputs(7117) <= '1';
    layer1_outputs(7118) <= b;
    layer1_outputs(7119) <= b and not a;
    layer1_outputs(7120) <= b and not a;
    layer1_outputs(7121) <= not b;
    layer1_outputs(7122) <= b and not a;
    layer1_outputs(7123) <= a or b;
    layer1_outputs(7124) <= not (a xor b);
    layer1_outputs(7125) <= a;
    layer1_outputs(7126) <= a and not b;
    layer1_outputs(7127) <= a and not b;
    layer1_outputs(7128) <= '0';
    layer1_outputs(7129) <= b;
    layer1_outputs(7130) <= not b;
    layer1_outputs(7131) <= b and not a;
    layer1_outputs(7132) <= a;
    layer1_outputs(7133) <= not b;
    layer1_outputs(7134) <= b;
    layer1_outputs(7135) <= not b;
    layer1_outputs(7136) <= not a or b;
    layer1_outputs(7137) <= '0';
    layer1_outputs(7138) <= a or b;
    layer1_outputs(7139) <= not a;
    layer1_outputs(7140) <= b;
    layer1_outputs(7141) <= b;
    layer1_outputs(7142) <= a xor b;
    layer1_outputs(7143) <= not a or b;
    layer1_outputs(7144) <= b and not a;
    layer1_outputs(7145) <= b;
    layer1_outputs(7146) <= b;
    layer1_outputs(7147) <= b;
    layer1_outputs(7148) <= not a;
    layer1_outputs(7149) <= '0';
    layer1_outputs(7150) <= not (a or b);
    layer1_outputs(7151) <= a and b;
    layer1_outputs(7152) <= not b;
    layer1_outputs(7153) <= '0';
    layer1_outputs(7154) <= b;
    layer1_outputs(7155) <= not b or a;
    layer1_outputs(7156) <= a;
    layer1_outputs(7157) <= not b;
    layer1_outputs(7158) <= '1';
    layer1_outputs(7159) <= '0';
    layer1_outputs(7160) <= not (a or b);
    layer1_outputs(7161) <= not b;
    layer1_outputs(7162) <= b;
    layer1_outputs(7163) <= b and not a;
    layer1_outputs(7164) <= not b;
    layer1_outputs(7165) <= b;
    layer1_outputs(7166) <= a and not b;
    layer1_outputs(7167) <= '1';
    layer1_outputs(7168) <= not a;
    layer1_outputs(7169) <= not b;
    layer1_outputs(7170) <= a or b;
    layer1_outputs(7171) <= '1';
    layer1_outputs(7172) <= b and not a;
    layer1_outputs(7173) <= not a;
    layer1_outputs(7174) <= not a;
    layer1_outputs(7175) <= not a or b;
    layer1_outputs(7176) <= not (a or b);
    layer1_outputs(7177) <= a and b;
    layer1_outputs(7178) <= '1';
    layer1_outputs(7179) <= b;
    layer1_outputs(7180) <= not a or b;
    layer1_outputs(7181) <= b;
    layer1_outputs(7182) <= not b;
    layer1_outputs(7183) <= not b or a;
    layer1_outputs(7184) <= '1';
    layer1_outputs(7185) <= not a;
    layer1_outputs(7186) <= not a;
    layer1_outputs(7187) <= not (a and b);
    layer1_outputs(7188) <= a or b;
    layer1_outputs(7189) <= a;
    layer1_outputs(7190) <= b and not a;
    layer1_outputs(7191) <= b and not a;
    layer1_outputs(7192) <= not (a and b);
    layer1_outputs(7193) <= not (a or b);
    layer1_outputs(7194) <= not (a and b);
    layer1_outputs(7195) <= '0';
    layer1_outputs(7196) <= '0';
    layer1_outputs(7197) <= a and b;
    layer1_outputs(7198) <= not (a xor b);
    layer1_outputs(7199) <= '0';
    layer1_outputs(7200) <= b;
    layer1_outputs(7201) <= not (a and b);
    layer1_outputs(7202) <= a;
    layer1_outputs(7203) <= '0';
    layer1_outputs(7204) <= not a or b;
    layer1_outputs(7205) <= not a or b;
    layer1_outputs(7206) <= '1';
    layer1_outputs(7207) <= a;
    layer1_outputs(7208) <= b;
    layer1_outputs(7209) <= not (a and b);
    layer1_outputs(7210) <= not (a xor b);
    layer1_outputs(7211) <= a;
    layer1_outputs(7212) <= a and b;
    layer1_outputs(7213) <= not b or a;
    layer1_outputs(7214) <= not a;
    layer1_outputs(7215) <= not b or a;
    layer1_outputs(7216) <= not a;
    layer1_outputs(7217) <= not (a or b);
    layer1_outputs(7218) <= '0';
    layer1_outputs(7219) <= b and not a;
    layer1_outputs(7220) <= b;
    layer1_outputs(7221) <= not b or a;
    layer1_outputs(7222) <= '1';
    layer1_outputs(7223) <= a;
    layer1_outputs(7224) <= '1';
    layer1_outputs(7225) <= not (a or b);
    layer1_outputs(7226) <= not a;
    layer1_outputs(7227) <= not a or b;
    layer1_outputs(7228) <= b and not a;
    layer1_outputs(7229) <= not a or b;
    layer1_outputs(7230) <= not b;
    layer1_outputs(7231) <= a and not b;
    layer1_outputs(7232) <= b and not a;
    layer1_outputs(7233) <= '1';
    layer1_outputs(7234) <= not a;
    layer1_outputs(7235) <= not a;
    layer1_outputs(7236) <= a;
    layer1_outputs(7237) <= not b or a;
    layer1_outputs(7238) <= a;
    layer1_outputs(7239) <= not b;
    layer1_outputs(7240) <= not b;
    layer1_outputs(7241) <= not a or b;
    layer1_outputs(7242) <= '1';
    layer1_outputs(7243) <= not (a or b);
    layer1_outputs(7244) <= b and not a;
    layer1_outputs(7245) <= a xor b;
    layer1_outputs(7246) <= a or b;
    layer1_outputs(7247) <= not (a xor b);
    layer1_outputs(7248) <= a;
    layer1_outputs(7249) <= not b;
    layer1_outputs(7250) <= not (a xor b);
    layer1_outputs(7251) <= a;
    layer1_outputs(7252) <= '1';
    layer1_outputs(7253) <= a and not b;
    layer1_outputs(7254) <= not a or b;
    layer1_outputs(7255) <= not (a xor b);
    layer1_outputs(7256) <= not a or b;
    layer1_outputs(7257) <= not (a and b);
    layer1_outputs(7258) <= b and not a;
    layer1_outputs(7259) <= a and not b;
    layer1_outputs(7260) <= a;
    layer1_outputs(7261) <= not a;
    layer1_outputs(7262) <= a xor b;
    layer1_outputs(7263) <= a and not b;
    layer1_outputs(7264) <= a and b;
    layer1_outputs(7265) <= b;
    layer1_outputs(7266) <= a and not b;
    layer1_outputs(7267) <= '1';
    layer1_outputs(7268) <= '1';
    layer1_outputs(7269) <= b;
    layer1_outputs(7270) <= not (a or b);
    layer1_outputs(7271) <= not b or a;
    layer1_outputs(7272) <= a or b;
    layer1_outputs(7273) <= not a;
    layer1_outputs(7274) <= not (a or b);
    layer1_outputs(7275) <= not a or b;
    layer1_outputs(7276) <= not (a xor b);
    layer1_outputs(7277) <= a or b;
    layer1_outputs(7278) <= not b;
    layer1_outputs(7279) <= not a or b;
    layer1_outputs(7280) <= not a or b;
    layer1_outputs(7281) <= a xor b;
    layer1_outputs(7282) <= b;
    layer1_outputs(7283) <= b and not a;
    layer1_outputs(7284) <= a and not b;
    layer1_outputs(7285) <= a xor b;
    layer1_outputs(7286) <= a or b;
    layer1_outputs(7287) <= a;
    layer1_outputs(7288) <= not a or b;
    layer1_outputs(7289) <= not (a xor b);
    layer1_outputs(7290) <= '1';
    layer1_outputs(7291) <= '0';
    layer1_outputs(7292) <= a;
    layer1_outputs(7293) <= not (a xor b);
    layer1_outputs(7294) <= not b;
    layer1_outputs(7295) <= a and b;
    layer1_outputs(7296) <= a or b;
    layer1_outputs(7297) <= b;
    layer1_outputs(7298) <= a and not b;
    layer1_outputs(7299) <= not (a and b);
    layer1_outputs(7300) <= not a;
    layer1_outputs(7301) <= not (a or b);
    layer1_outputs(7302) <= b and not a;
    layer1_outputs(7303) <= a and b;
    layer1_outputs(7304) <= a or b;
    layer1_outputs(7305) <= not (a or b);
    layer1_outputs(7306) <= not a or b;
    layer1_outputs(7307) <= not (a xor b);
    layer1_outputs(7308) <= a or b;
    layer1_outputs(7309) <= a and not b;
    layer1_outputs(7310) <= not b or a;
    layer1_outputs(7311) <= a;
    layer1_outputs(7312) <= a and not b;
    layer1_outputs(7313) <= not (a and b);
    layer1_outputs(7314) <= b and not a;
    layer1_outputs(7315) <= not (a xor b);
    layer1_outputs(7316) <= not (a or b);
    layer1_outputs(7317) <= a and not b;
    layer1_outputs(7318) <= not a or b;
    layer1_outputs(7319) <= not b or a;
    layer1_outputs(7320) <= not (a and b);
    layer1_outputs(7321) <= '1';
    layer1_outputs(7322) <= a xor b;
    layer1_outputs(7323) <= a;
    layer1_outputs(7324) <= a or b;
    layer1_outputs(7325) <= b;
    layer1_outputs(7326) <= not a or b;
    layer1_outputs(7327) <= a or b;
    layer1_outputs(7328) <= b;
    layer1_outputs(7329) <= not b;
    layer1_outputs(7330) <= a or b;
    layer1_outputs(7331) <= a xor b;
    layer1_outputs(7332) <= not a;
    layer1_outputs(7333) <= not b;
    layer1_outputs(7334) <= a or b;
    layer1_outputs(7335) <= a and b;
    layer1_outputs(7336) <= a or b;
    layer1_outputs(7337) <= not (a and b);
    layer1_outputs(7338) <= not (a or b);
    layer1_outputs(7339) <= not a;
    layer1_outputs(7340) <= not (a and b);
    layer1_outputs(7341) <= not b;
    layer1_outputs(7342) <= not a;
    layer1_outputs(7343) <= b;
    layer1_outputs(7344) <= not b or a;
    layer1_outputs(7345) <= '1';
    layer1_outputs(7346) <= a and not b;
    layer1_outputs(7347) <= not (a or b);
    layer1_outputs(7348) <= not a or b;
    layer1_outputs(7349) <= not b or a;
    layer1_outputs(7350) <= not (a and b);
    layer1_outputs(7351) <= b and not a;
    layer1_outputs(7352) <= not a or b;
    layer1_outputs(7353) <= '0';
    layer1_outputs(7354) <= a and b;
    layer1_outputs(7355) <= not a;
    layer1_outputs(7356) <= not (a or b);
    layer1_outputs(7357) <= not a;
    layer1_outputs(7358) <= a xor b;
    layer1_outputs(7359) <= not a or b;
    layer1_outputs(7360) <= not (a and b);
    layer1_outputs(7361) <= not b;
    layer1_outputs(7362) <= '0';
    layer1_outputs(7363) <= a or b;
    layer1_outputs(7364) <= a;
    layer1_outputs(7365) <= b;
    layer1_outputs(7366) <= not a or b;
    layer1_outputs(7367) <= not (a or b);
    layer1_outputs(7368) <= not a;
    layer1_outputs(7369) <= b and not a;
    layer1_outputs(7370) <= not b;
    layer1_outputs(7371) <= not a or b;
    layer1_outputs(7372) <= a and not b;
    layer1_outputs(7373) <= a or b;
    layer1_outputs(7374) <= a and not b;
    layer1_outputs(7375) <= not a or b;
    layer1_outputs(7376) <= b;
    layer1_outputs(7377) <= not (a or b);
    layer1_outputs(7378) <= not (a xor b);
    layer1_outputs(7379) <= '1';
    layer1_outputs(7380) <= b and not a;
    layer1_outputs(7381) <= '0';
    layer1_outputs(7382) <= not a;
    layer1_outputs(7383) <= b;
    layer1_outputs(7384) <= not b or a;
    layer1_outputs(7385) <= not (a xor b);
    layer1_outputs(7386) <= a and not b;
    layer1_outputs(7387) <= '1';
    layer1_outputs(7388) <= not a;
    layer1_outputs(7389) <= not (a xor b);
    layer1_outputs(7390) <= a or b;
    layer1_outputs(7391) <= a and not b;
    layer1_outputs(7392) <= not (a or b);
    layer1_outputs(7393) <= not (a or b);
    layer1_outputs(7394) <= b;
    layer1_outputs(7395) <= a and not b;
    layer1_outputs(7396) <= a and b;
    layer1_outputs(7397) <= a and not b;
    layer1_outputs(7398) <= not b or a;
    layer1_outputs(7399) <= b and not a;
    layer1_outputs(7400) <= not a or b;
    layer1_outputs(7401) <= a;
    layer1_outputs(7402) <= b;
    layer1_outputs(7403) <= not a or b;
    layer1_outputs(7404) <= a or b;
    layer1_outputs(7405) <= b and not a;
    layer1_outputs(7406) <= not (a and b);
    layer1_outputs(7407) <= b;
    layer1_outputs(7408) <= '1';
    layer1_outputs(7409) <= a and b;
    layer1_outputs(7410) <= not a or b;
    layer1_outputs(7411) <= not (a xor b);
    layer1_outputs(7412) <= '1';
    layer1_outputs(7413) <= not b or a;
    layer1_outputs(7414) <= a and not b;
    layer1_outputs(7415) <= not b or a;
    layer1_outputs(7416) <= not b;
    layer1_outputs(7417) <= '0';
    layer1_outputs(7418) <= not a;
    layer1_outputs(7419) <= b;
    layer1_outputs(7420) <= not (a xor b);
    layer1_outputs(7421) <= not (a and b);
    layer1_outputs(7422) <= not a;
    layer1_outputs(7423) <= not a;
    layer1_outputs(7424) <= not b;
    layer1_outputs(7425) <= a and b;
    layer1_outputs(7426) <= b and not a;
    layer1_outputs(7427) <= not b;
    layer1_outputs(7428) <= not a;
    layer1_outputs(7429) <= not (a xor b);
    layer1_outputs(7430) <= not a;
    layer1_outputs(7431) <= '0';
    layer1_outputs(7432) <= not b or a;
    layer1_outputs(7433) <= a;
    layer1_outputs(7434) <= a and b;
    layer1_outputs(7435) <= not (a or b);
    layer1_outputs(7436) <= b and not a;
    layer1_outputs(7437) <= b and not a;
    layer1_outputs(7438) <= a or b;
    layer1_outputs(7439) <= '0';
    layer1_outputs(7440) <= not a;
    layer1_outputs(7441) <= not (a or b);
    layer1_outputs(7442) <= not a;
    layer1_outputs(7443) <= a or b;
    layer1_outputs(7444) <= not b or a;
    layer1_outputs(7445) <= b;
    layer1_outputs(7446) <= not a or b;
    layer1_outputs(7447) <= not (a or b);
    layer1_outputs(7448) <= not a;
    layer1_outputs(7449) <= b and not a;
    layer1_outputs(7450) <= not (a and b);
    layer1_outputs(7451) <= '1';
    layer1_outputs(7452) <= b;
    layer1_outputs(7453) <= a xor b;
    layer1_outputs(7454) <= not b;
    layer1_outputs(7455) <= not (a and b);
    layer1_outputs(7456) <= b and not a;
    layer1_outputs(7457) <= a;
    layer1_outputs(7458) <= a and not b;
    layer1_outputs(7459) <= not b;
    layer1_outputs(7460) <= not b or a;
    layer1_outputs(7461) <= a or b;
    layer1_outputs(7462) <= a;
    layer1_outputs(7463) <= a or b;
    layer1_outputs(7464) <= '1';
    layer1_outputs(7465) <= a;
    layer1_outputs(7466) <= not b;
    layer1_outputs(7467) <= not (a or b);
    layer1_outputs(7468) <= '0';
    layer1_outputs(7469) <= not a or b;
    layer1_outputs(7470) <= not a;
    layer1_outputs(7471) <= not a;
    layer1_outputs(7472) <= a or b;
    layer1_outputs(7473) <= a or b;
    layer1_outputs(7474) <= not (a xor b);
    layer1_outputs(7475) <= '0';
    layer1_outputs(7476) <= not (a xor b);
    layer1_outputs(7477) <= not (a and b);
    layer1_outputs(7478) <= a or b;
    layer1_outputs(7479) <= not (a xor b);
    layer1_outputs(7480) <= a or b;
    layer1_outputs(7481) <= not a or b;
    layer1_outputs(7482) <= not (a and b);
    layer1_outputs(7483) <= b and not a;
    layer1_outputs(7484) <= not (a xor b);
    layer1_outputs(7485) <= b and not a;
    layer1_outputs(7486) <= not b;
    layer1_outputs(7487) <= not (a or b);
    layer1_outputs(7488) <= a;
    layer1_outputs(7489) <= b and not a;
    layer1_outputs(7490) <= b and not a;
    layer1_outputs(7491) <= '0';
    layer1_outputs(7492) <= not a;
    layer1_outputs(7493) <= a and not b;
    layer1_outputs(7494) <= a;
    layer1_outputs(7495) <= not b or a;
    layer1_outputs(7496) <= a and not b;
    layer1_outputs(7497) <= a;
    layer1_outputs(7498) <= a and b;
    layer1_outputs(7499) <= a xor b;
    layer1_outputs(7500) <= a or b;
    layer1_outputs(7501) <= not b or a;
    layer1_outputs(7502) <= not (a or b);
    layer1_outputs(7503) <= a and not b;
    layer1_outputs(7504) <= b and not a;
    layer1_outputs(7505) <= not (a and b);
    layer1_outputs(7506) <= not a;
    layer1_outputs(7507) <= b;
    layer1_outputs(7508) <= '1';
    layer1_outputs(7509) <= not a;
    layer1_outputs(7510) <= a;
    layer1_outputs(7511) <= not a or b;
    layer1_outputs(7512) <= a;
    layer1_outputs(7513) <= not a;
    layer1_outputs(7514) <= not a or b;
    layer1_outputs(7515) <= not b or a;
    layer1_outputs(7516) <= a;
    layer1_outputs(7517) <= '0';
    layer1_outputs(7518) <= not b;
    layer1_outputs(7519) <= a or b;
    layer1_outputs(7520) <= b and not a;
    layer1_outputs(7521) <= not a;
    layer1_outputs(7522) <= a or b;
    layer1_outputs(7523) <= b and not a;
    layer1_outputs(7524) <= not b or a;
    layer1_outputs(7525) <= not b or a;
    layer1_outputs(7526) <= not b;
    layer1_outputs(7527) <= a or b;
    layer1_outputs(7528) <= not a or b;
    layer1_outputs(7529) <= b;
    layer1_outputs(7530) <= a and b;
    layer1_outputs(7531) <= '0';
    layer1_outputs(7532) <= b and not a;
    layer1_outputs(7533) <= a or b;
    layer1_outputs(7534) <= b and not a;
    layer1_outputs(7535) <= '1';
    layer1_outputs(7536) <= not b or a;
    layer1_outputs(7537) <= a;
    layer1_outputs(7538) <= not a;
    layer1_outputs(7539) <= b and not a;
    layer1_outputs(7540) <= a or b;
    layer1_outputs(7541) <= b;
    layer1_outputs(7542) <= not a or b;
    layer1_outputs(7543) <= not b;
    layer1_outputs(7544) <= not a or b;
    layer1_outputs(7545) <= '0';
    layer1_outputs(7546) <= not (a and b);
    layer1_outputs(7547) <= not a;
    layer1_outputs(7548) <= a and not b;
    layer1_outputs(7549) <= not b or a;
    layer1_outputs(7550) <= b and not a;
    layer1_outputs(7551) <= not (a and b);
    layer1_outputs(7552) <= not a or b;
    layer1_outputs(7553) <= b and not a;
    layer1_outputs(7554) <= a and b;
    layer1_outputs(7555) <= not a or b;
    layer1_outputs(7556) <= '1';
    layer1_outputs(7557) <= '1';
    layer1_outputs(7558) <= a and b;
    layer1_outputs(7559) <= a and not b;
    layer1_outputs(7560) <= a and not b;
    layer1_outputs(7561) <= a and not b;
    layer1_outputs(7562) <= not a;
    layer1_outputs(7563) <= b;
    layer1_outputs(7564) <= a xor b;
    layer1_outputs(7565) <= a or b;
    layer1_outputs(7566) <= a;
    layer1_outputs(7567) <= '0';
    layer1_outputs(7568) <= a and b;
    layer1_outputs(7569) <= '0';
    layer1_outputs(7570) <= a;
    layer1_outputs(7571) <= not b or a;
    layer1_outputs(7572) <= not (a xor b);
    layer1_outputs(7573) <= b and not a;
    layer1_outputs(7574) <= a and not b;
    layer1_outputs(7575) <= '0';
    layer1_outputs(7576) <= a and not b;
    layer1_outputs(7577) <= a or b;
    layer1_outputs(7578) <= '0';
    layer1_outputs(7579) <= not a;
    layer1_outputs(7580) <= not b;
    layer1_outputs(7581) <= '0';
    layer1_outputs(7582) <= a and b;
    layer1_outputs(7583) <= a;
    layer1_outputs(7584) <= not b or a;
    layer1_outputs(7585) <= not (a and b);
    layer1_outputs(7586) <= a and b;
    layer1_outputs(7587) <= b and not a;
    layer1_outputs(7588) <= not (a xor b);
    layer1_outputs(7589) <= b;
    layer1_outputs(7590) <= a or b;
    layer1_outputs(7591) <= not (a and b);
    layer1_outputs(7592) <= a xor b;
    layer1_outputs(7593) <= not b or a;
    layer1_outputs(7594) <= not b or a;
    layer1_outputs(7595) <= not a or b;
    layer1_outputs(7596) <= b;
    layer1_outputs(7597) <= a;
    layer1_outputs(7598) <= not a or b;
    layer1_outputs(7599) <= a and b;
    layer1_outputs(7600) <= not (a or b);
    layer1_outputs(7601) <= not a;
    layer1_outputs(7602) <= a or b;
    layer1_outputs(7603) <= not a or b;
    layer1_outputs(7604) <= '0';
    layer1_outputs(7605) <= b and not a;
    layer1_outputs(7606) <= not a or b;
    layer1_outputs(7607) <= a and not b;
    layer1_outputs(7608) <= not a;
    layer1_outputs(7609) <= b;
    layer1_outputs(7610) <= a and b;
    layer1_outputs(7611) <= not a or b;
    layer1_outputs(7612) <= a;
    layer1_outputs(7613) <= '1';
    layer1_outputs(7614) <= not b;
    layer1_outputs(7615) <= not a;
    layer1_outputs(7616) <= a;
    layer1_outputs(7617) <= a or b;
    layer1_outputs(7618) <= not b;
    layer1_outputs(7619) <= '1';
    layer1_outputs(7620) <= not (a and b);
    layer1_outputs(7621) <= not b;
    layer1_outputs(7622) <= not (a and b);
    layer1_outputs(7623) <= not (a and b);
    layer1_outputs(7624) <= '1';
    layer1_outputs(7625) <= a or b;
    layer1_outputs(7626) <= b;
    layer1_outputs(7627) <= '1';
    layer1_outputs(7628) <= not b;
    layer1_outputs(7629) <= a and not b;
    layer1_outputs(7630) <= not (a and b);
    layer1_outputs(7631) <= not (a and b);
    layer1_outputs(7632) <= not a or b;
    layer1_outputs(7633) <= not a;
    layer1_outputs(7634) <= not a;
    layer1_outputs(7635) <= a and b;
    layer1_outputs(7636) <= '0';
    layer1_outputs(7637) <= not (a and b);
    layer1_outputs(7638) <= not b or a;
    layer1_outputs(7639) <= '1';
    layer1_outputs(7640) <= a and not b;
    layer1_outputs(7641) <= a or b;
    layer1_outputs(7642) <= a;
    layer1_outputs(7643) <= a;
    layer1_outputs(7644) <= a and not b;
    layer1_outputs(7645) <= a and b;
    layer1_outputs(7646) <= a and not b;
    layer1_outputs(7647) <= not b;
    layer1_outputs(7648) <= not b;
    layer1_outputs(7649) <= not a;
    layer1_outputs(7650) <= '0';
    layer1_outputs(7651) <= not b;
    layer1_outputs(7652) <= not a or b;
    layer1_outputs(7653) <= not b or a;
    layer1_outputs(7654) <= b;
    layer1_outputs(7655) <= '0';
    layer1_outputs(7656) <= not (a xor b);
    layer1_outputs(7657) <= a;
    layer1_outputs(7658) <= not (a and b);
    layer1_outputs(7659) <= not b;
    layer1_outputs(7660) <= b and not a;
    layer1_outputs(7661) <= a or b;
    layer1_outputs(7662) <= a;
    layer1_outputs(7663) <= not (a xor b);
    layer1_outputs(7664) <= not (a or b);
    layer1_outputs(7665) <= a or b;
    layer1_outputs(7666) <= not (a or b);
    layer1_outputs(7667) <= '1';
    layer1_outputs(7668) <= a xor b;
    layer1_outputs(7669) <= b;
    layer1_outputs(7670) <= a;
    layer1_outputs(7671) <= not (a and b);
    layer1_outputs(7672) <= '0';
    layer1_outputs(7673) <= a and not b;
    layer1_outputs(7674) <= a or b;
    layer1_outputs(7675) <= not b;
    layer1_outputs(7676) <= not (a or b);
    layer1_outputs(7677) <= a;
    layer1_outputs(7678) <= not b or a;
    layer1_outputs(7679) <= not b;
    layer1_outputs(7680) <= b;
    layer1_outputs(7681) <= not a;
    layer1_outputs(7682) <= not b;
    layer1_outputs(7683) <= '0';
    layer1_outputs(7684) <= '1';
    layer1_outputs(7685) <= '0';
    layer1_outputs(7686) <= not (a or b);
    layer1_outputs(7687) <= not a or b;
    layer1_outputs(7688) <= '1';
    layer1_outputs(7689) <= a xor b;
    layer1_outputs(7690) <= a and b;
    layer1_outputs(7691) <= b;
    layer1_outputs(7692) <= not (a or b);
    layer1_outputs(7693) <= not a or b;
    layer1_outputs(7694) <= '0';
    layer1_outputs(7695) <= a xor b;
    layer1_outputs(7696) <= b;
    layer1_outputs(7697) <= '0';
    layer1_outputs(7698) <= not a;
    layer1_outputs(7699) <= a or b;
    layer1_outputs(7700) <= not b or a;
    layer1_outputs(7701) <= a and b;
    layer1_outputs(7702) <= a or b;
    layer1_outputs(7703) <= b;
    layer1_outputs(7704) <= b;
    layer1_outputs(7705) <= not (a or b);
    layer1_outputs(7706) <= a or b;
    layer1_outputs(7707) <= '0';
    layer1_outputs(7708) <= not b;
    layer1_outputs(7709) <= not a or b;
    layer1_outputs(7710) <= not b;
    layer1_outputs(7711) <= b;
    layer1_outputs(7712) <= not (a or b);
    layer1_outputs(7713) <= not b or a;
    layer1_outputs(7714) <= b;
    layer1_outputs(7715) <= not a;
    layer1_outputs(7716) <= not b or a;
    layer1_outputs(7717) <= b and not a;
    layer1_outputs(7718) <= a and not b;
    layer1_outputs(7719) <= b;
    layer1_outputs(7720) <= b and not a;
    layer1_outputs(7721) <= not a or b;
    layer1_outputs(7722) <= a or b;
    layer1_outputs(7723) <= not b or a;
    layer1_outputs(7724) <= a and not b;
    layer1_outputs(7725) <= a and not b;
    layer1_outputs(7726) <= a and not b;
    layer1_outputs(7727) <= b and not a;
    layer1_outputs(7728) <= b;
    layer1_outputs(7729) <= a xor b;
    layer1_outputs(7730) <= not a;
    layer1_outputs(7731) <= not (a and b);
    layer1_outputs(7732) <= not a;
    layer1_outputs(7733) <= a and b;
    layer1_outputs(7734) <= a;
    layer1_outputs(7735) <= a;
    layer1_outputs(7736) <= not (a xor b);
    layer1_outputs(7737) <= not b;
    layer1_outputs(7738) <= b;
    layer1_outputs(7739) <= not (a and b);
    layer1_outputs(7740) <= a;
    layer1_outputs(7741) <= not b;
    layer1_outputs(7742) <= b and not a;
    layer1_outputs(7743) <= not (a and b);
    layer1_outputs(7744) <= a and not b;
    layer1_outputs(7745) <= a;
    layer1_outputs(7746) <= '1';
    layer1_outputs(7747) <= '1';
    layer1_outputs(7748) <= not (a xor b);
    layer1_outputs(7749) <= '0';
    layer1_outputs(7750) <= b;
    layer1_outputs(7751) <= b;
    layer1_outputs(7752) <= not (a and b);
    layer1_outputs(7753) <= not b or a;
    layer1_outputs(7754) <= '1';
    layer1_outputs(7755) <= b;
    layer1_outputs(7756) <= not a or b;
    layer1_outputs(7757) <= a and not b;
    layer1_outputs(7758) <= b and not a;
    layer1_outputs(7759) <= a or b;
    layer1_outputs(7760) <= a and not b;
    layer1_outputs(7761) <= not a or b;
    layer1_outputs(7762) <= not a;
    layer1_outputs(7763) <= b and not a;
    layer1_outputs(7764) <= a;
    layer1_outputs(7765) <= b and not a;
    layer1_outputs(7766) <= b and not a;
    layer1_outputs(7767) <= not b;
    layer1_outputs(7768) <= not (a and b);
    layer1_outputs(7769) <= not (a and b);
    layer1_outputs(7770) <= not (a or b);
    layer1_outputs(7771) <= not b;
    layer1_outputs(7772) <= a xor b;
    layer1_outputs(7773) <= a;
    layer1_outputs(7774) <= a xor b;
    layer1_outputs(7775) <= not a or b;
    layer1_outputs(7776) <= not (a and b);
    layer1_outputs(7777) <= a and b;
    layer1_outputs(7778) <= not a or b;
    layer1_outputs(7779) <= '1';
    layer1_outputs(7780) <= b and not a;
    layer1_outputs(7781) <= '0';
    layer1_outputs(7782) <= not a or b;
    layer1_outputs(7783) <= not b;
    layer1_outputs(7784) <= not b;
    layer1_outputs(7785) <= not b or a;
    layer1_outputs(7786) <= not b;
    layer1_outputs(7787) <= not (a or b);
    layer1_outputs(7788) <= not (a xor b);
    layer1_outputs(7789) <= not b or a;
    layer1_outputs(7790) <= not a or b;
    layer1_outputs(7791) <= not (a and b);
    layer1_outputs(7792) <= a xor b;
    layer1_outputs(7793) <= not (a and b);
    layer1_outputs(7794) <= a and not b;
    layer1_outputs(7795) <= not (a xor b);
    layer1_outputs(7796) <= a;
    layer1_outputs(7797) <= a or b;
    layer1_outputs(7798) <= a or b;
    layer1_outputs(7799) <= a xor b;
    layer1_outputs(7800) <= a or b;
    layer1_outputs(7801) <= a;
    layer1_outputs(7802) <= a and b;
    layer1_outputs(7803) <= a;
    layer1_outputs(7804) <= not (a and b);
    layer1_outputs(7805) <= not (a and b);
    layer1_outputs(7806) <= not b;
    layer1_outputs(7807) <= not (a or b);
    layer1_outputs(7808) <= a and b;
    layer1_outputs(7809) <= not b or a;
    layer1_outputs(7810) <= a and not b;
    layer1_outputs(7811) <= b;
    layer1_outputs(7812) <= '0';
    layer1_outputs(7813) <= not a;
    layer1_outputs(7814) <= not b;
    layer1_outputs(7815) <= not a or b;
    layer1_outputs(7816) <= not b or a;
    layer1_outputs(7817) <= not a;
    layer1_outputs(7818) <= '1';
    layer1_outputs(7819) <= not (a and b);
    layer1_outputs(7820) <= b;
    layer1_outputs(7821) <= a;
    layer1_outputs(7822) <= a or b;
    layer1_outputs(7823) <= b;
    layer1_outputs(7824) <= b;
    layer1_outputs(7825) <= not (a xor b);
    layer1_outputs(7826) <= not a;
    layer1_outputs(7827) <= not a or b;
    layer1_outputs(7828) <= not (a xor b);
    layer1_outputs(7829) <= not (a xor b);
    layer1_outputs(7830) <= a or b;
    layer1_outputs(7831) <= not b or a;
    layer1_outputs(7832) <= not b;
    layer1_outputs(7833) <= '0';
    layer1_outputs(7834) <= b;
    layer1_outputs(7835) <= a or b;
    layer1_outputs(7836) <= not (a and b);
    layer1_outputs(7837) <= a xor b;
    layer1_outputs(7838) <= not (a or b);
    layer1_outputs(7839) <= b;
    layer1_outputs(7840) <= a or b;
    layer1_outputs(7841) <= not (a or b);
    layer1_outputs(7842) <= not a;
    layer1_outputs(7843) <= not a or b;
    layer1_outputs(7844) <= not a;
    layer1_outputs(7845) <= not a or b;
    layer1_outputs(7846) <= '0';
    layer1_outputs(7847) <= b;
    layer1_outputs(7848) <= not (a xor b);
    layer1_outputs(7849) <= not (a or b);
    layer1_outputs(7850) <= b;
    layer1_outputs(7851) <= a and b;
    layer1_outputs(7852) <= not (a xor b);
    layer1_outputs(7853) <= a xor b;
    layer1_outputs(7854) <= b and not a;
    layer1_outputs(7855) <= not (a or b);
    layer1_outputs(7856) <= '1';
    layer1_outputs(7857) <= not (a and b);
    layer1_outputs(7858) <= a and not b;
    layer1_outputs(7859) <= b;
    layer1_outputs(7860) <= not b or a;
    layer1_outputs(7861) <= b and not a;
    layer1_outputs(7862) <= '0';
    layer1_outputs(7863) <= a xor b;
    layer1_outputs(7864) <= a;
    layer1_outputs(7865) <= not (a xor b);
    layer1_outputs(7866) <= '1';
    layer1_outputs(7867) <= not a;
    layer1_outputs(7868) <= a and not b;
    layer1_outputs(7869) <= b;
    layer1_outputs(7870) <= a or b;
    layer1_outputs(7871) <= not a or b;
    layer1_outputs(7872) <= a xor b;
    layer1_outputs(7873) <= not (a and b);
    layer1_outputs(7874) <= a;
    layer1_outputs(7875) <= a xor b;
    layer1_outputs(7876) <= '1';
    layer1_outputs(7877) <= not (a xor b);
    layer1_outputs(7878) <= a and b;
    layer1_outputs(7879) <= a or b;
    layer1_outputs(7880) <= not b or a;
    layer1_outputs(7881) <= not (a and b);
    layer1_outputs(7882) <= not (a or b);
    layer1_outputs(7883) <= b;
    layer1_outputs(7884) <= a or b;
    layer1_outputs(7885) <= a;
    layer1_outputs(7886) <= not b;
    layer1_outputs(7887) <= b and not a;
    layer1_outputs(7888) <= '1';
    layer1_outputs(7889) <= not b;
    layer1_outputs(7890) <= a and b;
    layer1_outputs(7891) <= not a;
    layer1_outputs(7892) <= '1';
    layer1_outputs(7893) <= not a or b;
    layer1_outputs(7894) <= b;
    layer1_outputs(7895) <= b and not a;
    layer1_outputs(7896) <= not a or b;
    layer1_outputs(7897) <= a or b;
    layer1_outputs(7898) <= a and not b;
    layer1_outputs(7899) <= b and not a;
    layer1_outputs(7900) <= not a or b;
    layer1_outputs(7901) <= a and not b;
    layer1_outputs(7902) <= not b;
    layer1_outputs(7903) <= not a or b;
    layer1_outputs(7904) <= a and b;
    layer1_outputs(7905) <= '0';
    layer1_outputs(7906) <= b and not a;
    layer1_outputs(7907) <= a xor b;
    layer1_outputs(7908) <= not b;
    layer1_outputs(7909) <= not (a xor b);
    layer1_outputs(7910) <= not (a and b);
    layer1_outputs(7911) <= b;
    layer1_outputs(7912) <= '1';
    layer1_outputs(7913) <= a;
    layer1_outputs(7914) <= b;
    layer1_outputs(7915) <= b;
    layer1_outputs(7916) <= a or b;
    layer1_outputs(7917) <= not a;
    layer1_outputs(7918) <= a and not b;
    layer1_outputs(7919) <= not a;
    layer1_outputs(7920) <= not (a or b);
    layer1_outputs(7921) <= a and not b;
    layer1_outputs(7922) <= not a;
    layer1_outputs(7923) <= '0';
    layer1_outputs(7924) <= not b or a;
    layer1_outputs(7925) <= not (a or b);
    layer1_outputs(7926) <= a;
    layer1_outputs(7927) <= a or b;
    layer1_outputs(7928) <= '0';
    layer1_outputs(7929) <= '0';
    layer1_outputs(7930) <= b and not a;
    layer1_outputs(7931) <= b;
    layer1_outputs(7932) <= '1';
    layer1_outputs(7933) <= not (a and b);
    layer1_outputs(7934) <= a;
    layer1_outputs(7935) <= '1';
    layer1_outputs(7936) <= not (a and b);
    layer1_outputs(7937) <= '1';
    layer1_outputs(7938) <= '1';
    layer1_outputs(7939) <= b;
    layer1_outputs(7940) <= not b or a;
    layer1_outputs(7941) <= a and not b;
    layer1_outputs(7942) <= a or b;
    layer1_outputs(7943) <= not (a and b);
    layer1_outputs(7944) <= not a;
    layer1_outputs(7945) <= not a;
    layer1_outputs(7946) <= a;
    layer1_outputs(7947) <= not (a and b);
    layer1_outputs(7948) <= a and not b;
    layer1_outputs(7949) <= b;
    layer1_outputs(7950) <= b and not a;
    layer1_outputs(7951) <= b;
    layer1_outputs(7952) <= a or b;
    layer1_outputs(7953) <= '1';
    layer1_outputs(7954) <= not a or b;
    layer1_outputs(7955) <= '0';
    layer1_outputs(7956) <= a and b;
    layer1_outputs(7957) <= '0';
    layer1_outputs(7958) <= b;
    layer1_outputs(7959) <= not b or a;
    layer1_outputs(7960) <= not (a and b);
    layer1_outputs(7961) <= a and not b;
    layer1_outputs(7962) <= '0';
    layer1_outputs(7963) <= b;
    layer1_outputs(7964) <= not b;
    layer1_outputs(7965) <= '0';
    layer1_outputs(7966) <= a or b;
    layer1_outputs(7967) <= not b or a;
    layer1_outputs(7968) <= b;
    layer1_outputs(7969) <= a and not b;
    layer1_outputs(7970) <= a and b;
    layer1_outputs(7971) <= a and not b;
    layer1_outputs(7972) <= a or b;
    layer1_outputs(7973) <= '1';
    layer1_outputs(7974) <= not (a and b);
    layer1_outputs(7975) <= '1';
    layer1_outputs(7976) <= a and b;
    layer1_outputs(7977) <= not b or a;
    layer1_outputs(7978) <= a and not b;
    layer1_outputs(7979) <= b;
    layer1_outputs(7980) <= '0';
    layer1_outputs(7981) <= not a or b;
    layer1_outputs(7982) <= not a;
    layer1_outputs(7983) <= a and b;
    layer1_outputs(7984) <= not (a and b);
    layer1_outputs(7985) <= a and b;
    layer1_outputs(7986) <= a;
    layer1_outputs(7987) <= b;
    layer1_outputs(7988) <= '0';
    layer1_outputs(7989) <= not a or b;
    layer1_outputs(7990) <= not a;
    layer1_outputs(7991) <= not b or a;
    layer1_outputs(7992) <= b;
    layer1_outputs(7993) <= a;
    layer1_outputs(7994) <= not (a xor b);
    layer1_outputs(7995) <= b and not a;
    layer1_outputs(7996) <= not b or a;
    layer1_outputs(7997) <= a and not b;
    layer1_outputs(7998) <= b;
    layer1_outputs(7999) <= a and b;
    layer1_outputs(8000) <= '0';
    layer1_outputs(8001) <= b;
    layer1_outputs(8002) <= not a;
    layer1_outputs(8003) <= not a or b;
    layer1_outputs(8004) <= not b or a;
    layer1_outputs(8005) <= a;
    layer1_outputs(8006) <= b;
    layer1_outputs(8007) <= not (a and b);
    layer1_outputs(8008) <= not (a xor b);
    layer1_outputs(8009) <= not a;
    layer1_outputs(8010) <= '1';
    layer1_outputs(8011) <= not b;
    layer1_outputs(8012) <= b and not a;
    layer1_outputs(8013) <= a and not b;
    layer1_outputs(8014) <= '1';
    layer1_outputs(8015) <= a and b;
    layer1_outputs(8016) <= a;
    layer1_outputs(8017) <= a and not b;
    layer1_outputs(8018) <= b;
    layer1_outputs(8019) <= b;
    layer1_outputs(8020) <= a or b;
    layer1_outputs(8021) <= '1';
    layer1_outputs(8022) <= not (a and b);
    layer1_outputs(8023) <= not b or a;
    layer1_outputs(8024) <= not a or b;
    layer1_outputs(8025) <= '1';
    layer1_outputs(8026) <= a;
    layer1_outputs(8027) <= a and b;
    layer1_outputs(8028) <= not a;
    layer1_outputs(8029) <= a;
    layer1_outputs(8030) <= b and not a;
    layer1_outputs(8031) <= a or b;
    layer1_outputs(8032) <= not a or b;
    layer1_outputs(8033) <= a and not b;
    layer1_outputs(8034) <= b and not a;
    layer1_outputs(8035) <= b;
    layer1_outputs(8036) <= not (a or b);
    layer1_outputs(8037) <= not (a and b);
    layer1_outputs(8038) <= not (a xor b);
    layer1_outputs(8039) <= not (a or b);
    layer1_outputs(8040) <= a and not b;
    layer1_outputs(8041) <= not a;
    layer1_outputs(8042) <= not a or b;
    layer1_outputs(8043) <= not (a xor b);
    layer1_outputs(8044) <= a and b;
    layer1_outputs(8045) <= b;
    layer1_outputs(8046) <= '1';
    layer1_outputs(8047) <= b;
    layer1_outputs(8048) <= a;
    layer1_outputs(8049) <= a or b;
    layer1_outputs(8050) <= a and b;
    layer1_outputs(8051) <= not (a or b);
    layer1_outputs(8052) <= a xor b;
    layer1_outputs(8053) <= not a or b;
    layer1_outputs(8054) <= a or b;
    layer1_outputs(8055) <= not a;
    layer1_outputs(8056) <= a or b;
    layer1_outputs(8057) <= not a or b;
    layer1_outputs(8058) <= not (a or b);
    layer1_outputs(8059) <= b;
    layer1_outputs(8060) <= a;
    layer1_outputs(8061) <= not a;
    layer1_outputs(8062) <= not a or b;
    layer1_outputs(8063) <= a or b;
    layer1_outputs(8064) <= not b;
    layer1_outputs(8065) <= not a or b;
    layer1_outputs(8066) <= '0';
    layer1_outputs(8067) <= b and not a;
    layer1_outputs(8068) <= not (a or b);
    layer1_outputs(8069) <= a;
    layer1_outputs(8070) <= a;
    layer1_outputs(8071) <= '1';
    layer1_outputs(8072) <= not b;
    layer1_outputs(8073) <= not a or b;
    layer1_outputs(8074) <= not a;
    layer1_outputs(8075) <= a and not b;
    layer1_outputs(8076) <= a and b;
    layer1_outputs(8077) <= b and not a;
    layer1_outputs(8078) <= b;
    layer1_outputs(8079) <= not (a and b);
    layer1_outputs(8080) <= not b or a;
    layer1_outputs(8081) <= not a or b;
    layer1_outputs(8082) <= b and not a;
    layer1_outputs(8083) <= a xor b;
    layer1_outputs(8084) <= not b or a;
    layer1_outputs(8085) <= not a or b;
    layer1_outputs(8086) <= not b;
    layer1_outputs(8087) <= b and not a;
    layer1_outputs(8088) <= b;
    layer1_outputs(8089) <= a and not b;
    layer1_outputs(8090) <= a;
    layer1_outputs(8091) <= not (a xor b);
    layer1_outputs(8092) <= not (a and b);
    layer1_outputs(8093) <= not a or b;
    layer1_outputs(8094) <= not a;
    layer1_outputs(8095) <= not (a or b);
    layer1_outputs(8096) <= a and b;
    layer1_outputs(8097) <= not (a and b);
    layer1_outputs(8098) <= b and not a;
    layer1_outputs(8099) <= a and not b;
    layer1_outputs(8100) <= not (a and b);
    layer1_outputs(8101) <= not (a and b);
    layer1_outputs(8102) <= not b;
    layer1_outputs(8103) <= not (a and b);
    layer1_outputs(8104) <= not b;
    layer1_outputs(8105) <= '1';
    layer1_outputs(8106) <= b;
    layer1_outputs(8107) <= b and not a;
    layer1_outputs(8108) <= a and not b;
    layer1_outputs(8109) <= a and not b;
    layer1_outputs(8110) <= a or b;
    layer1_outputs(8111) <= a xor b;
    layer1_outputs(8112) <= a and b;
    layer1_outputs(8113) <= not (a xor b);
    layer1_outputs(8114) <= b;
    layer1_outputs(8115) <= not a or b;
    layer1_outputs(8116) <= a and not b;
    layer1_outputs(8117) <= not (a xor b);
    layer1_outputs(8118) <= not (a and b);
    layer1_outputs(8119) <= b and not a;
    layer1_outputs(8120) <= not b;
    layer1_outputs(8121) <= a or b;
    layer1_outputs(8122) <= a and b;
    layer1_outputs(8123) <= a xor b;
    layer1_outputs(8124) <= not b;
    layer1_outputs(8125) <= not a or b;
    layer1_outputs(8126) <= not b or a;
    layer1_outputs(8127) <= '0';
    layer1_outputs(8128) <= not a or b;
    layer1_outputs(8129) <= a and b;
    layer1_outputs(8130) <= not (a or b);
    layer1_outputs(8131) <= '0';
    layer1_outputs(8132) <= a xor b;
    layer1_outputs(8133) <= b;
    layer1_outputs(8134) <= a and not b;
    layer1_outputs(8135) <= not a or b;
    layer1_outputs(8136) <= a or b;
    layer1_outputs(8137) <= not b;
    layer1_outputs(8138) <= not b or a;
    layer1_outputs(8139) <= not b or a;
    layer1_outputs(8140) <= not b;
    layer1_outputs(8141) <= not b or a;
    layer1_outputs(8142) <= not (a or b);
    layer1_outputs(8143) <= not (a and b);
    layer1_outputs(8144) <= b;
    layer1_outputs(8145) <= not b or a;
    layer1_outputs(8146) <= b and not a;
    layer1_outputs(8147) <= not a or b;
    layer1_outputs(8148) <= '0';
    layer1_outputs(8149) <= '0';
    layer1_outputs(8150) <= not a;
    layer1_outputs(8151) <= a and b;
    layer1_outputs(8152) <= b and not a;
    layer1_outputs(8153) <= a or b;
    layer1_outputs(8154) <= b;
    layer1_outputs(8155) <= not b or a;
    layer1_outputs(8156) <= not b or a;
    layer1_outputs(8157) <= a;
    layer1_outputs(8158) <= a and not b;
    layer1_outputs(8159) <= not (a or b);
    layer1_outputs(8160) <= a and b;
    layer1_outputs(8161) <= b and not a;
    layer1_outputs(8162) <= not (a or b);
    layer1_outputs(8163) <= '1';
    layer1_outputs(8164) <= '0';
    layer1_outputs(8165) <= not (a and b);
    layer1_outputs(8166) <= a and b;
    layer1_outputs(8167) <= not b or a;
    layer1_outputs(8168) <= b;
    layer1_outputs(8169) <= not (a xor b);
    layer1_outputs(8170) <= not b;
    layer1_outputs(8171) <= a and b;
    layer1_outputs(8172) <= a and not b;
    layer1_outputs(8173) <= b;
    layer1_outputs(8174) <= b and not a;
    layer1_outputs(8175) <= not b;
    layer1_outputs(8176) <= '0';
    layer1_outputs(8177) <= a or b;
    layer1_outputs(8178) <= b;
    layer1_outputs(8179) <= a and not b;
    layer1_outputs(8180) <= not b or a;
    layer1_outputs(8181) <= b;
    layer1_outputs(8182) <= not b;
    layer1_outputs(8183) <= a and b;
    layer1_outputs(8184) <= not a or b;
    layer1_outputs(8185) <= a or b;
    layer1_outputs(8186) <= b;
    layer1_outputs(8187) <= a;
    layer1_outputs(8188) <= not b;
    layer1_outputs(8189) <= '0';
    layer1_outputs(8190) <= a and b;
    layer1_outputs(8191) <= not b or a;
    layer1_outputs(8192) <= not b;
    layer1_outputs(8193) <= b and not a;
    layer1_outputs(8194) <= not a or b;
    layer1_outputs(8195) <= not a;
    layer1_outputs(8196) <= '1';
    layer1_outputs(8197) <= not a;
    layer1_outputs(8198) <= not a;
    layer1_outputs(8199) <= '1';
    layer1_outputs(8200) <= not (a or b);
    layer1_outputs(8201) <= not b or a;
    layer1_outputs(8202) <= '0';
    layer1_outputs(8203) <= '0';
    layer1_outputs(8204) <= not a or b;
    layer1_outputs(8205) <= not (a xor b);
    layer1_outputs(8206) <= not b;
    layer1_outputs(8207) <= '1';
    layer1_outputs(8208) <= a or b;
    layer1_outputs(8209) <= not b or a;
    layer1_outputs(8210) <= a or b;
    layer1_outputs(8211) <= a;
    layer1_outputs(8212) <= not a or b;
    layer1_outputs(8213) <= not (a and b);
    layer1_outputs(8214) <= b;
    layer1_outputs(8215) <= b and not a;
    layer1_outputs(8216) <= not b or a;
    layer1_outputs(8217) <= not b;
    layer1_outputs(8218) <= a xor b;
    layer1_outputs(8219) <= a;
    layer1_outputs(8220) <= b;
    layer1_outputs(8221) <= a;
    layer1_outputs(8222) <= not (a or b);
    layer1_outputs(8223) <= not b;
    layer1_outputs(8224) <= a;
    layer1_outputs(8225) <= '1';
    layer1_outputs(8226) <= '0';
    layer1_outputs(8227) <= not (a or b);
    layer1_outputs(8228) <= not b;
    layer1_outputs(8229) <= not (a xor b);
    layer1_outputs(8230) <= a and b;
    layer1_outputs(8231) <= not (a or b);
    layer1_outputs(8232) <= not b;
    layer1_outputs(8233) <= a and not b;
    layer1_outputs(8234) <= b;
    layer1_outputs(8235) <= not b or a;
    layer1_outputs(8236) <= a and not b;
    layer1_outputs(8237) <= not b;
    layer1_outputs(8238) <= not (a xor b);
    layer1_outputs(8239) <= not a;
    layer1_outputs(8240) <= not b;
    layer1_outputs(8241) <= b;
    layer1_outputs(8242) <= not a or b;
    layer1_outputs(8243) <= not b or a;
    layer1_outputs(8244) <= not a;
    layer1_outputs(8245) <= not b or a;
    layer1_outputs(8246) <= not b;
    layer1_outputs(8247) <= not (a or b);
    layer1_outputs(8248) <= not b or a;
    layer1_outputs(8249) <= not a;
    layer1_outputs(8250) <= not (a xor b);
    layer1_outputs(8251) <= a xor b;
    layer1_outputs(8252) <= not (a xor b);
    layer1_outputs(8253) <= not b;
    layer1_outputs(8254) <= a and not b;
    layer1_outputs(8255) <= a and not b;
    layer1_outputs(8256) <= a;
    layer1_outputs(8257) <= a;
    layer1_outputs(8258) <= a and b;
    layer1_outputs(8259) <= not a or b;
    layer1_outputs(8260) <= not b;
    layer1_outputs(8261) <= not b;
    layer1_outputs(8262) <= not b or a;
    layer1_outputs(8263) <= a and b;
    layer1_outputs(8264) <= not b or a;
    layer1_outputs(8265) <= a and b;
    layer1_outputs(8266) <= '0';
    layer1_outputs(8267) <= a and b;
    layer1_outputs(8268) <= a and b;
    layer1_outputs(8269) <= not (a or b);
    layer1_outputs(8270) <= '0';
    layer1_outputs(8271) <= b;
    layer1_outputs(8272) <= b and not a;
    layer1_outputs(8273) <= '1';
    layer1_outputs(8274) <= not b or a;
    layer1_outputs(8275) <= a or b;
    layer1_outputs(8276) <= a and not b;
    layer1_outputs(8277) <= not a;
    layer1_outputs(8278) <= b and not a;
    layer1_outputs(8279) <= not (a and b);
    layer1_outputs(8280) <= a or b;
    layer1_outputs(8281) <= not a;
    layer1_outputs(8282) <= not (a and b);
    layer1_outputs(8283) <= a;
    layer1_outputs(8284) <= not (a or b);
    layer1_outputs(8285) <= not (a and b);
    layer1_outputs(8286) <= a and not b;
    layer1_outputs(8287) <= '1';
    layer1_outputs(8288) <= b;
    layer1_outputs(8289) <= not b or a;
    layer1_outputs(8290) <= not (a and b);
    layer1_outputs(8291) <= not a or b;
    layer1_outputs(8292) <= not b or a;
    layer1_outputs(8293) <= not (a and b);
    layer1_outputs(8294) <= not (a and b);
    layer1_outputs(8295) <= '1';
    layer1_outputs(8296) <= not a;
    layer1_outputs(8297) <= a;
    layer1_outputs(8298) <= '0';
    layer1_outputs(8299) <= not a;
    layer1_outputs(8300) <= not b or a;
    layer1_outputs(8301) <= b and not a;
    layer1_outputs(8302) <= a and not b;
    layer1_outputs(8303) <= not a;
    layer1_outputs(8304) <= a and not b;
    layer1_outputs(8305) <= not b or a;
    layer1_outputs(8306) <= a and b;
    layer1_outputs(8307) <= not (a and b);
    layer1_outputs(8308) <= not b or a;
    layer1_outputs(8309) <= not a or b;
    layer1_outputs(8310) <= a or b;
    layer1_outputs(8311) <= '1';
    layer1_outputs(8312) <= a and b;
    layer1_outputs(8313) <= not (a or b);
    layer1_outputs(8314) <= not (a xor b);
    layer1_outputs(8315) <= a and b;
    layer1_outputs(8316) <= a and not b;
    layer1_outputs(8317) <= not a;
    layer1_outputs(8318) <= b;
    layer1_outputs(8319) <= '0';
    layer1_outputs(8320) <= '0';
    layer1_outputs(8321) <= not (a xor b);
    layer1_outputs(8322) <= b;
    layer1_outputs(8323) <= '0';
    layer1_outputs(8324) <= a;
    layer1_outputs(8325) <= not b;
    layer1_outputs(8326) <= a;
    layer1_outputs(8327) <= a;
    layer1_outputs(8328) <= not (a and b);
    layer1_outputs(8329) <= not a or b;
    layer1_outputs(8330) <= '0';
    layer1_outputs(8331) <= b;
    layer1_outputs(8332) <= not b;
    layer1_outputs(8333) <= not (a and b);
    layer1_outputs(8334) <= a;
    layer1_outputs(8335) <= not (a and b);
    layer1_outputs(8336) <= not (a or b);
    layer1_outputs(8337) <= not (a or b);
    layer1_outputs(8338) <= a and b;
    layer1_outputs(8339) <= b and not a;
    layer1_outputs(8340) <= '0';
    layer1_outputs(8341) <= '0';
    layer1_outputs(8342) <= a;
    layer1_outputs(8343) <= a and b;
    layer1_outputs(8344) <= a;
    layer1_outputs(8345) <= b;
    layer1_outputs(8346) <= a and b;
    layer1_outputs(8347) <= '1';
    layer1_outputs(8348) <= '1';
    layer1_outputs(8349) <= not a or b;
    layer1_outputs(8350) <= not b;
    layer1_outputs(8351) <= not (a and b);
    layer1_outputs(8352) <= a;
    layer1_outputs(8353) <= b;
    layer1_outputs(8354) <= a and not b;
    layer1_outputs(8355) <= a xor b;
    layer1_outputs(8356) <= a;
    layer1_outputs(8357) <= not a or b;
    layer1_outputs(8358) <= a or b;
    layer1_outputs(8359) <= a and b;
    layer1_outputs(8360) <= not b;
    layer1_outputs(8361) <= not (a xor b);
    layer1_outputs(8362) <= b;
    layer1_outputs(8363) <= a and not b;
    layer1_outputs(8364) <= b;
    layer1_outputs(8365) <= a and b;
    layer1_outputs(8366) <= '0';
    layer1_outputs(8367) <= a and not b;
    layer1_outputs(8368) <= not a or b;
    layer1_outputs(8369) <= not b or a;
    layer1_outputs(8370) <= a or b;
    layer1_outputs(8371) <= '1';
    layer1_outputs(8372) <= not b or a;
    layer1_outputs(8373) <= b;
    layer1_outputs(8374) <= not (a and b);
    layer1_outputs(8375) <= not a or b;
    layer1_outputs(8376) <= '0';
    layer1_outputs(8377) <= not (a and b);
    layer1_outputs(8378) <= not a;
    layer1_outputs(8379) <= not b;
    layer1_outputs(8380) <= b;
    layer1_outputs(8381) <= a and not b;
    layer1_outputs(8382) <= a xor b;
    layer1_outputs(8383) <= not b or a;
    layer1_outputs(8384) <= '1';
    layer1_outputs(8385) <= a or b;
    layer1_outputs(8386) <= b and not a;
    layer1_outputs(8387) <= not a;
    layer1_outputs(8388) <= not a or b;
    layer1_outputs(8389) <= not (a xor b);
    layer1_outputs(8390) <= not a;
    layer1_outputs(8391) <= b;
    layer1_outputs(8392) <= a and b;
    layer1_outputs(8393) <= b and not a;
    layer1_outputs(8394) <= not (a and b);
    layer1_outputs(8395) <= a or b;
    layer1_outputs(8396) <= '1';
    layer1_outputs(8397) <= '1';
    layer1_outputs(8398) <= a and not b;
    layer1_outputs(8399) <= not a;
    layer1_outputs(8400) <= not a or b;
    layer1_outputs(8401) <= not (a and b);
    layer1_outputs(8402) <= '1';
    layer1_outputs(8403) <= not a or b;
    layer1_outputs(8404) <= a and not b;
    layer1_outputs(8405) <= a and not b;
    layer1_outputs(8406) <= a and b;
    layer1_outputs(8407) <= a;
    layer1_outputs(8408) <= not a;
    layer1_outputs(8409) <= a;
    layer1_outputs(8410) <= b and not a;
    layer1_outputs(8411) <= a and not b;
    layer1_outputs(8412) <= a or b;
    layer1_outputs(8413) <= b and not a;
    layer1_outputs(8414) <= not b;
    layer1_outputs(8415) <= a and not b;
    layer1_outputs(8416) <= a;
    layer1_outputs(8417) <= a or b;
    layer1_outputs(8418) <= a and b;
    layer1_outputs(8419) <= not b or a;
    layer1_outputs(8420) <= not (a and b);
    layer1_outputs(8421) <= not b;
    layer1_outputs(8422) <= b and not a;
    layer1_outputs(8423) <= '1';
    layer1_outputs(8424) <= b;
    layer1_outputs(8425) <= not (a and b);
    layer1_outputs(8426) <= a and b;
    layer1_outputs(8427) <= not (a or b);
    layer1_outputs(8428) <= b;
    layer1_outputs(8429) <= b and not a;
    layer1_outputs(8430) <= '1';
    layer1_outputs(8431) <= a and b;
    layer1_outputs(8432) <= not (a xor b);
    layer1_outputs(8433) <= '1';
    layer1_outputs(8434) <= '1';
    layer1_outputs(8435) <= '0';
    layer1_outputs(8436) <= a and b;
    layer1_outputs(8437) <= a and b;
    layer1_outputs(8438) <= not a or b;
    layer1_outputs(8439) <= b and not a;
    layer1_outputs(8440) <= not b or a;
    layer1_outputs(8441) <= not (a and b);
    layer1_outputs(8442) <= b;
    layer1_outputs(8443) <= not (a or b);
    layer1_outputs(8444) <= a and b;
    layer1_outputs(8445) <= not a or b;
    layer1_outputs(8446) <= not a;
    layer1_outputs(8447) <= '0';
    layer1_outputs(8448) <= not (a or b);
    layer1_outputs(8449) <= not a or b;
    layer1_outputs(8450) <= '1';
    layer1_outputs(8451) <= not b;
    layer1_outputs(8452) <= a and not b;
    layer1_outputs(8453) <= b and not a;
    layer1_outputs(8454) <= not a or b;
    layer1_outputs(8455) <= b and not a;
    layer1_outputs(8456) <= not a;
    layer1_outputs(8457) <= not (a and b);
    layer1_outputs(8458) <= '0';
    layer1_outputs(8459) <= not (a or b);
    layer1_outputs(8460) <= b and not a;
    layer1_outputs(8461) <= not (a and b);
    layer1_outputs(8462) <= not b;
    layer1_outputs(8463) <= not b;
    layer1_outputs(8464) <= a;
    layer1_outputs(8465) <= not (a and b);
    layer1_outputs(8466) <= '0';
    layer1_outputs(8467) <= not a or b;
    layer1_outputs(8468) <= a xor b;
    layer1_outputs(8469) <= not b;
    layer1_outputs(8470) <= b;
    layer1_outputs(8471) <= a;
    layer1_outputs(8472) <= not a or b;
    layer1_outputs(8473) <= a and not b;
    layer1_outputs(8474) <= a or b;
    layer1_outputs(8475) <= not (a or b);
    layer1_outputs(8476) <= a and b;
    layer1_outputs(8477) <= '0';
    layer1_outputs(8478) <= not b;
    layer1_outputs(8479) <= not a;
    layer1_outputs(8480) <= not (a xor b);
    layer1_outputs(8481) <= '0';
    layer1_outputs(8482) <= a;
    layer1_outputs(8483) <= '0';
    layer1_outputs(8484) <= b and not a;
    layer1_outputs(8485) <= not b or a;
    layer1_outputs(8486) <= b and not a;
    layer1_outputs(8487) <= not (a or b);
    layer1_outputs(8488) <= not a;
    layer1_outputs(8489) <= not b or a;
    layer1_outputs(8490) <= '0';
    layer1_outputs(8491) <= b;
    layer1_outputs(8492) <= a and b;
    layer1_outputs(8493) <= a and not b;
    layer1_outputs(8494) <= not (a and b);
    layer1_outputs(8495) <= not (a and b);
    layer1_outputs(8496) <= not a;
    layer1_outputs(8497) <= '0';
    layer1_outputs(8498) <= not b;
    layer1_outputs(8499) <= '0';
    layer1_outputs(8500) <= not a or b;
    layer1_outputs(8501) <= not b or a;
    layer1_outputs(8502) <= a;
    layer1_outputs(8503) <= a xor b;
    layer1_outputs(8504) <= a and b;
    layer1_outputs(8505) <= not (a xor b);
    layer1_outputs(8506) <= b;
    layer1_outputs(8507) <= not a;
    layer1_outputs(8508) <= b;
    layer1_outputs(8509) <= not b;
    layer1_outputs(8510) <= not a;
    layer1_outputs(8511) <= '1';
    layer1_outputs(8512) <= a xor b;
    layer1_outputs(8513) <= b;
    layer1_outputs(8514) <= a or b;
    layer1_outputs(8515) <= a and b;
    layer1_outputs(8516) <= b and not a;
    layer1_outputs(8517) <= a xor b;
    layer1_outputs(8518) <= '1';
    layer1_outputs(8519) <= a and b;
    layer1_outputs(8520) <= not (a and b);
    layer1_outputs(8521) <= a or b;
    layer1_outputs(8522) <= not a or b;
    layer1_outputs(8523) <= b and not a;
    layer1_outputs(8524) <= not b or a;
    layer1_outputs(8525) <= '1';
    layer1_outputs(8526) <= b;
    layer1_outputs(8527) <= b;
    layer1_outputs(8528) <= b and not a;
    layer1_outputs(8529) <= b;
    layer1_outputs(8530) <= '0';
    layer1_outputs(8531) <= not a;
    layer1_outputs(8532) <= not a or b;
    layer1_outputs(8533) <= b and not a;
    layer1_outputs(8534) <= not (a and b);
    layer1_outputs(8535) <= a xor b;
    layer1_outputs(8536) <= not a;
    layer1_outputs(8537) <= a and not b;
    layer1_outputs(8538) <= a;
    layer1_outputs(8539) <= not a;
    layer1_outputs(8540) <= not b or a;
    layer1_outputs(8541) <= a and b;
    layer1_outputs(8542) <= a or b;
    layer1_outputs(8543) <= not a;
    layer1_outputs(8544) <= a;
    layer1_outputs(8545) <= '0';
    layer1_outputs(8546) <= '0';
    layer1_outputs(8547) <= a and b;
    layer1_outputs(8548) <= '1';
    layer1_outputs(8549) <= not (a or b);
    layer1_outputs(8550) <= a and b;
    layer1_outputs(8551) <= not a;
    layer1_outputs(8552) <= not a or b;
    layer1_outputs(8553) <= '0';
    layer1_outputs(8554) <= '0';
    layer1_outputs(8555) <= b;
    layer1_outputs(8556) <= a and not b;
    layer1_outputs(8557) <= not b or a;
    layer1_outputs(8558) <= a xor b;
    layer1_outputs(8559) <= b;
    layer1_outputs(8560) <= b;
    layer1_outputs(8561) <= not a or b;
    layer1_outputs(8562) <= a and not b;
    layer1_outputs(8563) <= not (a xor b);
    layer1_outputs(8564) <= not a or b;
    layer1_outputs(8565) <= b and not a;
    layer1_outputs(8566) <= b;
    layer1_outputs(8567) <= not (a or b);
    layer1_outputs(8568) <= not b or a;
    layer1_outputs(8569) <= not (a and b);
    layer1_outputs(8570) <= b and not a;
    layer1_outputs(8571) <= '1';
    layer1_outputs(8572) <= a xor b;
    layer1_outputs(8573) <= a;
    layer1_outputs(8574) <= a or b;
    layer1_outputs(8575) <= not b;
    layer1_outputs(8576) <= a and not b;
    layer1_outputs(8577) <= a and not b;
    layer1_outputs(8578) <= not (a and b);
    layer1_outputs(8579) <= not a or b;
    layer1_outputs(8580) <= not (a or b);
    layer1_outputs(8581) <= not a;
    layer1_outputs(8582) <= not a;
    layer1_outputs(8583) <= not (a and b);
    layer1_outputs(8584) <= not (a and b);
    layer1_outputs(8585) <= not (a or b);
    layer1_outputs(8586) <= a;
    layer1_outputs(8587) <= not b;
    layer1_outputs(8588) <= a xor b;
    layer1_outputs(8589) <= not (a or b);
    layer1_outputs(8590) <= a or b;
    layer1_outputs(8591) <= not (a and b);
    layer1_outputs(8592) <= not b;
    layer1_outputs(8593) <= '1';
    layer1_outputs(8594) <= a;
    layer1_outputs(8595) <= a and not b;
    layer1_outputs(8596) <= a and not b;
    layer1_outputs(8597) <= not (a or b);
    layer1_outputs(8598) <= b and not a;
    layer1_outputs(8599) <= a and b;
    layer1_outputs(8600) <= not b or a;
    layer1_outputs(8601) <= not b or a;
    layer1_outputs(8602) <= not a;
    layer1_outputs(8603) <= '0';
    layer1_outputs(8604) <= b;
    layer1_outputs(8605) <= a and not b;
    layer1_outputs(8606) <= a and b;
    layer1_outputs(8607) <= a and not b;
    layer1_outputs(8608) <= a or b;
    layer1_outputs(8609) <= a and b;
    layer1_outputs(8610) <= '1';
    layer1_outputs(8611) <= b and not a;
    layer1_outputs(8612) <= a and b;
    layer1_outputs(8613) <= a or b;
    layer1_outputs(8614) <= not a or b;
    layer1_outputs(8615) <= not (a and b);
    layer1_outputs(8616) <= not b or a;
    layer1_outputs(8617) <= not a;
    layer1_outputs(8618) <= b and not a;
    layer1_outputs(8619) <= not a;
    layer1_outputs(8620) <= not a;
    layer1_outputs(8621) <= '0';
    layer1_outputs(8622) <= a and not b;
    layer1_outputs(8623) <= '1';
    layer1_outputs(8624) <= not (a xor b);
    layer1_outputs(8625) <= '0';
    layer1_outputs(8626) <= a xor b;
    layer1_outputs(8627) <= not a or b;
    layer1_outputs(8628) <= b;
    layer1_outputs(8629) <= b;
    layer1_outputs(8630) <= a or b;
    layer1_outputs(8631) <= not (a and b);
    layer1_outputs(8632) <= a and b;
    layer1_outputs(8633) <= not a or b;
    layer1_outputs(8634) <= not a;
    layer1_outputs(8635) <= b and not a;
    layer1_outputs(8636) <= '1';
    layer1_outputs(8637) <= a and b;
    layer1_outputs(8638) <= a;
    layer1_outputs(8639) <= a and b;
    layer1_outputs(8640) <= not a;
    layer1_outputs(8641) <= '0';
    layer1_outputs(8642) <= not b or a;
    layer1_outputs(8643) <= not b;
    layer1_outputs(8644) <= a and b;
    layer1_outputs(8645) <= not b or a;
    layer1_outputs(8646) <= not b;
    layer1_outputs(8647) <= not a or b;
    layer1_outputs(8648) <= a;
    layer1_outputs(8649) <= a;
    layer1_outputs(8650) <= not a or b;
    layer1_outputs(8651) <= '0';
    layer1_outputs(8652) <= not b;
    layer1_outputs(8653) <= '0';
    layer1_outputs(8654) <= a;
    layer1_outputs(8655) <= not b or a;
    layer1_outputs(8656) <= a and not b;
    layer1_outputs(8657) <= a xor b;
    layer1_outputs(8658) <= not b;
    layer1_outputs(8659) <= not a;
    layer1_outputs(8660) <= a and not b;
    layer1_outputs(8661) <= not a;
    layer1_outputs(8662) <= not (a and b);
    layer1_outputs(8663) <= b and not a;
    layer1_outputs(8664) <= b and not a;
    layer1_outputs(8665) <= a;
    layer1_outputs(8666) <= not b;
    layer1_outputs(8667) <= not (a or b);
    layer1_outputs(8668) <= '0';
    layer1_outputs(8669) <= not b;
    layer1_outputs(8670) <= not a or b;
    layer1_outputs(8671) <= not a;
    layer1_outputs(8672) <= b and not a;
    layer1_outputs(8673) <= not a;
    layer1_outputs(8674) <= a and not b;
    layer1_outputs(8675) <= a;
    layer1_outputs(8676) <= not (a and b);
    layer1_outputs(8677) <= a and b;
    layer1_outputs(8678) <= '1';
    layer1_outputs(8679) <= b and not a;
    layer1_outputs(8680) <= not (a or b);
    layer1_outputs(8681) <= a xor b;
    layer1_outputs(8682) <= not b;
    layer1_outputs(8683) <= b and not a;
    layer1_outputs(8684) <= a or b;
    layer1_outputs(8685) <= not a;
    layer1_outputs(8686) <= a or b;
    layer1_outputs(8687) <= not a;
    layer1_outputs(8688) <= '0';
    layer1_outputs(8689) <= a and b;
    layer1_outputs(8690) <= '1';
    layer1_outputs(8691) <= a or b;
    layer1_outputs(8692) <= not b;
    layer1_outputs(8693) <= b and not a;
    layer1_outputs(8694) <= not (a xor b);
    layer1_outputs(8695) <= '1';
    layer1_outputs(8696) <= not (a xor b);
    layer1_outputs(8697) <= not (a and b);
    layer1_outputs(8698) <= b and not a;
    layer1_outputs(8699) <= not b or a;
    layer1_outputs(8700) <= not b;
    layer1_outputs(8701) <= a or b;
    layer1_outputs(8702) <= not a;
    layer1_outputs(8703) <= not (a xor b);
    layer1_outputs(8704) <= '0';
    layer1_outputs(8705) <= a and b;
    layer1_outputs(8706) <= b;
    layer1_outputs(8707) <= a and not b;
    layer1_outputs(8708) <= not a;
    layer1_outputs(8709) <= '0';
    layer1_outputs(8710) <= '1';
    layer1_outputs(8711) <= not (a and b);
    layer1_outputs(8712) <= not (a and b);
    layer1_outputs(8713) <= b;
    layer1_outputs(8714) <= not (a and b);
    layer1_outputs(8715) <= a or b;
    layer1_outputs(8716) <= not (a and b);
    layer1_outputs(8717) <= not (a and b);
    layer1_outputs(8718) <= not b or a;
    layer1_outputs(8719) <= '1';
    layer1_outputs(8720) <= '1';
    layer1_outputs(8721) <= a;
    layer1_outputs(8722) <= not a or b;
    layer1_outputs(8723) <= a and not b;
    layer1_outputs(8724) <= '0';
    layer1_outputs(8725) <= a or b;
    layer1_outputs(8726) <= not (a xor b);
    layer1_outputs(8727) <= '1';
    layer1_outputs(8728) <= not (a and b);
    layer1_outputs(8729) <= a and b;
    layer1_outputs(8730) <= b and not a;
    layer1_outputs(8731) <= a or b;
    layer1_outputs(8732) <= '1';
    layer1_outputs(8733) <= not b;
    layer1_outputs(8734) <= '0';
    layer1_outputs(8735) <= b;
    layer1_outputs(8736) <= not a;
    layer1_outputs(8737) <= b and not a;
    layer1_outputs(8738) <= not (a and b);
    layer1_outputs(8739) <= '1';
    layer1_outputs(8740) <= not (a or b);
    layer1_outputs(8741) <= a and not b;
    layer1_outputs(8742) <= a;
    layer1_outputs(8743) <= not (a and b);
    layer1_outputs(8744) <= not b;
    layer1_outputs(8745) <= a or b;
    layer1_outputs(8746) <= '0';
    layer1_outputs(8747) <= not (a xor b);
    layer1_outputs(8748) <= a and not b;
    layer1_outputs(8749) <= not (a xor b);
    layer1_outputs(8750) <= not b or a;
    layer1_outputs(8751) <= a and b;
    layer1_outputs(8752) <= not b or a;
    layer1_outputs(8753) <= '1';
    layer1_outputs(8754) <= not a;
    layer1_outputs(8755) <= '1';
    layer1_outputs(8756) <= a xor b;
    layer1_outputs(8757) <= '0';
    layer1_outputs(8758) <= not (a xor b);
    layer1_outputs(8759) <= '1';
    layer1_outputs(8760) <= a xor b;
    layer1_outputs(8761) <= not a;
    layer1_outputs(8762) <= a xor b;
    layer1_outputs(8763) <= b and not a;
    layer1_outputs(8764) <= b;
    layer1_outputs(8765) <= b;
    layer1_outputs(8766) <= b and not a;
    layer1_outputs(8767) <= not (a and b);
    layer1_outputs(8768) <= a and b;
    layer1_outputs(8769) <= not a;
    layer1_outputs(8770) <= not (a or b);
    layer1_outputs(8771) <= a and b;
    layer1_outputs(8772) <= not (a and b);
    layer1_outputs(8773) <= not (a and b);
    layer1_outputs(8774) <= not b or a;
    layer1_outputs(8775) <= '0';
    layer1_outputs(8776) <= a and b;
    layer1_outputs(8777) <= b and not a;
    layer1_outputs(8778) <= not (a and b);
    layer1_outputs(8779) <= a xor b;
    layer1_outputs(8780) <= b;
    layer1_outputs(8781) <= not a or b;
    layer1_outputs(8782) <= '1';
    layer1_outputs(8783) <= a xor b;
    layer1_outputs(8784) <= not b;
    layer1_outputs(8785) <= not a;
    layer1_outputs(8786) <= a or b;
    layer1_outputs(8787) <= not (a and b);
    layer1_outputs(8788) <= not (a and b);
    layer1_outputs(8789) <= not b or a;
    layer1_outputs(8790) <= a and not b;
    layer1_outputs(8791) <= a;
    layer1_outputs(8792) <= not (a and b);
    layer1_outputs(8793) <= a or b;
    layer1_outputs(8794) <= not (a or b);
    layer1_outputs(8795) <= not (a or b);
    layer1_outputs(8796) <= not b;
    layer1_outputs(8797) <= a xor b;
    layer1_outputs(8798) <= not (a xor b);
    layer1_outputs(8799) <= a and not b;
    layer1_outputs(8800) <= not (a or b);
    layer1_outputs(8801) <= '0';
    layer1_outputs(8802) <= not a;
    layer1_outputs(8803) <= not a;
    layer1_outputs(8804) <= not b;
    layer1_outputs(8805) <= a and not b;
    layer1_outputs(8806) <= b;
    layer1_outputs(8807) <= not b;
    layer1_outputs(8808) <= not (a or b);
    layer1_outputs(8809) <= not a or b;
    layer1_outputs(8810) <= not b;
    layer1_outputs(8811) <= not b;
    layer1_outputs(8812) <= b and not a;
    layer1_outputs(8813) <= '0';
    layer1_outputs(8814) <= a and b;
    layer1_outputs(8815) <= a and b;
    layer1_outputs(8816) <= a and not b;
    layer1_outputs(8817) <= not (a xor b);
    layer1_outputs(8818) <= a;
    layer1_outputs(8819) <= a and not b;
    layer1_outputs(8820) <= b and not a;
    layer1_outputs(8821) <= a or b;
    layer1_outputs(8822) <= '0';
    layer1_outputs(8823) <= not (a or b);
    layer1_outputs(8824) <= a;
    layer1_outputs(8825) <= not b;
    layer1_outputs(8826) <= a and not b;
    layer1_outputs(8827) <= b;
    layer1_outputs(8828) <= not b or a;
    layer1_outputs(8829) <= a and not b;
    layer1_outputs(8830) <= b and not a;
    layer1_outputs(8831) <= not b;
    layer1_outputs(8832) <= b;
    layer1_outputs(8833) <= not a;
    layer1_outputs(8834) <= a and b;
    layer1_outputs(8835) <= a or b;
    layer1_outputs(8836) <= a or b;
    layer1_outputs(8837) <= not a;
    layer1_outputs(8838) <= a or b;
    layer1_outputs(8839) <= not b or a;
    layer1_outputs(8840) <= not a or b;
    layer1_outputs(8841) <= not (a and b);
    layer1_outputs(8842) <= not b;
    layer1_outputs(8843) <= b and not a;
    layer1_outputs(8844) <= a and not b;
    layer1_outputs(8845) <= not (a and b);
    layer1_outputs(8846) <= not (a or b);
    layer1_outputs(8847) <= a and not b;
    layer1_outputs(8848) <= b;
    layer1_outputs(8849) <= '1';
    layer1_outputs(8850) <= b;
    layer1_outputs(8851) <= '0';
    layer1_outputs(8852) <= a and b;
    layer1_outputs(8853) <= not a or b;
    layer1_outputs(8854) <= a or b;
    layer1_outputs(8855) <= not (a or b);
    layer1_outputs(8856) <= a;
    layer1_outputs(8857) <= not a;
    layer1_outputs(8858) <= a xor b;
    layer1_outputs(8859) <= not b;
    layer1_outputs(8860) <= '0';
    layer1_outputs(8861) <= b and not a;
    layer1_outputs(8862) <= a;
    layer1_outputs(8863) <= '1';
    layer1_outputs(8864) <= a xor b;
    layer1_outputs(8865) <= not a or b;
    layer1_outputs(8866) <= a;
    layer1_outputs(8867) <= not (a xor b);
    layer1_outputs(8868) <= not b;
    layer1_outputs(8869) <= not a;
    layer1_outputs(8870) <= not b;
    layer1_outputs(8871) <= not a;
    layer1_outputs(8872) <= a xor b;
    layer1_outputs(8873) <= '1';
    layer1_outputs(8874) <= b;
    layer1_outputs(8875) <= a;
    layer1_outputs(8876) <= a and b;
    layer1_outputs(8877) <= a or b;
    layer1_outputs(8878) <= a or b;
    layer1_outputs(8879) <= a;
    layer1_outputs(8880) <= a;
    layer1_outputs(8881) <= not a or b;
    layer1_outputs(8882) <= a and not b;
    layer1_outputs(8883) <= not a;
    layer1_outputs(8884) <= not (a or b);
    layer1_outputs(8885) <= a xor b;
    layer1_outputs(8886) <= a or b;
    layer1_outputs(8887) <= not a;
    layer1_outputs(8888) <= not (a xor b);
    layer1_outputs(8889) <= a and b;
    layer1_outputs(8890) <= a and b;
    layer1_outputs(8891) <= not b;
    layer1_outputs(8892) <= a and not b;
    layer1_outputs(8893) <= not (a and b);
    layer1_outputs(8894) <= not b;
    layer1_outputs(8895) <= '0';
    layer1_outputs(8896) <= not (a and b);
    layer1_outputs(8897) <= not b or a;
    layer1_outputs(8898) <= a;
    layer1_outputs(8899) <= not (a or b);
    layer1_outputs(8900) <= b;
    layer1_outputs(8901) <= not a;
    layer1_outputs(8902) <= not (a and b);
    layer1_outputs(8903) <= not (a or b);
    layer1_outputs(8904) <= a;
    layer1_outputs(8905) <= b;
    layer1_outputs(8906) <= not b or a;
    layer1_outputs(8907) <= a or b;
    layer1_outputs(8908) <= a;
    layer1_outputs(8909) <= b;
    layer1_outputs(8910) <= b and not a;
    layer1_outputs(8911) <= not (a xor b);
    layer1_outputs(8912) <= '1';
    layer1_outputs(8913) <= b;
    layer1_outputs(8914) <= a and b;
    layer1_outputs(8915) <= b and not a;
    layer1_outputs(8916) <= not b;
    layer1_outputs(8917) <= not b;
    layer1_outputs(8918) <= '0';
    layer1_outputs(8919) <= a or b;
    layer1_outputs(8920) <= b and not a;
    layer1_outputs(8921) <= not b;
    layer1_outputs(8922) <= not b or a;
    layer1_outputs(8923) <= not a or b;
    layer1_outputs(8924) <= '0';
    layer1_outputs(8925) <= not b;
    layer1_outputs(8926) <= a;
    layer1_outputs(8927) <= not a or b;
    layer1_outputs(8928) <= not a;
    layer1_outputs(8929) <= '0';
    layer1_outputs(8930) <= not b or a;
    layer1_outputs(8931) <= not b;
    layer1_outputs(8932) <= not (a or b);
    layer1_outputs(8933) <= not (a or b);
    layer1_outputs(8934) <= not a;
    layer1_outputs(8935) <= not a;
    layer1_outputs(8936) <= a xor b;
    layer1_outputs(8937) <= a and b;
    layer1_outputs(8938) <= not b or a;
    layer1_outputs(8939) <= not (a and b);
    layer1_outputs(8940) <= b;
    layer1_outputs(8941) <= not (a xor b);
    layer1_outputs(8942) <= a and not b;
    layer1_outputs(8943) <= a;
    layer1_outputs(8944) <= not a;
    layer1_outputs(8945) <= not b or a;
    layer1_outputs(8946) <= not a or b;
    layer1_outputs(8947) <= not a or b;
    layer1_outputs(8948) <= a xor b;
    layer1_outputs(8949) <= not (a or b);
    layer1_outputs(8950) <= '0';
    layer1_outputs(8951) <= '1';
    layer1_outputs(8952) <= '0';
    layer1_outputs(8953) <= not b or a;
    layer1_outputs(8954) <= not b;
    layer1_outputs(8955) <= a;
    layer1_outputs(8956) <= b;
    layer1_outputs(8957) <= not b;
    layer1_outputs(8958) <= not b;
    layer1_outputs(8959) <= not (a xor b);
    layer1_outputs(8960) <= a xor b;
    layer1_outputs(8961) <= '0';
    layer1_outputs(8962) <= a;
    layer1_outputs(8963) <= not (a and b);
    layer1_outputs(8964) <= a and not b;
    layer1_outputs(8965) <= b and not a;
    layer1_outputs(8966) <= not a or b;
    layer1_outputs(8967) <= '1';
    layer1_outputs(8968) <= '0';
    layer1_outputs(8969) <= not b or a;
    layer1_outputs(8970) <= a and b;
    layer1_outputs(8971) <= not a;
    layer1_outputs(8972) <= a xor b;
    layer1_outputs(8973) <= not a or b;
    layer1_outputs(8974) <= a and b;
    layer1_outputs(8975) <= a and b;
    layer1_outputs(8976) <= a and b;
    layer1_outputs(8977) <= not (a xor b);
    layer1_outputs(8978) <= not (a or b);
    layer1_outputs(8979) <= not a or b;
    layer1_outputs(8980) <= not b;
    layer1_outputs(8981) <= b;
    layer1_outputs(8982) <= not a;
    layer1_outputs(8983) <= not (a or b);
    layer1_outputs(8984) <= not a or b;
    layer1_outputs(8985) <= not b;
    layer1_outputs(8986) <= not a or b;
    layer1_outputs(8987) <= a and not b;
    layer1_outputs(8988) <= b;
    layer1_outputs(8989) <= a and b;
    layer1_outputs(8990) <= not (a xor b);
    layer1_outputs(8991) <= a or b;
    layer1_outputs(8992) <= not (a and b);
    layer1_outputs(8993) <= a and b;
    layer1_outputs(8994) <= a;
    layer1_outputs(8995) <= a or b;
    layer1_outputs(8996) <= not b or a;
    layer1_outputs(8997) <= b and not a;
    layer1_outputs(8998) <= a xor b;
    layer1_outputs(8999) <= a;
    layer1_outputs(9000) <= a xor b;
    layer1_outputs(9001) <= '1';
    layer1_outputs(9002) <= not b or a;
    layer1_outputs(9003) <= a and not b;
    layer1_outputs(9004) <= '1';
    layer1_outputs(9005) <= not b;
    layer1_outputs(9006) <= not a;
    layer1_outputs(9007) <= a or b;
    layer1_outputs(9008) <= not b;
    layer1_outputs(9009) <= '0';
    layer1_outputs(9010) <= a or b;
    layer1_outputs(9011) <= not b or a;
    layer1_outputs(9012) <= not (a and b);
    layer1_outputs(9013) <= not a;
    layer1_outputs(9014) <= b;
    layer1_outputs(9015) <= not a or b;
    layer1_outputs(9016) <= a;
    layer1_outputs(9017) <= not a;
    layer1_outputs(9018) <= not (a or b);
    layer1_outputs(9019) <= not b;
    layer1_outputs(9020) <= a xor b;
    layer1_outputs(9021) <= not b;
    layer1_outputs(9022) <= not a;
    layer1_outputs(9023) <= b and not a;
    layer1_outputs(9024) <= b and not a;
    layer1_outputs(9025) <= b;
    layer1_outputs(9026) <= not (a and b);
    layer1_outputs(9027) <= a and not b;
    layer1_outputs(9028) <= not b or a;
    layer1_outputs(9029) <= not (a xor b);
    layer1_outputs(9030) <= a;
    layer1_outputs(9031) <= not b;
    layer1_outputs(9032) <= not a;
    layer1_outputs(9033) <= b and not a;
    layer1_outputs(9034) <= b;
    layer1_outputs(9035) <= b and not a;
    layer1_outputs(9036) <= b;
    layer1_outputs(9037) <= a xor b;
    layer1_outputs(9038) <= a;
    layer1_outputs(9039) <= not a;
    layer1_outputs(9040) <= a and not b;
    layer1_outputs(9041) <= b and not a;
    layer1_outputs(9042) <= a or b;
    layer1_outputs(9043) <= b;
    layer1_outputs(9044) <= not a;
    layer1_outputs(9045) <= not b;
    layer1_outputs(9046) <= not a;
    layer1_outputs(9047) <= a or b;
    layer1_outputs(9048) <= a and not b;
    layer1_outputs(9049) <= not b;
    layer1_outputs(9050) <= not b or a;
    layer1_outputs(9051) <= a xor b;
    layer1_outputs(9052) <= not a;
    layer1_outputs(9053) <= a and b;
    layer1_outputs(9054) <= b and not a;
    layer1_outputs(9055) <= a;
    layer1_outputs(9056) <= a xor b;
    layer1_outputs(9057) <= a and b;
    layer1_outputs(9058) <= a;
    layer1_outputs(9059) <= a or b;
    layer1_outputs(9060) <= b;
    layer1_outputs(9061) <= '1';
    layer1_outputs(9062) <= '1';
    layer1_outputs(9063) <= not b;
    layer1_outputs(9064) <= '1';
    layer1_outputs(9065) <= not (a and b);
    layer1_outputs(9066) <= a or b;
    layer1_outputs(9067) <= a xor b;
    layer1_outputs(9068) <= b;
    layer1_outputs(9069) <= '0';
    layer1_outputs(9070) <= not b;
    layer1_outputs(9071) <= a and b;
    layer1_outputs(9072) <= not b;
    layer1_outputs(9073) <= not a or b;
    layer1_outputs(9074) <= not b;
    layer1_outputs(9075) <= not a;
    layer1_outputs(9076) <= a and b;
    layer1_outputs(9077) <= b;
    layer1_outputs(9078) <= not a;
    layer1_outputs(9079) <= not a or b;
    layer1_outputs(9080) <= a and not b;
    layer1_outputs(9081) <= not a;
    layer1_outputs(9082) <= not a;
    layer1_outputs(9083) <= a and b;
    layer1_outputs(9084) <= not b or a;
    layer1_outputs(9085) <= '1';
    layer1_outputs(9086) <= b and not a;
    layer1_outputs(9087) <= b and not a;
    layer1_outputs(9088) <= a and b;
    layer1_outputs(9089) <= not a or b;
    layer1_outputs(9090) <= a or b;
    layer1_outputs(9091) <= a or b;
    layer1_outputs(9092) <= not (a and b);
    layer1_outputs(9093) <= b;
    layer1_outputs(9094) <= b;
    layer1_outputs(9095) <= not b;
    layer1_outputs(9096) <= a and not b;
    layer1_outputs(9097) <= not a;
    layer1_outputs(9098) <= a and b;
    layer1_outputs(9099) <= not b or a;
    layer1_outputs(9100) <= not b;
    layer1_outputs(9101) <= not (a and b);
    layer1_outputs(9102) <= a;
    layer1_outputs(9103) <= a and not b;
    layer1_outputs(9104) <= b and not a;
    layer1_outputs(9105) <= not (a and b);
    layer1_outputs(9106) <= a xor b;
    layer1_outputs(9107) <= not a;
    layer1_outputs(9108) <= a and not b;
    layer1_outputs(9109) <= a or b;
    layer1_outputs(9110) <= a and not b;
    layer1_outputs(9111) <= not b;
    layer1_outputs(9112) <= not a;
    layer1_outputs(9113) <= not b or a;
    layer1_outputs(9114) <= a and b;
    layer1_outputs(9115) <= not a or b;
    layer1_outputs(9116) <= b;
    layer1_outputs(9117) <= b;
    layer1_outputs(9118) <= b;
    layer1_outputs(9119) <= not a;
    layer1_outputs(9120) <= not a;
    layer1_outputs(9121) <= not a or b;
    layer1_outputs(9122) <= '1';
    layer1_outputs(9123) <= not b or a;
    layer1_outputs(9124) <= b and not a;
    layer1_outputs(9125) <= b;
    layer1_outputs(9126) <= not b or a;
    layer1_outputs(9127) <= a and not b;
    layer1_outputs(9128) <= not (a xor b);
    layer1_outputs(9129) <= a and b;
    layer1_outputs(9130) <= '0';
    layer1_outputs(9131) <= b and not a;
    layer1_outputs(9132) <= not a;
    layer1_outputs(9133) <= not (a or b);
    layer1_outputs(9134) <= not (a xor b);
    layer1_outputs(9135) <= a;
    layer1_outputs(9136) <= not a or b;
    layer1_outputs(9137) <= a and b;
    layer1_outputs(9138) <= not a or b;
    layer1_outputs(9139) <= not (a or b);
    layer1_outputs(9140) <= '1';
    layer1_outputs(9141) <= a and not b;
    layer1_outputs(9142) <= b and not a;
    layer1_outputs(9143) <= not a;
    layer1_outputs(9144) <= a;
    layer1_outputs(9145) <= '0';
    layer1_outputs(9146) <= not a;
    layer1_outputs(9147) <= a;
    layer1_outputs(9148) <= b and not a;
    layer1_outputs(9149) <= '1';
    layer1_outputs(9150) <= a;
    layer1_outputs(9151) <= a and not b;
    layer1_outputs(9152) <= a xor b;
    layer1_outputs(9153) <= not a;
    layer1_outputs(9154) <= not (a and b);
    layer1_outputs(9155) <= not (a xor b);
    layer1_outputs(9156) <= '0';
    layer1_outputs(9157) <= a or b;
    layer1_outputs(9158) <= not b;
    layer1_outputs(9159) <= b and not a;
    layer1_outputs(9160) <= a or b;
    layer1_outputs(9161) <= not b or a;
    layer1_outputs(9162) <= a or b;
    layer1_outputs(9163) <= not a or b;
    layer1_outputs(9164) <= a and b;
    layer1_outputs(9165) <= not b or a;
    layer1_outputs(9166) <= not (a or b);
    layer1_outputs(9167) <= not b or a;
    layer1_outputs(9168) <= not (a and b);
    layer1_outputs(9169) <= a and not b;
    layer1_outputs(9170) <= b;
    layer1_outputs(9171) <= not (a and b);
    layer1_outputs(9172) <= not (a and b);
    layer1_outputs(9173) <= not a;
    layer1_outputs(9174) <= not b;
    layer1_outputs(9175) <= not a or b;
    layer1_outputs(9176) <= '1';
    layer1_outputs(9177) <= '0';
    layer1_outputs(9178) <= b;
    layer1_outputs(9179) <= not (a and b);
    layer1_outputs(9180) <= not (a xor b);
    layer1_outputs(9181) <= not a;
    layer1_outputs(9182) <= not b or a;
    layer1_outputs(9183) <= '0';
    layer1_outputs(9184) <= not a or b;
    layer1_outputs(9185) <= not (a or b);
    layer1_outputs(9186) <= not (a or b);
    layer1_outputs(9187) <= not (a or b);
    layer1_outputs(9188) <= not a or b;
    layer1_outputs(9189) <= a xor b;
    layer1_outputs(9190) <= a and not b;
    layer1_outputs(9191) <= '0';
    layer1_outputs(9192) <= '1';
    layer1_outputs(9193) <= b;
    layer1_outputs(9194) <= not (a xor b);
    layer1_outputs(9195) <= b;
    layer1_outputs(9196) <= '0';
    layer1_outputs(9197) <= b;
    layer1_outputs(9198) <= a xor b;
    layer1_outputs(9199) <= not (a and b);
    layer1_outputs(9200) <= '0';
    layer1_outputs(9201) <= '0';
    layer1_outputs(9202) <= a;
    layer1_outputs(9203) <= not a;
    layer1_outputs(9204) <= not (a and b);
    layer1_outputs(9205) <= not (a and b);
    layer1_outputs(9206) <= a and not b;
    layer1_outputs(9207) <= not b or a;
    layer1_outputs(9208) <= a;
    layer1_outputs(9209) <= not a;
    layer1_outputs(9210) <= b;
    layer1_outputs(9211) <= b and not a;
    layer1_outputs(9212) <= b;
    layer1_outputs(9213) <= a xor b;
    layer1_outputs(9214) <= a and not b;
    layer1_outputs(9215) <= a and b;
    layer1_outputs(9216) <= not b or a;
    layer1_outputs(9217) <= a or b;
    layer1_outputs(9218) <= not b or a;
    layer1_outputs(9219) <= a or b;
    layer1_outputs(9220) <= '0';
    layer1_outputs(9221) <= not a or b;
    layer1_outputs(9222) <= '0';
    layer1_outputs(9223) <= not (a and b);
    layer1_outputs(9224) <= not a or b;
    layer1_outputs(9225) <= a xor b;
    layer1_outputs(9226) <= b;
    layer1_outputs(9227) <= not a;
    layer1_outputs(9228) <= not a;
    layer1_outputs(9229) <= a and not b;
    layer1_outputs(9230) <= a or b;
    layer1_outputs(9231) <= not b;
    layer1_outputs(9232) <= a;
    layer1_outputs(9233) <= '0';
    layer1_outputs(9234) <= '1';
    layer1_outputs(9235) <= a and b;
    layer1_outputs(9236) <= a;
    layer1_outputs(9237) <= a or b;
    layer1_outputs(9238) <= a;
    layer1_outputs(9239) <= not (a xor b);
    layer1_outputs(9240) <= a and not b;
    layer1_outputs(9241) <= not a or b;
    layer1_outputs(9242) <= not a or b;
    layer1_outputs(9243) <= b and not a;
    layer1_outputs(9244) <= not a;
    layer1_outputs(9245) <= b and not a;
    layer1_outputs(9246) <= not b or a;
    layer1_outputs(9247) <= not b;
    layer1_outputs(9248) <= b;
    layer1_outputs(9249) <= '0';
    layer1_outputs(9250) <= not (a xor b);
    layer1_outputs(9251) <= '0';
    layer1_outputs(9252) <= not b;
    layer1_outputs(9253) <= '0';
    layer1_outputs(9254) <= not (a and b);
    layer1_outputs(9255) <= '1';
    layer1_outputs(9256) <= b and not a;
    layer1_outputs(9257) <= not (a or b);
    layer1_outputs(9258) <= a or b;
    layer1_outputs(9259) <= '0';
    layer1_outputs(9260) <= not (a or b);
    layer1_outputs(9261) <= not b or a;
    layer1_outputs(9262) <= '0';
    layer1_outputs(9263) <= a;
    layer1_outputs(9264) <= a xor b;
    layer1_outputs(9265) <= not b or a;
    layer1_outputs(9266) <= b;
    layer1_outputs(9267) <= a xor b;
    layer1_outputs(9268) <= not a;
    layer1_outputs(9269) <= b;
    layer1_outputs(9270) <= not a or b;
    layer1_outputs(9271) <= '1';
    layer1_outputs(9272) <= not b;
    layer1_outputs(9273) <= not (a or b);
    layer1_outputs(9274) <= b;
    layer1_outputs(9275) <= a or b;
    layer1_outputs(9276) <= '0';
    layer1_outputs(9277) <= not b or a;
    layer1_outputs(9278) <= not (a and b);
    layer1_outputs(9279) <= '1';
    layer1_outputs(9280) <= not (a xor b);
    layer1_outputs(9281) <= a and b;
    layer1_outputs(9282) <= b;
    layer1_outputs(9283) <= not b or a;
    layer1_outputs(9284) <= a and not b;
    layer1_outputs(9285) <= '0';
    layer1_outputs(9286) <= not b;
    layer1_outputs(9287) <= not b or a;
    layer1_outputs(9288) <= a and not b;
    layer1_outputs(9289) <= not (a and b);
    layer1_outputs(9290) <= not (a xor b);
    layer1_outputs(9291) <= b;
    layer1_outputs(9292) <= a and not b;
    layer1_outputs(9293) <= not a or b;
    layer1_outputs(9294) <= a;
    layer1_outputs(9295) <= '1';
    layer1_outputs(9296) <= not a;
    layer1_outputs(9297) <= not (a and b);
    layer1_outputs(9298) <= b;
    layer1_outputs(9299) <= not a or b;
    layer1_outputs(9300) <= '0';
    layer1_outputs(9301) <= b and not a;
    layer1_outputs(9302) <= not a;
    layer1_outputs(9303) <= '0';
    layer1_outputs(9304) <= not (a xor b);
    layer1_outputs(9305) <= '0';
    layer1_outputs(9306) <= b and not a;
    layer1_outputs(9307) <= '0';
    layer1_outputs(9308) <= b and not a;
    layer1_outputs(9309) <= not (a and b);
    layer1_outputs(9310) <= not a or b;
    layer1_outputs(9311) <= not (a or b);
    layer1_outputs(9312) <= not b or a;
    layer1_outputs(9313) <= a and not b;
    layer1_outputs(9314) <= not b or a;
    layer1_outputs(9315) <= a or b;
    layer1_outputs(9316) <= b and not a;
    layer1_outputs(9317) <= not b;
    layer1_outputs(9318) <= '0';
    layer1_outputs(9319) <= a or b;
    layer1_outputs(9320) <= a or b;
    layer1_outputs(9321) <= not (a and b);
    layer1_outputs(9322) <= a and b;
    layer1_outputs(9323) <= not (a or b);
    layer1_outputs(9324) <= '0';
    layer1_outputs(9325) <= not b;
    layer1_outputs(9326) <= '1';
    layer1_outputs(9327) <= not (a and b);
    layer1_outputs(9328) <= a and not b;
    layer1_outputs(9329) <= not (a xor b);
    layer1_outputs(9330) <= not b;
    layer1_outputs(9331) <= a;
    layer1_outputs(9332) <= not b;
    layer1_outputs(9333) <= a and not b;
    layer1_outputs(9334) <= not (a and b);
    layer1_outputs(9335) <= not (a or b);
    layer1_outputs(9336) <= not (a and b);
    layer1_outputs(9337) <= not (a or b);
    layer1_outputs(9338) <= '0';
    layer1_outputs(9339) <= not b;
    layer1_outputs(9340) <= not a or b;
    layer1_outputs(9341) <= '1';
    layer1_outputs(9342) <= a;
    layer1_outputs(9343) <= '1';
    layer1_outputs(9344) <= not (a and b);
    layer1_outputs(9345) <= b;
    layer1_outputs(9346) <= b and not a;
    layer1_outputs(9347) <= not (a and b);
    layer1_outputs(9348) <= not (a and b);
    layer1_outputs(9349) <= '1';
    layer1_outputs(9350) <= '1';
    layer1_outputs(9351) <= a xor b;
    layer1_outputs(9352) <= '0';
    layer1_outputs(9353) <= a or b;
    layer1_outputs(9354) <= '0';
    layer1_outputs(9355) <= '1';
    layer1_outputs(9356) <= b and not a;
    layer1_outputs(9357) <= not a or b;
    layer1_outputs(9358) <= not (a xor b);
    layer1_outputs(9359) <= a or b;
    layer1_outputs(9360) <= not a;
    layer1_outputs(9361) <= b;
    layer1_outputs(9362) <= b and not a;
    layer1_outputs(9363) <= a and b;
    layer1_outputs(9364) <= not a or b;
    layer1_outputs(9365) <= '0';
    layer1_outputs(9366) <= a and not b;
    layer1_outputs(9367) <= not (a xor b);
    layer1_outputs(9368) <= b and not a;
    layer1_outputs(9369) <= not b or a;
    layer1_outputs(9370) <= b and not a;
    layer1_outputs(9371) <= not b;
    layer1_outputs(9372) <= b and not a;
    layer1_outputs(9373) <= '0';
    layer1_outputs(9374) <= not (a and b);
    layer1_outputs(9375) <= a and b;
    layer1_outputs(9376) <= not b;
    layer1_outputs(9377) <= a and not b;
    layer1_outputs(9378) <= a and b;
    layer1_outputs(9379) <= a xor b;
    layer1_outputs(9380) <= not a;
    layer1_outputs(9381) <= a and not b;
    layer1_outputs(9382) <= b;
    layer1_outputs(9383) <= a;
    layer1_outputs(9384) <= not a;
    layer1_outputs(9385) <= not b or a;
    layer1_outputs(9386) <= a or b;
    layer1_outputs(9387) <= b;
    layer1_outputs(9388) <= a;
    layer1_outputs(9389) <= not a or b;
    layer1_outputs(9390) <= not (a and b);
    layer1_outputs(9391) <= not (a or b);
    layer1_outputs(9392) <= a or b;
    layer1_outputs(9393) <= not (a or b);
    layer1_outputs(9394) <= a and b;
    layer1_outputs(9395) <= not a or b;
    layer1_outputs(9396) <= a;
    layer1_outputs(9397) <= '1';
    layer1_outputs(9398) <= '0';
    layer1_outputs(9399) <= not b;
    layer1_outputs(9400) <= not (a and b);
    layer1_outputs(9401) <= b;
    layer1_outputs(9402) <= not (a and b);
    layer1_outputs(9403) <= b;
    layer1_outputs(9404) <= '0';
    layer1_outputs(9405) <= not b or a;
    layer1_outputs(9406) <= a xor b;
    layer1_outputs(9407) <= not b;
    layer1_outputs(9408) <= not (a xor b);
    layer1_outputs(9409) <= a xor b;
    layer1_outputs(9410) <= a;
    layer1_outputs(9411) <= not b;
    layer1_outputs(9412) <= a and b;
    layer1_outputs(9413) <= not b;
    layer1_outputs(9414) <= a and b;
    layer1_outputs(9415) <= b;
    layer1_outputs(9416) <= b and not a;
    layer1_outputs(9417) <= a and not b;
    layer1_outputs(9418) <= not b or a;
    layer1_outputs(9419) <= b;
    layer1_outputs(9420) <= '0';
    layer1_outputs(9421) <= not a or b;
    layer1_outputs(9422) <= not (a or b);
    layer1_outputs(9423) <= '0';
    layer1_outputs(9424) <= a and b;
    layer1_outputs(9425) <= a xor b;
    layer1_outputs(9426) <= not a or b;
    layer1_outputs(9427) <= a or b;
    layer1_outputs(9428) <= a or b;
    layer1_outputs(9429) <= '0';
    layer1_outputs(9430) <= a;
    layer1_outputs(9431) <= not a;
    layer1_outputs(9432) <= b;
    layer1_outputs(9433) <= b;
    layer1_outputs(9434) <= a or b;
    layer1_outputs(9435) <= b;
    layer1_outputs(9436) <= a or b;
    layer1_outputs(9437) <= b and not a;
    layer1_outputs(9438) <= not (a or b);
    layer1_outputs(9439) <= '0';
    layer1_outputs(9440) <= b;
    layer1_outputs(9441) <= a and not b;
    layer1_outputs(9442) <= '0';
    layer1_outputs(9443) <= '1';
    layer1_outputs(9444) <= not b;
    layer1_outputs(9445) <= a and b;
    layer1_outputs(9446) <= not (a xor b);
    layer1_outputs(9447) <= '0';
    layer1_outputs(9448) <= a xor b;
    layer1_outputs(9449) <= '0';
    layer1_outputs(9450) <= not b;
    layer1_outputs(9451) <= not b;
    layer1_outputs(9452) <= not (a xor b);
    layer1_outputs(9453) <= not b or a;
    layer1_outputs(9454) <= not a or b;
    layer1_outputs(9455) <= not (a and b);
    layer1_outputs(9456) <= not (a or b);
    layer1_outputs(9457) <= not a or b;
    layer1_outputs(9458) <= not b;
    layer1_outputs(9459) <= a and not b;
    layer1_outputs(9460) <= '1';
    layer1_outputs(9461) <= not b or a;
    layer1_outputs(9462) <= b and not a;
    layer1_outputs(9463) <= a and not b;
    layer1_outputs(9464) <= b and not a;
    layer1_outputs(9465) <= a and not b;
    layer1_outputs(9466) <= a or b;
    layer1_outputs(9467) <= a and b;
    layer1_outputs(9468) <= '1';
    layer1_outputs(9469) <= not (a or b);
    layer1_outputs(9470) <= '1';
    layer1_outputs(9471) <= a and not b;
    layer1_outputs(9472) <= a;
    layer1_outputs(9473) <= a and b;
    layer1_outputs(9474) <= not (a and b);
    layer1_outputs(9475) <= '0';
    layer1_outputs(9476) <= b;
    layer1_outputs(9477) <= b;
    layer1_outputs(9478) <= not a;
    layer1_outputs(9479) <= b and not a;
    layer1_outputs(9480) <= a and b;
    layer1_outputs(9481) <= not b;
    layer1_outputs(9482) <= not b;
    layer1_outputs(9483) <= b;
    layer1_outputs(9484) <= a and not b;
    layer1_outputs(9485) <= a and b;
    layer1_outputs(9486) <= not a or b;
    layer1_outputs(9487) <= not a;
    layer1_outputs(9488) <= not b or a;
    layer1_outputs(9489) <= a or b;
    layer1_outputs(9490) <= '0';
    layer1_outputs(9491) <= not a or b;
    layer1_outputs(9492) <= not a;
    layer1_outputs(9493) <= not b;
    layer1_outputs(9494) <= not (a and b);
    layer1_outputs(9495) <= not (a xor b);
    layer1_outputs(9496) <= not b;
    layer1_outputs(9497) <= not (a or b);
    layer1_outputs(9498) <= a and not b;
    layer1_outputs(9499) <= a xor b;
    layer1_outputs(9500) <= a or b;
    layer1_outputs(9501) <= not (a or b);
    layer1_outputs(9502) <= not a or b;
    layer1_outputs(9503) <= not a;
    layer1_outputs(9504) <= not b;
    layer1_outputs(9505) <= not a;
    layer1_outputs(9506) <= b and not a;
    layer1_outputs(9507) <= not b;
    layer1_outputs(9508) <= not (a and b);
    layer1_outputs(9509) <= a and b;
    layer1_outputs(9510) <= '1';
    layer1_outputs(9511) <= a;
    layer1_outputs(9512) <= not a;
    layer1_outputs(9513) <= '1';
    layer1_outputs(9514) <= not b;
    layer1_outputs(9515) <= not b;
    layer1_outputs(9516) <= not b or a;
    layer1_outputs(9517) <= not (a or b);
    layer1_outputs(9518) <= not b;
    layer1_outputs(9519) <= a and b;
    layer1_outputs(9520) <= not (a or b);
    layer1_outputs(9521) <= not b or a;
    layer1_outputs(9522) <= a;
    layer1_outputs(9523) <= b;
    layer1_outputs(9524) <= not b or a;
    layer1_outputs(9525) <= a;
    layer1_outputs(9526) <= '0';
    layer1_outputs(9527) <= a and b;
    layer1_outputs(9528) <= not a;
    layer1_outputs(9529) <= not b;
    layer1_outputs(9530) <= '1';
    layer1_outputs(9531) <= a;
    layer1_outputs(9532) <= a and not b;
    layer1_outputs(9533) <= a or b;
    layer1_outputs(9534) <= not b or a;
    layer1_outputs(9535) <= b;
    layer1_outputs(9536) <= not a;
    layer1_outputs(9537) <= a and b;
    layer1_outputs(9538) <= '1';
    layer1_outputs(9539) <= not b;
    layer1_outputs(9540) <= a;
    layer1_outputs(9541) <= not (a xor b);
    layer1_outputs(9542) <= a;
    layer1_outputs(9543) <= a and not b;
    layer1_outputs(9544) <= not (a and b);
    layer1_outputs(9545) <= not (a and b);
    layer1_outputs(9546) <= not (a and b);
    layer1_outputs(9547) <= a and b;
    layer1_outputs(9548) <= not a;
    layer1_outputs(9549) <= not a;
    layer1_outputs(9550) <= not b or a;
    layer1_outputs(9551) <= not (a or b);
    layer1_outputs(9552) <= a;
    layer1_outputs(9553) <= not (a xor b);
    layer1_outputs(9554) <= not (a xor b);
    layer1_outputs(9555) <= not (a or b);
    layer1_outputs(9556) <= not b;
    layer1_outputs(9557) <= not (a and b);
    layer1_outputs(9558) <= b;
    layer1_outputs(9559) <= not a or b;
    layer1_outputs(9560) <= b and not a;
    layer1_outputs(9561) <= not a or b;
    layer1_outputs(9562) <= a or b;
    layer1_outputs(9563) <= not a;
    layer1_outputs(9564) <= a and b;
    layer1_outputs(9565) <= b;
    layer1_outputs(9566) <= '1';
    layer1_outputs(9567) <= '1';
    layer1_outputs(9568) <= not b or a;
    layer1_outputs(9569) <= not (a xor b);
    layer1_outputs(9570) <= '1';
    layer1_outputs(9571) <= '1';
    layer1_outputs(9572) <= not a or b;
    layer1_outputs(9573) <= a or b;
    layer1_outputs(9574) <= not (a and b);
    layer1_outputs(9575) <= a and not b;
    layer1_outputs(9576) <= '0';
    layer1_outputs(9577) <= not a;
    layer1_outputs(9578) <= not (a and b);
    layer1_outputs(9579) <= not b;
    layer1_outputs(9580) <= not a or b;
    layer1_outputs(9581) <= '1';
    layer1_outputs(9582) <= not (a or b);
    layer1_outputs(9583) <= a and not b;
    layer1_outputs(9584) <= a or b;
    layer1_outputs(9585) <= b and not a;
    layer1_outputs(9586) <= not b or a;
    layer1_outputs(9587) <= not a or b;
    layer1_outputs(9588) <= a and not b;
    layer1_outputs(9589) <= not b or a;
    layer1_outputs(9590) <= '1';
    layer1_outputs(9591) <= a and not b;
    layer1_outputs(9592) <= a and b;
    layer1_outputs(9593) <= not a or b;
    layer1_outputs(9594) <= b and not a;
    layer1_outputs(9595) <= not a or b;
    layer1_outputs(9596) <= not (a and b);
    layer1_outputs(9597) <= not b;
    layer1_outputs(9598) <= a or b;
    layer1_outputs(9599) <= b;
    layer1_outputs(9600) <= '0';
    layer1_outputs(9601) <= not (a xor b);
    layer1_outputs(9602) <= not b;
    layer1_outputs(9603) <= '0';
    layer1_outputs(9604) <= a or b;
    layer1_outputs(9605) <= not b;
    layer1_outputs(9606) <= a xor b;
    layer1_outputs(9607) <= a and not b;
    layer1_outputs(9608) <= not (a and b);
    layer1_outputs(9609) <= not b;
    layer1_outputs(9610) <= a and b;
    layer1_outputs(9611) <= b and not a;
    layer1_outputs(9612) <= not a;
    layer1_outputs(9613) <= a;
    layer1_outputs(9614) <= a;
    layer1_outputs(9615) <= a or b;
    layer1_outputs(9616) <= '0';
    layer1_outputs(9617) <= not (a and b);
    layer1_outputs(9618) <= not b;
    layer1_outputs(9619) <= a or b;
    layer1_outputs(9620) <= not a or b;
    layer1_outputs(9621) <= not b or a;
    layer1_outputs(9622) <= not a or b;
    layer1_outputs(9623) <= a and not b;
    layer1_outputs(9624) <= a;
    layer1_outputs(9625) <= a and b;
    layer1_outputs(9626) <= not (a and b);
    layer1_outputs(9627) <= not a or b;
    layer1_outputs(9628) <= a and not b;
    layer1_outputs(9629) <= not a or b;
    layer1_outputs(9630) <= not b or a;
    layer1_outputs(9631) <= '1';
    layer1_outputs(9632) <= a and not b;
    layer1_outputs(9633) <= not a;
    layer1_outputs(9634) <= not b or a;
    layer1_outputs(9635) <= not (a xor b);
    layer1_outputs(9636) <= a;
    layer1_outputs(9637) <= '0';
    layer1_outputs(9638) <= a xor b;
    layer1_outputs(9639) <= '1';
    layer1_outputs(9640) <= not (a xor b);
    layer1_outputs(9641) <= not (a and b);
    layer1_outputs(9642) <= b and not a;
    layer1_outputs(9643) <= a and b;
    layer1_outputs(9644) <= '0';
    layer1_outputs(9645) <= b and not a;
    layer1_outputs(9646) <= '0';
    layer1_outputs(9647) <= a and b;
    layer1_outputs(9648) <= not (a or b);
    layer1_outputs(9649) <= a and not b;
    layer1_outputs(9650) <= not a or b;
    layer1_outputs(9651) <= '1';
    layer1_outputs(9652) <= a;
    layer1_outputs(9653) <= not a or b;
    layer1_outputs(9654) <= not b;
    layer1_outputs(9655) <= not (a or b);
    layer1_outputs(9656) <= not (a and b);
    layer1_outputs(9657) <= not a or b;
    layer1_outputs(9658) <= not (a or b);
    layer1_outputs(9659) <= b and not a;
    layer1_outputs(9660) <= not a or b;
    layer1_outputs(9661) <= a;
    layer1_outputs(9662) <= '0';
    layer1_outputs(9663) <= not (a and b);
    layer1_outputs(9664) <= not b or a;
    layer1_outputs(9665) <= a and not b;
    layer1_outputs(9666) <= not a;
    layer1_outputs(9667) <= not b or a;
    layer1_outputs(9668) <= not (a or b);
    layer1_outputs(9669) <= a;
    layer1_outputs(9670) <= not a;
    layer1_outputs(9671) <= not (a and b);
    layer1_outputs(9672) <= not a or b;
    layer1_outputs(9673) <= a;
    layer1_outputs(9674) <= not (a or b);
    layer1_outputs(9675) <= b;
    layer1_outputs(9676) <= not (a and b);
    layer1_outputs(9677) <= '0';
    layer1_outputs(9678) <= not (a or b);
    layer1_outputs(9679) <= not (a xor b);
    layer1_outputs(9680) <= not a;
    layer1_outputs(9681) <= b and not a;
    layer1_outputs(9682) <= a xor b;
    layer1_outputs(9683) <= not (a or b);
    layer1_outputs(9684) <= '1';
    layer1_outputs(9685) <= a;
    layer1_outputs(9686) <= a and not b;
    layer1_outputs(9687) <= not (a or b);
    layer1_outputs(9688) <= b;
    layer1_outputs(9689) <= not (a and b);
    layer1_outputs(9690) <= b and not a;
    layer1_outputs(9691) <= b and not a;
    layer1_outputs(9692) <= not a or b;
    layer1_outputs(9693) <= a and b;
    layer1_outputs(9694) <= '0';
    layer1_outputs(9695) <= a and not b;
    layer1_outputs(9696) <= not a or b;
    layer1_outputs(9697) <= not (a or b);
    layer1_outputs(9698) <= '0';
    layer1_outputs(9699) <= not (a or b);
    layer1_outputs(9700) <= not b;
    layer1_outputs(9701) <= a and b;
    layer1_outputs(9702) <= a or b;
    layer1_outputs(9703) <= not a or b;
    layer1_outputs(9704) <= b;
    layer1_outputs(9705) <= a;
    layer1_outputs(9706) <= not (a or b);
    layer1_outputs(9707) <= a and b;
    layer1_outputs(9708) <= not (a or b);
    layer1_outputs(9709) <= a and b;
    layer1_outputs(9710) <= not (a and b);
    layer1_outputs(9711) <= not (a and b);
    layer1_outputs(9712) <= not b;
    layer1_outputs(9713) <= b and not a;
    layer1_outputs(9714) <= a and not b;
    layer1_outputs(9715) <= not (a and b);
    layer1_outputs(9716) <= not b;
    layer1_outputs(9717) <= a xor b;
    layer1_outputs(9718) <= b;
    layer1_outputs(9719) <= not a;
    layer1_outputs(9720) <= not (a and b);
    layer1_outputs(9721) <= not a;
    layer1_outputs(9722) <= a and b;
    layer1_outputs(9723) <= b and not a;
    layer1_outputs(9724) <= b and not a;
    layer1_outputs(9725) <= not a;
    layer1_outputs(9726) <= not b;
    layer1_outputs(9727) <= '1';
    layer1_outputs(9728) <= not (a xor b);
    layer1_outputs(9729) <= b and not a;
    layer1_outputs(9730) <= a xor b;
    layer1_outputs(9731) <= '0';
    layer1_outputs(9732) <= a and b;
    layer1_outputs(9733) <= b and not a;
    layer1_outputs(9734) <= a;
    layer1_outputs(9735) <= a and b;
    layer1_outputs(9736) <= not (a or b);
    layer1_outputs(9737) <= a and not b;
    layer1_outputs(9738) <= not (a or b);
    layer1_outputs(9739) <= a and b;
    layer1_outputs(9740) <= a;
    layer1_outputs(9741) <= a;
    layer1_outputs(9742) <= not b;
    layer1_outputs(9743) <= b;
    layer1_outputs(9744) <= not b or a;
    layer1_outputs(9745) <= not (a and b);
    layer1_outputs(9746) <= a and not b;
    layer1_outputs(9747) <= not (a and b);
    layer1_outputs(9748) <= not b;
    layer1_outputs(9749) <= b;
    layer1_outputs(9750) <= not b;
    layer1_outputs(9751) <= b;
    layer1_outputs(9752) <= not a or b;
    layer1_outputs(9753) <= a or b;
    layer1_outputs(9754) <= not (a xor b);
    layer1_outputs(9755) <= not (a or b);
    layer1_outputs(9756) <= a xor b;
    layer1_outputs(9757) <= '1';
    layer1_outputs(9758) <= a and b;
    layer1_outputs(9759) <= not b or a;
    layer1_outputs(9760) <= not b;
    layer1_outputs(9761) <= b;
    layer1_outputs(9762) <= not b or a;
    layer1_outputs(9763) <= not (a and b);
    layer1_outputs(9764) <= b;
    layer1_outputs(9765) <= not a;
    layer1_outputs(9766) <= not b or a;
    layer1_outputs(9767) <= b;
    layer1_outputs(9768) <= a or b;
    layer1_outputs(9769) <= not b;
    layer1_outputs(9770) <= not a;
    layer1_outputs(9771) <= b;
    layer1_outputs(9772) <= '1';
    layer1_outputs(9773) <= not (a xor b);
    layer1_outputs(9774) <= not a;
    layer1_outputs(9775) <= '0';
    layer1_outputs(9776) <= a and b;
    layer1_outputs(9777) <= a;
    layer1_outputs(9778) <= not (a and b);
    layer1_outputs(9779) <= not a;
    layer1_outputs(9780) <= '0';
    layer1_outputs(9781) <= not a or b;
    layer1_outputs(9782) <= a and not b;
    layer1_outputs(9783) <= b and not a;
    layer1_outputs(9784) <= '1';
    layer1_outputs(9785) <= not (a xor b);
    layer1_outputs(9786) <= not (a or b);
    layer1_outputs(9787) <= not (a or b);
    layer1_outputs(9788) <= not (a and b);
    layer1_outputs(9789) <= not (a xor b);
    layer1_outputs(9790) <= b and not a;
    layer1_outputs(9791) <= a;
    layer1_outputs(9792) <= a and not b;
    layer1_outputs(9793) <= a and not b;
    layer1_outputs(9794) <= a;
    layer1_outputs(9795) <= not (a or b);
    layer1_outputs(9796) <= a;
    layer1_outputs(9797) <= a or b;
    layer1_outputs(9798) <= not (a xor b);
    layer1_outputs(9799) <= b and not a;
    layer1_outputs(9800) <= not b or a;
    layer1_outputs(9801) <= a and not b;
    layer1_outputs(9802) <= not b or a;
    layer1_outputs(9803) <= a;
    layer1_outputs(9804) <= not a or b;
    layer1_outputs(9805) <= not b or a;
    layer1_outputs(9806) <= b;
    layer1_outputs(9807) <= a xor b;
    layer1_outputs(9808) <= not b or a;
    layer1_outputs(9809) <= not (a and b);
    layer1_outputs(9810) <= not b;
    layer1_outputs(9811) <= a;
    layer1_outputs(9812) <= b and not a;
    layer1_outputs(9813) <= not (a and b);
    layer1_outputs(9814) <= '1';
    layer1_outputs(9815) <= a and not b;
    layer1_outputs(9816) <= a xor b;
    layer1_outputs(9817) <= a and b;
    layer1_outputs(9818) <= not b;
    layer1_outputs(9819) <= a;
    layer1_outputs(9820) <= a or b;
    layer1_outputs(9821) <= not b;
    layer1_outputs(9822) <= not (a xor b);
    layer1_outputs(9823) <= a;
    layer1_outputs(9824) <= b and not a;
    layer1_outputs(9825) <= not (a xor b);
    layer1_outputs(9826) <= a;
    layer1_outputs(9827) <= not a or b;
    layer1_outputs(9828) <= not a;
    layer1_outputs(9829) <= not (a or b);
    layer1_outputs(9830) <= a and b;
    layer1_outputs(9831) <= not (a or b);
    layer1_outputs(9832) <= not a;
    layer1_outputs(9833) <= not a or b;
    layer1_outputs(9834) <= not b;
    layer1_outputs(9835) <= '1';
    layer1_outputs(9836) <= not a or b;
    layer1_outputs(9837) <= b;
    layer1_outputs(9838) <= not b or a;
    layer1_outputs(9839) <= '1';
    layer1_outputs(9840) <= '1';
    layer1_outputs(9841) <= a and not b;
    layer1_outputs(9842) <= not a or b;
    layer1_outputs(9843) <= not b or a;
    layer1_outputs(9844) <= not a or b;
    layer1_outputs(9845) <= not a;
    layer1_outputs(9846) <= a and b;
    layer1_outputs(9847) <= a;
    layer1_outputs(9848) <= a or b;
    layer1_outputs(9849) <= a or b;
    layer1_outputs(9850) <= not a or b;
    layer1_outputs(9851) <= not b or a;
    layer1_outputs(9852) <= not b;
    layer1_outputs(9853) <= a;
    layer1_outputs(9854) <= a;
    layer1_outputs(9855) <= a;
    layer1_outputs(9856) <= not b;
    layer1_outputs(9857) <= not (a or b);
    layer1_outputs(9858) <= '0';
    layer1_outputs(9859) <= not a;
    layer1_outputs(9860) <= a and not b;
    layer1_outputs(9861) <= not b or a;
    layer1_outputs(9862) <= not a or b;
    layer1_outputs(9863) <= not b;
    layer1_outputs(9864) <= a xor b;
    layer1_outputs(9865) <= a;
    layer1_outputs(9866) <= b;
    layer1_outputs(9867) <= a xor b;
    layer1_outputs(9868) <= not b;
    layer1_outputs(9869) <= a or b;
    layer1_outputs(9870) <= a and not b;
    layer1_outputs(9871) <= a;
    layer1_outputs(9872) <= '1';
    layer1_outputs(9873) <= not b or a;
    layer1_outputs(9874) <= a;
    layer1_outputs(9875) <= not b;
    layer1_outputs(9876) <= not b;
    layer1_outputs(9877) <= '0';
    layer1_outputs(9878) <= b and not a;
    layer1_outputs(9879) <= not b;
    layer1_outputs(9880) <= not b or a;
    layer1_outputs(9881) <= not (a or b);
    layer1_outputs(9882) <= not a;
    layer1_outputs(9883) <= not a;
    layer1_outputs(9884) <= a or b;
    layer1_outputs(9885) <= not a;
    layer1_outputs(9886) <= a;
    layer1_outputs(9887) <= a and b;
    layer1_outputs(9888) <= not b;
    layer1_outputs(9889) <= a xor b;
    layer1_outputs(9890) <= a or b;
    layer1_outputs(9891) <= a or b;
    layer1_outputs(9892) <= a or b;
    layer1_outputs(9893) <= a and not b;
    layer1_outputs(9894) <= not a;
    layer1_outputs(9895) <= a or b;
    layer1_outputs(9896) <= not (a and b);
    layer1_outputs(9897) <= a and b;
    layer1_outputs(9898) <= b;
    layer1_outputs(9899) <= not (a or b);
    layer1_outputs(9900) <= '1';
    layer1_outputs(9901) <= b;
    layer1_outputs(9902) <= not a;
    layer1_outputs(9903) <= b;
    layer1_outputs(9904) <= not a;
    layer1_outputs(9905) <= not (a or b);
    layer1_outputs(9906) <= a or b;
    layer1_outputs(9907) <= a xor b;
    layer1_outputs(9908) <= b;
    layer1_outputs(9909) <= not b;
    layer1_outputs(9910) <= b;
    layer1_outputs(9911) <= b;
    layer1_outputs(9912) <= '1';
    layer1_outputs(9913) <= a or b;
    layer1_outputs(9914) <= not b or a;
    layer1_outputs(9915) <= not a;
    layer1_outputs(9916) <= not a or b;
    layer1_outputs(9917) <= not (a or b);
    layer1_outputs(9918) <= not b or a;
    layer1_outputs(9919) <= a and b;
    layer1_outputs(9920) <= not a or b;
    layer1_outputs(9921) <= not (a or b);
    layer1_outputs(9922) <= '1';
    layer1_outputs(9923) <= a and b;
    layer1_outputs(9924) <= b;
    layer1_outputs(9925) <= a xor b;
    layer1_outputs(9926) <= a xor b;
    layer1_outputs(9927) <= '0';
    layer1_outputs(9928) <= not a;
    layer1_outputs(9929) <= b and not a;
    layer1_outputs(9930) <= a xor b;
    layer1_outputs(9931) <= not b or a;
    layer1_outputs(9932) <= '0';
    layer1_outputs(9933) <= not b or a;
    layer1_outputs(9934) <= b and not a;
    layer1_outputs(9935) <= not a or b;
    layer1_outputs(9936) <= not b;
    layer1_outputs(9937) <= '1';
    layer1_outputs(9938) <= a and not b;
    layer1_outputs(9939) <= not b;
    layer1_outputs(9940) <= a and b;
    layer1_outputs(9941) <= '0';
    layer1_outputs(9942) <= not (a and b);
    layer1_outputs(9943) <= b and not a;
    layer1_outputs(9944) <= a xor b;
    layer1_outputs(9945) <= not a;
    layer1_outputs(9946) <= not (a or b);
    layer1_outputs(9947) <= a or b;
    layer1_outputs(9948) <= a xor b;
    layer1_outputs(9949) <= a xor b;
    layer1_outputs(9950) <= a or b;
    layer1_outputs(9951) <= not a or b;
    layer1_outputs(9952) <= a or b;
    layer1_outputs(9953) <= not a;
    layer1_outputs(9954) <= a xor b;
    layer1_outputs(9955) <= not a;
    layer1_outputs(9956) <= a and not b;
    layer1_outputs(9957) <= b;
    layer1_outputs(9958) <= not b;
    layer1_outputs(9959) <= a and not b;
    layer1_outputs(9960) <= not (a xor b);
    layer1_outputs(9961) <= not (a and b);
    layer1_outputs(9962) <= b;
    layer1_outputs(9963) <= not b;
    layer1_outputs(9964) <= a;
    layer1_outputs(9965) <= a;
    layer1_outputs(9966) <= a and not b;
    layer1_outputs(9967) <= a and b;
    layer1_outputs(9968) <= b and not a;
    layer1_outputs(9969) <= a and not b;
    layer1_outputs(9970) <= b;
    layer1_outputs(9971) <= not (a and b);
    layer1_outputs(9972) <= not b;
    layer1_outputs(9973) <= '1';
    layer1_outputs(9974) <= '0';
    layer1_outputs(9975) <= a and b;
    layer1_outputs(9976) <= '1';
    layer1_outputs(9977) <= a and b;
    layer1_outputs(9978) <= '1';
    layer1_outputs(9979) <= not (a or b);
    layer1_outputs(9980) <= b and not a;
    layer1_outputs(9981) <= not b;
    layer1_outputs(9982) <= a and not b;
    layer1_outputs(9983) <= a;
    layer1_outputs(9984) <= a;
    layer1_outputs(9985) <= not b;
    layer1_outputs(9986) <= b;
    layer1_outputs(9987) <= not b or a;
    layer1_outputs(9988) <= '1';
    layer1_outputs(9989) <= a and not b;
    layer1_outputs(9990) <= a and b;
    layer1_outputs(9991) <= not b or a;
    layer1_outputs(9992) <= not a;
    layer1_outputs(9993) <= a;
    layer1_outputs(9994) <= b;
    layer1_outputs(9995) <= not (a xor b);
    layer1_outputs(9996) <= not (a or b);
    layer1_outputs(9997) <= not a;
    layer1_outputs(9998) <= a or b;
    layer1_outputs(9999) <= b and not a;
    layer1_outputs(10000) <= not (a or b);
    layer1_outputs(10001) <= not b or a;
    layer1_outputs(10002) <= b;
    layer1_outputs(10003) <= not (a or b);
    layer1_outputs(10004) <= a and b;
    layer1_outputs(10005) <= a;
    layer1_outputs(10006) <= b and not a;
    layer1_outputs(10007) <= not a;
    layer1_outputs(10008) <= not b;
    layer1_outputs(10009) <= a or b;
    layer1_outputs(10010) <= '1';
    layer1_outputs(10011) <= b and not a;
    layer1_outputs(10012) <= not a or b;
    layer1_outputs(10013) <= '0';
    layer1_outputs(10014) <= a or b;
    layer1_outputs(10015) <= '0';
    layer1_outputs(10016) <= a;
    layer1_outputs(10017) <= b;
    layer1_outputs(10018) <= not (a or b);
    layer1_outputs(10019) <= not (a xor b);
    layer1_outputs(10020) <= a;
    layer1_outputs(10021) <= not (a and b);
    layer1_outputs(10022) <= not (a xor b);
    layer1_outputs(10023) <= not a;
    layer1_outputs(10024) <= not b or a;
    layer1_outputs(10025) <= not (a xor b);
    layer1_outputs(10026) <= '1';
    layer1_outputs(10027) <= b;
    layer1_outputs(10028) <= not (a xor b);
    layer1_outputs(10029) <= not b;
    layer1_outputs(10030) <= not a;
    layer1_outputs(10031) <= b and not a;
    layer1_outputs(10032) <= not a or b;
    layer1_outputs(10033) <= a and b;
    layer1_outputs(10034) <= '0';
    layer1_outputs(10035) <= a;
    layer1_outputs(10036) <= a;
    layer1_outputs(10037) <= b;
    layer1_outputs(10038) <= a xor b;
    layer1_outputs(10039) <= b and not a;
    layer1_outputs(10040) <= a or b;
    layer1_outputs(10041) <= not b or a;
    layer1_outputs(10042) <= not b;
    layer1_outputs(10043) <= a and b;
    layer1_outputs(10044) <= not (a or b);
    layer1_outputs(10045) <= a or b;
    layer1_outputs(10046) <= a;
    layer1_outputs(10047) <= b;
    layer1_outputs(10048) <= not (a and b);
    layer1_outputs(10049) <= not b;
    layer1_outputs(10050) <= b and not a;
    layer1_outputs(10051) <= a;
    layer1_outputs(10052) <= not b;
    layer1_outputs(10053) <= a and not b;
    layer1_outputs(10054) <= a xor b;
    layer1_outputs(10055) <= not (a or b);
    layer1_outputs(10056) <= not a or b;
    layer1_outputs(10057) <= not b or a;
    layer1_outputs(10058) <= not (a xor b);
    layer1_outputs(10059) <= not (a xor b);
    layer1_outputs(10060) <= not b;
    layer1_outputs(10061) <= a and not b;
    layer1_outputs(10062) <= a and b;
    layer1_outputs(10063) <= not (a xor b);
    layer1_outputs(10064) <= '0';
    layer1_outputs(10065) <= b;
    layer1_outputs(10066) <= not b or a;
    layer1_outputs(10067) <= '0';
    layer1_outputs(10068) <= not (a and b);
    layer1_outputs(10069) <= a and b;
    layer1_outputs(10070) <= not a;
    layer1_outputs(10071) <= a;
    layer1_outputs(10072) <= not a;
    layer1_outputs(10073) <= not b or a;
    layer1_outputs(10074) <= a xor b;
    layer1_outputs(10075) <= not b;
    layer1_outputs(10076) <= not b;
    layer1_outputs(10077) <= a;
    layer1_outputs(10078) <= b;
    layer1_outputs(10079) <= b;
    layer1_outputs(10080) <= '0';
    layer1_outputs(10081) <= not (a and b);
    layer1_outputs(10082) <= '0';
    layer1_outputs(10083) <= a and not b;
    layer1_outputs(10084) <= b and not a;
    layer1_outputs(10085) <= '1';
    layer1_outputs(10086) <= b and not a;
    layer1_outputs(10087) <= '0';
    layer1_outputs(10088) <= '1';
    layer1_outputs(10089) <= not (a and b);
    layer1_outputs(10090) <= '0';
    layer1_outputs(10091) <= a;
    layer1_outputs(10092) <= not a or b;
    layer1_outputs(10093) <= not a;
    layer1_outputs(10094) <= not a;
    layer1_outputs(10095) <= not (a xor b);
    layer1_outputs(10096) <= not (a or b);
    layer1_outputs(10097) <= not a;
    layer1_outputs(10098) <= not b;
    layer1_outputs(10099) <= a and not b;
    layer1_outputs(10100) <= not a or b;
    layer1_outputs(10101) <= not a or b;
    layer1_outputs(10102) <= b and not a;
    layer1_outputs(10103) <= b;
    layer1_outputs(10104) <= a;
    layer1_outputs(10105) <= a and not b;
    layer1_outputs(10106) <= b;
    layer1_outputs(10107) <= b;
    layer1_outputs(10108) <= a;
    layer1_outputs(10109) <= a xor b;
    layer1_outputs(10110) <= a and not b;
    layer1_outputs(10111) <= not (a or b);
    layer1_outputs(10112) <= '0';
    layer1_outputs(10113) <= b;
    layer1_outputs(10114) <= not a;
    layer1_outputs(10115) <= not b;
    layer1_outputs(10116) <= not (a and b);
    layer1_outputs(10117) <= not (a or b);
    layer1_outputs(10118) <= b and not a;
    layer1_outputs(10119) <= a and b;
    layer1_outputs(10120) <= not b or a;
    layer1_outputs(10121) <= '0';
    layer1_outputs(10122) <= '1';
    layer1_outputs(10123) <= a and b;
    layer1_outputs(10124) <= b;
    layer1_outputs(10125) <= '0';
    layer1_outputs(10126) <= a and b;
    layer1_outputs(10127) <= a or b;
    layer1_outputs(10128) <= a or b;
    layer1_outputs(10129) <= a;
    layer1_outputs(10130) <= b and not a;
    layer1_outputs(10131) <= a and b;
    layer1_outputs(10132) <= not b;
    layer1_outputs(10133) <= not b;
    layer1_outputs(10134) <= a or b;
    layer1_outputs(10135) <= not a;
    layer1_outputs(10136) <= '1';
    layer1_outputs(10137) <= a xor b;
    layer1_outputs(10138) <= b;
    layer1_outputs(10139) <= not a or b;
    layer1_outputs(10140) <= not b;
    layer1_outputs(10141) <= not b;
    layer1_outputs(10142) <= not (a or b);
    layer1_outputs(10143) <= not a or b;
    layer1_outputs(10144) <= not b;
    layer1_outputs(10145) <= not (a and b);
    layer1_outputs(10146) <= a;
    layer1_outputs(10147) <= not (a or b);
    layer1_outputs(10148) <= not b or a;
    layer1_outputs(10149) <= b and not a;
    layer1_outputs(10150) <= b;
    layer1_outputs(10151) <= a or b;
    layer1_outputs(10152) <= a or b;
    layer1_outputs(10153) <= a and not b;
    layer1_outputs(10154) <= not a or b;
    layer1_outputs(10155) <= not (a xor b);
    layer1_outputs(10156) <= '0';
    layer1_outputs(10157) <= a xor b;
    layer1_outputs(10158) <= not a or b;
    layer1_outputs(10159) <= not a or b;
    layer1_outputs(10160) <= b and not a;
    layer1_outputs(10161) <= not b or a;
    layer1_outputs(10162) <= a or b;
    layer1_outputs(10163) <= a and not b;
    layer1_outputs(10164) <= not (a xor b);
    layer1_outputs(10165) <= not a;
    layer1_outputs(10166) <= not (a and b);
    layer1_outputs(10167) <= '1';
    layer1_outputs(10168) <= a;
    layer1_outputs(10169) <= not a or b;
    layer1_outputs(10170) <= '1';
    layer1_outputs(10171) <= not b or a;
    layer1_outputs(10172) <= a;
    layer1_outputs(10173) <= '0';
    layer1_outputs(10174) <= not (a xor b);
    layer1_outputs(10175) <= '1';
    layer1_outputs(10176) <= a;
    layer1_outputs(10177) <= not (a and b);
    layer1_outputs(10178) <= not b;
    layer1_outputs(10179) <= b and not a;
    layer1_outputs(10180) <= not b;
    layer1_outputs(10181) <= '1';
    layer1_outputs(10182) <= a xor b;
    layer1_outputs(10183) <= not a or b;
    layer1_outputs(10184) <= b;
    layer1_outputs(10185) <= '0';
    layer1_outputs(10186) <= a and b;
    layer1_outputs(10187) <= a and not b;
    layer1_outputs(10188) <= not (a and b);
    layer1_outputs(10189) <= b;
    layer1_outputs(10190) <= a or b;
    layer1_outputs(10191) <= b;
    layer1_outputs(10192) <= not a;
    layer1_outputs(10193) <= a or b;
    layer1_outputs(10194) <= not a;
    layer1_outputs(10195) <= a;
    layer1_outputs(10196) <= not (a and b);
    layer1_outputs(10197) <= not a;
    layer1_outputs(10198) <= not (a xor b);
    layer1_outputs(10199) <= b and not a;
    layer1_outputs(10200) <= a and b;
    layer1_outputs(10201) <= a or b;
    layer1_outputs(10202) <= not b;
    layer1_outputs(10203) <= not a or b;
    layer1_outputs(10204) <= a and b;
    layer1_outputs(10205) <= a;
    layer1_outputs(10206) <= a and b;
    layer1_outputs(10207) <= a and b;
    layer1_outputs(10208) <= not b;
    layer1_outputs(10209) <= a and b;
    layer1_outputs(10210) <= not b;
    layer1_outputs(10211) <= not (a and b);
    layer1_outputs(10212) <= not a;
    layer1_outputs(10213) <= '1';
    layer1_outputs(10214) <= a;
    layer1_outputs(10215) <= not b or a;
    layer1_outputs(10216) <= not (a xor b);
    layer1_outputs(10217) <= a;
    layer1_outputs(10218) <= not (a and b);
    layer1_outputs(10219) <= '0';
    layer1_outputs(10220) <= a and b;
    layer1_outputs(10221) <= not (a xor b);
    layer1_outputs(10222) <= a and not b;
    layer1_outputs(10223) <= not (a or b);
    layer1_outputs(10224) <= not (a or b);
    layer1_outputs(10225) <= a and not b;
    layer1_outputs(10226) <= a and b;
    layer1_outputs(10227) <= not a or b;
    layer1_outputs(10228) <= a;
    layer1_outputs(10229) <= not a;
    layer1_outputs(10230) <= a or b;
    layer1_outputs(10231) <= not a or b;
    layer1_outputs(10232) <= b and not a;
    layer1_outputs(10233) <= a and b;
    layer1_outputs(10234) <= b and not a;
    layer1_outputs(10235) <= not (a and b);
    layer1_outputs(10236) <= a and not b;
    layer1_outputs(10237) <= a;
    layer1_outputs(10238) <= not b or a;
    layer1_outputs(10239) <= '1';
    layer2_outputs(0) <= '1';
    layer2_outputs(1) <= a;
    layer2_outputs(2) <= b;
    layer2_outputs(3) <= not (a xor b);
    layer2_outputs(4) <= not a or b;
    layer2_outputs(5) <= not (a and b);
    layer2_outputs(6) <= '1';
    layer2_outputs(7) <= a;
    layer2_outputs(8) <= a and b;
    layer2_outputs(9) <= b;
    layer2_outputs(10) <= not (a and b);
    layer2_outputs(11) <= not b or a;
    layer2_outputs(12) <= not b;
    layer2_outputs(13) <= a;
    layer2_outputs(14) <= not (a xor b);
    layer2_outputs(15) <= not a or b;
    layer2_outputs(16) <= a;
    layer2_outputs(17) <= b and not a;
    layer2_outputs(18) <= not b;
    layer2_outputs(19) <= a and b;
    layer2_outputs(20) <= not b or a;
    layer2_outputs(21) <= not b or a;
    layer2_outputs(22) <= not a or b;
    layer2_outputs(23) <= '0';
    layer2_outputs(24) <= not b;
    layer2_outputs(25) <= a or b;
    layer2_outputs(26) <= not b;
    layer2_outputs(27) <= a and not b;
    layer2_outputs(28) <= '1';
    layer2_outputs(29) <= b;
    layer2_outputs(30) <= not (a xor b);
    layer2_outputs(31) <= not (a and b);
    layer2_outputs(32) <= not (a and b);
    layer2_outputs(33) <= not (a xor b);
    layer2_outputs(34) <= not b;
    layer2_outputs(35) <= a;
    layer2_outputs(36) <= '0';
    layer2_outputs(37) <= not b;
    layer2_outputs(38) <= not b or a;
    layer2_outputs(39) <= not b;
    layer2_outputs(40) <= not a;
    layer2_outputs(41) <= a xor b;
    layer2_outputs(42) <= b;
    layer2_outputs(43) <= not a;
    layer2_outputs(44) <= a xor b;
    layer2_outputs(45) <= b and not a;
    layer2_outputs(46) <= a;
    layer2_outputs(47) <= not a or b;
    layer2_outputs(48) <= not (a or b);
    layer2_outputs(49) <= not (a or b);
    layer2_outputs(50) <= a;
    layer2_outputs(51) <= a and b;
    layer2_outputs(52) <= not (a and b);
    layer2_outputs(53) <= not a or b;
    layer2_outputs(54) <= not (a or b);
    layer2_outputs(55) <= a and b;
    layer2_outputs(56) <= b;
    layer2_outputs(57) <= b;
    layer2_outputs(58) <= not (a or b);
    layer2_outputs(59) <= b;
    layer2_outputs(60) <= a xor b;
    layer2_outputs(61) <= not (a or b);
    layer2_outputs(62) <= b and not a;
    layer2_outputs(63) <= not b or a;
    layer2_outputs(64) <= not b;
    layer2_outputs(65) <= a and b;
    layer2_outputs(66) <= b;
    layer2_outputs(67) <= not b;
    layer2_outputs(68) <= not b;
    layer2_outputs(69) <= b and not a;
    layer2_outputs(70) <= b;
    layer2_outputs(71) <= not (a and b);
    layer2_outputs(72) <= not a;
    layer2_outputs(73) <= a and not b;
    layer2_outputs(74) <= not (a and b);
    layer2_outputs(75) <= b and not a;
    layer2_outputs(76) <= a and b;
    layer2_outputs(77) <= not (a and b);
    layer2_outputs(78) <= a or b;
    layer2_outputs(79) <= a or b;
    layer2_outputs(80) <= not b;
    layer2_outputs(81) <= a xor b;
    layer2_outputs(82) <= '1';
    layer2_outputs(83) <= b;
    layer2_outputs(84) <= not b;
    layer2_outputs(85) <= not a or b;
    layer2_outputs(86) <= not a or b;
    layer2_outputs(87) <= not (a xor b);
    layer2_outputs(88) <= not a or b;
    layer2_outputs(89) <= not b or a;
    layer2_outputs(90) <= not a or b;
    layer2_outputs(91) <= '1';
    layer2_outputs(92) <= a and b;
    layer2_outputs(93) <= a or b;
    layer2_outputs(94) <= '1';
    layer2_outputs(95) <= a;
    layer2_outputs(96) <= '1';
    layer2_outputs(97) <= not (a and b);
    layer2_outputs(98) <= a and not b;
    layer2_outputs(99) <= a;
    layer2_outputs(100) <= a;
    layer2_outputs(101) <= '0';
    layer2_outputs(102) <= not b;
    layer2_outputs(103) <= '1';
    layer2_outputs(104) <= not (a and b);
    layer2_outputs(105) <= a;
    layer2_outputs(106) <= a and b;
    layer2_outputs(107) <= b and not a;
    layer2_outputs(108) <= not b;
    layer2_outputs(109) <= '1';
    layer2_outputs(110) <= a and b;
    layer2_outputs(111) <= not b;
    layer2_outputs(112) <= not b or a;
    layer2_outputs(113) <= not a or b;
    layer2_outputs(114) <= not a;
    layer2_outputs(115) <= not a or b;
    layer2_outputs(116) <= not a or b;
    layer2_outputs(117) <= a;
    layer2_outputs(118) <= a;
    layer2_outputs(119) <= a and b;
    layer2_outputs(120) <= not (a and b);
    layer2_outputs(121) <= a and b;
    layer2_outputs(122) <= a and b;
    layer2_outputs(123) <= '1';
    layer2_outputs(124) <= a or b;
    layer2_outputs(125) <= not a;
    layer2_outputs(126) <= b;
    layer2_outputs(127) <= a and not b;
    layer2_outputs(128) <= not (a or b);
    layer2_outputs(129) <= not a or b;
    layer2_outputs(130) <= a and not b;
    layer2_outputs(131) <= a or b;
    layer2_outputs(132) <= not b;
    layer2_outputs(133) <= not a;
    layer2_outputs(134) <= b;
    layer2_outputs(135) <= not (a or b);
    layer2_outputs(136) <= a xor b;
    layer2_outputs(137) <= a xor b;
    layer2_outputs(138) <= a and b;
    layer2_outputs(139) <= a and not b;
    layer2_outputs(140) <= a or b;
    layer2_outputs(141) <= not (a or b);
    layer2_outputs(142) <= b and not a;
    layer2_outputs(143) <= not (a and b);
    layer2_outputs(144) <= b;
    layer2_outputs(145) <= b and not a;
    layer2_outputs(146) <= '1';
    layer2_outputs(147) <= not b;
    layer2_outputs(148) <= not (a and b);
    layer2_outputs(149) <= a xor b;
    layer2_outputs(150) <= b and not a;
    layer2_outputs(151) <= not (a and b);
    layer2_outputs(152) <= not a or b;
    layer2_outputs(153) <= not (a or b);
    layer2_outputs(154) <= a and b;
    layer2_outputs(155) <= not (a or b);
    layer2_outputs(156) <= a and not b;
    layer2_outputs(157) <= not a or b;
    layer2_outputs(158) <= a and not b;
    layer2_outputs(159) <= a;
    layer2_outputs(160) <= a and b;
    layer2_outputs(161) <= b;
    layer2_outputs(162) <= '1';
    layer2_outputs(163) <= not a;
    layer2_outputs(164) <= a or b;
    layer2_outputs(165) <= b;
    layer2_outputs(166) <= a or b;
    layer2_outputs(167) <= not a or b;
    layer2_outputs(168) <= '0';
    layer2_outputs(169) <= a and b;
    layer2_outputs(170) <= not (a and b);
    layer2_outputs(171) <= not (a and b);
    layer2_outputs(172) <= a;
    layer2_outputs(173) <= a and not b;
    layer2_outputs(174) <= a and b;
    layer2_outputs(175) <= '0';
    layer2_outputs(176) <= not a or b;
    layer2_outputs(177) <= b;
    layer2_outputs(178) <= b;
    layer2_outputs(179) <= '0';
    layer2_outputs(180) <= not b;
    layer2_outputs(181) <= not a;
    layer2_outputs(182) <= b;
    layer2_outputs(183) <= not a;
    layer2_outputs(184) <= not b;
    layer2_outputs(185) <= not b;
    layer2_outputs(186) <= not a;
    layer2_outputs(187) <= not b or a;
    layer2_outputs(188) <= not b;
    layer2_outputs(189) <= not (a and b);
    layer2_outputs(190) <= not a or b;
    layer2_outputs(191) <= '0';
    layer2_outputs(192) <= a or b;
    layer2_outputs(193) <= a;
    layer2_outputs(194) <= '1';
    layer2_outputs(195) <= a or b;
    layer2_outputs(196) <= b;
    layer2_outputs(197) <= a or b;
    layer2_outputs(198) <= not a;
    layer2_outputs(199) <= not b or a;
    layer2_outputs(200) <= b;
    layer2_outputs(201) <= a or b;
    layer2_outputs(202) <= not b or a;
    layer2_outputs(203) <= not a;
    layer2_outputs(204) <= not a;
    layer2_outputs(205) <= b and not a;
    layer2_outputs(206) <= not (a xor b);
    layer2_outputs(207) <= a;
    layer2_outputs(208) <= not b;
    layer2_outputs(209) <= b;
    layer2_outputs(210) <= '0';
    layer2_outputs(211) <= a or b;
    layer2_outputs(212) <= a;
    layer2_outputs(213) <= a;
    layer2_outputs(214) <= a xor b;
    layer2_outputs(215) <= not (a or b);
    layer2_outputs(216) <= not a or b;
    layer2_outputs(217) <= '1';
    layer2_outputs(218) <= a or b;
    layer2_outputs(219) <= '1';
    layer2_outputs(220) <= '0';
    layer2_outputs(221) <= not b;
    layer2_outputs(222) <= not (a or b);
    layer2_outputs(223) <= a;
    layer2_outputs(224) <= b;
    layer2_outputs(225) <= not a or b;
    layer2_outputs(226) <= b and not a;
    layer2_outputs(227) <= a and b;
    layer2_outputs(228) <= b;
    layer2_outputs(229) <= b;
    layer2_outputs(230) <= not b;
    layer2_outputs(231) <= not b or a;
    layer2_outputs(232) <= not b or a;
    layer2_outputs(233) <= b;
    layer2_outputs(234) <= not b or a;
    layer2_outputs(235) <= '1';
    layer2_outputs(236) <= a;
    layer2_outputs(237) <= not (a or b);
    layer2_outputs(238) <= '1';
    layer2_outputs(239) <= b;
    layer2_outputs(240) <= b;
    layer2_outputs(241) <= b;
    layer2_outputs(242) <= not (a xor b);
    layer2_outputs(243) <= a and b;
    layer2_outputs(244) <= a;
    layer2_outputs(245) <= a and not b;
    layer2_outputs(246) <= not (a or b);
    layer2_outputs(247) <= a and not b;
    layer2_outputs(248) <= '1';
    layer2_outputs(249) <= a xor b;
    layer2_outputs(250) <= a xor b;
    layer2_outputs(251) <= a;
    layer2_outputs(252) <= a or b;
    layer2_outputs(253) <= a xor b;
    layer2_outputs(254) <= a or b;
    layer2_outputs(255) <= not (a or b);
    layer2_outputs(256) <= not b;
    layer2_outputs(257) <= b and not a;
    layer2_outputs(258) <= a xor b;
    layer2_outputs(259) <= a and not b;
    layer2_outputs(260) <= '0';
    layer2_outputs(261) <= a xor b;
    layer2_outputs(262) <= '0';
    layer2_outputs(263) <= not b or a;
    layer2_outputs(264) <= not a or b;
    layer2_outputs(265) <= not (a and b);
    layer2_outputs(266) <= not (a and b);
    layer2_outputs(267) <= not b;
    layer2_outputs(268) <= not b or a;
    layer2_outputs(269) <= not (a or b);
    layer2_outputs(270) <= '1';
    layer2_outputs(271) <= not (a and b);
    layer2_outputs(272) <= a and b;
    layer2_outputs(273) <= not a;
    layer2_outputs(274) <= a;
    layer2_outputs(275) <= not a;
    layer2_outputs(276) <= not (a or b);
    layer2_outputs(277) <= not a;
    layer2_outputs(278) <= not a;
    layer2_outputs(279) <= not b;
    layer2_outputs(280) <= not (a xor b);
    layer2_outputs(281) <= b;
    layer2_outputs(282) <= not a;
    layer2_outputs(283) <= not a or b;
    layer2_outputs(284) <= not b or a;
    layer2_outputs(285) <= a and b;
    layer2_outputs(286) <= a and b;
    layer2_outputs(287) <= not b;
    layer2_outputs(288) <= b and not a;
    layer2_outputs(289) <= not b or a;
    layer2_outputs(290) <= not (a and b);
    layer2_outputs(291) <= a and b;
    layer2_outputs(292) <= not b or a;
    layer2_outputs(293) <= not b;
    layer2_outputs(294) <= not b;
    layer2_outputs(295) <= b and not a;
    layer2_outputs(296) <= a;
    layer2_outputs(297) <= not a;
    layer2_outputs(298) <= '0';
    layer2_outputs(299) <= not (a or b);
    layer2_outputs(300) <= not a;
    layer2_outputs(301) <= '1';
    layer2_outputs(302) <= not b or a;
    layer2_outputs(303) <= not b or a;
    layer2_outputs(304) <= b and not a;
    layer2_outputs(305) <= '1';
    layer2_outputs(306) <= not (a or b);
    layer2_outputs(307) <= a and not b;
    layer2_outputs(308) <= not (a and b);
    layer2_outputs(309) <= b;
    layer2_outputs(310) <= not a or b;
    layer2_outputs(311) <= not b;
    layer2_outputs(312) <= a or b;
    layer2_outputs(313) <= not a;
    layer2_outputs(314) <= a;
    layer2_outputs(315) <= not a;
    layer2_outputs(316) <= a;
    layer2_outputs(317) <= not (a and b);
    layer2_outputs(318) <= not b;
    layer2_outputs(319) <= a and b;
    layer2_outputs(320) <= a or b;
    layer2_outputs(321) <= b and not a;
    layer2_outputs(322) <= b;
    layer2_outputs(323) <= a or b;
    layer2_outputs(324) <= not a or b;
    layer2_outputs(325) <= a and not b;
    layer2_outputs(326) <= not (a or b);
    layer2_outputs(327) <= a xor b;
    layer2_outputs(328) <= a or b;
    layer2_outputs(329) <= not (a or b);
    layer2_outputs(330) <= not a;
    layer2_outputs(331) <= not a or b;
    layer2_outputs(332) <= b;
    layer2_outputs(333) <= a and not b;
    layer2_outputs(334) <= b;
    layer2_outputs(335) <= not (a or b);
    layer2_outputs(336) <= a or b;
    layer2_outputs(337) <= a and not b;
    layer2_outputs(338) <= '0';
    layer2_outputs(339) <= not b;
    layer2_outputs(340) <= not (a xor b);
    layer2_outputs(341) <= a and not b;
    layer2_outputs(342) <= not (a or b);
    layer2_outputs(343) <= not (a xor b);
    layer2_outputs(344) <= a;
    layer2_outputs(345) <= a;
    layer2_outputs(346) <= b and not a;
    layer2_outputs(347) <= not (a or b);
    layer2_outputs(348) <= a;
    layer2_outputs(349) <= '0';
    layer2_outputs(350) <= not b;
    layer2_outputs(351) <= not a or b;
    layer2_outputs(352) <= not (a xor b);
    layer2_outputs(353) <= a and not b;
    layer2_outputs(354) <= a;
    layer2_outputs(355) <= '0';
    layer2_outputs(356) <= not a or b;
    layer2_outputs(357) <= b;
    layer2_outputs(358) <= not a or b;
    layer2_outputs(359) <= b;
    layer2_outputs(360) <= b;
    layer2_outputs(361) <= b;
    layer2_outputs(362) <= not a;
    layer2_outputs(363) <= not b;
    layer2_outputs(364) <= not b;
    layer2_outputs(365) <= '0';
    layer2_outputs(366) <= not (a xor b);
    layer2_outputs(367) <= not b;
    layer2_outputs(368) <= '0';
    layer2_outputs(369) <= b;
    layer2_outputs(370) <= a;
    layer2_outputs(371) <= a xor b;
    layer2_outputs(372) <= b;
    layer2_outputs(373) <= not (a or b);
    layer2_outputs(374) <= a;
    layer2_outputs(375) <= not (a and b);
    layer2_outputs(376) <= a;
    layer2_outputs(377) <= b;
    layer2_outputs(378) <= '1';
    layer2_outputs(379) <= b;
    layer2_outputs(380) <= '1';
    layer2_outputs(381) <= b and not a;
    layer2_outputs(382) <= not a;
    layer2_outputs(383) <= not (a or b);
    layer2_outputs(384) <= not (a or b);
    layer2_outputs(385) <= b and not a;
    layer2_outputs(386) <= a;
    layer2_outputs(387) <= a;
    layer2_outputs(388) <= a and b;
    layer2_outputs(389) <= not a;
    layer2_outputs(390) <= a or b;
    layer2_outputs(391) <= not a;
    layer2_outputs(392) <= not (a xor b);
    layer2_outputs(393) <= not b or a;
    layer2_outputs(394) <= a and b;
    layer2_outputs(395) <= not b;
    layer2_outputs(396) <= not (a xor b);
    layer2_outputs(397) <= not a or b;
    layer2_outputs(398) <= not a;
    layer2_outputs(399) <= not (a and b);
    layer2_outputs(400) <= '0';
    layer2_outputs(401) <= a or b;
    layer2_outputs(402) <= a and b;
    layer2_outputs(403) <= '1';
    layer2_outputs(404) <= b;
    layer2_outputs(405) <= not a;
    layer2_outputs(406) <= not (a xor b);
    layer2_outputs(407) <= a;
    layer2_outputs(408) <= not a;
    layer2_outputs(409) <= '0';
    layer2_outputs(410) <= not b or a;
    layer2_outputs(411) <= a and not b;
    layer2_outputs(412) <= a or b;
    layer2_outputs(413) <= not b or a;
    layer2_outputs(414) <= not a;
    layer2_outputs(415) <= b and not a;
    layer2_outputs(416) <= not (a or b);
    layer2_outputs(417) <= '0';
    layer2_outputs(418) <= a or b;
    layer2_outputs(419) <= a;
    layer2_outputs(420) <= not a;
    layer2_outputs(421) <= b and not a;
    layer2_outputs(422) <= not b or a;
    layer2_outputs(423) <= b and not a;
    layer2_outputs(424) <= a and not b;
    layer2_outputs(425) <= not b;
    layer2_outputs(426) <= a and b;
    layer2_outputs(427) <= not b;
    layer2_outputs(428) <= a and b;
    layer2_outputs(429) <= '1';
    layer2_outputs(430) <= not b or a;
    layer2_outputs(431) <= not b;
    layer2_outputs(432) <= b;
    layer2_outputs(433) <= not (a or b);
    layer2_outputs(434) <= not b;
    layer2_outputs(435) <= not b;
    layer2_outputs(436) <= not (a or b);
    layer2_outputs(437) <= b;
    layer2_outputs(438) <= not (a or b);
    layer2_outputs(439) <= a and not b;
    layer2_outputs(440) <= '1';
    layer2_outputs(441) <= a or b;
    layer2_outputs(442) <= b;
    layer2_outputs(443) <= not b;
    layer2_outputs(444) <= not a or b;
    layer2_outputs(445) <= '0';
    layer2_outputs(446) <= not b;
    layer2_outputs(447) <= not a;
    layer2_outputs(448) <= not (a or b);
    layer2_outputs(449) <= '0';
    layer2_outputs(450) <= a;
    layer2_outputs(451) <= '0';
    layer2_outputs(452) <= not b or a;
    layer2_outputs(453) <= b;
    layer2_outputs(454) <= a or b;
    layer2_outputs(455) <= a and b;
    layer2_outputs(456) <= a and not b;
    layer2_outputs(457) <= a and b;
    layer2_outputs(458) <= not a;
    layer2_outputs(459) <= b;
    layer2_outputs(460) <= '1';
    layer2_outputs(461) <= not a or b;
    layer2_outputs(462) <= a xor b;
    layer2_outputs(463) <= not (a and b);
    layer2_outputs(464) <= not a;
    layer2_outputs(465) <= '0';
    layer2_outputs(466) <= not a or b;
    layer2_outputs(467) <= a or b;
    layer2_outputs(468) <= not b;
    layer2_outputs(469) <= not (a or b);
    layer2_outputs(470) <= a;
    layer2_outputs(471) <= a or b;
    layer2_outputs(472) <= not b or a;
    layer2_outputs(473) <= not b or a;
    layer2_outputs(474) <= b;
    layer2_outputs(475) <= not a;
    layer2_outputs(476) <= a xor b;
    layer2_outputs(477) <= b;
    layer2_outputs(478) <= not b;
    layer2_outputs(479) <= not (a or b);
    layer2_outputs(480) <= not (a and b);
    layer2_outputs(481) <= not a;
    layer2_outputs(482) <= a;
    layer2_outputs(483) <= not b;
    layer2_outputs(484) <= '0';
    layer2_outputs(485) <= not b;
    layer2_outputs(486) <= '0';
    layer2_outputs(487) <= a and b;
    layer2_outputs(488) <= a and b;
    layer2_outputs(489) <= not (a or b);
    layer2_outputs(490) <= not (a and b);
    layer2_outputs(491) <= a and b;
    layer2_outputs(492) <= not a or b;
    layer2_outputs(493) <= a and b;
    layer2_outputs(494) <= '1';
    layer2_outputs(495) <= b;
    layer2_outputs(496) <= not (a and b);
    layer2_outputs(497) <= not b;
    layer2_outputs(498) <= not a;
    layer2_outputs(499) <= not a or b;
    layer2_outputs(500) <= not b or a;
    layer2_outputs(501) <= not (a and b);
    layer2_outputs(502) <= a and b;
    layer2_outputs(503) <= not a or b;
    layer2_outputs(504) <= not (a and b);
    layer2_outputs(505) <= '0';
    layer2_outputs(506) <= '0';
    layer2_outputs(507) <= b;
    layer2_outputs(508) <= a;
    layer2_outputs(509) <= not b;
    layer2_outputs(510) <= not b or a;
    layer2_outputs(511) <= a;
    layer2_outputs(512) <= a;
    layer2_outputs(513) <= not (a and b);
    layer2_outputs(514) <= not b or a;
    layer2_outputs(515) <= a xor b;
    layer2_outputs(516) <= b and not a;
    layer2_outputs(517) <= a and not b;
    layer2_outputs(518) <= a or b;
    layer2_outputs(519) <= not a;
    layer2_outputs(520) <= not a;
    layer2_outputs(521) <= not (a or b);
    layer2_outputs(522) <= b;
    layer2_outputs(523) <= '0';
    layer2_outputs(524) <= a;
    layer2_outputs(525) <= not a or b;
    layer2_outputs(526) <= not (a or b);
    layer2_outputs(527) <= not a;
    layer2_outputs(528) <= a xor b;
    layer2_outputs(529) <= not (a xor b);
    layer2_outputs(530) <= '1';
    layer2_outputs(531) <= not a;
    layer2_outputs(532) <= not (a and b);
    layer2_outputs(533) <= a or b;
    layer2_outputs(534) <= not (a or b);
    layer2_outputs(535) <= not a;
    layer2_outputs(536) <= a and not b;
    layer2_outputs(537) <= '1';
    layer2_outputs(538) <= not b;
    layer2_outputs(539) <= not a or b;
    layer2_outputs(540) <= b;
    layer2_outputs(541) <= '0';
    layer2_outputs(542) <= not a or b;
    layer2_outputs(543) <= not (a xor b);
    layer2_outputs(544) <= not (a xor b);
    layer2_outputs(545) <= not (a or b);
    layer2_outputs(546) <= not b or a;
    layer2_outputs(547) <= a or b;
    layer2_outputs(548) <= b;
    layer2_outputs(549) <= '1';
    layer2_outputs(550) <= not b or a;
    layer2_outputs(551) <= not a;
    layer2_outputs(552) <= a and b;
    layer2_outputs(553) <= a and not b;
    layer2_outputs(554) <= b and not a;
    layer2_outputs(555) <= not b;
    layer2_outputs(556) <= not b or a;
    layer2_outputs(557) <= '1';
    layer2_outputs(558) <= not (a and b);
    layer2_outputs(559) <= '1';
    layer2_outputs(560) <= a and b;
    layer2_outputs(561) <= not (a and b);
    layer2_outputs(562) <= not a or b;
    layer2_outputs(563) <= not a;
    layer2_outputs(564) <= b and not a;
    layer2_outputs(565) <= not (a or b);
    layer2_outputs(566) <= '0';
    layer2_outputs(567) <= not b or a;
    layer2_outputs(568) <= a xor b;
    layer2_outputs(569) <= a;
    layer2_outputs(570) <= b;
    layer2_outputs(571) <= not (a and b);
    layer2_outputs(572) <= not (a or b);
    layer2_outputs(573) <= b;
    layer2_outputs(574) <= b;
    layer2_outputs(575) <= not b or a;
    layer2_outputs(576) <= '0';
    layer2_outputs(577) <= b;
    layer2_outputs(578) <= '0';
    layer2_outputs(579) <= b and not a;
    layer2_outputs(580) <= not a;
    layer2_outputs(581) <= not b;
    layer2_outputs(582) <= not b or a;
    layer2_outputs(583) <= b and not a;
    layer2_outputs(584) <= not a;
    layer2_outputs(585) <= not b;
    layer2_outputs(586) <= a or b;
    layer2_outputs(587) <= not b;
    layer2_outputs(588) <= not (a or b);
    layer2_outputs(589) <= '1';
    layer2_outputs(590) <= not b or a;
    layer2_outputs(591) <= not a or b;
    layer2_outputs(592) <= a or b;
    layer2_outputs(593) <= a or b;
    layer2_outputs(594) <= a;
    layer2_outputs(595) <= not b or a;
    layer2_outputs(596) <= not a or b;
    layer2_outputs(597) <= a and b;
    layer2_outputs(598) <= a or b;
    layer2_outputs(599) <= not (a or b);
    layer2_outputs(600) <= '1';
    layer2_outputs(601) <= not a;
    layer2_outputs(602) <= a and b;
    layer2_outputs(603) <= '1';
    layer2_outputs(604) <= not a or b;
    layer2_outputs(605) <= not b;
    layer2_outputs(606) <= '0';
    layer2_outputs(607) <= a;
    layer2_outputs(608) <= a and b;
    layer2_outputs(609) <= not (a and b);
    layer2_outputs(610) <= not a or b;
    layer2_outputs(611) <= b and not a;
    layer2_outputs(612) <= not (a and b);
    layer2_outputs(613) <= not b or a;
    layer2_outputs(614) <= not a or b;
    layer2_outputs(615) <= '1';
    layer2_outputs(616) <= a and not b;
    layer2_outputs(617) <= a;
    layer2_outputs(618) <= not b or a;
    layer2_outputs(619) <= not (a and b);
    layer2_outputs(620) <= not (a and b);
    layer2_outputs(621) <= '1';
    layer2_outputs(622) <= not b or a;
    layer2_outputs(623) <= a;
    layer2_outputs(624) <= not b or a;
    layer2_outputs(625) <= b and not a;
    layer2_outputs(626) <= '1';
    layer2_outputs(627) <= b;
    layer2_outputs(628) <= b;
    layer2_outputs(629) <= a and b;
    layer2_outputs(630) <= not (a and b);
    layer2_outputs(631) <= a and not b;
    layer2_outputs(632) <= '1';
    layer2_outputs(633) <= not a or b;
    layer2_outputs(634) <= not b;
    layer2_outputs(635) <= not b or a;
    layer2_outputs(636) <= '1';
    layer2_outputs(637) <= not b or a;
    layer2_outputs(638) <= not (a or b);
    layer2_outputs(639) <= not b;
    layer2_outputs(640) <= a or b;
    layer2_outputs(641) <= not b or a;
    layer2_outputs(642) <= not (a xor b);
    layer2_outputs(643) <= a and not b;
    layer2_outputs(644) <= not b;
    layer2_outputs(645) <= b;
    layer2_outputs(646) <= '1';
    layer2_outputs(647) <= a and not b;
    layer2_outputs(648) <= a or b;
    layer2_outputs(649) <= '1';
    layer2_outputs(650) <= not a;
    layer2_outputs(651) <= not (a or b);
    layer2_outputs(652) <= not (a and b);
    layer2_outputs(653) <= a;
    layer2_outputs(654) <= not a;
    layer2_outputs(655) <= not a or b;
    layer2_outputs(656) <= a;
    layer2_outputs(657) <= not b;
    layer2_outputs(658) <= not b or a;
    layer2_outputs(659) <= not a;
    layer2_outputs(660) <= a and not b;
    layer2_outputs(661) <= not b or a;
    layer2_outputs(662) <= '1';
    layer2_outputs(663) <= '1';
    layer2_outputs(664) <= a or b;
    layer2_outputs(665) <= a and b;
    layer2_outputs(666) <= not b or a;
    layer2_outputs(667) <= not (a and b);
    layer2_outputs(668) <= not (a xor b);
    layer2_outputs(669) <= not (a xor b);
    layer2_outputs(670) <= not (a xor b);
    layer2_outputs(671) <= not b or a;
    layer2_outputs(672) <= not (a xor b);
    layer2_outputs(673) <= not a;
    layer2_outputs(674) <= not a;
    layer2_outputs(675) <= not a or b;
    layer2_outputs(676) <= not b;
    layer2_outputs(677) <= a and not b;
    layer2_outputs(678) <= not b;
    layer2_outputs(679) <= not b;
    layer2_outputs(680) <= b;
    layer2_outputs(681) <= a;
    layer2_outputs(682) <= not b;
    layer2_outputs(683) <= a;
    layer2_outputs(684) <= not (a or b);
    layer2_outputs(685) <= not b or a;
    layer2_outputs(686) <= a;
    layer2_outputs(687) <= '1';
    layer2_outputs(688) <= not (a xor b);
    layer2_outputs(689) <= b;
    layer2_outputs(690) <= a;
    layer2_outputs(691) <= not (a and b);
    layer2_outputs(692) <= '0';
    layer2_outputs(693) <= a and not b;
    layer2_outputs(694) <= not a or b;
    layer2_outputs(695) <= '1';
    layer2_outputs(696) <= not a or b;
    layer2_outputs(697) <= not (a and b);
    layer2_outputs(698) <= not a or b;
    layer2_outputs(699) <= not a;
    layer2_outputs(700) <= not b or a;
    layer2_outputs(701) <= not b;
    layer2_outputs(702) <= a or b;
    layer2_outputs(703) <= '1';
    layer2_outputs(704) <= not a;
    layer2_outputs(705) <= b;
    layer2_outputs(706) <= '1';
    layer2_outputs(707) <= b;
    layer2_outputs(708) <= a;
    layer2_outputs(709) <= a;
    layer2_outputs(710) <= not a;
    layer2_outputs(711) <= '1';
    layer2_outputs(712) <= b;
    layer2_outputs(713) <= a and b;
    layer2_outputs(714) <= b;
    layer2_outputs(715) <= a or b;
    layer2_outputs(716) <= not b or a;
    layer2_outputs(717) <= b;
    layer2_outputs(718) <= not b or a;
    layer2_outputs(719) <= not a or b;
    layer2_outputs(720) <= b and not a;
    layer2_outputs(721) <= not a or b;
    layer2_outputs(722) <= not b;
    layer2_outputs(723) <= not a;
    layer2_outputs(724) <= not (a and b);
    layer2_outputs(725) <= b;
    layer2_outputs(726) <= b and not a;
    layer2_outputs(727) <= a;
    layer2_outputs(728) <= not (a and b);
    layer2_outputs(729) <= a or b;
    layer2_outputs(730) <= not a;
    layer2_outputs(731) <= a;
    layer2_outputs(732) <= a and b;
    layer2_outputs(733) <= '0';
    layer2_outputs(734) <= a or b;
    layer2_outputs(735) <= b;
    layer2_outputs(736) <= b and not a;
    layer2_outputs(737) <= a;
    layer2_outputs(738) <= not b;
    layer2_outputs(739) <= b;
    layer2_outputs(740) <= a or b;
    layer2_outputs(741) <= not (a and b);
    layer2_outputs(742) <= b;
    layer2_outputs(743) <= a xor b;
    layer2_outputs(744) <= a or b;
    layer2_outputs(745) <= not b;
    layer2_outputs(746) <= not a;
    layer2_outputs(747) <= not (a and b);
    layer2_outputs(748) <= not a;
    layer2_outputs(749) <= not b or a;
    layer2_outputs(750) <= not (a and b);
    layer2_outputs(751) <= b;
    layer2_outputs(752) <= '0';
    layer2_outputs(753) <= not (a and b);
    layer2_outputs(754) <= a xor b;
    layer2_outputs(755) <= b and not a;
    layer2_outputs(756) <= b;
    layer2_outputs(757) <= not a or b;
    layer2_outputs(758) <= '1';
    layer2_outputs(759) <= a xor b;
    layer2_outputs(760) <= a;
    layer2_outputs(761) <= not a;
    layer2_outputs(762) <= not a;
    layer2_outputs(763) <= a or b;
    layer2_outputs(764) <= a xor b;
    layer2_outputs(765) <= b;
    layer2_outputs(766) <= not a;
    layer2_outputs(767) <= not a or b;
    layer2_outputs(768) <= not a;
    layer2_outputs(769) <= a and b;
    layer2_outputs(770) <= a xor b;
    layer2_outputs(771) <= not (a xor b);
    layer2_outputs(772) <= a and b;
    layer2_outputs(773) <= a and b;
    layer2_outputs(774) <= a xor b;
    layer2_outputs(775) <= a or b;
    layer2_outputs(776) <= b and not a;
    layer2_outputs(777) <= not a;
    layer2_outputs(778) <= '1';
    layer2_outputs(779) <= b and not a;
    layer2_outputs(780) <= not b;
    layer2_outputs(781) <= a and not b;
    layer2_outputs(782) <= not b or a;
    layer2_outputs(783) <= b and not a;
    layer2_outputs(784) <= not b;
    layer2_outputs(785) <= not (a xor b);
    layer2_outputs(786) <= b and not a;
    layer2_outputs(787) <= '0';
    layer2_outputs(788) <= not b or a;
    layer2_outputs(789) <= a and not b;
    layer2_outputs(790) <= not (a or b);
    layer2_outputs(791) <= not b or a;
    layer2_outputs(792) <= '0';
    layer2_outputs(793) <= not (a or b);
    layer2_outputs(794) <= a;
    layer2_outputs(795) <= not (a or b);
    layer2_outputs(796) <= not (a and b);
    layer2_outputs(797) <= b;
    layer2_outputs(798) <= a and not b;
    layer2_outputs(799) <= b and not a;
    layer2_outputs(800) <= a and b;
    layer2_outputs(801) <= not a;
    layer2_outputs(802) <= not (a xor b);
    layer2_outputs(803) <= '1';
    layer2_outputs(804) <= a xor b;
    layer2_outputs(805) <= a or b;
    layer2_outputs(806) <= a and not b;
    layer2_outputs(807) <= not (a and b);
    layer2_outputs(808) <= '0';
    layer2_outputs(809) <= a and b;
    layer2_outputs(810) <= a;
    layer2_outputs(811) <= '1';
    layer2_outputs(812) <= not b;
    layer2_outputs(813) <= '1';
    layer2_outputs(814) <= not a;
    layer2_outputs(815) <= a or b;
    layer2_outputs(816) <= '0';
    layer2_outputs(817) <= a and not b;
    layer2_outputs(818) <= b and not a;
    layer2_outputs(819) <= b;
    layer2_outputs(820) <= not b;
    layer2_outputs(821) <= '1';
    layer2_outputs(822) <= a;
    layer2_outputs(823) <= not a;
    layer2_outputs(824) <= '0';
    layer2_outputs(825) <= b and not a;
    layer2_outputs(826) <= '0';
    layer2_outputs(827) <= a;
    layer2_outputs(828) <= a;
    layer2_outputs(829) <= '1';
    layer2_outputs(830) <= '1';
    layer2_outputs(831) <= not a or b;
    layer2_outputs(832) <= a or b;
    layer2_outputs(833) <= b;
    layer2_outputs(834) <= not a;
    layer2_outputs(835) <= b and not a;
    layer2_outputs(836) <= a;
    layer2_outputs(837) <= not b or a;
    layer2_outputs(838) <= a;
    layer2_outputs(839) <= a or b;
    layer2_outputs(840) <= not b;
    layer2_outputs(841) <= a;
    layer2_outputs(842) <= not a;
    layer2_outputs(843) <= not b or a;
    layer2_outputs(844) <= not (a or b);
    layer2_outputs(845) <= not (a and b);
    layer2_outputs(846) <= a xor b;
    layer2_outputs(847) <= a and b;
    layer2_outputs(848) <= not b or a;
    layer2_outputs(849) <= b and not a;
    layer2_outputs(850) <= b and not a;
    layer2_outputs(851) <= not a or b;
    layer2_outputs(852) <= b and not a;
    layer2_outputs(853) <= '0';
    layer2_outputs(854) <= not b;
    layer2_outputs(855) <= '0';
    layer2_outputs(856) <= a;
    layer2_outputs(857) <= a;
    layer2_outputs(858) <= not b or a;
    layer2_outputs(859) <= '0';
    layer2_outputs(860) <= not (a or b);
    layer2_outputs(861) <= a and not b;
    layer2_outputs(862) <= not a;
    layer2_outputs(863) <= not a;
    layer2_outputs(864) <= b and not a;
    layer2_outputs(865) <= a or b;
    layer2_outputs(866) <= a;
    layer2_outputs(867) <= b;
    layer2_outputs(868) <= b and not a;
    layer2_outputs(869) <= a and b;
    layer2_outputs(870) <= not b;
    layer2_outputs(871) <= not (a xor b);
    layer2_outputs(872) <= not (a xor b);
    layer2_outputs(873) <= not (a xor b);
    layer2_outputs(874) <= not b;
    layer2_outputs(875) <= not a or b;
    layer2_outputs(876) <= not (a or b);
    layer2_outputs(877) <= a and b;
    layer2_outputs(878) <= not a;
    layer2_outputs(879) <= b;
    layer2_outputs(880) <= b;
    layer2_outputs(881) <= '1';
    layer2_outputs(882) <= b;
    layer2_outputs(883) <= b;
    layer2_outputs(884) <= not b;
    layer2_outputs(885) <= not b;
    layer2_outputs(886) <= not (a xor b);
    layer2_outputs(887) <= not a or b;
    layer2_outputs(888) <= not b;
    layer2_outputs(889) <= a;
    layer2_outputs(890) <= b;
    layer2_outputs(891) <= a and b;
    layer2_outputs(892) <= b;
    layer2_outputs(893) <= '1';
    layer2_outputs(894) <= a;
    layer2_outputs(895) <= a;
    layer2_outputs(896) <= '0';
    layer2_outputs(897) <= '0';
    layer2_outputs(898) <= '0';
    layer2_outputs(899) <= '1';
    layer2_outputs(900) <= not b or a;
    layer2_outputs(901) <= a and b;
    layer2_outputs(902) <= a and not b;
    layer2_outputs(903) <= a or b;
    layer2_outputs(904) <= not (a and b);
    layer2_outputs(905) <= not a or b;
    layer2_outputs(906) <= not b;
    layer2_outputs(907) <= a xor b;
    layer2_outputs(908) <= not (a and b);
    layer2_outputs(909) <= a and not b;
    layer2_outputs(910) <= a or b;
    layer2_outputs(911) <= a xor b;
    layer2_outputs(912) <= not (a or b);
    layer2_outputs(913) <= not (a and b);
    layer2_outputs(914) <= '1';
    layer2_outputs(915) <= a and b;
    layer2_outputs(916) <= not (a or b);
    layer2_outputs(917) <= not a or b;
    layer2_outputs(918) <= not b;
    layer2_outputs(919) <= '1';
    layer2_outputs(920) <= b;
    layer2_outputs(921) <= not (a or b);
    layer2_outputs(922) <= a;
    layer2_outputs(923) <= not b;
    layer2_outputs(924) <= not b or a;
    layer2_outputs(925) <= not (a or b);
    layer2_outputs(926) <= not a;
    layer2_outputs(927) <= not b or a;
    layer2_outputs(928) <= a;
    layer2_outputs(929) <= not a;
    layer2_outputs(930) <= a;
    layer2_outputs(931) <= a;
    layer2_outputs(932) <= a and not b;
    layer2_outputs(933) <= not (a xor b);
    layer2_outputs(934) <= a and b;
    layer2_outputs(935) <= not (a or b);
    layer2_outputs(936) <= a;
    layer2_outputs(937) <= a;
    layer2_outputs(938) <= a xor b;
    layer2_outputs(939) <= not a;
    layer2_outputs(940) <= not b;
    layer2_outputs(941) <= b;
    layer2_outputs(942) <= not a;
    layer2_outputs(943) <= a and not b;
    layer2_outputs(944) <= not a;
    layer2_outputs(945) <= not (a xor b);
    layer2_outputs(946) <= a and b;
    layer2_outputs(947) <= not a or b;
    layer2_outputs(948) <= not b;
    layer2_outputs(949) <= a and b;
    layer2_outputs(950) <= not a;
    layer2_outputs(951) <= '0';
    layer2_outputs(952) <= b and not a;
    layer2_outputs(953) <= not (a or b);
    layer2_outputs(954) <= '1';
    layer2_outputs(955) <= a and not b;
    layer2_outputs(956) <= '0';
    layer2_outputs(957) <= not a;
    layer2_outputs(958) <= a and b;
    layer2_outputs(959) <= not b or a;
    layer2_outputs(960) <= a;
    layer2_outputs(961) <= not b;
    layer2_outputs(962) <= '0';
    layer2_outputs(963) <= '0';
    layer2_outputs(964) <= not (a and b);
    layer2_outputs(965) <= a xor b;
    layer2_outputs(966) <= a and b;
    layer2_outputs(967) <= a;
    layer2_outputs(968) <= not (a and b);
    layer2_outputs(969) <= not (a and b);
    layer2_outputs(970) <= not b;
    layer2_outputs(971) <= not b;
    layer2_outputs(972) <= not a;
    layer2_outputs(973) <= not (a and b);
    layer2_outputs(974) <= a;
    layer2_outputs(975) <= not a or b;
    layer2_outputs(976) <= a;
    layer2_outputs(977) <= a and b;
    layer2_outputs(978) <= not (a and b);
    layer2_outputs(979) <= not a;
    layer2_outputs(980) <= not a;
    layer2_outputs(981) <= not (a xor b);
    layer2_outputs(982) <= b and not a;
    layer2_outputs(983) <= not b;
    layer2_outputs(984) <= a;
    layer2_outputs(985) <= not a;
    layer2_outputs(986) <= not (a xor b);
    layer2_outputs(987) <= a and not b;
    layer2_outputs(988) <= '1';
    layer2_outputs(989) <= '1';
    layer2_outputs(990) <= not b or a;
    layer2_outputs(991) <= not a;
    layer2_outputs(992) <= b and not a;
    layer2_outputs(993) <= not (a and b);
    layer2_outputs(994) <= '1';
    layer2_outputs(995) <= a or b;
    layer2_outputs(996) <= '0';
    layer2_outputs(997) <= not a or b;
    layer2_outputs(998) <= b and not a;
    layer2_outputs(999) <= a and b;
    layer2_outputs(1000) <= a;
    layer2_outputs(1001) <= not b or a;
    layer2_outputs(1002) <= not (a xor b);
    layer2_outputs(1003) <= b;
    layer2_outputs(1004) <= not a or b;
    layer2_outputs(1005) <= '0';
    layer2_outputs(1006) <= b and not a;
    layer2_outputs(1007) <= a xor b;
    layer2_outputs(1008) <= a and not b;
    layer2_outputs(1009) <= a and b;
    layer2_outputs(1010) <= not b or a;
    layer2_outputs(1011) <= b and not a;
    layer2_outputs(1012) <= a;
    layer2_outputs(1013) <= not a or b;
    layer2_outputs(1014) <= a or b;
    layer2_outputs(1015) <= not a;
    layer2_outputs(1016) <= not b or a;
    layer2_outputs(1017) <= not b or a;
    layer2_outputs(1018) <= a and not b;
    layer2_outputs(1019) <= not (a xor b);
    layer2_outputs(1020) <= '0';
    layer2_outputs(1021) <= not a or b;
    layer2_outputs(1022) <= not b;
    layer2_outputs(1023) <= not b or a;
    layer2_outputs(1024) <= a or b;
    layer2_outputs(1025) <= a xor b;
    layer2_outputs(1026) <= '0';
    layer2_outputs(1027) <= b;
    layer2_outputs(1028) <= not b;
    layer2_outputs(1029) <= a xor b;
    layer2_outputs(1030) <= b and not a;
    layer2_outputs(1031) <= not b;
    layer2_outputs(1032) <= '0';
    layer2_outputs(1033) <= '0';
    layer2_outputs(1034) <= not b or a;
    layer2_outputs(1035) <= not a;
    layer2_outputs(1036) <= '1';
    layer2_outputs(1037) <= not b or a;
    layer2_outputs(1038) <= a and not b;
    layer2_outputs(1039) <= not a;
    layer2_outputs(1040) <= not (a or b);
    layer2_outputs(1041) <= not (a xor b);
    layer2_outputs(1042) <= b;
    layer2_outputs(1043) <= not a;
    layer2_outputs(1044) <= b and not a;
    layer2_outputs(1045) <= a;
    layer2_outputs(1046) <= a and not b;
    layer2_outputs(1047) <= a;
    layer2_outputs(1048) <= not (a xor b);
    layer2_outputs(1049) <= not (a and b);
    layer2_outputs(1050) <= not (a and b);
    layer2_outputs(1051) <= not a or b;
    layer2_outputs(1052) <= a xor b;
    layer2_outputs(1053) <= not b or a;
    layer2_outputs(1054) <= not a;
    layer2_outputs(1055) <= a and not b;
    layer2_outputs(1056) <= '1';
    layer2_outputs(1057) <= a;
    layer2_outputs(1058) <= '0';
    layer2_outputs(1059) <= a or b;
    layer2_outputs(1060) <= not a or b;
    layer2_outputs(1061) <= '1';
    layer2_outputs(1062) <= '0';
    layer2_outputs(1063) <= not (a xor b);
    layer2_outputs(1064) <= b;
    layer2_outputs(1065) <= not (a and b);
    layer2_outputs(1066) <= not b;
    layer2_outputs(1067) <= not (a xor b);
    layer2_outputs(1068) <= not b or a;
    layer2_outputs(1069) <= '1';
    layer2_outputs(1070) <= b and not a;
    layer2_outputs(1071) <= not b;
    layer2_outputs(1072) <= '1';
    layer2_outputs(1073) <= '1';
    layer2_outputs(1074) <= b and not a;
    layer2_outputs(1075) <= a;
    layer2_outputs(1076) <= a and b;
    layer2_outputs(1077) <= not (a xor b);
    layer2_outputs(1078) <= a;
    layer2_outputs(1079) <= not a or b;
    layer2_outputs(1080) <= not a;
    layer2_outputs(1081) <= b;
    layer2_outputs(1082) <= not b;
    layer2_outputs(1083) <= b;
    layer2_outputs(1084) <= a and b;
    layer2_outputs(1085) <= not a;
    layer2_outputs(1086) <= a or b;
    layer2_outputs(1087) <= a and b;
    layer2_outputs(1088) <= not b or a;
    layer2_outputs(1089) <= not (a and b);
    layer2_outputs(1090) <= a and b;
    layer2_outputs(1091) <= a xor b;
    layer2_outputs(1092) <= '1';
    layer2_outputs(1093) <= not (a and b);
    layer2_outputs(1094) <= '1';
    layer2_outputs(1095) <= not (a and b);
    layer2_outputs(1096) <= a xor b;
    layer2_outputs(1097) <= b;
    layer2_outputs(1098) <= a and b;
    layer2_outputs(1099) <= a or b;
    layer2_outputs(1100) <= not (a or b);
    layer2_outputs(1101) <= a;
    layer2_outputs(1102) <= a and b;
    layer2_outputs(1103) <= not b or a;
    layer2_outputs(1104) <= b;
    layer2_outputs(1105) <= '1';
    layer2_outputs(1106) <= not b or a;
    layer2_outputs(1107) <= b;
    layer2_outputs(1108) <= a and not b;
    layer2_outputs(1109) <= b;
    layer2_outputs(1110) <= b;
    layer2_outputs(1111) <= not (a xor b);
    layer2_outputs(1112) <= not (a or b);
    layer2_outputs(1113) <= a xor b;
    layer2_outputs(1114) <= b and not a;
    layer2_outputs(1115) <= not (a and b);
    layer2_outputs(1116) <= a and b;
    layer2_outputs(1117) <= not b;
    layer2_outputs(1118) <= b;
    layer2_outputs(1119) <= not a;
    layer2_outputs(1120) <= b and not a;
    layer2_outputs(1121) <= '1';
    layer2_outputs(1122) <= b and not a;
    layer2_outputs(1123) <= not b;
    layer2_outputs(1124) <= not a;
    layer2_outputs(1125) <= a xor b;
    layer2_outputs(1126) <= '1';
    layer2_outputs(1127) <= b;
    layer2_outputs(1128) <= a and b;
    layer2_outputs(1129) <= not a;
    layer2_outputs(1130) <= not b;
    layer2_outputs(1131) <= a and b;
    layer2_outputs(1132) <= not b or a;
    layer2_outputs(1133) <= not (a or b);
    layer2_outputs(1134) <= not (a and b);
    layer2_outputs(1135) <= a;
    layer2_outputs(1136) <= a;
    layer2_outputs(1137) <= not (a or b);
    layer2_outputs(1138) <= not (a or b);
    layer2_outputs(1139) <= not (a or b);
    layer2_outputs(1140) <= not (a or b);
    layer2_outputs(1141) <= not a;
    layer2_outputs(1142) <= a and not b;
    layer2_outputs(1143) <= '1';
    layer2_outputs(1144) <= a and b;
    layer2_outputs(1145) <= not (a or b);
    layer2_outputs(1146) <= a;
    layer2_outputs(1147) <= not b or a;
    layer2_outputs(1148) <= a and b;
    layer2_outputs(1149) <= not (a and b);
    layer2_outputs(1150) <= '1';
    layer2_outputs(1151) <= not a;
    layer2_outputs(1152) <= a;
    layer2_outputs(1153) <= not a;
    layer2_outputs(1154) <= a or b;
    layer2_outputs(1155) <= a and b;
    layer2_outputs(1156) <= a or b;
    layer2_outputs(1157) <= not (a and b);
    layer2_outputs(1158) <= not (a or b);
    layer2_outputs(1159) <= a;
    layer2_outputs(1160) <= a and b;
    layer2_outputs(1161) <= not (a or b);
    layer2_outputs(1162) <= not b;
    layer2_outputs(1163) <= a or b;
    layer2_outputs(1164) <= not (a and b);
    layer2_outputs(1165) <= a and b;
    layer2_outputs(1166) <= a or b;
    layer2_outputs(1167) <= b;
    layer2_outputs(1168) <= a xor b;
    layer2_outputs(1169) <= a and b;
    layer2_outputs(1170) <= b;
    layer2_outputs(1171) <= a;
    layer2_outputs(1172) <= a;
    layer2_outputs(1173) <= a or b;
    layer2_outputs(1174) <= a;
    layer2_outputs(1175) <= '0';
    layer2_outputs(1176) <= b;
    layer2_outputs(1177) <= not (a and b);
    layer2_outputs(1178) <= a;
    layer2_outputs(1179) <= a or b;
    layer2_outputs(1180) <= not (a and b);
    layer2_outputs(1181) <= b;
    layer2_outputs(1182) <= not (a or b);
    layer2_outputs(1183) <= b;
    layer2_outputs(1184) <= b and not a;
    layer2_outputs(1185) <= not a;
    layer2_outputs(1186) <= a;
    layer2_outputs(1187) <= a and not b;
    layer2_outputs(1188) <= not b or a;
    layer2_outputs(1189) <= not (a xor b);
    layer2_outputs(1190) <= not a or b;
    layer2_outputs(1191) <= '0';
    layer2_outputs(1192) <= not (a or b);
    layer2_outputs(1193) <= '1';
    layer2_outputs(1194) <= b;
    layer2_outputs(1195) <= a or b;
    layer2_outputs(1196) <= '0';
    layer2_outputs(1197) <= not b or a;
    layer2_outputs(1198) <= b;
    layer2_outputs(1199) <= not (a and b);
    layer2_outputs(1200) <= a;
    layer2_outputs(1201) <= not a;
    layer2_outputs(1202) <= not (a or b);
    layer2_outputs(1203) <= not (a and b);
    layer2_outputs(1204) <= b;
    layer2_outputs(1205) <= a;
    layer2_outputs(1206) <= not b;
    layer2_outputs(1207) <= b;
    layer2_outputs(1208) <= not b;
    layer2_outputs(1209) <= not b;
    layer2_outputs(1210) <= not b;
    layer2_outputs(1211) <= '0';
    layer2_outputs(1212) <= a and not b;
    layer2_outputs(1213) <= not a or b;
    layer2_outputs(1214) <= not (a and b);
    layer2_outputs(1215) <= a;
    layer2_outputs(1216) <= not b;
    layer2_outputs(1217) <= a and not b;
    layer2_outputs(1218) <= a or b;
    layer2_outputs(1219) <= b;
    layer2_outputs(1220) <= a;
    layer2_outputs(1221) <= a;
    layer2_outputs(1222) <= a and b;
    layer2_outputs(1223) <= a or b;
    layer2_outputs(1224) <= not b or a;
    layer2_outputs(1225) <= not a;
    layer2_outputs(1226) <= not a or b;
    layer2_outputs(1227) <= not a;
    layer2_outputs(1228) <= b;
    layer2_outputs(1229) <= '0';
    layer2_outputs(1230) <= b and not a;
    layer2_outputs(1231) <= not (a or b);
    layer2_outputs(1232) <= b;
    layer2_outputs(1233) <= not a;
    layer2_outputs(1234) <= '0';
    layer2_outputs(1235) <= not (a or b);
    layer2_outputs(1236) <= not (a and b);
    layer2_outputs(1237) <= not (a or b);
    layer2_outputs(1238) <= a;
    layer2_outputs(1239) <= a;
    layer2_outputs(1240) <= '1';
    layer2_outputs(1241) <= not a;
    layer2_outputs(1242) <= not b;
    layer2_outputs(1243) <= '1';
    layer2_outputs(1244) <= a or b;
    layer2_outputs(1245) <= a and b;
    layer2_outputs(1246) <= not a;
    layer2_outputs(1247) <= a;
    layer2_outputs(1248) <= not (a and b);
    layer2_outputs(1249) <= '0';
    layer2_outputs(1250) <= a;
    layer2_outputs(1251) <= a xor b;
    layer2_outputs(1252) <= '1';
    layer2_outputs(1253) <= not (a and b);
    layer2_outputs(1254) <= a or b;
    layer2_outputs(1255) <= b and not a;
    layer2_outputs(1256) <= not (a and b);
    layer2_outputs(1257) <= b and not a;
    layer2_outputs(1258) <= not a;
    layer2_outputs(1259) <= b;
    layer2_outputs(1260) <= a and not b;
    layer2_outputs(1261) <= a and not b;
    layer2_outputs(1262) <= a;
    layer2_outputs(1263) <= '0';
    layer2_outputs(1264) <= b and not a;
    layer2_outputs(1265) <= a;
    layer2_outputs(1266) <= b;
    layer2_outputs(1267) <= a or b;
    layer2_outputs(1268) <= not (a or b);
    layer2_outputs(1269) <= not (a xor b);
    layer2_outputs(1270) <= a and not b;
    layer2_outputs(1271) <= '1';
    layer2_outputs(1272) <= not (a or b);
    layer2_outputs(1273) <= not b or a;
    layer2_outputs(1274) <= a or b;
    layer2_outputs(1275) <= not (a or b);
    layer2_outputs(1276) <= a or b;
    layer2_outputs(1277) <= a xor b;
    layer2_outputs(1278) <= '0';
    layer2_outputs(1279) <= not b;
    layer2_outputs(1280) <= not b;
    layer2_outputs(1281) <= a and not b;
    layer2_outputs(1282) <= not a;
    layer2_outputs(1283) <= a and b;
    layer2_outputs(1284) <= b;
    layer2_outputs(1285) <= b;
    layer2_outputs(1286) <= b;
    layer2_outputs(1287) <= a and b;
    layer2_outputs(1288) <= a and b;
    layer2_outputs(1289) <= a;
    layer2_outputs(1290) <= not a or b;
    layer2_outputs(1291) <= a and not b;
    layer2_outputs(1292) <= a xor b;
    layer2_outputs(1293) <= not a or b;
    layer2_outputs(1294) <= not (a xor b);
    layer2_outputs(1295) <= b;
    layer2_outputs(1296) <= b;
    layer2_outputs(1297) <= not a or b;
    layer2_outputs(1298) <= '1';
    layer2_outputs(1299) <= a xor b;
    layer2_outputs(1300) <= b;
    layer2_outputs(1301) <= '1';
    layer2_outputs(1302) <= not b;
    layer2_outputs(1303) <= not a or b;
    layer2_outputs(1304) <= not a or b;
    layer2_outputs(1305) <= not a;
    layer2_outputs(1306) <= not b;
    layer2_outputs(1307) <= not (a and b);
    layer2_outputs(1308) <= not b or a;
    layer2_outputs(1309) <= not b or a;
    layer2_outputs(1310) <= not b;
    layer2_outputs(1311) <= a;
    layer2_outputs(1312) <= a or b;
    layer2_outputs(1313) <= a or b;
    layer2_outputs(1314) <= a;
    layer2_outputs(1315) <= a and b;
    layer2_outputs(1316) <= a;
    layer2_outputs(1317) <= a xor b;
    layer2_outputs(1318) <= b and not a;
    layer2_outputs(1319) <= a;
    layer2_outputs(1320) <= b and not a;
    layer2_outputs(1321) <= a and b;
    layer2_outputs(1322) <= a;
    layer2_outputs(1323) <= not (a and b);
    layer2_outputs(1324) <= b;
    layer2_outputs(1325) <= a;
    layer2_outputs(1326) <= not (a and b);
    layer2_outputs(1327) <= not b;
    layer2_outputs(1328) <= not a or b;
    layer2_outputs(1329) <= '0';
    layer2_outputs(1330) <= b;
    layer2_outputs(1331) <= not (a xor b);
    layer2_outputs(1332) <= '1';
    layer2_outputs(1333) <= not a or b;
    layer2_outputs(1334) <= '0';
    layer2_outputs(1335) <= not b;
    layer2_outputs(1336) <= a and not b;
    layer2_outputs(1337) <= not a or b;
    layer2_outputs(1338) <= not b;
    layer2_outputs(1339) <= a;
    layer2_outputs(1340) <= not a;
    layer2_outputs(1341) <= not (a xor b);
    layer2_outputs(1342) <= b;
    layer2_outputs(1343) <= not a;
    layer2_outputs(1344) <= not (a or b);
    layer2_outputs(1345) <= a;
    layer2_outputs(1346) <= a and b;
    layer2_outputs(1347) <= a or b;
    layer2_outputs(1348) <= not (a or b);
    layer2_outputs(1349) <= '0';
    layer2_outputs(1350) <= b;
    layer2_outputs(1351) <= not b or a;
    layer2_outputs(1352) <= not (a or b);
    layer2_outputs(1353) <= not b;
    layer2_outputs(1354) <= not b;
    layer2_outputs(1355) <= '1';
    layer2_outputs(1356) <= a;
    layer2_outputs(1357) <= b;
    layer2_outputs(1358) <= not (a or b);
    layer2_outputs(1359) <= b;
    layer2_outputs(1360) <= a;
    layer2_outputs(1361) <= not (a xor b);
    layer2_outputs(1362) <= a and not b;
    layer2_outputs(1363) <= '0';
    layer2_outputs(1364) <= a or b;
    layer2_outputs(1365) <= not (a and b);
    layer2_outputs(1366) <= not (a or b);
    layer2_outputs(1367) <= a or b;
    layer2_outputs(1368) <= a and not b;
    layer2_outputs(1369) <= a xor b;
    layer2_outputs(1370) <= b and not a;
    layer2_outputs(1371) <= a and b;
    layer2_outputs(1372) <= a and not b;
    layer2_outputs(1373) <= not b or a;
    layer2_outputs(1374) <= a and b;
    layer2_outputs(1375) <= a;
    layer2_outputs(1376) <= not a;
    layer2_outputs(1377) <= not a or b;
    layer2_outputs(1378) <= not b or a;
    layer2_outputs(1379) <= a;
    layer2_outputs(1380) <= not (a or b);
    layer2_outputs(1381) <= not b;
    layer2_outputs(1382) <= a and b;
    layer2_outputs(1383) <= a or b;
    layer2_outputs(1384) <= '1';
    layer2_outputs(1385) <= not (a or b);
    layer2_outputs(1386) <= not b;
    layer2_outputs(1387) <= '1';
    layer2_outputs(1388) <= b and not a;
    layer2_outputs(1389) <= a and b;
    layer2_outputs(1390) <= '1';
    layer2_outputs(1391) <= not a or b;
    layer2_outputs(1392) <= not (a or b);
    layer2_outputs(1393) <= a and not b;
    layer2_outputs(1394) <= '1';
    layer2_outputs(1395) <= b and not a;
    layer2_outputs(1396) <= a xor b;
    layer2_outputs(1397) <= b;
    layer2_outputs(1398) <= b;
    layer2_outputs(1399) <= a or b;
    layer2_outputs(1400) <= a and not b;
    layer2_outputs(1401) <= '0';
    layer2_outputs(1402) <= a;
    layer2_outputs(1403) <= '0';
    layer2_outputs(1404) <= '1';
    layer2_outputs(1405) <= a xor b;
    layer2_outputs(1406) <= not a;
    layer2_outputs(1407) <= a;
    layer2_outputs(1408) <= not a;
    layer2_outputs(1409) <= not a or b;
    layer2_outputs(1410) <= b;
    layer2_outputs(1411) <= a;
    layer2_outputs(1412) <= not b or a;
    layer2_outputs(1413) <= a and b;
    layer2_outputs(1414) <= not (a or b);
    layer2_outputs(1415) <= b;
    layer2_outputs(1416) <= not b;
    layer2_outputs(1417) <= a or b;
    layer2_outputs(1418) <= not (a or b);
    layer2_outputs(1419) <= a or b;
    layer2_outputs(1420) <= a xor b;
    layer2_outputs(1421) <= not a;
    layer2_outputs(1422) <= a;
    layer2_outputs(1423) <= not a or b;
    layer2_outputs(1424) <= not a or b;
    layer2_outputs(1425) <= a and b;
    layer2_outputs(1426) <= not b;
    layer2_outputs(1427) <= not a;
    layer2_outputs(1428) <= a;
    layer2_outputs(1429) <= a;
    layer2_outputs(1430) <= a or b;
    layer2_outputs(1431) <= a or b;
    layer2_outputs(1432) <= a;
    layer2_outputs(1433) <= a or b;
    layer2_outputs(1434) <= b;
    layer2_outputs(1435) <= a and b;
    layer2_outputs(1436) <= not (a or b);
    layer2_outputs(1437) <= a or b;
    layer2_outputs(1438) <= not (a and b);
    layer2_outputs(1439) <= not a or b;
    layer2_outputs(1440) <= b and not a;
    layer2_outputs(1441) <= a xor b;
    layer2_outputs(1442) <= not (a and b);
    layer2_outputs(1443) <= a and b;
    layer2_outputs(1444) <= '0';
    layer2_outputs(1445) <= not a;
    layer2_outputs(1446) <= not b;
    layer2_outputs(1447) <= a xor b;
    layer2_outputs(1448) <= a and b;
    layer2_outputs(1449) <= not (a or b);
    layer2_outputs(1450) <= a xor b;
    layer2_outputs(1451) <= not (a and b);
    layer2_outputs(1452) <= not b;
    layer2_outputs(1453) <= not b or a;
    layer2_outputs(1454) <= a and b;
    layer2_outputs(1455) <= not (a and b);
    layer2_outputs(1456) <= a xor b;
    layer2_outputs(1457) <= not b;
    layer2_outputs(1458) <= b and not a;
    layer2_outputs(1459) <= '0';
    layer2_outputs(1460) <= a;
    layer2_outputs(1461) <= a and b;
    layer2_outputs(1462) <= b;
    layer2_outputs(1463) <= '1';
    layer2_outputs(1464) <= a;
    layer2_outputs(1465) <= not b;
    layer2_outputs(1466) <= '1';
    layer2_outputs(1467) <= a or b;
    layer2_outputs(1468) <= a and not b;
    layer2_outputs(1469) <= not (a or b);
    layer2_outputs(1470) <= a;
    layer2_outputs(1471) <= not (a and b);
    layer2_outputs(1472) <= not a or b;
    layer2_outputs(1473) <= not (a or b);
    layer2_outputs(1474) <= a and not b;
    layer2_outputs(1475) <= a and b;
    layer2_outputs(1476) <= b;
    layer2_outputs(1477) <= a xor b;
    layer2_outputs(1478) <= '1';
    layer2_outputs(1479) <= not b or a;
    layer2_outputs(1480) <= a;
    layer2_outputs(1481) <= a and b;
    layer2_outputs(1482) <= b;
    layer2_outputs(1483) <= not a;
    layer2_outputs(1484) <= a and not b;
    layer2_outputs(1485) <= b;
    layer2_outputs(1486) <= not b;
    layer2_outputs(1487) <= b and not a;
    layer2_outputs(1488) <= b;
    layer2_outputs(1489) <= b and not a;
    layer2_outputs(1490) <= a and not b;
    layer2_outputs(1491) <= '1';
    layer2_outputs(1492) <= not a or b;
    layer2_outputs(1493) <= a;
    layer2_outputs(1494) <= a or b;
    layer2_outputs(1495) <= b and not a;
    layer2_outputs(1496) <= not b;
    layer2_outputs(1497) <= not a or b;
    layer2_outputs(1498) <= a xor b;
    layer2_outputs(1499) <= not a or b;
    layer2_outputs(1500) <= not b or a;
    layer2_outputs(1501) <= not b or a;
    layer2_outputs(1502) <= '1';
    layer2_outputs(1503) <= a;
    layer2_outputs(1504) <= not a or b;
    layer2_outputs(1505) <= b and not a;
    layer2_outputs(1506) <= not a or b;
    layer2_outputs(1507) <= '0';
    layer2_outputs(1508) <= a;
    layer2_outputs(1509) <= '1';
    layer2_outputs(1510) <= not b or a;
    layer2_outputs(1511) <= a xor b;
    layer2_outputs(1512) <= b;
    layer2_outputs(1513) <= a or b;
    layer2_outputs(1514) <= not b or a;
    layer2_outputs(1515) <= '1';
    layer2_outputs(1516) <= '1';
    layer2_outputs(1517) <= not b;
    layer2_outputs(1518) <= b and not a;
    layer2_outputs(1519) <= not b;
    layer2_outputs(1520) <= not a or b;
    layer2_outputs(1521) <= a or b;
    layer2_outputs(1522) <= '0';
    layer2_outputs(1523) <= a or b;
    layer2_outputs(1524) <= a;
    layer2_outputs(1525) <= not (a and b);
    layer2_outputs(1526) <= a xor b;
    layer2_outputs(1527) <= not b or a;
    layer2_outputs(1528) <= a and b;
    layer2_outputs(1529) <= a and b;
    layer2_outputs(1530) <= not (a and b);
    layer2_outputs(1531) <= '0';
    layer2_outputs(1532) <= a and not b;
    layer2_outputs(1533) <= b;
    layer2_outputs(1534) <= a xor b;
    layer2_outputs(1535) <= not a;
    layer2_outputs(1536) <= a and not b;
    layer2_outputs(1537) <= a;
    layer2_outputs(1538) <= b and not a;
    layer2_outputs(1539) <= a and b;
    layer2_outputs(1540) <= not b;
    layer2_outputs(1541) <= not b or a;
    layer2_outputs(1542) <= a or b;
    layer2_outputs(1543) <= not (a and b);
    layer2_outputs(1544) <= not b;
    layer2_outputs(1545) <= not (a and b);
    layer2_outputs(1546) <= a;
    layer2_outputs(1547) <= a or b;
    layer2_outputs(1548) <= '1';
    layer2_outputs(1549) <= a and not b;
    layer2_outputs(1550) <= '0';
    layer2_outputs(1551) <= a and not b;
    layer2_outputs(1552) <= a;
    layer2_outputs(1553) <= a and not b;
    layer2_outputs(1554) <= a and b;
    layer2_outputs(1555) <= not a;
    layer2_outputs(1556) <= a and b;
    layer2_outputs(1557) <= '0';
    layer2_outputs(1558) <= b;
    layer2_outputs(1559) <= not (a or b);
    layer2_outputs(1560) <= not b;
    layer2_outputs(1561) <= not b;
    layer2_outputs(1562) <= not b or a;
    layer2_outputs(1563) <= a;
    layer2_outputs(1564) <= not (a xor b);
    layer2_outputs(1565) <= not a;
    layer2_outputs(1566) <= not a;
    layer2_outputs(1567) <= a and not b;
    layer2_outputs(1568) <= b and not a;
    layer2_outputs(1569) <= b and not a;
    layer2_outputs(1570) <= a;
    layer2_outputs(1571) <= not a;
    layer2_outputs(1572) <= not (a and b);
    layer2_outputs(1573) <= not a;
    layer2_outputs(1574) <= not b or a;
    layer2_outputs(1575) <= not a;
    layer2_outputs(1576) <= b;
    layer2_outputs(1577) <= not b;
    layer2_outputs(1578) <= not b or a;
    layer2_outputs(1579) <= '1';
    layer2_outputs(1580) <= not a or b;
    layer2_outputs(1581) <= '1';
    layer2_outputs(1582) <= not a or b;
    layer2_outputs(1583) <= not b or a;
    layer2_outputs(1584) <= a;
    layer2_outputs(1585) <= a and not b;
    layer2_outputs(1586) <= b and not a;
    layer2_outputs(1587) <= '0';
    layer2_outputs(1588) <= not a or b;
    layer2_outputs(1589) <= a or b;
    layer2_outputs(1590) <= a;
    layer2_outputs(1591) <= not a or b;
    layer2_outputs(1592) <= a and not b;
    layer2_outputs(1593) <= b;
    layer2_outputs(1594) <= '1';
    layer2_outputs(1595) <= b and not a;
    layer2_outputs(1596) <= b;
    layer2_outputs(1597) <= not (a xor b);
    layer2_outputs(1598) <= not (a xor b);
    layer2_outputs(1599) <= not b or a;
    layer2_outputs(1600) <= not a;
    layer2_outputs(1601) <= b;
    layer2_outputs(1602) <= a and not b;
    layer2_outputs(1603) <= a and not b;
    layer2_outputs(1604) <= b and not a;
    layer2_outputs(1605) <= not a or b;
    layer2_outputs(1606) <= not (a and b);
    layer2_outputs(1607) <= not b or a;
    layer2_outputs(1608) <= a or b;
    layer2_outputs(1609) <= b;
    layer2_outputs(1610) <= not b;
    layer2_outputs(1611) <= not a;
    layer2_outputs(1612) <= a and not b;
    layer2_outputs(1613) <= b and not a;
    layer2_outputs(1614) <= not a or b;
    layer2_outputs(1615) <= a and b;
    layer2_outputs(1616) <= a xor b;
    layer2_outputs(1617) <= not (a or b);
    layer2_outputs(1618) <= not a;
    layer2_outputs(1619) <= not a;
    layer2_outputs(1620) <= not a or b;
    layer2_outputs(1621) <= b and not a;
    layer2_outputs(1622) <= a xor b;
    layer2_outputs(1623) <= b and not a;
    layer2_outputs(1624) <= a;
    layer2_outputs(1625) <= not b;
    layer2_outputs(1626) <= not (a or b);
    layer2_outputs(1627) <= a;
    layer2_outputs(1628) <= a or b;
    layer2_outputs(1629) <= not b;
    layer2_outputs(1630) <= not b;
    layer2_outputs(1631) <= '0';
    layer2_outputs(1632) <= a or b;
    layer2_outputs(1633) <= not a;
    layer2_outputs(1634) <= not a;
    layer2_outputs(1635) <= not a;
    layer2_outputs(1636) <= '1';
    layer2_outputs(1637) <= not (a or b);
    layer2_outputs(1638) <= a and not b;
    layer2_outputs(1639) <= not a or b;
    layer2_outputs(1640) <= b;
    layer2_outputs(1641) <= not (a and b);
    layer2_outputs(1642) <= not (a or b);
    layer2_outputs(1643) <= not a;
    layer2_outputs(1644) <= not (a or b);
    layer2_outputs(1645) <= a or b;
    layer2_outputs(1646) <= not (a or b);
    layer2_outputs(1647) <= not (a and b);
    layer2_outputs(1648) <= a or b;
    layer2_outputs(1649) <= a and not b;
    layer2_outputs(1650) <= not a;
    layer2_outputs(1651) <= not a or b;
    layer2_outputs(1652) <= not (a and b);
    layer2_outputs(1653) <= '1';
    layer2_outputs(1654) <= '1';
    layer2_outputs(1655) <= not (a xor b);
    layer2_outputs(1656) <= b;
    layer2_outputs(1657) <= a and not b;
    layer2_outputs(1658) <= not b;
    layer2_outputs(1659) <= b;
    layer2_outputs(1660) <= a and not b;
    layer2_outputs(1661) <= a or b;
    layer2_outputs(1662) <= '0';
    layer2_outputs(1663) <= b;
    layer2_outputs(1664) <= not (a and b);
    layer2_outputs(1665) <= a;
    layer2_outputs(1666) <= '0';
    layer2_outputs(1667) <= not b or a;
    layer2_outputs(1668) <= not b;
    layer2_outputs(1669) <= a xor b;
    layer2_outputs(1670) <= not a or b;
    layer2_outputs(1671) <= not a or b;
    layer2_outputs(1672) <= not (a and b);
    layer2_outputs(1673) <= '0';
    layer2_outputs(1674) <= b and not a;
    layer2_outputs(1675) <= not a or b;
    layer2_outputs(1676) <= a;
    layer2_outputs(1677) <= not b;
    layer2_outputs(1678) <= not (a or b);
    layer2_outputs(1679) <= not (a or b);
    layer2_outputs(1680) <= not a or b;
    layer2_outputs(1681) <= not (a and b);
    layer2_outputs(1682) <= '1';
    layer2_outputs(1683) <= not b or a;
    layer2_outputs(1684) <= not a;
    layer2_outputs(1685) <= not a;
    layer2_outputs(1686) <= a;
    layer2_outputs(1687) <= b;
    layer2_outputs(1688) <= not b or a;
    layer2_outputs(1689) <= not b;
    layer2_outputs(1690) <= '1';
    layer2_outputs(1691) <= not (a and b);
    layer2_outputs(1692) <= a and not b;
    layer2_outputs(1693) <= a;
    layer2_outputs(1694) <= not b;
    layer2_outputs(1695) <= not (a and b);
    layer2_outputs(1696) <= not (a and b);
    layer2_outputs(1697) <= '0';
    layer2_outputs(1698) <= '1';
    layer2_outputs(1699) <= a xor b;
    layer2_outputs(1700) <= not b;
    layer2_outputs(1701) <= not b;
    layer2_outputs(1702) <= not a;
    layer2_outputs(1703) <= not (a or b);
    layer2_outputs(1704) <= a and b;
    layer2_outputs(1705) <= not a;
    layer2_outputs(1706) <= not (a xor b);
    layer2_outputs(1707) <= b;
    layer2_outputs(1708) <= b and not a;
    layer2_outputs(1709) <= a and not b;
    layer2_outputs(1710) <= not (a and b);
    layer2_outputs(1711) <= '1';
    layer2_outputs(1712) <= '0';
    layer2_outputs(1713) <= b and not a;
    layer2_outputs(1714) <= not a or b;
    layer2_outputs(1715) <= not b;
    layer2_outputs(1716) <= not a or b;
    layer2_outputs(1717) <= not b;
    layer2_outputs(1718) <= a or b;
    layer2_outputs(1719) <= not a;
    layer2_outputs(1720) <= a and not b;
    layer2_outputs(1721) <= b and not a;
    layer2_outputs(1722) <= not a;
    layer2_outputs(1723) <= not (a or b);
    layer2_outputs(1724) <= a and b;
    layer2_outputs(1725) <= not b or a;
    layer2_outputs(1726) <= '1';
    layer2_outputs(1727) <= not b;
    layer2_outputs(1728) <= b and not a;
    layer2_outputs(1729) <= not a or b;
    layer2_outputs(1730) <= not a;
    layer2_outputs(1731) <= not a or b;
    layer2_outputs(1732) <= a and not b;
    layer2_outputs(1733) <= not a;
    layer2_outputs(1734) <= a;
    layer2_outputs(1735) <= a;
    layer2_outputs(1736) <= not (a xor b);
    layer2_outputs(1737) <= not a;
    layer2_outputs(1738) <= a;
    layer2_outputs(1739) <= b;
    layer2_outputs(1740) <= '0';
    layer2_outputs(1741) <= a and b;
    layer2_outputs(1742) <= a or b;
    layer2_outputs(1743) <= a and not b;
    layer2_outputs(1744) <= not (a or b);
    layer2_outputs(1745) <= a or b;
    layer2_outputs(1746) <= b;
    layer2_outputs(1747) <= not (a or b);
    layer2_outputs(1748) <= not b;
    layer2_outputs(1749) <= not (a or b);
    layer2_outputs(1750) <= a;
    layer2_outputs(1751) <= '1';
    layer2_outputs(1752) <= not (a and b);
    layer2_outputs(1753) <= a and not b;
    layer2_outputs(1754) <= a and b;
    layer2_outputs(1755) <= a and not b;
    layer2_outputs(1756) <= not b;
    layer2_outputs(1757) <= a or b;
    layer2_outputs(1758) <= a;
    layer2_outputs(1759) <= '1';
    layer2_outputs(1760) <= not a or b;
    layer2_outputs(1761) <= a or b;
    layer2_outputs(1762) <= a;
    layer2_outputs(1763) <= '1';
    layer2_outputs(1764) <= a xor b;
    layer2_outputs(1765) <= not a or b;
    layer2_outputs(1766) <= '0';
    layer2_outputs(1767) <= not (a or b);
    layer2_outputs(1768) <= b and not a;
    layer2_outputs(1769) <= not (a and b);
    layer2_outputs(1770) <= not (a and b);
    layer2_outputs(1771) <= not a;
    layer2_outputs(1772) <= '1';
    layer2_outputs(1773) <= a xor b;
    layer2_outputs(1774) <= a;
    layer2_outputs(1775) <= not (a and b);
    layer2_outputs(1776) <= not (a and b);
    layer2_outputs(1777) <= a;
    layer2_outputs(1778) <= not a or b;
    layer2_outputs(1779) <= b and not a;
    layer2_outputs(1780) <= not a or b;
    layer2_outputs(1781) <= a and not b;
    layer2_outputs(1782) <= a xor b;
    layer2_outputs(1783) <= '0';
    layer2_outputs(1784) <= b and not a;
    layer2_outputs(1785) <= a and b;
    layer2_outputs(1786) <= a and not b;
    layer2_outputs(1787) <= not (a xor b);
    layer2_outputs(1788) <= not a;
    layer2_outputs(1789) <= b and not a;
    layer2_outputs(1790) <= not a or b;
    layer2_outputs(1791) <= '1';
    layer2_outputs(1792) <= not a or b;
    layer2_outputs(1793) <= '0';
    layer2_outputs(1794) <= not b or a;
    layer2_outputs(1795) <= not b or a;
    layer2_outputs(1796) <= not (a or b);
    layer2_outputs(1797) <= not a or b;
    layer2_outputs(1798) <= not a;
    layer2_outputs(1799) <= not (a and b);
    layer2_outputs(1800) <= not b or a;
    layer2_outputs(1801) <= b;
    layer2_outputs(1802) <= a or b;
    layer2_outputs(1803) <= not b or a;
    layer2_outputs(1804) <= '0';
    layer2_outputs(1805) <= a or b;
    layer2_outputs(1806) <= a and b;
    layer2_outputs(1807) <= not a;
    layer2_outputs(1808) <= a;
    layer2_outputs(1809) <= not (a and b);
    layer2_outputs(1810) <= not b;
    layer2_outputs(1811) <= a or b;
    layer2_outputs(1812) <= not b or a;
    layer2_outputs(1813) <= not (a xor b);
    layer2_outputs(1814) <= a or b;
    layer2_outputs(1815) <= a or b;
    layer2_outputs(1816) <= not (a and b);
    layer2_outputs(1817) <= '1';
    layer2_outputs(1818) <= b;
    layer2_outputs(1819) <= not b or a;
    layer2_outputs(1820) <= not a or b;
    layer2_outputs(1821) <= a and not b;
    layer2_outputs(1822) <= a;
    layer2_outputs(1823) <= a or b;
    layer2_outputs(1824) <= b and not a;
    layer2_outputs(1825) <= b;
    layer2_outputs(1826) <= not a;
    layer2_outputs(1827) <= '0';
    layer2_outputs(1828) <= not a or b;
    layer2_outputs(1829) <= a xor b;
    layer2_outputs(1830) <= a xor b;
    layer2_outputs(1831) <= not (a or b);
    layer2_outputs(1832) <= a and not b;
    layer2_outputs(1833) <= a xor b;
    layer2_outputs(1834) <= b;
    layer2_outputs(1835) <= a or b;
    layer2_outputs(1836) <= not a;
    layer2_outputs(1837) <= not a or b;
    layer2_outputs(1838) <= '1';
    layer2_outputs(1839) <= not (a or b);
    layer2_outputs(1840) <= not a;
    layer2_outputs(1841) <= '0';
    layer2_outputs(1842) <= a;
    layer2_outputs(1843) <= '0';
    layer2_outputs(1844) <= not b;
    layer2_outputs(1845) <= b and not a;
    layer2_outputs(1846) <= b;
    layer2_outputs(1847) <= not b or a;
    layer2_outputs(1848) <= a and b;
    layer2_outputs(1849) <= a;
    layer2_outputs(1850) <= a and not b;
    layer2_outputs(1851) <= a xor b;
    layer2_outputs(1852) <= not (a and b);
    layer2_outputs(1853) <= not (a and b);
    layer2_outputs(1854) <= b;
    layer2_outputs(1855) <= a;
    layer2_outputs(1856) <= a;
    layer2_outputs(1857) <= a xor b;
    layer2_outputs(1858) <= a and b;
    layer2_outputs(1859) <= not b or a;
    layer2_outputs(1860) <= not (a and b);
    layer2_outputs(1861) <= b and not a;
    layer2_outputs(1862) <= a and b;
    layer2_outputs(1863) <= a and not b;
    layer2_outputs(1864) <= '1';
    layer2_outputs(1865) <= b and not a;
    layer2_outputs(1866) <= a;
    layer2_outputs(1867) <= b;
    layer2_outputs(1868) <= a xor b;
    layer2_outputs(1869) <= a xor b;
    layer2_outputs(1870) <= not (a or b);
    layer2_outputs(1871) <= b and not a;
    layer2_outputs(1872) <= not b;
    layer2_outputs(1873) <= a and not b;
    layer2_outputs(1874) <= '0';
    layer2_outputs(1875) <= a and not b;
    layer2_outputs(1876) <= '0';
    layer2_outputs(1877) <= b and not a;
    layer2_outputs(1878) <= not (a and b);
    layer2_outputs(1879) <= not (a and b);
    layer2_outputs(1880) <= a;
    layer2_outputs(1881) <= not b or a;
    layer2_outputs(1882) <= not a;
    layer2_outputs(1883) <= not (a or b);
    layer2_outputs(1884) <= '1';
    layer2_outputs(1885) <= a and not b;
    layer2_outputs(1886) <= b;
    layer2_outputs(1887) <= a xor b;
    layer2_outputs(1888) <= not a;
    layer2_outputs(1889) <= not a;
    layer2_outputs(1890) <= '0';
    layer2_outputs(1891) <= a;
    layer2_outputs(1892) <= a and b;
    layer2_outputs(1893) <= a and b;
    layer2_outputs(1894) <= not b or a;
    layer2_outputs(1895) <= a;
    layer2_outputs(1896) <= not (a and b);
    layer2_outputs(1897) <= not a;
    layer2_outputs(1898) <= b and not a;
    layer2_outputs(1899) <= not a or b;
    layer2_outputs(1900) <= not b or a;
    layer2_outputs(1901) <= not (a or b);
    layer2_outputs(1902) <= not a;
    layer2_outputs(1903) <= not a;
    layer2_outputs(1904) <= not (a or b);
    layer2_outputs(1905) <= not a;
    layer2_outputs(1906) <= b;
    layer2_outputs(1907) <= b;
    layer2_outputs(1908) <= '1';
    layer2_outputs(1909) <= not a or b;
    layer2_outputs(1910) <= not a;
    layer2_outputs(1911) <= not (a or b);
    layer2_outputs(1912) <= a or b;
    layer2_outputs(1913) <= not (a or b);
    layer2_outputs(1914) <= not a or b;
    layer2_outputs(1915) <= not b;
    layer2_outputs(1916) <= '1';
    layer2_outputs(1917) <= b;
    layer2_outputs(1918) <= a and b;
    layer2_outputs(1919) <= a or b;
    layer2_outputs(1920) <= b;
    layer2_outputs(1921) <= a and not b;
    layer2_outputs(1922) <= b and not a;
    layer2_outputs(1923) <= not (a xor b);
    layer2_outputs(1924) <= a;
    layer2_outputs(1925) <= b;
    layer2_outputs(1926) <= a and not b;
    layer2_outputs(1927) <= not a;
    layer2_outputs(1928) <= b and not a;
    layer2_outputs(1929) <= a or b;
    layer2_outputs(1930) <= not b;
    layer2_outputs(1931) <= not b;
    layer2_outputs(1932) <= a or b;
    layer2_outputs(1933) <= a;
    layer2_outputs(1934) <= not (a or b);
    layer2_outputs(1935) <= a and b;
    layer2_outputs(1936) <= not b or a;
    layer2_outputs(1937) <= b and not a;
    layer2_outputs(1938) <= a and b;
    layer2_outputs(1939) <= a and not b;
    layer2_outputs(1940) <= a and b;
    layer2_outputs(1941) <= a or b;
    layer2_outputs(1942) <= b and not a;
    layer2_outputs(1943) <= not b or a;
    layer2_outputs(1944) <= a and b;
    layer2_outputs(1945) <= b;
    layer2_outputs(1946) <= b;
    layer2_outputs(1947) <= a;
    layer2_outputs(1948) <= a;
    layer2_outputs(1949) <= '0';
    layer2_outputs(1950) <= a and b;
    layer2_outputs(1951) <= a and b;
    layer2_outputs(1952) <= not a;
    layer2_outputs(1953) <= not (a or b);
    layer2_outputs(1954) <= a xor b;
    layer2_outputs(1955) <= not a or b;
    layer2_outputs(1956) <= not a;
    layer2_outputs(1957) <= b;
    layer2_outputs(1958) <= b;
    layer2_outputs(1959) <= not (a or b);
    layer2_outputs(1960) <= not (a or b);
    layer2_outputs(1961) <= a and b;
    layer2_outputs(1962) <= '0';
    layer2_outputs(1963) <= not (a or b);
    layer2_outputs(1964) <= not (a xor b);
    layer2_outputs(1965) <= '0';
    layer2_outputs(1966) <= not (a or b);
    layer2_outputs(1967) <= b;
    layer2_outputs(1968) <= b;
    layer2_outputs(1969) <= not b or a;
    layer2_outputs(1970) <= not b or a;
    layer2_outputs(1971) <= a xor b;
    layer2_outputs(1972) <= a;
    layer2_outputs(1973) <= not (a xor b);
    layer2_outputs(1974) <= not b;
    layer2_outputs(1975) <= a or b;
    layer2_outputs(1976) <= a;
    layer2_outputs(1977) <= a and b;
    layer2_outputs(1978) <= b;
    layer2_outputs(1979) <= not b or a;
    layer2_outputs(1980) <= not a;
    layer2_outputs(1981) <= not b;
    layer2_outputs(1982) <= a;
    layer2_outputs(1983) <= not a;
    layer2_outputs(1984) <= a and b;
    layer2_outputs(1985) <= not a;
    layer2_outputs(1986) <= not b;
    layer2_outputs(1987) <= a and not b;
    layer2_outputs(1988) <= not a or b;
    layer2_outputs(1989) <= not b;
    layer2_outputs(1990) <= b and not a;
    layer2_outputs(1991) <= not a or b;
    layer2_outputs(1992) <= a xor b;
    layer2_outputs(1993) <= not (a and b);
    layer2_outputs(1994) <= not (a and b);
    layer2_outputs(1995) <= '1';
    layer2_outputs(1996) <= not b;
    layer2_outputs(1997) <= a and not b;
    layer2_outputs(1998) <= not (a or b);
    layer2_outputs(1999) <= a;
    layer2_outputs(2000) <= a and not b;
    layer2_outputs(2001) <= a and b;
    layer2_outputs(2002) <= not a;
    layer2_outputs(2003) <= not b;
    layer2_outputs(2004) <= '1';
    layer2_outputs(2005) <= '0';
    layer2_outputs(2006) <= a and not b;
    layer2_outputs(2007) <= not (a and b);
    layer2_outputs(2008) <= '0';
    layer2_outputs(2009) <= not a;
    layer2_outputs(2010) <= a and b;
    layer2_outputs(2011) <= not (a and b);
    layer2_outputs(2012) <= not a;
    layer2_outputs(2013) <= not (a and b);
    layer2_outputs(2014) <= not a or b;
    layer2_outputs(2015) <= a;
    layer2_outputs(2016) <= not a;
    layer2_outputs(2017) <= not (a and b);
    layer2_outputs(2018) <= '0';
    layer2_outputs(2019) <= not (a or b);
    layer2_outputs(2020) <= not (a xor b);
    layer2_outputs(2021) <= a and not b;
    layer2_outputs(2022) <= '0';
    layer2_outputs(2023) <= not b;
    layer2_outputs(2024) <= not a;
    layer2_outputs(2025) <= '0';
    layer2_outputs(2026) <= not (a or b);
    layer2_outputs(2027) <= a and b;
    layer2_outputs(2028) <= b;
    layer2_outputs(2029) <= a and not b;
    layer2_outputs(2030) <= not (a and b);
    layer2_outputs(2031) <= not b;
    layer2_outputs(2032) <= b and not a;
    layer2_outputs(2033) <= a and b;
    layer2_outputs(2034) <= not b;
    layer2_outputs(2035) <= '0';
    layer2_outputs(2036) <= a or b;
    layer2_outputs(2037) <= not b or a;
    layer2_outputs(2038) <= not a or b;
    layer2_outputs(2039) <= not a or b;
    layer2_outputs(2040) <= not (a and b);
    layer2_outputs(2041) <= not a;
    layer2_outputs(2042) <= a;
    layer2_outputs(2043) <= not (a xor b);
    layer2_outputs(2044) <= not (a or b);
    layer2_outputs(2045) <= a;
    layer2_outputs(2046) <= not (a or b);
    layer2_outputs(2047) <= '0';
    layer2_outputs(2048) <= a and b;
    layer2_outputs(2049) <= a and not b;
    layer2_outputs(2050) <= b;
    layer2_outputs(2051) <= '0';
    layer2_outputs(2052) <= not b or a;
    layer2_outputs(2053) <= not (a xor b);
    layer2_outputs(2054) <= not b or a;
    layer2_outputs(2055) <= '0';
    layer2_outputs(2056) <= a and not b;
    layer2_outputs(2057) <= a or b;
    layer2_outputs(2058) <= not b or a;
    layer2_outputs(2059) <= b and not a;
    layer2_outputs(2060) <= '1';
    layer2_outputs(2061) <= not (a xor b);
    layer2_outputs(2062) <= a or b;
    layer2_outputs(2063) <= a or b;
    layer2_outputs(2064) <= a or b;
    layer2_outputs(2065) <= not a or b;
    layer2_outputs(2066) <= b;
    layer2_outputs(2067) <= not (a or b);
    layer2_outputs(2068) <= a;
    layer2_outputs(2069) <= a and b;
    layer2_outputs(2070) <= not (a or b);
    layer2_outputs(2071) <= a and not b;
    layer2_outputs(2072) <= a and not b;
    layer2_outputs(2073) <= a;
    layer2_outputs(2074) <= '1';
    layer2_outputs(2075) <= b;
    layer2_outputs(2076) <= b and not a;
    layer2_outputs(2077) <= a;
    layer2_outputs(2078) <= not a;
    layer2_outputs(2079) <= '0';
    layer2_outputs(2080) <= b and not a;
    layer2_outputs(2081) <= not (a or b);
    layer2_outputs(2082) <= not (a and b);
    layer2_outputs(2083) <= not b or a;
    layer2_outputs(2084) <= a and b;
    layer2_outputs(2085) <= not b;
    layer2_outputs(2086) <= b;
    layer2_outputs(2087) <= a;
    layer2_outputs(2088) <= a and not b;
    layer2_outputs(2089) <= b;
    layer2_outputs(2090) <= a xor b;
    layer2_outputs(2091) <= not (a or b);
    layer2_outputs(2092) <= '0';
    layer2_outputs(2093) <= '0';
    layer2_outputs(2094) <= not (a or b);
    layer2_outputs(2095) <= not a or b;
    layer2_outputs(2096) <= a xor b;
    layer2_outputs(2097) <= b and not a;
    layer2_outputs(2098) <= not a;
    layer2_outputs(2099) <= not a or b;
    layer2_outputs(2100) <= not b or a;
    layer2_outputs(2101) <= b;
    layer2_outputs(2102) <= '0';
    layer2_outputs(2103) <= not b or a;
    layer2_outputs(2104) <= a and b;
    layer2_outputs(2105) <= not a or b;
    layer2_outputs(2106) <= not b;
    layer2_outputs(2107) <= a and b;
    layer2_outputs(2108) <= not (a or b);
    layer2_outputs(2109) <= not (a or b);
    layer2_outputs(2110) <= not b;
    layer2_outputs(2111) <= b and not a;
    layer2_outputs(2112) <= not (a xor b);
    layer2_outputs(2113) <= a;
    layer2_outputs(2114) <= a or b;
    layer2_outputs(2115) <= not (a or b);
    layer2_outputs(2116) <= a or b;
    layer2_outputs(2117) <= a;
    layer2_outputs(2118) <= not a or b;
    layer2_outputs(2119) <= a and b;
    layer2_outputs(2120) <= a and b;
    layer2_outputs(2121) <= b;
    layer2_outputs(2122) <= a or b;
    layer2_outputs(2123) <= not (a xor b);
    layer2_outputs(2124) <= not a or b;
    layer2_outputs(2125) <= not b;
    layer2_outputs(2126) <= not (a and b);
    layer2_outputs(2127) <= b;
    layer2_outputs(2128) <= not (a and b);
    layer2_outputs(2129) <= not b or a;
    layer2_outputs(2130) <= '0';
    layer2_outputs(2131) <= a and not b;
    layer2_outputs(2132) <= a and b;
    layer2_outputs(2133) <= a;
    layer2_outputs(2134) <= not b;
    layer2_outputs(2135) <= not b or a;
    layer2_outputs(2136) <= not b;
    layer2_outputs(2137) <= not b;
    layer2_outputs(2138) <= not b;
    layer2_outputs(2139) <= not b;
    layer2_outputs(2140) <= not a;
    layer2_outputs(2141) <= a or b;
    layer2_outputs(2142) <= '0';
    layer2_outputs(2143) <= not a or b;
    layer2_outputs(2144) <= not a or b;
    layer2_outputs(2145) <= '0';
    layer2_outputs(2146) <= not a or b;
    layer2_outputs(2147) <= '0';
    layer2_outputs(2148) <= a;
    layer2_outputs(2149) <= not (a and b);
    layer2_outputs(2150) <= a xor b;
    layer2_outputs(2151) <= not (a or b);
    layer2_outputs(2152) <= not b or a;
    layer2_outputs(2153) <= a and not b;
    layer2_outputs(2154) <= a or b;
    layer2_outputs(2155) <= not a or b;
    layer2_outputs(2156) <= not a or b;
    layer2_outputs(2157) <= a;
    layer2_outputs(2158) <= a and b;
    layer2_outputs(2159) <= b;
    layer2_outputs(2160) <= '1';
    layer2_outputs(2161) <= not a;
    layer2_outputs(2162) <= not (a and b);
    layer2_outputs(2163) <= a and b;
    layer2_outputs(2164) <= '1';
    layer2_outputs(2165) <= b and not a;
    layer2_outputs(2166) <= not a;
    layer2_outputs(2167) <= a;
    layer2_outputs(2168) <= a and b;
    layer2_outputs(2169) <= b;
    layer2_outputs(2170) <= a xor b;
    layer2_outputs(2171) <= not b or a;
    layer2_outputs(2172) <= not (a xor b);
    layer2_outputs(2173) <= a xor b;
    layer2_outputs(2174) <= a;
    layer2_outputs(2175) <= '1';
    layer2_outputs(2176) <= a or b;
    layer2_outputs(2177) <= a or b;
    layer2_outputs(2178) <= a and not b;
    layer2_outputs(2179) <= a or b;
    layer2_outputs(2180) <= a and b;
    layer2_outputs(2181) <= b;
    layer2_outputs(2182) <= not (a and b);
    layer2_outputs(2183) <= not b or a;
    layer2_outputs(2184) <= a and not b;
    layer2_outputs(2185) <= b and not a;
    layer2_outputs(2186) <= not b or a;
    layer2_outputs(2187) <= a and not b;
    layer2_outputs(2188) <= not a;
    layer2_outputs(2189) <= a xor b;
    layer2_outputs(2190) <= a and not b;
    layer2_outputs(2191) <= not (a or b);
    layer2_outputs(2192) <= not a;
    layer2_outputs(2193) <= not a;
    layer2_outputs(2194) <= '0';
    layer2_outputs(2195) <= not a;
    layer2_outputs(2196) <= a;
    layer2_outputs(2197) <= b;
    layer2_outputs(2198) <= b and not a;
    layer2_outputs(2199) <= a or b;
    layer2_outputs(2200) <= '0';
    layer2_outputs(2201) <= not a or b;
    layer2_outputs(2202) <= not (a and b);
    layer2_outputs(2203) <= a;
    layer2_outputs(2204) <= a and not b;
    layer2_outputs(2205) <= a xor b;
    layer2_outputs(2206) <= not a or b;
    layer2_outputs(2207) <= '1';
    layer2_outputs(2208) <= not b or a;
    layer2_outputs(2209) <= not (a or b);
    layer2_outputs(2210) <= not (a xor b);
    layer2_outputs(2211) <= not (a or b);
    layer2_outputs(2212) <= '1';
    layer2_outputs(2213) <= not (a and b);
    layer2_outputs(2214) <= not b or a;
    layer2_outputs(2215) <= a xor b;
    layer2_outputs(2216) <= not (a and b);
    layer2_outputs(2217) <= '1';
    layer2_outputs(2218) <= b;
    layer2_outputs(2219) <= not b;
    layer2_outputs(2220) <= a;
    layer2_outputs(2221) <= not (a and b);
    layer2_outputs(2222) <= '0';
    layer2_outputs(2223) <= b and not a;
    layer2_outputs(2224) <= a or b;
    layer2_outputs(2225) <= '1';
    layer2_outputs(2226) <= a or b;
    layer2_outputs(2227) <= not (a xor b);
    layer2_outputs(2228) <= '0';
    layer2_outputs(2229) <= a;
    layer2_outputs(2230) <= not b or a;
    layer2_outputs(2231) <= a;
    layer2_outputs(2232) <= not a;
    layer2_outputs(2233) <= b and not a;
    layer2_outputs(2234) <= not (a and b);
    layer2_outputs(2235) <= b;
    layer2_outputs(2236) <= not b or a;
    layer2_outputs(2237) <= not a or b;
    layer2_outputs(2238) <= a or b;
    layer2_outputs(2239) <= a and b;
    layer2_outputs(2240) <= not (a or b);
    layer2_outputs(2241) <= b and not a;
    layer2_outputs(2242) <= a xor b;
    layer2_outputs(2243) <= '0';
    layer2_outputs(2244) <= not (a xor b);
    layer2_outputs(2245) <= not (a or b);
    layer2_outputs(2246) <= not b;
    layer2_outputs(2247) <= a or b;
    layer2_outputs(2248) <= '0';
    layer2_outputs(2249) <= b and not a;
    layer2_outputs(2250) <= not b or a;
    layer2_outputs(2251) <= b;
    layer2_outputs(2252) <= not a;
    layer2_outputs(2253) <= b and not a;
    layer2_outputs(2254) <= a and b;
    layer2_outputs(2255) <= not (a and b);
    layer2_outputs(2256) <= a and not b;
    layer2_outputs(2257) <= a;
    layer2_outputs(2258) <= not a;
    layer2_outputs(2259) <= not a;
    layer2_outputs(2260) <= not b;
    layer2_outputs(2261) <= not (a and b);
    layer2_outputs(2262) <= not a or b;
    layer2_outputs(2263) <= b;
    layer2_outputs(2264) <= not (a and b);
    layer2_outputs(2265) <= not (a and b);
    layer2_outputs(2266) <= not a or b;
    layer2_outputs(2267) <= a and b;
    layer2_outputs(2268) <= not a or b;
    layer2_outputs(2269) <= not b;
    layer2_outputs(2270) <= not b;
    layer2_outputs(2271) <= not (a and b);
    layer2_outputs(2272) <= not a;
    layer2_outputs(2273) <= a;
    layer2_outputs(2274) <= not (a or b);
    layer2_outputs(2275) <= '1';
    layer2_outputs(2276) <= '0';
    layer2_outputs(2277) <= not b or a;
    layer2_outputs(2278) <= a and not b;
    layer2_outputs(2279) <= not (a and b);
    layer2_outputs(2280) <= not b;
    layer2_outputs(2281) <= '0';
    layer2_outputs(2282) <= a;
    layer2_outputs(2283) <= a and not b;
    layer2_outputs(2284) <= a xor b;
    layer2_outputs(2285) <= a;
    layer2_outputs(2286) <= not b;
    layer2_outputs(2287) <= not b;
    layer2_outputs(2288) <= not b or a;
    layer2_outputs(2289) <= not a;
    layer2_outputs(2290) <= a;
    layer2_outputs(2291) <= a and not b;
    layer2_outputs(2292) <= not (a and b);
    layer2_outputs(2293) <= not (a and b);
    layer2_outputs(2294) <= not b or a;
    layer2_outputs(2295) <= not (a or b);
    layer2_outputs(2296) <= not a;
    layer2_outputs(2297) <= not b;
    layer2_outputs(2298) <= a or b;
    layer2_outputs(2299) <= not b or a;
    layer2_outputs(2300) <= a;
    layer2_outputs(2301) <= not (a and b);
    layer2_outputs(2302) <= not (a xor b);
    layer2_outputs(2303) <= b;
    layer2_outputs(2304) <= a or b;
    layer2_outputs(2305) <= not (a or b);
    layer2_outputs(2306) <= not b;
    layer2_outputs(2307) <= a or b;
    layer2_outputs(2308) <= not (a and b);
    layer2_outputs(2309) <= b;
    layer2_outputs(2310) <= '0';
    layer2_outputs(2311) <= a and not b;
    layer2_outputs(2312) <= b;
    layer2_outputs(2313) <= not b or a;
    layer2_outputs(2314) <= '0';
    layer2_outputs(2315) <= not (a or b);
    layer2_outputs(2316) <= b;
    layer2_outputs(2317) <= not (a or b);
    layer2_outputs(2318) <= not a;
    layer2_outputs(2319) <= '1';
    layer2_outputs(2320) <= not a or b;
    layer2_outputs(2321) <= not a;
    layer2_outputs(2322) <= not b;
    layer2_outputs(2323) <= a and b;
    layer2_outputs(2324) <= a and not b;
    layer2_outputs(2325) <= a;
    layer2_outputs(2326) <= a or b;
    layer2_outputs(2327) <= '0';
    layer2_outputs(2328) <= not a;
    layer2_outputs(2329) <= not b;
    layer2_outputs(2330) <= '0';
    layer2_outputs(2331) <= not a;
    layer2_outputs(2332) <= not b;
    layer2_outputs(2333) <= '1';
    layer2_outputs(2334) <= a;
    layer2_outputs(2335) <= a;
    layer2_outputs(2336) <= not (a and b);
    layer2_outputs(2337) <= a;
    layer2_outputs(2338) <= b;
    layer2_outputs(2339) <= not b;
    layer2_outputs(2340) <= not b or a;
    layer2_outputs(2341) <= not (a or b);
    layer2_outputs(2342) <= '0';
    layer2_outputs(2343) <= b and not a;
    layer2_outputs(2344) <= b and not a;
    layer2_outputs(2345) <= not a;
    layer2_outputs(2346) <= b;
    layer2_outputs(2347) <= not (a or b);
    layer2_outputs(2348) <= not (a or b);
    layer2_outputs(2349) <= a or b;
    layer2_outputs(2350) <= '0';
    layer2_outputs(2351) <= not (a or b);
    layer2_outputs(2352) <= not a or b;
    layer2_outputs(2353) <= '0';
    layer2_outputs(2354) <= '1';
    layer2_outputs(2355) <= a or b;
    layer2_outputs(2356) <= not (a xor b);
    layer2_outputs(2357) <= b;
    layer2_outputs(2358) <= b and not a;
    layer2_outputs(2359) <= not (a or b);
    layer2_outputs(2360) <= '0';
    layer2_outputs(2361) <= a and b;
    layer2_outputs(2362) <= not b or a;
    layer2_outputs(2363) <= not (a and b);
    layer2_outputs(2364) <= a;
    layer2_outputs(2365) <= '0';
    layer2_outputs(2366) <= not b or a;
    layer2_outputs(2367) <= b;
    layer2_outputs(2368) <= not (a and b);
    layer2_outputs(2369) <= a;
    layer2_outputs(2370) <= a or b;
    layer2_outputs(2371) <= a and b;
    layer2_outputs(2372) <= b;
    layer2_outputs(2373) <= a;
    layer2_outputs(2374) <= not a;
    layer2_outputs(2375) <= b and not a;
    layer2_outputs(2376) <= a;
    layer2_outputs(2377) <= not (a and b);
    layer2_outputs(2378) <= a and b;
    layer2_outputs(2379) <= not a;
    layer2_outputs(2380) <= not (a and b);
    layer2_outputs(2381) <= b;
    layer2_outputs(2382) <= not (a xor b);
    layer2_outputs(2383) <= b;
    layer2_outputs(2384) <= a or b;
    layer2_outputs(2385) <= not a;
    layer2_outputs(2386) <= not a;
    layer2_outputs(2387) <= a;
    layer2_outputs(2388) <= b and not a;
    layer2_outputs(2389) <= b;
    layer2_outputs(2390) <= a or b;
    layer2_outputs(2391) <= a;
    layer2_outputs(2392) <= b and not a;
    layer2_outputs(2393) <= not b;
    layer2_outputs(2394) <= not (a or b);
    layer2_outputs(2395) <= not a;
    layer2_outputs(2396) <= '0';
    layer2_outputs(2397) <= a or b;
    layer2_outputs(2398) <= not (a or b);
    layer2_outputs(2399) <= a and not b;
    layer2_outputs(2400) <= b and not a;
    layer2_outputs(2401) <= b;
    layer2_outputs(2402) <= a and b;
    layer2_outputs(2403) <= not a;
    layer2_outputs(2404) <= a;
    layer2_outputs(2405) <= a;
    layer2_outputs(2406) <= a xor b;
    layer2_outputs(2407) <= a and not b;
    layer2_outputs(2408) <= a;
    layer2_outputs(2409) <= a and not b;
    layer2_outputs(2410) <= not b;
    layer2_outputs(2411) <= '1';
    layer2_outputs(2412) <= b and not a;
    layer2_outputs(2413) <= a and b;
    layer2_outputs(2414) <= '1';
    layer2_outputs(2415) <= b;
    layer2_outputs(2416) <= '1';
    layer2_outputs(2417) <= not a or b;
    layer2_outputs(2418) <= b;
    layer2_outputs(2419) <= not (a and b);
    layer2_outputs(2420) <= not (a or b);
    layer2_outputs(2421) <= a and not b;
    layer2_outputs(2422) <= b;
    layer2_outputs(2423) <= not (a or b);
    layer2_outputs(2424) <= a and b;
    layer2_outputs(2425) <= a xor b;
    layer2_outputs(2426) <= a or b;
    layer2_outputs(2427) <= not b;
    layer2_outputs(2428) <= not a;
    layer2_outputs(2429) <= not a or b;
    layer2_outputs(2430) <= b;
    layer2_outputs(2431) <= not b or a;
    layer2_outputs(2432) <= a or b;
    layer2_outputs(2433) <= not (a xor b);
    layer2_outputs(2434) <= b;
    layer2_outputs(2435) <= a;
    layer2_outputs(2436) <= not b;
    layer2_outputs(2437) <= b;
    layer2_outputs(2438) <= a xor b;
    layer2_outputs(2439) <= not b or a;
    layer2_outputs(2440) <= a and b;
    layer2_outputs(2441) <= b;
    layer2_outputs(2442) <= not a;
    layer2_outputs(2443) <= not (a or b);
    layer2_outputs(2444) <= '0';
    layer2_outputs(2445) <= a and b;
    layer2_outputs(2446) <= not a;
    layer2_outputs(2447) <= b;
    layer2_outputs(2448) <= b and not a;
    layer2_outputs(2449) <= a and not b;
    layer2_outputs(2450) <= not a or b;
    layer2_outputs(2451) <= '1';
    layer2_outputs(2452) <= b;
    layer2_outputs(2453) <= not b;
    layer2_outputs(2454) <= not (a or b);
    layer2_outputs(2455) <= not a or b;
    layer2_outputs(2456) <= b;
    layer2_outputs(2457) <= a;
    layer2_outputs(2458) <= a and b;
    layer2_outputs(2459) <= b;
    layer2_outputs(2460) <= a;
    layer2_outputs(2461) <= not b or a;
    layer2_outputs(2462) <= a or b;
    layer2_outputs(2463) <= not a or b;
    layer2_outputs(2464) <= b;
    layer2_outputs(2465) <= not a;
    layer2_outputs(2466) <= a or b;
    layer2_outputs(2467) <= '1';
    layer2_outputs(2468) <= not a;
    layer2_outputs(2469) <= '0';
    layer2_outputs(2470) <= b and not a;
    layer2_outputs(2471) <= a;
    layer2_outputs(2472) <= not b;
    layer2_outputs(2473) <= a xor b;
    layer2_outputs(2474) <= not a;
    layer2_outputs(2475) <= b;
    layer2_outputs(2476) <= b;
    layer2_outputs(2477) <= '1';
    layer2_outputs(2478) <= not b;
    layer2_outputs(2479) <= a or b;
    layer2_outputs(2480) <= b;
    layer2_outputs(2481) <= a or b;
    layer2_outputs(2482) <= not a;
    layer2_outputs(2483) <= not (a or b);
    layer2_outputs(2484) <= '0';
    layer2_outputs(2485) <= not (a and b);
    layer2_outputs(2486) <= a;
    layer2_outputs(2487) <= not b or a;
    layer2_outputs(2488) <= not b;
    layer2_outputs(2489) <= not b;
    layer2_outputs(2490) <= not (a xor b);
    layer2_outputs(2491) <= a;
    layer2_outputs(2492) <= a and not b;
    layer2_outputs(2493) <= a;
    layer2_outputs(2494) <= a and b;
    layer2_outputs(2495) <= a and not b;
    layer2_outputs(2496) <= not (a or b);
    layer2_outputs(2497) <= '1';
    layer2_outputs(2498) <= '0';
    layer2_outputs(2499) <= not b;
    layer2_outputs(2500) <= not b;
    layer2_outputs(2501) <= not a;
    layer2_outputs(2502) <= not a;
    layer2_outputs(2503) <= '0';
    layer2_outputs(2504) <= a or b;
    layer2_outputs(2505) <= not b;
    layer2_outputs(2506) <= b and not a;
    layer2_outputs(2507) <= not b or a;
    layer2_outputs(2508) <= b;
    layer2_outputs(2509) <= b and not a;
    layer2_outputs(2510) <= a and not b;
    layer2_outputs(2511) <= b;
    layer2_outputs(2512) <= '1';
    layer2_outputs(2513) <= '0';
    layer2_outputs(2514) <= b;
    layer2_outputs(2515) <= not (a or b);
    layer2_outputs(2516) <= not a;
    layer2_outputs(2517) <= a or b;
    layer2_outputs(2518) <= b;
    layer2_outputs(2519) <= a or b;
    layer2_outputs(2520) <= b;
    layer2_outputs(2521) <= not a or b;
    layer2_outputs(2522) <= a;
    layer2_outputs(2523) <= '0';
    layer2_outputs(2524) <= a and b;
    layer2_outputs(2525) <= a and not b;
    layer2_outputs(2526) <= not b;
    layer2_outputs(2527) <= not a;
    layer2_outputs(2528) <= not b;
    layer2_outputs(2529) <= not (a and b);
    layer2_outputs(2530) <= '1';
    layer2_outputs(2531) <= '0';
    layer2_outputs(2532) <= '1';
    layer2_outputs(2533) <= not a or b;
    layer2_outputs(2534) <= not (a or b);
    layer2_outputs(2535) <= not a;
    layer2_outputs(2536) <= a;
    layer2_outputs(2537) <= '0';
    layer2_outputs(2538) <= a;
    layer2_outputs(2539) <= a and b;
    layer2_outputs(2540) <= a and b;
    layer2_outputs(2541) <= a or b;
    layer2_outputs(2542) <= not b;
    layer2_outputs(2543) <= a;
    layer2_outputs(2544) <= not a or b;
    layer2_outputs(2545) <= not b;
    layer2_outputs(2546) <= b;
    layer2_outputs(2547) <= a;
    layer2_outputs(2548) <= b;
    layer2_outputs(2549) <= b and not a;
    layer2_outputs(2550) <= a and not b;
    layer2_outputs(2551) <= not b;
    layer2_outputs(2552) <= a and not b;
    layer2_outputs(2553) <= b and not a;
    layer2_outputs(2554) <= b and not a;
    layer2_outputs(2555) <= a and not b;
    layer2_outputs(2556) <= not b or a;
    layer2_outputs(2557) <= a;
    layer2_outputs(2558) <= not (a or b);
    layer2_outputs(2559) <= '1';
    layer2_outputs(2560) <= a xor b;
    layer2_outputs(2561) <= a or b;
    layer2_outputs(2562) <= a or b;
    layer2_outputs(2563) <= b and not a;
    layer2_outputs(2564) <= not a or b;
    layer2_outputs(2565) <= a or b;
    layer2_outputs(2566) <= b;
    layer2_outputs(2567) <= b and not a;
    layer2_outputs(2568) <= a and not b;
    layer2_outputs(2569) <= b;
    layer2_outputs(2570) <= not a or b;
    layer2_outputs(2571) <= a xor b;
    layer2_outputs(2572) <= not a;
    layer2_outputs(2573) <= a;
    layer2_outputs(2574) <= a;
    layer2_outputs(2575) <= b and not a;
    layer2_outputs(2576) <= a;
    layer2_outputs(2577) <= not (a and b);
    layer2_outputs(2578) <= '1';
    layer2_outputs(2579) <= not b;
    layer2_outputs(2580) <= not (a or b);
    layer2_outputs(2581) <= b;
    layer2_outputs(2582) <= not (a or b);
    layer2_outputs(2583) <= b and not a;
    layer2_outputs(2584) <= b;
    layer2_outputs(2585) <= a xor b;
    layer2_outputs(2586) <= a or b;
    layer2_outputs(2587) <= a;
    layer2_outputs(2588) <= not (a and b);
    layer2_outputs(2589) <= not b;
    layer2_outputs(2590) <= not a or b;
    layer2_outputs(2591) <= a or b;
    layer2_outputs(2592) <= a and not b;
    layer2_outputs(2593) <= not a;
    layer2_outputs(2594) <= '0';
    layer2_outputs(2595) <= a and not b;
    layer2_outputs(2596) <= a;
    layer2_outputs(2597) <= '1';
    layer2_outputs(2598) <= '1';
    layer2_outputs(2599) <= b;
    layer2_outputs(2600) <= a and not b;
    layer2_outputs(2601) <= b;
    layer2_outputs(2602) <= '0';
    layer2_outputs(2603) <= b;
    layer2_outputs(2604) <= a xor b;
    layer2_outputs(2605) <= not (a and b);
    layer2_outputs(2606) <= not (a xor b);
    layer2_outputs(2607) <= a and not b;
    layer2_outputs(2608) <= not a;
    layer2_outputs(2609) <= b and not a;
    layer2_outputs(2610) <= a and b;
    layer2_outputs(2611) <= '1';
    layer2_outputs(2612) <= not (a or b);
    layer2_outputs(2613) <= not a;
    layer2_outputs(2614) <= not a or b;
    layer2_outputs(2615) <= a and b;
    layer2_outputs(2616) <= not (a or b);
    layer2_outputs(2617) <= b;
    layer2_outputs(2618) <= b;
    layer2_outputs(2619) <= a or b;
    layer2_outputs(2620) <= '1';
    layer2_outputs(2621) <= '1';
    layer2_outputs(2622) <= not a or b;
    layer2_outputs(2623) <= b and not a;
    layer2_outputs(2624) <= not b or a;
    layer2_outputs(2625) <= b and not a;
    layer2_outputs(2626) <= a or b;
    layer2_outputs(2627) <= not a;
    layer2_outputs(2628) <= not (a and b);
    layer2_outputs(2629) <= not a;
    layer2_outputs(2630) <= '1';
    layer2_outputs(2631) <= a and not b;
    layer2_outputs(2632) <= not a;
    layer2_outputs(2633) <= b;
    layer2_outputs(2634) <= a;
    layer2_outputs(2635) <= a and not b;
    layer2_outputs(2636) <= '0';
    layer2_outputs(2637) <= b and not a;
    layer2_outputs(2638) <= not a;
    layer2_outputs(2639) <= a;
    layer2_outputs(2640) <= b and not a;
    layer2_outputs(2641) <= a and not b;
    layer2_outputs(2642) <= a;
    layer2_outputs(2643) <= not a or b;
    layer2_outputs(2644) <= not (a and b);
    layer2_outputs(2645) <= not (a xor b);
    layer2_outputs(2646) <= a xor b;
    layer2_outputs(2647) <= a;
    layer2_outputs(2648) <= a;
    layer2_outputs(2649) <= '0';
    layer2_outputs(2650) <= not (a or b);
    layer2_outputs(2651) <= a or b;
    layer2_outputs(2652) <= not b;
    layer2_outputs(2653) <= not a;
    layer2_outputs(2654) <= not a;
    layer2_outputs(2655) <= a xor b;
    layer2_outputs(2656) <= b;
    layer2_outputs(2657) <= a or b;
    layer2_outputs(2658) <= a and b;
    layer2_outputs(2659) <= not a;
    layer2_outputs(2660) <= not b;
    layer2_outputs(2661) <= a and not b;
    layer2_outputs(2662) <= not a;
    layer2_outputs(2663) <= b and not a;
    layer2_outputs(2664) <= not b or a;
    layer2_outputs(2665) <= not (a or b);
    layer2_outputs(2666) <= not (a or b);
    layer2_outputs(2667) <= '1';
    layer2_outputs(2668) <= a and b;
    layer2_outputs(2669) <= not (a and b);
    layer2_outputs(2670) <= not b or a;
    layer2_outputs(2671) <= not b;
    layer2_outputs(2672) <= a and b;
    layer2_outputs(2673) <= a;
    layer2_outputs(2674) <= a;
    layer2_outputs(2675) <= b;
    layer2_outputs(2676) <= b and not a;
    layer2_outputs(2677) <= b and not a;
    layer2_outputs(2678) <= not (a and b);
    layer2_outputs(2679) <= '0';
    layer2_outputs(2680) <= '1';
    layer2_outputs(2681) <= b;
    layer2_outputs(2682) <= '1';
    layer2_outputs(2683) <= not (a or b);
    layer2_outputs(2684) <= b;
    layer2_outputs(2685) <= a or b;
    layer2_outputs(2686) <= not (a or b);
    layer2_outputs(2687) <= b and not a;
    layer2_outputs(2688) <= '1';
    layer2_outputs(2689) <= a and not b;
    layer2_outputs(2690) <= not (a or b);
    layer2_outputs(2691) <= b and not a;
    layer2_outputs(2692) <= not a;
    layer2_outputs(2693) <= b and not a;
    layer2_outputs(2694) <= not (a and b);
    layer2_outputs(2695) <= '0';
    layer2_outputs(2696) <= not b;
    layer2_outputs(2697) <= b;
    layer2_outputs(2698) <= not a;
    layer2_outputs(2699) <= a and b;
    layer2_outputs(2700) <= not a;
    layer2_outputs(2701) <= b;
    layer2_outputs(2702) <= b and not a;
    layer2_outputs(2703) <= a and not b;
    layer2_outputs(2704) <= b and not a;
    layer2_outputs(2705) <= b;
    layer2_outputs(2706) <= not a;
    layer2_outputs(2707) <= a and not b;
    layer2_outputs(2708) <= not (a and b);
    layer2_outputs(2709) <= not a or b;
    layer2_outputs(2710) <= not (a and b);
    layer2_outputs(2711) <= a;
    layer2_outputs(2712) <= b and not a;
    layer2_outputs(2713) <= a or b;
    layer2_outputs(2714) <= a xor b;
    layer2_outputs(2715) <= a or b;
    layer2_outputs(2716) <= '1';
    layer2_outputs(2717) <= not a or b;
    layer2_outputs(2718) <= b and not a;
    layer2_outputs(2719) <= not b;
    layer2_outputs(2720) <= a and not b;
    layer2_outputs(2721) <= not (a and b);
    layer2_outputs(2722) <= not b;
    layer2_outputs(2723) <= a or b;
    layer2_outputs(2724) <= b and not a;
    layer2_outputs(2725) <= not a;
    layer2_outputs(2726) <= not a;
    layer2_outputs(2727) <= b and not a;
    layer2_outputs(2728) <= not b;
    layer2_outputs(2729) <= a and b;
    layer2_outputs(2730) <= not a;
    layer2_outputs(2731) <= a;
    layer2_outputs(2732) <= not a;
    layer2_outputs(2733) <= a;
    layer2_outputs(2734) <= '0';
    layer2_outputs(2735) <= a and b;
    layer2_outputs(2736) <= not b;
    layer2_outputs(2737) <= a and b;
    layer2_outputs(2738) <= a or b;
    layer2_outputs(2739) <= a or b;
    layer2_outputs(2740) <= a;
    layer2_outputs(2741) <= a;
    layer2_outputs(2742) <= a and not b;
    layer2_outputs(2743) <= a or b;
    layer2_outputs(2744) <= a or b;
    layer2_outputs(2745) <= not a;
    layer2_outputs(2746) <= a or b;
    layer2_outputs(2747) <= a and not b;
    layer2_outputs(2748) <= b;
    layer2_outputs(2749) <= a and b;
    layer2_outputs(2750) <= a or b;
    layer2_outputs(2751) <= a or b;
    layer2_outputs(2752) <= not b;
    layer2_outputs(2753) <= not (a and b);
    layer2_outputs(2754) <= a;
    layer2_outputs(2755) <= not b or a;
    layer2_outputs(2756) <= a and not b;
    layer2_outputs(2757) <= not b or a;
    layer2_outputs(2758) <= b;
    layer2_outputs(2759) <= not (a or b);
    layer2_outputs(2760) <= b and not a;
    layer2_outputs(2761) <= a and b;
    layer2_outputs(2762) <= a or b;
    layer2_outputs(2763) <= b and not a;
    layer2_outputs(2764) <= b and not a;
    layer2_outputs(2765) <= '1';
    layer2_outputs(2766) <= not (a and b);
    layer2_outputs(2767) <= b;
    layer2_outputs(2768) <= not b or a;
    layer2_outputs(2769) <= not a;
    layer2_outputs(2770) <= a and b;
    layer2_outputs(2771) <= not b or a;
    layer2_outputs(2772) <= '1';
    layer2_outputs(2773) <= '1';
    layer2_outputs(2774) <= '0';
    layer2_outputs(2775) <= not b;
    layer2_outputs(2776) <= a and b;
    layer2_outputs(2777) <= a and b;
    layer2_outputs(2778) <= not a;
    layer2_outputs(2779) <= b;
    layer2_outputs(2780) <= '0';
    layer2_outputs(2781) <= '1';
    layer2_outputs(2782) <= not b;
    layer2_outputs(2783) <= b;
    layer2_outputs(2784) <= not a or b;
    layer2_outputs(2785) <= b;
    layer2_outputs(2786) <= a;
    layer2_outputs(2787) <= b and not a;
    layer2_outputs(2788) <= not (a and b);
    layer2_outputs(2789) <= b and not a;
    layer2_outputs(2790) <= not a or b;
    layer2_outputs(2791) <= not (a or b);
    layer2_outputs(2792) <= b;
    layer2_outputs(2793) <= b and not a;
    layer2_outputs(2794) <= '0';
    layer2_outputs(2795) <= a;
    layer2_outputs(2796) <= a and not b;
    layer2_outputs(2797) <= not b or a;
    layer2_outputs(2798) <= not b;
    layer2_outputs(2799) <= a or b;
    layer2_outputs(2800) <= not (a or b);
    layer2_outputs(2801) <= '1';
    layer2_outputs(2802) <= not b;
    layer2_outputs(2803) <= not (a or b);
    layer2_outputs(2804) <= a and b;
    layer2_outputs(2805) <= a;
    layer2_outputs(2806) <= not b or a;
    layer2_outputs(2807) <= a or b;
    layer2_outputs(2808) <= a;
    layer2_outputs(2809) <= a and b;
    layer2_outputs(2810) <= a and not b;
    layer2_outputs(2811) <= a and b;
    layer2_outputs(2812) <= not b or a;
    layer2_outputs(2813) <= b;
    layer2_outputs(2814) <= a xor b;
    layer2_outputs(2815) <= not b;
    layer2_outputs(2816) <= not a;
    layer2_outputs(2817) <= not a or b;
    layer2_outputs(2818) <= not b;
    layer2_outputs(2819) <= not b;
    layer2_outputs(2820) <= b;
    layer2_outputs(2821) <= not a;
    layer2_outputs(2822) <= a xor b;
    layer2_outputs(2823) <= a or b;
    layer2_outputs(2824) <= a and not b;
    layer2_outputs(2825) <= not a or b;
    layer2_outputs(2826) <= not b or a;
    layer2_outputs(2827) <= not a;
    layer2_outputs(2828) <= not a or b;
    layer2_outputs(2829) <= a;
    layer2_outputs(2830) <= not b;
    layer2_outputs(2831) <= a;
    layer2_outputs(2832) <= '1';
    layer2_outputs(2833) <= a or b;
    layer2_outputs(2834) <= a or b;
    layer2_outputs(2835) <= not (a or b);
    layer2_outputs(2836) <= not (a or b);
    layer2_outputs(2837) <= a and b;
    layer2_outputs(2838) <= not a or b;
    layer2_outputs(2839) <= not b;
    layer2_outputs(2840) <= '1';
    layer2_outputs(2841) <= not b;
    layer2_outputs(2842) <= a and not b;
    layer2_outputs(2843) <= '1';
    layer2_outputs(2844) <= not (a or b);
    layer2_outputs(2845) <= not a;
    layer2_outputs(2846) <= a or b;
    layer2_outputs(2847) <= a or b;
    layer2_outputs(2848) <= a or b;
    layer2_outputs(2849) <= '0';
    layer2_outputs(2850) <= b;
    layer2_outputs(2851) <= a;
    layer2_outputs(2852) <= a and not b;
    layer2_outputs(2853) <= not b;
    layer2_outputs(2854) <= not a;
    layer2_outputs(2855) <= not b or a;
    layer2_outputs(2856) <= not b;
    layer2_outputs(2857) <= b;
    layer2_outputs(2858) <= a and not b;
    layer2_outputs(2859) <= not b or a;
    layer2_outputs(2860) <= b;
    layer2_outputs(2861) <= not a or b;
    layer2_outputs(2862) <= b;
    layer2_outputs(2863) <= a and b;
    layer2_outputs(2864) <= a xor b;
    layer2_outputs(2865) <= a;
    layer2_outputs(2866) <= a or b;
    layer2_outputs(2867) <= '0';
    layer2_outputs(2868) <= not a or b;
    layer2_outputs(2869) <= a or b;
    layer2_outputs(2870) <= not a;
    layer2_outputs(2871) <= a and b;
    layer2_outputs(2872) <= a and b;
    layer2_outputs(2873) <= b and not a;
    layer2_outputs(2874) <= a or b;
    layer2_outputs(2875) <= '1';
    layer2_outputs(2876) <= a and b;
    layer2_outputs(2877) <= not b or a;
    layer2_outputs(2878) <= b;
    layer2_outputs(2879) <= not (a or b);
    layer2_outputs(2880) <= not a;
    layer2_outputs(2881) <= a and not b;
    layer2_outputs(2882) <= '0';
    layer2_outputs(2883) <= a or b;
    layer2_outputs(2884) <= not a;
    layer2_outputs(2885) <= not (a or b);
    layer2_outputs(2886) <= a xor b;
    layer2_outputs(2887) <= not (a xor b);
    layer2_outputs(2888) <= a and not b;
    layer2_outputs(2889) <= not a;
    layer2_outputs(2890) <= a and b;
    layer2_outputs(2891) <= not b or a;
    layer2_outputs(2892) <= a and not b;
    layer2_outputs(2893) <= not (a xor b);
    layer2_outputs(2894) <= a and b;
    layer2_outputs(2895) <= a or b;
    layer2_outputs(2896) <= '1';
    layer2_outputs(2897) <= b;
    layer2_outputs(2898) <= a and not b;
    layer2_outputs(2899) <= not (a xor b);
    layer2_outputs(2900) <= a or b;
    layer2_outputs(2901) <= '0';
    layer2_outputs(2902) <= not (a and b);
    layer2_outputs(2903) <= a and b;
    layer2_outputs(2904) <= a or b;
    layer2_outputs(2905) <= b;
    layer2_outputs(2906) <= '1';
    layer2_outputs(2907) <= not a or b;
    layer2_outputs(2908) <= a or b;
    layer2_outputs(2909) <= not a;
    layer2_outputs(2910) <= not b or a;
    layer2_outputs(2911) <= not b or a;
    layer2_outputs(2912) <= not b;
    layer2_outputs(2913) <= a;
    layer2_outputs(2914) <= not b;
    layer2_outputs(2915) <= not a or b;
    layer2_outputs(2916) <= '1';
    layer2_outputs(2917) <= a;
    layer2_outputs(2918) <= not b;
    layer2_outputs(2919) <= not a;
    layer2_outputs(2920) <= not a;
    layer2_outputs(2921) <= a and not b;
    layer2_outputs(2922) <= not a;
    layer2_outputs(2923) <= b;
    layer2_outputs(2924) <= '0';
    layer2_outputs(2925) <= '1';
    layer2_outputs(2926) <= b and not a;
    layer2_outputs(2927) <= b;
    layer2_outputs(2928) <= '1';
    layer2_outputs(2929) <= not a;
    layer2_outputs(2930) <= not b or a;
    layer2_outputs(2931) <= '1';
    layer2_outputs(2932) <= b;
    layer2_outputs(2933) <= not b;
    layer2_outputs(2934) <= not (a and b);
    layer2_outputs(2935) <= '0';
    layer2_outputs(2936) <= not (a or b);
    layer2_outputs(2937) <= not (a xor b);
    layer2_outputs(2938) <= not b or a;
    layer2_outputs(2939) <= not b or a;
    layer2_outputs(2940) <= not b;
    layer2_outputs(2941) <= not b or a;
    layer2_outputs(2942) <= b and not a;
    layer2_outputs(2943) <= a xor b;
    layer2_outputs(2944) <= not b;
    layer2_outputs(2945) <= not b or a;
    layer2_outputs(2946) <= a and not b;
    layer2_outputs(2947) <= '0';
    layer2_outputs(2948) <= a and b;
    layer2_outputs(2949) <= '1';
    layer2_outputs(2950) <= a and b;
    layer2_outputs(2951) <= not b;
    layer2_outputs(2952) <= not (a and b);
    layer2_outputs(2953) <= a;
    layer2_outputs(2954) <= not b or a;
    layer2_outputs(2955) <= b;
    layer2_outputs(2956) <= b;
    layer2_outputs(2957) <= a;
    layer2_outputs(2958) <= b;
    layer2_outputs(2959) <= not b;
    layer2_outputs(2960) <= not b or a;
    layer2_outputs(2961) <= not a;
    layer2_outputs(2962) <= b and not a;
    layer2_outputs(2963) <= not (a xor b);
    layer2_outputs(2964) <= not a;
    layer2_outputs(2965) <= not b;
    layer2_outputs(2966) <= b;
    layer2_outputs(2967) <= '1';
    layer2_outputs(2968) <= b;
    layer2_outputs(2969) <= a or b;
    layer2_outputs(2970) <= not a;
    layer2_outputs(2971) <= a;
    layer2_outputs(2972) <= b;
    layer2_outputs(2973) <= not b;
    layer2_outputs(2974) <= not b;
    layer2_outputs(2975) <= not (a and b);
    layer2_outputs(2976) <= not (a xor b);
    layer2_outputs(2977) <= not (a xor b);
    layer2_outputs(2978) <= a and not b;
    layer2_outputs(2979) <= b;
    layer2_outputs(2980) <= not b;
    layer2_outputs(2981) <= not b or a;
    layer2_outputs(2982) <= not a or b;
    layer2_outputs(2983) <= not a;
    layer2_outputs(2984) <= '0';
    layer2_outputs(2985) <= not b;
    layer2_outputs(2986) <= b and not a;
    layer2_outputs(2987) <= b;
    layer2_outputs(2988) <= a and not b;
    layer2_outputs(2989) <= not (a xor b);
    layer2_outputs(2990) <= '1';
    layer2_outputs(2991) <= a;
    layer2_outputs(2992) <= '0';
    layer2_outputs(2993) <= a and not b;
    layer2_outputs(2994) <= a and not b;
    layer2_outputs(2995) <= a;
    layer2_outputs(2996) <= a or b;
    layer2_outputs(2997) <= not b or a;
    layer2_outputs(2998) <= a;
    layer2_outputs(2999) <= a and b;
    layer2_outputs(3000) <= not (a xor b);
    layer2_outputs(3001) <= '0';
    layer2_outputs(3002) <= a and not b;
    layer2_outputs(3003) <= not (a or b);
    layer2_outputs(3004) <= not (a and b);
    layer2_outputs(3005) <= not (a and b);
    layer2_outputs(3006) <= not b or a;
    layer2_outputs(3007) <= not (a and b);
    layer2_outputs(3008) <= not (a or b);
    layer2_outputs(3009) <= a;
    layer2_outputs(3010) <= not a or b;
    layer2_outputs(3011) <= not b or a;
    layer2_outputs(3012) <= a;
    layer2_outputs(3013) <= not (a or b);
    layer2_outputs(3014) <= not b or a;
    layer2_outputs(3015) <= b and not a;
    layer2_outputs(3016) <= b and not a;
    layer2_outputs(3017) <= not (a and b);
    layer2_outputs(3018) <= b;
    layer2_outputs(3019) <= not a or b;
    layer2_outputs(3020) <= not (a or b);
    layer2_outputs(3021) <= not (a and b);
    layer2_outputs(3022) <= a and not b;
    layer2_outputs(3023) <= b and not a;
    layer2_outputs(3024) <= b and not a;
    layer2_outputs(3025) <= not (a xor b);
    layer2_outputs(3026) <= b;
    layer2_outputs(3027) <= b;
    layer2_outputs(3028) <= '1';
    layer2_outputs(3029) <= '0';
    layer2_outputs(3030) <= a and not b;
    layer2_outputs(3031) <= a and b;
    layer2_outputs(3032) <= b and not a;
    layer2_outputs(3033) <= a and b;
    layer2_outputs(3034) <= a and b;
    layer2_outputs(3035) <= a;
    layer2_outputs(3036) <= b and not a;
    layer2_outputs(3037) <= not b or a;
    layer2_outputs(3038) <= b and not a;
    layer2_outputs(3039) <= b;
    layer2_outputs(3040) <= not b;
    layer2_outputs(3041) <= '1';
    layer2_outputs(3042) <= a;
    layer2_outputs(3043) <= '1';
    layer2_outputs(3044) <= not b or a;
    layer2_outputs(3045) <= not b;
    layer2_outputs(3046) <= b;
    layer2_outputs(3047) <= not b;
    layer2_outputs(3048) <= b;
    layer2_outputs(3049) <= not b;
    layer2_outputs(3050) <= b and not a;
    layer2_outputs(3051) <= not a;
    layer2_outputs(3052) <= a or b;
    layer2_outputs(3053) <= not b;
    layer2_outputs(3054) <= b;
    layer2_outputs(3055) <= '1';
    layer2_outputs(3056) <= '0';
    layer2_outputs(3057) <= not b or a;
    layer2_outputs(3058) <= not (a and b);
    layer2_outputs(3059) <= '1';
    layer2_outputs(3060) <= not a or b;
    layer2_outputs(3061) <= not b;
    layer2_outputs(3062) <= '1';
    layer2_outputs(3063) <= a;
    layer2_outputs(3064) <= not a;
    layer2_outputs(3065) <= b and not a;
    layer2_outputs(3066) <= b;
    layer2_outputs(3067) <= a xor b;
    layer2_outputs(3068) <= a;
    layer2_outputs(3069) <= a or b;
    layer2_outputs(3070) <= a and b;
    layer2_outputs(3071) <= '1';
    layer2_outputs(3072) <= not (a or b);
    layer2_outputs(3073) <= not a or b;
    layer2_outputs(3074) <= a;
    layer2_outputs(3075) <= b;
    layer2_outputs(3076) <= a and not b;
    layer2_outputs(3077) <= not (a or b);
    layer2_outputs(3078) <= b;
    layer2_outputs(3079) <= not b;
    layer2_outputs(3080) <= b and not a;
    layer2_outputs(3081) <= '1';
    layer2_outputs(3082) <= b and not a;
    layer2_outputs(3083) <= not a;
    layer2_outputs(3084) <= a and b;
    layer2_outputs(3085) <= '1';
    layer2_outputs(3086) <= not a or b;
    layer2_outputs(3087) <= a and not b;
    layer2_outputs(3088) <= not b;
    layer2_outputs(3089) <= not (a or b);
    layer2_outputs(3090) <= b and not a;
    layer2_outputs(3091) <= '1';
    layer2_outputs(3092) <= not (a and b);
    layer2_outputs(3093) <= not a or b;
    layer2_outputs(3094) <= not b or a;
    layer2_outputs(3095) <= '0';
    layer2_outputs(3096) <= '1';
    layer2_outputs(3097) <= not b;
    layer2_outputs(3098) <= not (a and b);
    layer2_outputs(3099) <= '0';
    layer2_outputs(3100) <= not (a and b);
    layer2_outputs(3101) <= a and not b;
    layer2_outputs(3102) <= not b or a;
    layer2_outputs(3103) <= '0';
    layer2_outputs(3104) <= a and not b;
    layer2_outputs(3105) <= not b or a;
    layer2_outputs(3106) <= not b;
    layer2_outputs(3107) <= not a;
    layer2_outputs(3108) <= not b;
    layer2_outputs(3109) <= a or b;
    layer2_outputs(3110) <= '0';
    layer2_outputs(3111) <= b and not a;
    layer2_outputs(3112) <= not a;
    layer2_outputs(3113) <= a or b;
    layer2_outputs(3114) <= b;
    layer2_outputs(3115) <= b and not a;
    layer2_outputs(3116) <= not b;
    layer2_outputs(3117) <= a;
    layer2_outputs(3118) <= not (a and b);
    layer2_outputs(3119) <= a and not b;
    layer2_outputs(3120) <= not b;
    layer2_outputs(3121) <= not (a and b);
    layer2_outputs(3122) <= a;
    layer2_outputs(3123) <= a;
    layer2_outputs(3124) <= not (a xor b);
    layer2_outputs(3125) <= '0';
    layer2_outputs(3126) <= b and not a;
    layer2_outputs(3127) <= a;
    layer2_outputs(3128) <= not (a and b);
    layer2_outputs(3129) <= '0';
    layer2_outputs(3130) <= not b or a;
    layer2_outputs(3131) <= not a;
    layer2_outputs(3132) <= not a;
    layer2_outputs(3133) <= b;
    layer2_outputs(3134) <= not a;
    layer2_outputs(3135) <= not a or b;
    layer2_outputs(3136) <= a;
    layer2_outputs(3137) <= b;
    layer2_outputs(3138) <= not a;
    layer2_outputs(3139) <= not a or b;
    layer2_outputs(3140) <= not b or a;
    layer2_outputs(3141) <= b and not a;
    layer2_outputs(3142) <= not (a or b);
    layer2_outputs(3143) <= b;
    layer2_outputs(3144) <= b and not a;
    layer2_outputs(3145) <= a;
    layer2_outputs(3146) <= not a;
    layer2_outputs(3147) <= not b;
    layer2_outputs(3148) <= a;
    layer2_outputs(3149) <= b;
    layer2_outputs(3150) <= not (a xor b);
    layer2_outputs(3151) <= a or b;
    layer2_outputs(3152) <= not a;
    layer2_outputs(3153) <= b;
    layer2_outputs(3154) <= a;
    layer2_outputs(3155) <= not (a and b);
    layer2_outputs(3156) <= a or b;
    layer2_outputs(3157) <= '1';
    layer2_outputs(3158) <= '1';
    layer2_outputs(3159) <= not a;
    layer2_outputs(3160) <= a;
    layer2_outputs(3161) <= a;
    layer2_outputs(3162) <= a;
    layer2_outputs(3163) <= a and b;
    layer2_outputs(3164) <= '1';
    layer2_outputs(3165) <= '1';
    layer2_outputs(3166) <= not (a xor b);
    layer2_outputs(3167) <= a and not b;
    layer2_outputs(3168) <= not b;
    layer2_outputs(3169) <= not a;
    layer2_outputs(3170) <= b and not a;
    layer2_outputs(3171) <= not a;
    layer2_outputs(3172) <= a and b;
    layer2_outputs(3173) <= not a;
    layer2_outputs(3174) <= b and not a;
    layer2_outputs(3175) <= not (a or b);
    layer2_outputs(3176) <= a and not b;
    layer2_outputs(3177) <= b and not a;
    layer2_outputs(3178) <= '0';
    layer2_outputs(3179) <= a and b;
    layer2_outputs(3180) <= not (a and b);
    layer2_outputs(3181) <= not a;
    layer2_outputs(3182) <= not b;
    layer2_outputs(3183) <= '1';
    layer2_outputs(3184) <= b and not a;
    layer2_outputs(3185) <= a and not b;
    layer2_outputs(3186) <= not (a xor b);
    layer2_outputs(3187) <= not b;
    layer2_outputs(3188) <= b;
    layer2_outputs(3189) <= a and b;
    layer2_outputs(3190) <= a;
    layer2_outputs(3191) <= not b or a;
    layer2_outputs(3192) <= not b or a;
    layer2_outputs(3193) <= a and b;
    layer2_outputs(3194) <= not (a or b);
    layer2_outputs(3195) <= not b;
    layer2_outputs(3196) <= a;
    layer2_outputs(3197) <= '0';
    layer2_outputs(3198) <= not b;
    layer2_outputs(3199) <= a or b;
    layer2_outputs(3200) <= a and b;
    layer2_outputs(3201) <= a and not b;
    layer2_outputs(3202) <= a or b;
    layer2_outputs(3203) <= b and not a;
    layer2_outputs(3204) <= b;
    layer2_outputs(3205) <= not a or b;
    layer2_outputs(3206) <= not (a and b);
    layer2_outputs(3207) <= not b;
    layer2_outputs(3208) <= a xor b;
    layer2_outputs(3209) <= not a or b;
    layer2_outputs(3210) <= a xor b;
    layer2_outputs(3211) <= b;
    layer2_outputs(3212) <= a and not b;
    layer2_outputs(3213) <= a and b;
    layer2_outputs(3214) <= not a or b;
    layer2_outputs(3215) <= a xor b;
    layer2_outputs(3216) <= a and not b;
    layer2_outputs(3217) <= not (a xor b);
    layer2_outputs(3218) <= '0';
    layer2_outputs(3219) <= not a or b;
    layer2_outputs(3220) <= a;
    layer2_outputs(3221) <= not (a or b);
    layer2_outputs(3222) <= '0';
    layer2_outputs(3223) <= not (a or b);
    layer2_outputs(3224) <= b;
    layer2_outputs(3225) <= not a or b;
    layer2_outputs(3226) <= a or b;
    layer2_outputs(3227) <= a or b;
    layer2_outputs(3228) <= not a;
    layer2_outputs(3229) <= not a or b;
    layer2_outputs(3230) <= a or b;
    layer2_outputs(3231) <= not a;
    layer2_outputs(3232) <= not (a xor b);
    layer2_outputs(3233) <= a;
    layer2_outputs(3234) <= a xor b;
    layer2_outputs(3235) <= a and not b;
    layer2_outputs(3236) <= a and b;
    layer2_outputs(3237) <= '1';
    layer2_outputs(3238) <= '0';
    layer2_outputs(3239) <= '1';
    layer2_outputs(3240) <= not b or a;
    layer2_outputs(3241) <= not a;
    layer2_outputs(3242) <= not a;
    layer2_outputs(3243) <= not b or a;
    layer2_outputs(3244) <= b and not a;
    layer2_outputs(3245) <= b and not a;
    layer2_outputs(3246) <= a or b;
    layer2_outputs(3247) <= not (a or b);
    layer2_outputs(3248) <= not a;
    layer2_outputs(3249) <= not a or b;
    layer2_outputs(3250) <= a;
    layer2_outputs(3251) <= not b;
    layer2_outputs(3252) <= a;
    layer2_outputs(3253) <= b;
    layer2_outputs(3254) <= not a or b;
    layer2_outputs(3255) <= not (a and b);
    layer2_outputs(3256) <= b;
    layer2_outputs(3257) <= b and not a;
    layer2_outputs(3258) <= not b or a;
    layer2_outputs(3259) <= not b;
    layer2_outputs(3260) <= a xor b;
    layer2_outputs(3261) <= not (a xor b);
    layer2_outputs(3262) <= not b;
    layer2_outputs(3263) <= b and not a;
    layer2_outputs(3264) <= '0';
    layer2_outputs(3265) <= not (a and b);
    layer2_outputs(3266) <= not b;
    layer2_outputs(3267) <= not a or b;
    layer2_outputs(3268) <= a and b;
    layer2_outputs(3269) <= b and not a;
    layer2_outputs(3270) <= '0';
    layer2_outputs(3271) <= a and b;
    layer2_outputs(3272) <= not b or a;
    layer2_outputs(3273) <= not b;
    layer2_outputs(3274) <= a or b;
    layer2_outputs(3275) <= a;
    layer2_outputs(3276) <= a or b;
    layer2_outputs(3277) <= b;
    layer2_outputs(3278) <= a xor b;
    layer2_outputs(3279) <= '1';
    layer2_outputs(3280) <= not a or b;
    layer2_outputs(3281) <= not (a and b);
    layer2_outputs(3282) <= not b;
    layer2_outputs(3283) <= not a;
    layer2_outputs(3284) <= a or b;
    layer2_outputs(3285) <= not (a xor b);
    layer2_outputs(3286) <= not (a and b);
    layer2_outputs(3287) <= not b or a;
    layer2_outputs(3288) <= not b;
    layer2_outputs(3289) <= a;
    layer2_outputs(3290) <= a or b;
    layer2_outputs(3291) <= a and not b;
    layer2_outputs(3292) <= not a;
    layer2_outputs(3293) <= not (a or b);
    layer2_outputs(3294) <= not (a and b);
    layer2_outputs(3295) <= a and b;
    layer2_outputs(3296) <= not (a and b);
    layer2_outputs(3297) <= not (a or b);
    layer2_outputs(3298) <= a and b;
    layer2_outputs(3299) <= a and b;
    layer2_outputs(3300) <= a and not b;
    layer2_outputs(3301) <= a or b;
    layer2_outputs(3302) <= not b or a;
    layer2_outputs(3303) <= not a;
    layer2_outputs(3304) <= b and not a;
    layer2_outputs(3305) <= a or b;
    layer2_outputs(3306) <= '0';
    layer2_outputs(3307) <= not b;
    layer2_outputs(3308) <= b;
    layer2_outputs(3309) <= a and not b;
    layer2_outputs(3310) <= not a or b;
    layer2_outputs(3311) <= not (a and b);
    layer2_outputs(3312) <= a and b;
    layer2_outputs(3313) <= a and not b;
    layer2_outputs(3314) <= '0';
    layer2_outputs(3315) <= not a or b;
    layer2_outputs(3316) <= a xor b;
    layer2_outputs(3317) <= b;
    layer2_outputs(3318) <= not a;
    layer2_outputs(3319) <= not a or b;
    layer2_outputs(3320) <= not (a xor b);
    layer2_outputs(3321) <= a or b;
    layer2_outputs(3322) <= not b;
    layer2_outputs(3323) <= '1';
    layer2_outputs(3324) <= not (a and b);
    layer2_outputs(3325) <= '1';
    layer2_outputs(3326) <= a or b;
    layer2_outputs(3327) <= not a or b;
    layer2_outputs(3328) <= not (a and b);
    layer2_outputs(3329) <= not b;
    layer2_outputs(3330) <= '1';
    layer2_outputs(3331) <= a and b;
    layer2_outputs(3332) <= not b or a;
    layer2_outputs(3333) <= '0';
    layer2_outputs(3334) <= a and not b;
    layer2_outputs(3335) <= not (a or b);
    layer2_outputs(3336) <= b and not a;
    layer2_outputs(3337) <= not (a or b);
    layer2_outputs(3338) <= a;
    layer2_outputs(3339) <= not b;
    layer2_outputs(3340) <= a;
    layer2_outputs(3341) <= not (a xor b);
    layer2_outputs(3342) <= not b;
    layer2_outputs(3343) <= a and b;
    layer2_outputs(3344) <= a;
    layer2_outputs(3345) <= not (a xor b);
    layer2_outputs(3346) <= not a;
    layer2_outputs(3347) <= a;
    layer2_outputs(3348) <= '0';
    layer2_outputs(3349) <= b;
    layer2_outputs(3350) <= not a;
    layer2_outputs(3351) <= b;
    layer2_outputs(3352) <= a and not b;
    layer2_outputs(3353) <= a and b;
    layer2_outputs(3354) <= a;
    layer2_outputs(3355) <= not a or b;
    layer2_outputs(3356) <= '0';
    layer2_outputs(3357) <= a;
    layer2_outputs(3358) <= not b;
    layer2_outputs(3359) <= not (a and b);
    layer2_outputs(3360) <= a and b;
    layer2_outputs(3361) <= b;
    layer2_outputs(3362) <= not a;
    layer2_outputs(3363) <= a xor b;
    layer2_outputs(3364) <= not (a xor b);
    layer2_outputs(3365) <= not (a and b);
    layer2_outputs(3366) <= '0';
    layer2_outputs(3367) <= not b;
    layer2_outputs(3368) <= '1';
    layer2_outputs(3369) <= not (a or b);
    layer2_outputs(3370) <= not (a or b);
    layer2_outputs(3371) <= b and not a;
    layer2_outputs(3372) <= '0';
    layer2_outputs(3373) <= not a or b;
    layer2_outputs(3374) <= a and b;
    layer2_outputs(3375) <= a;
    layer2_outputs(3376) <= not a or b;
    layer2_outputs(3377) <= a or b;
    layer2_outputs(3378) <= a;
    layer2_outputs(3379) <= b and not a;
    layer2_outputs(3380) <= a and not b;
    layer2_outputs(3381) <= not a;
    layer2_outputs(3382) <= not (a or b);
    layer2_outputs(3383) <= not b or a;
    layer2_outputs(3384) <= '1';
    layer2_outputs(3385) <= not (a or b);
    layer2_outputs(3386) <= b and not a;
    layer2_outputs(3387) <= a and b;
    layer2_outputs(3388) <= a and not b;
    layer2_outputs(3389) <= a and b;
    layer2_outputs(3390) <= not b;
    layer2_outputs(3391) <= b and not a;
    layer2_outputs(3392) <= not (a and b);
    layer2_outputs(3393) <= a or b;
    layer2_outputs(3394) <= b and not a;
    layer2_outputs(3395) <= b and not a;
    layer2_outputs(3396) <= a;
    layer2_outputs(3397) <= a xor b;
    layer2_outputs(3398) <= b and not a;
    layer2_outputs(3399) <= not a;
    layer2_outputs(3400) <= not b;
    layer2_outputs(3401) <= not a;
    layer2_outputs(3402) <= not (a or b);
    layer2_outputs(3403) <= not (a and b);
    layer2_outputs(3404) <= a;
    layer2_outputs(3405) <= a;
    layer2_outputs(3406) <= b and not a;
    layer2_outputs(3407) <= not a;
    layer2_outputs(3408) <= not b;
    layer2_outputs(3409) <= not (a and b);
    layer2_outputs(3410) <= b;
    layer2_outputs(3411) <= not b or a;
    layer2_outputs(3412) <= not b;
    layer2_outputs(3413) <= b;
    layer2_outputs(3414) <= b;
    layer2_outputs(3415) <= not (a xor b);
    layer2_outputs(3416) <= a and not b;
    layer2_outputs(3417) <= not b or a;
    layer2_outputs(3418) <= not b or a;
    layer2_outputs(3419) <= a xor b;
    layer2_outputs(3420) <= a or b;
    layer2_outputs(3421) <= not (a and b);
    layer2_outputs(3422) <= '0';
    layer2_outputs(3423) <= a or b;
    layer2_outputs(3424) <= b;
    layer2_outputs(3425) <= not b;
    layer2_outputs(3426) <= not (a xor b);
    layer2_outputs(3427) <= not b;
    layer2_outputs(3428) <= not b;
    layer2_outputs(3429) <= not a or b;
    layer2_outputs(3430) <= not b;
    layer2_outputs(3431) <= a;
    layer2_outputs(3432) <= not (a and b);
    layer2_outputs(3433) <= not (a or b);
    layer2_outputs(3434) <= not b;
    layer2_outputs(3435) <= b;
    layer2_outputs(3436) <= b;
    layer2_outputs(3437) <= a or b;
    layer2_outputs(3438) <= b and not a;
    layer2_outputs(3439) <= '0';
    layer2_outputs(3440) <= b;
    layer2_outputs(3441) <= '0';
    layer2_outputs(3442) <= a or b;
    layer2_outputs(3443) <= a;
    layer2_outputs(3444) <= '1';
    layer2_outputs(3445) <= not (a or b);
    layer2_outputs(3446) <= a and not b;
    layer2_outputs(3447) <= a and b;
    layer2_outputs(3448) <= a and b;
    layer2_outputs(3449) <= '1';
    layer2_outputs(3450) <= a and b;
    layer2_outputs(3451) <= a and not b;
    layer2_outputs(3452) <= a and not b;
    layer2_outputs(3453) <= not a or b;
    layer2_outputs(3454) <= not b or a;
    layer2_outputs(3455) <= not (a and b);
    layer2_outputs(3456) <= not (a and b);
    layer2_outputs(3457) <= a or b;
    layer2_outputs(3458) <= not b;
    layer2_outputs(3459) <= '0';
    layer2_outputs(3460) <= a;
    layer2_outputs(3461) <= not (a and b);
    layer2_outputs(3462) <= not b;
    layer2_outputs(3463) <= not b;
    layer2_outputs(3464) <= '1';
    layer2_outputs(3465) <= b;
    layer2_outputs(3466) <= not (a or b);
    layer2_outputs(3467) <= not b;
    layer2_outputs(3468) <= not b;
    layer2_outputs(3469) <= not (a and b);
    layer2_outputs(3470) <= not (a and b);
    layer2_outputs(3471) <= not (a xor b);
    layer2_outputs(3472) <= a and not b;
    layer2_outputs(3473) <= '0';
    layer2_outputs(3474) <= not b;
    layer2_outputs(3475) <= not (a and b);
    layer2_outputs(3476) <= a and b;
    layer2_outputs(3477) <= not a;
    layer2_outputs(3478) <= not a or b;
    layer2_outputs(3479) <= a and not b;
    layer2_outputs(3480) <= not b;
    layer2_outputs(3481) <= b;
    layer2_outputs(3482) <= '0';
    layer2_outputs(3483) <= not a or b;
    layer2_outputs(3484) <= a and not b;
    layer2_outputs(3485) <= b and not a;
    layer2_outputs(3486) <= not b or a;
    layer2_outputs(3487) <= '1';
    layer2_outputs(3488) <= not a;
    layer2_outputs(3489) <= not (a and b);
    layer2_outputs(3490) <= a;
    layer2_outputs(3491) <= a xor b;
    layer2_outputs(3492) <= a xor b;
    layer2_outputs(3493) <= '0';
    layer2_outputs(3494) <= a;
    layer2_outputs(3495) <= not b or a;
    layer2_outputs(3496) <= a and not b;
    layer2_outputs(3497) <= a;
    layer2_outputs(3498) <= a xor b;
    layer2_outputs(3499) <= not (a and b);
    layer2_outputs(3500) <= not (a and b);
    layer2_outputs(3501) <= a;
    layer2_outputs(3502) <= not b;
    layer2_outputs(3503) <= b and not a;
    layer2_outputs(3504) <= not b;
    layer2_outputs(3505) <= a xor b;
    layer2_outputs(3506) <= not b;
    layer2_outputs(3507) <= not (a and b);
    layer2_outputs(3508) <= not b;
    layer2_outputs(3509) <= not (a or b);
    layer2_outputs(3510) <= not b or a;
    layer2_outputs(3511) <= '1';
    layer2_outputs(3512) <= not b;
    layer2_outputs(3513) <= a and not b;
    layer2_outputs(3514) <= b and not a;
    layer2_outputs(3515) <= '0';
    layer2_outputs(3516) <= a and not b;
    layer2_outputs(3517) <= b;
    layer2_outputs(3518) <= a and not b;
    layer2_outputs(3519) <= a;
    layer2_outputs(3520) <= not a;
    layer2_outputs(3521) <= not b;
    layer2_outputs(3522) <= not (a and b);
    layer2_outputs(3523) <= a and b;
    layer2_outputs(3524) <= '0';
    layer2_outputs(3525) <= not a or b;
    layer2_outputs(3526) <= not b or a;
    layer2_outputs(3527) <= b;
    layer2_outputs(3528) <= not (a xor b);
    layer2_outputs(3529) <= not b or a;
    layer2_outputs(3530) <= '0';
    layer2_outputs(3531) <= not a;
    layer2_outputs(3532) <= not (a or b);
    layer2_outputs(3533) <= b and not a;
    layer2_outputs(3534) <= not (a xor b);
    layer2_outputs(3535) <= '0';
    layer2_outputs(3536) <= not (a or b);
    layer2_outputs(3537) <= b;
    layer2_outputs(3538) <= '0';
    layer2_outputs(3539) <= not (a and b);
    layer2_outputs(3540) <= a and not b;
    layer2_outputs(3541) <= not b;
    layer2_outputs(3542) <= not a;
    layer2_outputs(3543) <= a and b;
    layer2_outputs(3544) <= b and not a;
    layer2_outputs(3545) <= not b or a;
    layer2_outputs(3546) <= b;
    layer2_outputs(3547) <= a and b;
    layer2_outputs(3548) <= not a;
    layer2_outputs(3549) <= not (a xor b);
    layer2_outputs(3550) <= b and not a;
    layer2_outputs(3551) <= not a or b;
    layer2_outputs(3552) <= a or b;
    layer2_outputs(3553) <= not a or b;
    layer2_outputs(3554) <= a or b;
    layer2_outputs(3555) <= '0';
    layer2_outputs(3556) <= a and not b;
    layer2_outputs(3557) <= not a;
    layer2_outputs(3558) <= not b or a;
    layer2_outputs(3559) <= a and not b;
    layer2_outputs(3560) <= not b;
    layer2_outputs(3561) <= a and not b;
    layer2_outputs(3562) <= b and not a;
    layer2_outputs(3563) <= a and not b;
    layer2_outputs(3564) <= a xor b;
    layer2_outputs(3565) <= a;
    layer2_outputs(3566) <= a and b;
    layer2_outputs(3567) <= a;
    layer2_outputs(3568) <= not (a and b);
    layer2_outputs(3569) <= a or b;
    layer2_outputs(3570) <= not b or a;
    layer2_outputs(3571) <= not (a and b);
    layer2_outputs(3572) <= not a;
    layer2_outputs(3573) <= '1';
    layer2_outputs(3574) <= b and not a;
    layer2_outputs(3575) <= not b;
    layer2_outputs(3576) <= not a;
    layer2_outputs(3577) <= '1';
    layer2_outputs(3578) <= not a;
    layer2_outputs(3579) <= a or b;
    layer2_outputs(3580) <= not (a or b);
    layer2_outputs(3581) <= a;
    layer2_outputs(3582) <= b and not a;
    layer2_outputs(3583) <= b and not a;
    layer2_outputs(3584) <= b and not a;
    layer2_outputs(3585) <= a and b;
    layer2_outputs(3586) <= not b;
    layer2_outputs(3587) <= b and not a;
    layer2_outputs(3588) <= not b or a;
    layer2_outputs(3589) <= not (a and b);
    layer2_outputs(3590) <= b;
    layer2_outputs(3591) <= not (a or b);
    layer2_outputs(3592) <= not (a and b);
    layer2_outputs(3593) <= not (a and b);
    layer2_outputs(3594) <= a xor b;
    layer2_outputs(3595) <= a or b;
    layer2_outputs(3596) <= not a or b;
    layer2_outputs(3597) <= not (a and b);
    layer2_outputs(3598) <= not a;
    layer2_outputs(3599) <= not b or a;
    layer2_outputs(3600) <= not (a or b);
    layer2_outputs(3601) <= not (a and b);
    layer2_outputs(3602) <= a or b;
    layer2_outputs(3603) <= '0';
    layer2_outputs(3604) <= not a or b;
    layer2_outputs(3605) <= not (a or b);
    layer2_outputs(3606) <= b and not a;
    layer2_outputs(3607) <= not a or b;
    layer2_outputs(3608) <= not (a and b);
    layer2_outputs(3609) <= b;
    layer2_outputs(3610) <= not a;
    layer2_outputs(3611) <= b;
    layer2_outputs(3612) <= not a or b;
    layer2_outputs(3613) <= not a;
    layer2_outputs(3614) <= b;
    layer2_outputs(3615) <= not b;
    layer2_outputs(3616) <= '1';
    layer2_outputs(3617) <= a;
    layer2_outputs(3618) <= not a or b;
    layer2_outputs(3619) <= a;
    layer2_outputs(3620) <= not b or a;
    layer2_outputs(3621) <= a or b;
    layer2_outputs(3622) <= '1';
    layer2_outputs(3623) <= not (a xor b);
    layer2_outputs(3624) <= b;
    layer2_outputs(3625) <= a and not b;
    layer2_outputs(3626) <= not a;
    layer2_outputs(3627) <= not (a xor b);
    layer2_outputs(3628) <= not b or a;
    layer2_outputs(3629) <= not b;
    layer2_outputs(3630) <= not b;
    layer2_outputs(3631) <= not a;
    layer2_outputs(3632) <= not (a or b);
    layer2_outputs(3633) <= a;
    layer2_outputs(3634) <= a and not b;
    layer2_outputs(3635) <= not (a or b);
    layer2_outputs(3636) <= '0';
    layer2_outputs(3637) <= not a;
    layer2_outputs(3638) <= not (a or b);
    layer2_outputs(3639) <= b;
    layer2_outputs(3640) <= not b or a;
    layer2_outputs(3641) <= '0';
    layer2_outputs(3642) <= not a;
    layer2_outputs(3643) <= a and not b;
    layer2_outputs(3644) <= a or b;
    layer2_outputs(3645) <= not b;
    layer2_outputs(3646) <= a and b;
    layer2_outputs(3647) <= not (a or b);
    layer2_outputs(3648) <= not a;
    layer2_outputs(3649) <= not b;
    layer2_outputs(3650) <= a or b;
    layer2_outputs(3651) <= not a or b;
    layer2_outputs(3652) <= not (a and b);
    layer2_outputs(3653) <= '1';
    layer2_outputs(3654) <= not b;
    layer2_outputs(3655) <= not a;
    layer2_outputs(3656) <= a;
    layer2_outputs(3657) <= not (a and b);
    layer2_outputs(3658) <= not b;
    layer2_outputs(3659) <= a;
    layer2_outputs(3660) <= '0';
    layer2_outputs(3661) <= not (a xor b);
    layer2_outputs(3662) <= not (a or b);
    layer2_outputs(3663) <= not b or a;
    layer2_outputs(3664) <= not a or b;
    layer2_outputs(3665) <= not a;
    layer2_outputs(3666) <= a xor b;
    layer2_outputs(3667) <= b;
    layer2_outputs(3668) <= a and not b;
    layer2_outputs(3669) <= not (a and b);
    layer2_outputs(3670) <= a and not b;
    layer2_outputs(3671) <= not (a and b);
    layer2_outputs(3672) <= b;
    layer2_outputs(3673) <= b and not a;
    layer2_outputs(3674) <= '0';
    layer2_outputs(3675) <= a;
    layer2_outputs(3676) <= not b;
    layer2_outputs(3677) <= not b;
    layer2_outputs(3678) <= b and not a;
    layer2_outputs(3679) <= not b;
    layer2_outputs(3680) <= not (a or b);
    layer2_outputs(3681) <= not a;
    layer2_outputs(3682) <= not b or a;
    layer2_outputs(3683) <= not a;
    layer2_outputs(3684) <= not (a or b);
    layer2_outputs(3685) <= a;
    layer2_outputs(3686) <= not (a and b);
    layer2_outputs(3687) <= b;
    layer2_outputs(3688) <= a or b;
    layer2_outputs(3689) <= not a or b;
    layer2_outputs(3690) <= '1';
    layer2_outputs(3691) <= not b or a;
    layer2_outputs(3692) <= not a;
    layer2_outputs(3693) <= a or b;
    layer2_outputs(3694) <= not a or b;
    layer2_outputs(3695) <= b;
    layer2_outputs(3696) <= a and not b;
    layer2_outputs(3697) <= not b;
    layer2_outputs(3698) <= b;
    layer2_outputs(3699) <= not a;
    layer2_outputs(3700) <= a and not b;
    layer2_outputs(3701) <= not b;
    layer2_outputs(3702) <= a or b;
    layer2_outputs(3703) <= not a or b;
    layer2_outputs(3704) <= not (a xor b);
    layer2_outputs(3705) <= a or b;
    layer2_outputs(3706) <= b;
    layer2_outputs(3707) <= not b;
    layer2_outputs(3708) <= b and not a;
    layer2_outputs(3709) <= a and not b;
    layer2_outputs(3710) <= not b or a;
    layer2_outputs(3711) <= not a;
    layer2_outputs(3712) <= '1';
    layer2_outputs(3713) <= not b;
    layer2_outputs(3714) <= '1';
    layer2_outputs(3715) <= b;
    layer2_outputs(3716) <= not b;
    layer2_outputs(3717) <= a and not b;
    layer2_outputs(3718) <= not (a and b);
    layer2_outputs(3719) <= '1';
    layer2_outputs(3720) <= a xor b;
    layer2_outputs(3721) <= not (a and b);
    layer2_outputs(3722) <= not b or a;
    layer2_outputs(3723) <= b and not a;
    layer2_outputs(3724) <= not (a xor b);
    layer2_outputs(3725) <= a and not b;
    layer2_outputs(3726) <= not (a and b);
    layer2_outputs(3727) <= not b or a;
    layer2_outputs(3728) <= not b;
    layer2_outputs(3729) <= '0';
    layer2_outputs(3730) <= a;
    layer2_outputs(3731) <= a;
    layer2_outputs(3732) <= a or b;
    layer2_outputs(3733) <= not a;
    layer2_outputs(3734) <= not b or a;
    layer2_outputs(3735) <= b;
    layer2_outputs(3736) <= b and not a;
    layer2_outputs(3737) <= not (a or b);
    layer2_outputs(3738) <= not b or a;
    layer2_outputs(3739) <= not a;
    layer2_outputs(3740) <= '1';
    layer2_outputs(3741) <= '0';
    layer2_outputs(3742) <= not b;
    layer2_outputs(3743) <= '1';
    layer2_outputs(3744) <= not (a or b);
    layer2_outputs(3745) <= a;
    layer2_outputs(3746) <= a and b;
    layer2_outputs(3747) <= not (a or b);
    layer2_outputs(3748) <= not a or b;
    layer2_outputs(3749) <= not a or b;
    layer2_outputs(3750) <= not b;
    layer2_outputs(3751) <= not b;
    layer2_outputs(3752) <= a xor b;
    layer2_outputs(3753) <= not a;
    layer2_outputs(3754) <= a;
    layer2_outputs(3755) <= '1';
    layer2_outputs(3756) <= not (a xor b);
    layer2_outputs(3757) <= not b;
    layer2_outputs(3758) <= a;
    layer2_outputs(3759) <= a and b;
    layer2_outputs(3760) <= a xor b;
    layer2_outputs(3761) <= a and not b;
    layer2_outputs(3762) <= not a or b;
    layer2_outputs(3763) <= a and b;
    layer2_outputs(3764) <= not b;
    layer2_outputs(3765) <= a;
    layer2_outputs(3766) <= b;
    layer2_outputs(3767) <= not (a xor b);
    layer2_outputs(3768) <= b;
    layer2_outputs(3769) <= b and not a;
    layer2_outputs(3770) <= not a;
    layer2_outputs(3771) <= a and b;
    layer2_outputs(3772) <= a or b;
    layer2_outputs(3773) <= not a or b;
    layer2_outputs(3774) <= not (a and b);
    layer2_outputs(3775) <= b;
    layer2_outputs(3776) <= b and not a;
    layer2_outputs(3777) <= '0';
    layer2_outputs(3778) <= a and b;
    layer2_outputs(3779) <= not (a or b);
    layer2_outputs(3780) <= a and b;
    layer2_outputs(3781) <= '1';
    layer2_outputs(3782) <= a;
    layer2_outputs(3783) <= not b or a;
    layer2_outputs(3784) <= a and b;
    layer2_outputs(3785) <= not (a xor b);
    layer2_outputs(3786) <= not b or a;
    layer2_outputs(3787) <= b and not a;
    layer2_outputs(3788) <= a;
    layer2_outputs(3789) <= a;
    layer2_outputs(3790) <= b;
    layer2_outputs(3791) <= a;
    layer2_outputs(3792) <= not (a xor b);
    layer2_outputs(3793) <= a and b;
    layer2_outputs(3794) <= b and not a;
    layer2_outputs(3795) <= b;
    layer2_outputs(3796) <= not (a and b);
    layer2_outputs(3797) <= b and not a;
    layer2_outputs(3798) <= a and not b;
    layer2_outputs(3799) <= '0';
    layer2_outputs(3800) <= a;
    layer2_outputs(3801) <= not (a xor b);
    layer2_outputs(3802) <= not b;
    layer2_outputs(3803) <= not b or a;
    layer2_outputs(3804) <= not (a and b);
    layer2_outputs(3805) <= not (a xor b);
    layer2_outputs(3806) <= a or b;
    layer2_outputs(3807) <= not a;
    layer2_outputs(3808) <= a or b;
    layer2_outputs(3809) <= a or b;
    layer2_outputs(3810) <= not (a and b);
    layer2_outputs(3811) <= not b;
    layer2_outputs(3812) <= a or b;
    layer2_outputs(3813) <= '0';
    layer2_outputs(3814) <= b;
    layer2_outputs(3815) <= a and not b;
    layer2_outputs(3816) <= not (a or b);
    layer2_outputs(3817) <= '1';
    layer2_outputs(3818) <= a and not b;
    layer2_outputs(3819) <= not a or b;
    layer2_outputs(3820) <= a or b;
    layer2_outputs(3821) <= a and not b;
    layer2_outputs(3822) <= a and b;
    layer2_outputs(3823) <= b;
    layer2_outputs(3824) <= not b;
    layer2_outputs(3825) <= a;
    layer2_outputs(3826) <= b;
    layer2_outputs(3827) <= not b or a;
    layer2_outputs(3828) <= not b;
    layer2_outputs(3829) <= a;
    layer2_outputs(3830) <= not b;
    layer2_outputs(3831) <= b;
    layer2_outputs(3832) <= a and not b;
    layer2_outputs(3833) <= b and not a;
    layer2_outputs(3834) <= b and not a;
    layer2_outputs(3835) <= '0';
    layer2_outputs(3836) <= a;
    layer2_outputs(3837) <= '1';
    layer2_outputs(3838) <= a or b;
    layer2_outputs(3839) <= not a;
    layer2_outputs(3840) <= '1';
    layer2_outputs(3841) <= not b;
    layer2_outputs(3842) <= not b;
    layer2_outputs(3843) <= a xor b;
    layer2_outputs(3844) <= a;
    layer2_outputs(3845) <= not b or a;
    layer2_outputs(3846) <= a and not b;
    layer2_outputs(3847) <= not (a and b);
    layer2_outputs(3848) <= a;
    layer2_outputs(3849) <= a and b;
    layer2_outputs(3850) <= b;
    layer2_outputs(3851) <= not a;
    layer2_outputs(3852) <= not a or b;
    layer2_outputs(3853) <= a;
    layer2_outputs(3854) <= a and b;
    layer2_outputs(3855) <= not (a xor b);
    layer2_outputs(3856) <= a or b;
    layer2_outputs(3857) <= b and not a;
    layer2_outputs(3858) <= not a;
    layer2_outputs(3859) <= b and not a;
    layer2_outputs(3860) <= a;
    layer2_outputs(3861) <= '1';
    layer2_outputs(3862) <= not a;
    layer2_outputs(3863) <= a or b;
    layer2_outputs(3864) <= not (a xor b);
    layer2_outputs(3865) <= b;
    layer2_outputs(3866) <= a or b;
    layer2_outputs(3867) <= not b;
    layer2_outputs(3868) <= '0';
    layer2_outputs(3869) <= '1';
    layer2_outputs(3870) <= not b;
    layer2_outputs(3871) <= a and not b;
    layer2_outputs(3872) <= a and not b;
    layer2_outputs(3873) <= not b;
    layer2_outputs(3874) <= '0';
    layer2_outputs(3875) <= a and b;
    layer2_outputs(3876) <= not a or b;
    layer2_outputs(3877) <= a;
    layer2_outputs(3878) <= not (a or b);
    layer2_outputs(3879) <= '0';
    layer2_outputs(3880) <= b and not a;
    layer2_outputs(3881) <= a xor b;
    layer2_outputs(3882) <= a;
    layer2_outputs(3883) <= a and not b;
    layer2_outputs(3884) <= b;
    layer2_outputs(3885) <= a and not b;
    layer2_outputs(3886) <= a and b;
    layer2_outputs(3887) <= a or b;
    layer2_outputs(3888) <= not (a xor b);
    layer2_outputs(3889) <= a xor b;
    layer2_outputs(3890) <= a and b;
    layer2_outputs(3891) <= a and not b;
    layer2_outputs(3892) <= b and not a;
    layer2_outputs(3893) <= a xor b;
    layer2_outputs(3894) <= not (a xor b);
    layer2_outputs(3895) <= '0';
    layer2_outputs(3896) <= a or b;
    layer2_outputs(3897) <= not b;
    layer2_outputs(3898) <= not (a or b);
    layer2_outputs(3899) <= a;
    layer2_outputs(3900) <= not a or b;
    layer2_outputs(3901) <= a and b;
    layer2_outputs(3902) <= not a or b;
    layer2_outputs(3903) <= a and not b;
    layer2_outputs(3904) <= '0';
    layer2_outputs(3905) <= a and b;
    layer2_outputs(3906) <= not a;
    layer2_outputs(3907) <= not b or a;
    layer2_outputs(3908) <= not b;
    layer2_outputs(3909) <= a and b;
    layer2_outputs(3910) <= not b or a;
    layer2_outputs(3911) <= not a;
    layer2_outputs(3912) <= not a or b;
    layer2_outputs(3913) <= not a or b;
    layer2_outputs(3914) <= not (a or b);
    layer2_outputs(3915) <= not b;
    layer2_outputs(3916) <= '1';
    layer2_outputs(3917) <= not a or b;
    layer2_outputs(3918) <= a;
    layer2_outputs(3919) <= not b;
    layer2_outputs(3920) <= a;
    layer2_outputs(3921) <= not b;
    layer2_outputs(3922) <= not a or b;
    layer2_outputs(3923) <= not b or a;
    layer2_outputs(3924) <= b;
    layer2_outputs(3925) <= not a;
    layer2_outputs(3926) <= a and b;
    layer2_outputs(3927) <= b and not a;
    layer2_outputs(3928) <= a and b;
    layer2_outputs(3929) <= not (a and b);
    layer2_outputs(3930) <= b and not a;
    layer2_outputs(3931) <= b;
    layer2_outputs(3932) <= not (a or b);
    layer2_outputs(3933) <= not (a and b);
    layer2_outputs(3934) <= b;
    layer2_outputs(3935) <= not a;
    layer2_outputs(3936) <= not (a or b);
    layer2_outputs(3937) <= not b;
    layer2_outputs(3938) <= not (a or b);
    layer2_outputs(3939) <= a;
    layer2_outputs(3940) <= not (a and b);
    layer2_outputs(3941) <= not b or a;
    layer2_outputs(3942) <= not b or a;
    layer2_outputs(3943) <= not (a xor b);
    layer2_outputs(3944) <= not a;
    layer2_outputs(3945) <= not b or a;
    layer2_outputs(3946) <= a and not b;
    layer2_outputs(3947) <= not a or b;
    layer2_outputs(3948) <= a and not b;
    layer2_outputs(3949) <= a;
    layer2_outputs(3950) <= a and b;
    layer2_outputs(3951) <= not b;
    layer2_outputs(3952) <= not a;
    layer2_outputs(3953) <= not a;
    layer2_outputs(3954) <= not (a or b);
    layer2_outputs(3955) <= '1';
    layer2_outputs(3956) <= a;
    layer2_outputs(3957) <= b and not a;
    layer2_outputs(3958) <= not a;
    layer2_outputs(3959) <= a;
    layer2_outputs(3960) <= '0';
    layer2_outputs(3961) <= a and b;
    layer2_outputs(3962) <= not (a or b);
    layer2_outputs(3963) <= b;
    layer2_outputs(3964) <= '1';
    layer2_outputs(3965) <= '0';
    layer2_outputs(3966) <= a;
    layer2_outputs(3967) <= b;
    layer2_outputs(3968) <= b and not a;
    layer2_outputs(3969) <= not b;
    layer2_outputs(3970) <= a and b;
    layer2_outputs(3971) <= a and not b;
    layer2_outputs(3972) <= not a or b;
    layer2_outputs(3973) <= not (a and b);
    layer2_outputs(3974) <= b;
    layer2_outputs(3975) <= a and b;
    layer2_outputs(3976) <= not a;
    layer2_outputs(3977) <= a and b;
    layer2_outputs(3978) <= not (a or b);
    layer2_outputs(3979) <= a or b;
    layer2_outputs(3980) <= a;
    layer2_outputs(3981) <= not b or a;
    layer2_outputs(3982) <= a or b;
    layer2_outputs(3983) <= b and not a;
    layer2_outputs(3984) <= not (a and b);
    layer2_outputs(3985) <= '0';
    layer2_outputs(3986) <= not (a and b);
    layer2_outputs(3987) <= a;
    layer2_outputs(3988) <= not b;
    layer2_outputs(3989) <= not (a and b);
    layer2_outputs(3990) <= '0';
    layer2_outputs(3991) <= '1';
    layer2_outputs(3992) <= a and not b;
    layer2_outputs(3993) <= not (a xor b);
    layer2_outputs(3994) <= not a or b;
    layer2_outputs(3995) <= not b or a;
    layer2_outputs(3996) <= '0';
    layer2_outputs(3997) <= b and not a;
    layer2_outputs(3998) <= a or b;
    layer2_outputs(3999) <= not b or a;
    layer2_outputs(4000) <= a;
    layer2_outputs(4001) <= a and not b;
    layer2_outputs(4002) <= not (a or b);
    layer2_outputs(4003) <= a and b;
    layer2_outputs(4004) <= not (a or b);
    layer2_outputs(4005) <= a;
    layer2_outputs(4006) <= not a;
    layer2_outputs(4007) <= '0';
    layer2_outputs(4008) <= a and b;
    layer2_outputs(4009) <= '0';
    layer2_outputs(4010) <= a;
    layer2_outputs(4011) <= '1';
    layer2_outputs(4012) <= not a or b;
    layer2_outputs(4013) <= not b or a;
    layer2_outputs(4014) <= a;
    layer2_outputs(4015) <= b and not a;
    layer2_outputs(4016) <= not (a xor b);
    layer2_outputs(4017) <= b and not a;
    layer2_outputs(4018) <= not (a or b);
    layer2_outputs(4019) <= not a;
    layer2_outputs(4020) <= '0';
    layer2_outputs(4021) <= a or b;
    layer2_outputs(4022) <= a xor b;
    layer2_outputs(4023) <= a xor b;
    layer2_outputs(4024) <= a;
    layer2_outputs(4025) <= not (a or b);
    layer2_outputs(4026) <= a or b;
    layer2_outputs(4027) <= b;
    layer2_outputs(4028) <= not (a xor b);
    layer2_outputs(4029) <= a xor b;
    layer2_outputs(4030) <= not a or b;
    layer2_outputs(4031) <= a or b;
    layer2_outputs(4032) <= a and not b;
    layer2_outputs(4033) <= a;
    layer2_outputs(4034) <= not b or a;
    layer2_outputs(4035) <= not (a or b);
    layer2_outputs(4036) <= a and not b;
    layer2_outputs(4037) <= not (a or b);
    layer2_outputs(4038) <= a;
    layer2_outputs(4039) <= '0';
    layer2_outputs(4040) <= '1';
    layer2_outputs(4041) <= not (a and b);
    layer2_outputs(4042) <= b and not a;
    layer2_outputs(4043) <= not (a or b);
    layer2_outputs(4044) <= not b;
    layer2_outputs(4045) <= not a or b;
    layer2_outputs(4046) <= a xor b;
    layer2_outputs(4047) <= a and b;
    layer2_outputs(4048) <= not (a and b);
    layer2_outputs(4049) <= not b;
    layer2_outputs(4050) <= not (a or b);
    layer2_outputs(4051) <= a;
    layer2_outputs(4052) <= not (a and b);
    layer2_outputs(4053) <= a or b;
    layer2_outputs(4054) <= not a;
    layer2_outputs(4055) <= not (a and b);
    layer2_outputs(4056) <= a;
    layer2_outputs(4057) <= a or b;
    layer2_outputs(4058) <= a and b;
    layer2_outputs(4059) <= b;
    layer2_outputs(4060) <= not a;
    layer2_outputs(4061) <= not b;
    layer2_outputs(4062) <= not (a and b);
    layer2_outputs(4063) <= a and not b;
    layer2_outputs(4064) <= '0';
    layer2_outputs(4065) <= b and not a;
    layer2_outputs(4066) <= not a or b;
    layer2_outputs(4067) <= not a;
    layer2_outputs(4068) <= not (a xor b);
    layer2_outputs(4069) <= a or b;
    layer2_outputs(4070) <= a xor b;
    layer2_outputs(4071) <= not (a or b);
    layer2_outputs(4072) <= '0';
    layer2_outputs(4073) <= a;
    layer2_outputs(4074) <= a and not b;
    layer2_outputs(4075) <= a and not b;
    layer2_outputs(4076) <= a;
    layer2_outputs(4077) <= not b;
    layer2_outputs(4078) <= not a;
    layer2_outputs(4079) <= a or b;
    layer2_outputs(4080) <= '1';
    layer2_outputs(4081) <= a and not b;
    layer2_outputs(4082) <= a and not b;
    layer2_outputs(4083) <= b;
    layer2_outputs(4084) <= b and not a;
    layer2_outputs(4085) <= not a;
    layer2_outputs(4086) <= not a;
    layer2_outputs(4087) <= '0';
    layer2_outputs(4088) <= not (a xor b);
    layer2_outputs(4089) <= '0';
    layer2_outputs(4090) <= not (a and b);
    layer2_outputs(4091) <= not b or a;
    layer2_outputs(4092) <= not a or b;
    layer2_outputs(4093) <= a or b;
    layer2_outputs(4094) <= b;
    layer2_outputs(4095) <= a or b;
    layer2_outputs(4096) <= a and not b;
    layer2_outputs(4097) <= '1';
    layer2_outputs(4098) <= not a;
    layer2_outputs(4099) <= not (a and b);
    layer2_outputs(4100) <= not a or b;
    layer2_outputs(4101) <= not (a or b);
    layer2_outputs(4102) <= '1';
    layer2_outputs(4103) <= a and not b;
    layer2_outputs(4104) <= not b;
    layer2_outputs(4105) <= not a;
    layer2_outputs(4106) <= not (a or b);
    layer2_outputs(4107) <= a;
    layer2_outputs(4108) <= a;
    layer2_outputs(4109) <= not (a and b);
    layer2_outputs(4110) <= a or b;
    layer2_outputs(4111) <= a and b;
    layer2_outputs(4112) <= not b;
    layer2_outputs(4113) <= a;
    layer2_outputs(4114) <= a and b;
    layer2_outputs(4115) <= not a;
    layer2_outputs(4116) <= a xor b;
    layer2_outputs(4117) <= not (a xor b);
    layer2_outputs(4118) <= b and not a;
    layer2_outputs(4119) <= a xor b;
    layer2_outputs(4120) <= a and b;
    layer2_outputs(4121) <= not a;
    layer2_outputs(4122) <= '1';
    layer2_outputs(4123) <= a;
    layer2_outputs(4124) <= '1';
    layer2_outputs(4125) <= not b;
    layer2_outputs(4126) <= not (a and b);
    layer2_outputs(4127) <= not a;
    layer2_outputs(4128) <= a;
    layer2_outputs(4129) <= not (a or b);
    layer2_outputs(4130) <= '0';
    layer2_outputs(4131) <= not (a or b);
    layer2_outputs(4132) <= a;
    layer2_outputs(4133) <= not (a or b);
    layer2_outputs(4134) <= not (a xor b);
    layer2_outputs(4135) <= not a;
    layer2_outputs(4136) <= a and not b;
    layer2_outputs(4137) <= b;
    layer2_outputs(4138) <= not b;
    layer2_outputs(4139) <= a and not b;
    layer2_outputs(4140) <= not a or b;
    layer2_outputs(4141) <= b and not a;
    layer2_outputs(4142) <= a;
    layer2_outputs(4143) <= b;
    layer2_outputs(4144) <= not (a xor b);
    layer2_outputs(4145) <= '0';
    layer2_outputs(4146) <= b and not a;
    layer2_outputs(4147) <= a or b;
    layer2_outputs(4148) <= a;
    layer2_outputs(4149) <= '0';
    layer2_outputs(4150) <= a;
    layer2_outputs(4151) <= a;
    layer2_outputs(4152) <= not a or b;
    layer2_outputs(4153) <= '0';
    layer2_outputs(4154) <= not b or a;
    layer2_outputs(4155) <= '1';
    layer2_outputs(4156) <= not (a and b);
    layer2_outputs(4157) <= b and not a;
    layer2_outputs(4158) <= not b or a;
    layer2_outputs(4159) <= a and not b;
    layer2_outputs(4160) <= not (a or b);
    layer2_outputs(4161) <= b and not a;
    layer2_outputs(4162) <= not (a and b);
    layer2_outputs(4163) <= a xor b;
    layer2_outputs(4164) <= not b;
    layer2_outputs(4165) <= a;
    layer2_outputs(4166) <= b and not a;
    layer2_outputs(4167) <= not b;
    layer2_outputs(4168) <= a and not b;
    layer2_outputs(4169) <= not b or a;
    layer2_outputs(4170) <= a and b;
    layer2_outputs(4171) <= not a;
    layer2_outputs(4172) <= not b;
    layer2_outputs(4173) <= a and b;
    layer2_outputs(4174) <= b;
    layer2_outputs(4175) <= not a or b;
    layer2_outputs(4176) <= not a or b;
    layer2_outputs(4177) <= not b or a;
    layer2_outputs(4178) <= a and not b;
    layer2_outputs(4179) <= not b or a;
    layer2_outputs(4180) <= a;
    layer2_outputs(4181) <= b;
    layer2_outputs(4182) <= b;
    layer2_outputs(4183) <= b and not a;
    layer2_outputs(4184) <= a xor b;
    layer2_outputs(4185) <= a;
    layer2_outputs(4186) <= a and b;
    layer2_outputs(4187) <= '0';
    layer2_outputs(4188) <= not a or b;
    layer2_outputs(4189) <= not b;
    layer2_outputs(4190) <= not b;
    layer2_outputs(4191) <= a and not b;
    layer2_outputs(4192) <= a and not b;
    layer2_outputs(4193) <= not (a and b);
    layer2_outputs(4194) <= not (a or b);
    layer2_outputs(4195) <= not (a or b);
    layer2_outputs(4196) <= b and not a;
    layer2_outputs(4197) <= not b;
    layer2_outputs(4198) <= a;
    layer2_outputs(4199) <= a or b;
    layer2_outputs(4200) <= not a or b;
    layer2_outputs(4201) <= not a;
    layer2_outputs(4202) <= a and b;
    layer2_outputs(4203) <= a;
    layer2_outputs(4204) <= not a;
    layer2_outputs(4205) <= not a or b;
    layer2_outputs(4206) <= b and not a;
    layer2_outputs(4207) <= a and b;
    layer2_outputs(4208) <= not (a and b);
    layer2_outputs(4209) <= a and b;
    layer2_outputs(4210) <= not b or a;
    layer2_outputs(4211) <= not a;
    layer2_outputs(4212) <= not (a xor b);
    layer2_outputs(4213) <= b and not a;
    layer2_outputs(4214) <= '0';
    layer2_outputs(4215) <= b;
    layer2_outputs(4216) <= b and not a;
    layer2_outputs(4217) <= a xor b;
    layer2_outputs(4218) <= b;
    layer2_outputs(4219) <= not (a and b);
    layer2_outputs(4220) <= a;
    layer2_outputs(4221) <= not b;
    layer2_outputs(4222) <= b and not a;
    layer2_outputs(4223) <= not a or b;
    layer2_outputs(4224) <= not a;
    layer2_outputs(4225) <= a and not b;
    layer2_outputs(4226) <= a or b;
    layer2_outputs(4227) <= a and not b;
    layer2_outputs(4228) <= '1';
    layer2_outputs(4229) <= not (a and b);
    layer2_outputs(4230) <= a and b;
    layer2_outputs(4231) <= '0';
    layer2_outputs(4232) <= not a;
    layer2_outputs(4233) <= a and not b;
    layer2_outputs(4234) <= a and b;
    layer2_outputs(4235) <= not b;
    layer2_outputs(4236) <= a;
    layer2_outputs(4237) <= a and b;
    layer2_outputs(4238) <= a or b;
    layer2_outputs(4239) <= b and not a;
    layer2_outputs(4240) <= not b or a;
    layer2_outputs(4241) <= b;
    layer2_outputs(4242) <= not b;
    layer2_outputs(4243) <= b and not a;
    layer2_outputs(4244) <= '1';
    layer2_outputs(4245) <= not (a or b);
    layer2_outputs(4246) <= not (a and b);
    layer2_outputs(4247) <= not (a and b);
    layer2_outputs(4248) <= not (a or b);
    layer2_outputs(4249) <= b;
    layer2_outputs(4250) <= not a or b;
    layer2_outputs(4251) <= not a or b;
    layer2_outputs(4252) <= a and b;
    layer2_outputs(4253) <= not b;
    layer2_outputs(4254) <= b and not a;
    layer2_outputs(4255) <= '1';
    layer2_outputs(4256) <= not b;
    layer2_outputs(4257) <= b and not a;
    layer2_outputs(4258) <= not b or a;
    layer2_outputs(4259) <= not (a and b);
    layer2_outputs(4260) <= '1';
    layer2_outputs(4261) <= not a;
    layer2_outputs(4262) <= a;
    layer2_outputs(4263) <= '0';
    layer2_outputs(4264) <= '1';
    layer2_outputs(4265) <= not (a and b);
    layer2_outputs(4266) <= not a;
    layer2_outputs(4267) <= a and b;
    layer2_outputs(4268) <= '1';
    layer2_outputs(4269) <= b;
    layer2_outputs(4270) <= not a or b;
    layer2_outputs(4271) <= not a;
    layer2_outputs(4272) <= not a or b;
    layer2_outputs(4273) <= b;
    layer2_outputs(4274) <= a and not b;
    layer2_outputs(4275) <= a;
    layer2_outputs(4276) <= a or b;
    layer2_outputs(4277) <= a or b;
    layer2_outputs(4278) <= '1';
    layer2_outputs(4279) <= '0';
    layer2_outputs(4280) <= b;
    layer2_outputs(4281) <= '1';
    layer2_outputs(4282) <= not a;
    layer2_outputs(4283) <= not (a or b);
    layer2_outputs(4284) <= a and not b;
    layer2_outputs(4285) <= not a;
    layer2_outputs(4286) <= not a;
    layer2_outputs(4287) <= b and not a;
    layer2_outputs(4288) <= b and not a;
    layer2_outputs(4289) <= not a or b;
    layer2_outputs(4290) <= not (a and b);
    layer2_outputs(4291) <= b;
    layer2_outputs(4292) <= not b or a;
    layer2_outputs(4293) <= '0';
    layer2_outputs(4294) <= a or b;
    layer2_outputs(4295) <= a and not b;
    layer2_outputs(4296) <= b and not a;
    layer2_outputs(4297) <= a;
    layer2_outputs(4298) <= not a;
    layer2_outputs(4299) <= a and b;
    layer2_outputs(4300) <= '1';
    layer2_outputs(4301) <= a or b;
    layer2_outputs(4302) <= b;
    layer2_outputs(4303) <= b;
    layer2_outputs(4304) <= not (a and b);
    layer2_outputs(4305) <= '1';
    layer2_outputs(4306) <= not a or b;
    layer2_outputs(4307) <= b;
    layer2_outputs(4308) <= not a;
    layer2_outputs(4309) <= a;
    layer2_outputs(4310) <= not b;
    layer2_outputs(4311) <= '1';
    layer2_outputs(4312) <= a or b;
    layer2_outputs(4313) <= not b or a;
    layer2_outputs(4314) <= a or b;
    layer2_outputs(4315) <= a and b;
    layer2_outputs(4316) <= '0';
    layer2_outputs(4317) <= a or b;
    layer2_outputs(4318) <= not b;
    layer2_outputs(4319) <= not (a and b);
    layer2_outputs(4320) <= not a or b;
    layer2_outputs(4321) <= not (a xor b);
    layer2_outputs(4322) <= a and b;
    layer2_outputs(4323) <= '1';
    layer2_outputs(4324) <= a or b;
    layer2_outputs(4325) <= a or b;
    layer2_outputs(4326) <= not b;
    layer2_outputs(4327) <= a and not b;
    layer2_outputs(4328) <= a and b;
    layer2_outputs(4329) <= not a;
    layer2_outputs(4330) <= not (a or b);
    layer2_outputs(4331) <= not (a xor b);
    layer2_outputs(4332) <= '0';
    layer2_outputs(4333) <= not b;
    layer2_outputs(4334) <= not (a or b);
    layer2_outputs(4335) <= b and not a;
    layer2_outputs(4336) <= not (a xor b);
    layer2_outputs(4337) <= b;
    layer2_outputs(4338) <= b and not a;
    layer2_outputs(4339) <= '1';
    layer2_outputs(4340) <= not a;
    layer2_outputs(4341) <= a or b;
    layer2_outputs(4342) <= a and b;
    layer2_outputs(4343) <= a and not b;
    layer2_outputs(4344) <= not a;
    layer2_outputs(4345) <= a;
    layer2_outputs(4346) <= not (a or b);
    layer2_outputs(4347) <= not (a and b);
    layer2_outputs(4348) <= a and not b;
    layer2_outputs(4349) <= a or b;
    layer2_outputs(4350) <= a or b;
    layer2_outputs(4351) <= not b or a;
    layer2_outputs(4352) <= not a or b;
    layer2_outputs(4353) <= b and not a;
    layer2_outputs(4354) <= a;
    layer2_outputs(4355) <= '1';
    layer2_outputs(4356) <= a;
    layer2_outputs(4357) <= not (a and b);
    layer2_outputs(4358) <= '1';
    layer2_outputs(4359) <= not b;
    layer2_outputs(4360) <= b;
    layer2_outputs(4361) <= b;
    layer2_outputs(4362) <= not (a or b);
    layer2_outputs(4363) <= b and not a;
    layer2_outputs(4364) <= not b or a;
    layer2_outputs(4365) <= not b;
    layer2_outputs(4366) <= not b or a;
    layer2_outputs(4367) <= '0';
    layer2_outputs(4368) <= b and not a;
    layer2_outputs(4369) <= a;
    layer2_outputs(4370) <= not a;
    layer2_outputs(4371) <= not a;
    layer2_outputs(4372) <= a;
    layer2_outputs(4373) <= a and b;
    layer2_outputs(4374) <= not a or b;
    layer2_outputs(4375) <= not a or b;
    layer2_outputs(4376) <= b and not a;
    layer2_outputs(4377) <= not (a or b);
    layer2_outputs(4378) <= not b;
    layer2_outputs(4379) <= a;
    layer2_outputs(4380) <= a and b;
    layer2_outputs(4381) <= b;
    layer2_outputs(4382) <= not a;
    layer2_outputs(4383) <= '1';
    layer2_outputs(4384) <= not (a or b);
    layer2_outputs(4385) <= a;
    layer2_outputs(4386) <= '0';
    layer2_outputs(4387) <= a and not b;
    layer2_outputs(4388) <= not b;
    layer2_outputs(4389) <= not b;
    layer2_outputs(4390) <= not a;
    layer2_outputs(4391) <= not a or b;
    layer2_outputs(4392) <= a and not b;
    layer2_outputs(4393) <= b and not a;
    layer2_outputs(4394) <= not b;
    layer2_outputs(4395) <= not (a and b);
    layer2_outputs(4396) <= not (a or b);
    layer2_outputs(4397) <= a and b;
    layer2_outputs(4398) <= a;
    layer2_outputs(4399) <= not (a or b);
    layer2_outputs(4400) <= not a;
    layer2_outputs(4401) <= b;
    layer2_outputs(4402) <= a and b;
    layer2_outputs(4403) <= b and not a;
    layer2_outputs(4404) <= not (a or b);
    layer2_outputs(4405) <= not b;
    layer2_outputs(4406) <= not a or b;
    layer2_outputs(4407) <= a and b;
    layer2_outputs(4408) <= a;
    layer2_outputs(4409) <= b;
    layer2_outputs(4410) <= a or b;
    layer2_outputs(4411) <= '0';
    layer2_outputs(4412) <= '1';
    layer2_outputs(4413) <= a and b;
    layer2_outputs(4414) <= b;
    layer2_outputs(4415) <= b;
    layer2_outputs(4416) <= a and not b;
    layer2_outputs(4417) <= b;
    layer2_outputs(4418) <= '1';
    layer2_outputs(4419) <= not a;
    layer2_outputs(4420) <= b and not a;
    layer2_outputs(4421) <= not (a or b);
    layer2_outputs(4422) <= not a or b;
    layer2_outputs(4423) <= a and b;
    layer2_outputs(4424) <= '0';
    layer2_outputs(4425) <= a xor b;
    layer2_outputs(4426) <= b;
    layer2_outputs(4427) <= a or b;
    layer2_outputs(4428) <= '0';
    layer2_outputs(4429) <= a;
    layer2_outputs(4430) <= '1';
    layer2_outputs(4431) <= not a;
    layer2_outputs(4432) <= a xor b;
    layer2_outputs(4433) <= b;
    layer2_outputs(4434) <= b;
    layer2_outputs(4435) <= a or b;
    layer2_outputs(4436) <= b;
    layer2_outputs(4437) <= a;
    layer2_outputs(4438) <= b;
    layer2_outputs(4439) <= not (a and b);
    layer2_outputs(4440) <= not a;
    layer2_outputs(4441) <= not (a or b);
    layer2_outputs(4442) <= '0';
    layer2_outputs(4443) <= b;
    layer2_outputs(4444) <= not a or b;
    layer2_outputs(4445) <= not (a xor b);
    layer2_outputs(4446) <= '1';
    layer2_outputs(4447) <= not (a and b);
    layer2_outputs(4448) <= b;
    layer2_outputs(4449) <= not a;
    layer2_outputs(4450) <= a;
    layer2_outputs(4451) <= not b or a;
    layer2_outputs(4452) <= not (a xor b);
    layer2_outputs(4453) <= not b;
    layer2_outputs(4454) <= a and b;
    layer2_outputs(4455) <= not (a and b);
    layer2_outputs(4456) <= a and not b;
    layer2_outputs(4457) <= a and not b;
    layer2_outputs(4458) <= a and not b;
    layer2_outputs(4459) <= not (a or b);
    layer2_outputs(4460) <= not a or b;
    layer2_outputs(4461) <= a and not b;
    layer2_outputs(4462) <= b and not a;
    layer2_outputs(4463) <= b and not a;
    layer2_outputs(4464) <= a and not b;
    layer2_outputs(4465) <= not (a xor b);
    layer2_outputs(4466) <= a or b;
    layer2_outputs(4467) <= '0';
    layer2_outputs(4468) <= not a;
    layer2_outputs(4469) <= not (a and b);
    layer2_outputs(4470) <= not b;
    layer2_outputs(4471) <= not (a and b);
    layer2_outputs(4472) <= '0';
    layer2_outputs(4473) <= a and not b;
    layer2_outputs(4474) <= not (a or b);
    layer2_outputs(4475) <= not a or b;
    layer2_outputs(4476) <= b;
    layer2_outputs(4477) <= not (a and b);
    layer2_outputs(4478) <= not (a or b);
    layer2_outputs(4479) <= b and not a;
    layer2_outputs(4480) <= b and not a;
    layer2_outputs(4481) <= not (a xor b);
    layer2_outputs(4482) <= a and not b;
    layer2_outputs(4483) <= '1';
    layer2_outputs(4484) <= not (a and b);
    layer2_outputs(4485) <= a or b;
    layer2_outputs(4486) <= not (a or b);
    layer2_outputs(4487) <= a;
    layer2_outputs(4488) <= b;
    layer2_outputs(4489) <= a xor b;
    layer2_outputs(4490) <= not (a and b);
    layer2_outputs(4491) <= not (a or b);
    layer2_outputs(4492) <= a and b;
    layer2_outputs(4493) <= a;
    layer2_outputs(4494) <= not b or a;
    layer2_outputs(4495) <= not (a and b);
    layer2_outputs(4496) <= not a or b;
    layer2_outputs(4497) <= not b;
    layer2_outputs(4498) <= a and not b;
    layer2_outputs(4499) <= '1';
    layer2_outputs(4500) <= not a;
    layer2_outputs(4501) <= not (a and b);
    layer2_outputs(4502) <= b and not a;
    layer2_outputs(4503) <= not (a xor b);
    layer2_outputs(4504) <= a and not b;
    layer2_outputs(4505) <= a and not b;
    layer2_outputs(4506) <= not b or a;
    layer2_outputs(4507) <= not b or a;
    layer2_outputs(4508) <= not b;
    layer2_outputs(4509) <= not a or b;
    layer2_outputs(4510) <= '0';
    layer2_outputs(4511) <= a and not b;
    layer2_outputs(4512) <= not (a or b);
    layer2_outputs(4513) <= not (a or b);
    layer2_outputs(4514) <= not (a and b);
    layer2_outputs(4515) <= a and not b;
    layer2_outputs(4516) <= not b or a;
    layer2_outputs(4517) <= not (a or b);
    layer2_outputs(4518) <= not (a and b);
    layer2_outputs(4519) <= not a or b;
    layer2_outputs(4520) <= a;
    layer2_outputs(4521) <= not b;
    layer2_outputs(4522) <= not (a xor b);
    layer2_outputs(4523) <= b;
    layer2_outputs(4524) <= a xor b;
    layer2_outputs(4525) <= not a or b;
    layer2_outputs(4526) <= '1';
    layer2_outputs(4527) <= b;
    layer2_outputs(4528) <= a;
    layer2_outputs(4529) <= not a;
    layer2_outputs(4530) <= b and not a;
    layer2_outputs(4531) <= b;
    layer2_outputs(4532) <= a xor b;
    layer2_outputs(4533) <= a;
    layer2_outputs(4534) <= a and b;
    layer2_outputs(4535) <= '1';
    layer2_outputs(4536) <= not (a and b);
    layer2_outputs(4537) <= b and not a;
    layer2_outputs(4538) <= a or b;
    layer2_outputs(4539) <= not (a or b);
    layer2_outputs(4540) <= a;
    layer2_outputs(4541) <= not a;
    layer2_outputs(4542) <= a and b;
    layer2_outputs(4543) <= a or b;
    layer2_outputs(4544) <= not a;
    layer2_outputs(4545) <= a;
    layer2_outputs(4546) <= a or b;
    layer2_outputs(4547) <= '0';
    layer2_outputs(4548) <= '1';
    layer2_outputs(4549) <= a and not b;
    layer2_outputs(4550) <= a and not b;
    layer2_outputs(4551) <= a or b;
    layer2_outputs(4552) <= not (a or b);
    layer2_outputs(4553) <= not (a or b);
    layer2_outputs(4554) <= b;
    layer2_outputs(4555) <= not (a xor b);
    layer2_outputs(4556) <= not b;
    layer2_outputs(4557) <= not (a or b);
    layer2_outputs(4558) <= b;
    layer2_outputs(4559) <= not a;
    layer2_outputs(4560) <= not a;
    layer2_outputs(4561) <= not b or a;
    layer2_outputs(4562) <= not (a xor b);
    layer2_outputs(4563) <= b;
    layer2_outputs(4564) <= not (a or b);
    layer2_outputs(4565) <= b;
    layer2_outputs(4566) <= not b;
    layer2_outputs(4567) <= not a or b;
    layer2_outputs(4568) <= not (a and b);
    layer2_outputs(4569) <= not a or b;
    layer2_outputs(4570) <= not (a or b);
    layer2_outputs(4571) <= b;
    layer2_outputs(4572) <= not a;
    layer2_outputs(4573) <= a or b;
    layer2_outputs(4574) <= '1';
    layer2_outputs(4575) <= not a;
    layer2_outputs(4576) <= '1';
    layer2_outputs(4577) <= not a or b;
    layer2_outputs(4578) <= not a or b;
    layer2_outputs(4579) <= a or b;
    layer2_outputs(4580) <= not b;
    layer2_outputs(4581) <= a and not b;
    layer2_outputs(4582) <= a xor b;
    layer2_outputs(4583) <= not (a and b);
    layer2_outputs(4584) <= not (a or b);
    layer2_outputs(4585) <= not a or b;
    layer2_outputs(4586) <= not b;
    layer2_outputs(4587) <= a and not b;
    layer2_outputs(4588) <= not b;
    layer2_outputs(4589) <= a xor b;
    layer2_outputs(4590) <= not b;
    layer2_outputs(4591) <= not a;
    layer2_outputs(4592) <= b and not a;
    layer2_outputs(4593) <= '0';
    layer2_outputs(4594) <= not b or a;
    layer2_outputs(4595) <= not b;
    layer2_outputs(4596) <= '1';
    layer2_outputs(4597) <= not b;
    layer2_outputs(4598) <= a;
    layer2_outputs(4599) <= '1';
    layer2_outputs(4600) <= not b;
    layer2_outputs(4601) <= a and not b;
    layer2_outputs(4602) <= not (a or b);
    layer2_outputs(4603) <= b;
    layer2_outputs(4604) <= not (a xor b);
    layer2_outputs(4605) <= not b or a;
    layer2_outputs(4606) <= a and not b;
    layer2_outputs(4607) <= b;
    layer2_outputs(4608) <= a xor b;
    layer2_outputs(4609) <= not b;
    layer2_outputs(4610) <= '0';
    layer2_outputs(4611) <= not b;
    layer2_outputs(4612) <= not (a xor b);
    layer2_outputs(4613) <= not b or a;
    layer2_outputs(4614) <= b;
    layer2_outputs(4615) <= a;
    layer2_outputs(4616) <= '0';
    layer2_outputs(4617) <= not b or a;
    layer2_outputs(4618) <= not b or a;
    layer2_outputs(4619) <= not a;
    layer2_outputs(4620) <= b;
    layer2_outputs(4621) <= not a or b;
    layer2_outputs(4622) <= not b or a;
    layer2_outputs(4623) <= a and b;
    layer2_outputs(4624) <= not b or a;
    layer2_outputs(4625) <= a xor b;
    layer2_outputs(4626) <= a xor b;
    layer2_outputs(4627) <= a;
    layer2_outputs(4628) <= b and not a;
    layer2_outputs(4629) <= not (a or b);
    layer2_outputs(4630) <= '1';
    layer2_outputs(4631) <= a;
    layer2_outputs(4632) <= a and b;
    layer2_outputs(4633) <= not a or b;
    layer2_outputs(4634) <= '1';
    layer2_outputs(4635) <= not b or a;
    layer2_outputs(4636) <= not (a or b);
    layer2_outputs(4637) <= not (a and b);
    layer2_outputs(4638) <= a or b;
    layer2_outputs(4639) <= '0';
    layer2_outputs(4640) <= a;
    layer2_outputs(4641) <= a and b;
    layer2_outputs(4642) <= not b;
    layer2_outputs(4643) <= b;
    layer2_outputs(4644) <= not a;
    layer2_outputs(4645) <= a or b;
    layer2_outputs(4646) <= '1';
    layer2_outputs(4647) <= not a;
    layer2_outputs(4648) <= not (a and b);
    layer2_outputs(4649) <= not b or a;
    layer2_outputs(4650) <= a and not b;
    layer2_outputs(4651) <= a and not b;
    layer2_outputs(4652) <= not b;
    layer2_outputs(4653) <= not (a and b);
    layer2_outputs(4654) <= a and b;
    layer2_outputs(4655) <= not a or b;
    layer2_outputs(4656) <= b and not a;
    layer2_outputs(4657) <= not b;
    layer2_outputs(4658) <= a xor b;
    layer2_outputs(4659) <= not a or b;
    layer2_outputs(4660) <= '0';
    layer2_outputs(4661) <= not (a or b);
    layer2_outputs(4662) <= not (a and b);
    layer2_outputs(4663) <= a and b;
    layer2_outputs(4664) <= a;
    layer2_outputs(4665) <= not (a and b);
    layer2_outputs(4666) <= a and b;
    layer2_outputs(4667) <= not (a or b);
    layer2_outputs(4668) <= '0';
    layer2_outputs(4669) <= a;
    layer2_outputs(4670) <= not b;
    layer2_outputs(4671) <= not b or a;
    layer2_outputs(4672) <= b and not a;
    layer2_outputs(4673) <= not a or b;
    layer2_outputs(4674) <= '0';
    layer2_outputs(4675) <= a and not b;
    layer2_outputs(4676) <= '0';
    layer2_outputs(4677) <= not a;
    layer2_outputs(4678) <= a;
    layer2_outputs(4679) <= a and b;
    layer2_outputs(4680) <= a or b;
    layer2_outputs(4681) <= a or b;
    layer2_outputs(4682) <= not a;
    layer2_outputs(4683) <= a or b;
    layer2_outputs(4684) <= not (a and b);
    layer2_outputs(4685) <= not a;
    layer2_outputs(4686) <= not b;
    layer2_outputs(4687) <= a;
    layer2_outputs(4688) <= not b or a;
    layer2_outputs(4689) <= not b or a;
    layer2_outputs(4690) <= b and not a;
    layer2_outputs(4691) <= a and not b;
    layer2_outputs(4692) <= '1';
    layer2_outputs(4693) <= not (a and b);
    layer2_outputs(4694) <= not (a and b);
    layer2_outputs(4695) <= a;
    layer2_outputs(4696) <= '0';
    layer2_outputs(4697) <= b;
    layer2_outputs(4698) <= a and not b;
    layer2_outputs(4699) <= not b or a;
    layer2_outputs(4700) <= a or b;
    layer2_outputs(4701) <= not (a or b);
    layer2_outputs(4702) <= not b or a;
    layer2_outputs(4703) <= not a or b;
    layer2_outputs(4704) <= not a;
    layer2_outputs(4705) <= not a or b;
    layer2_outputs(4706) <= a;
    layer2_outputs(4707) <= a and b;
    layer2_outputs(4708) <= not a or b;
    layer2_outputs(4709) <= a and not b;
    layer2_outputs(4710) <= not (a or b);
    layer2_outputs(4711) <= not b or a;
    layer2_outputs(4712) <= not (a and b);
    layer2_outputs(4713) <= not b;
    layer2_outputs(4714) <= not (a or b);
    layer2_outputs(4715) <= not b;
    layer2_outputs(4716) <= not (a or b);
    layer2_outputs(4717) <= a or b;
    layer2_outputs(4718) <= '1';
    layer2_outputs(4719) <= a xor b;
    layer2_outputs(4720) <= a;
    layer2_outputs(4721) <= not b;
    layer2_outputs(4722) <= not (a and b);
    layer2_outputs(4723) <= a;
    layer2_outputs(4724) <= a and not b;
    layer2_outputs(4725) <= not a or b;
    layer2_outputs(4726) <= not b or a;
    layer2_outputs(4727) <= a or b;
    layer2_outputs(4728) <= a and b;
    layer2_outputs(4729) <= not b or a;
    layer2_outputs(4730) <= not (a and b);
    layer2_outputs(4731) <= not b or a;
    layer2_outputs(4732) <= b;
    layer2_outputs(4733) <= a;
    layer2_outputs(4734) <= not (a xor b);
    layer2_outputs(4735) <= a and not b;
    layer2_outputs(4736) <= b and not a;
    layer2_outputs(4737) <= a and b;
    layer2_outputs(4738) <= not b or a;
    layer2_outputs(4739) <= a;
    layer2_outputs(4740) <= b and not a;
    layer2_outputs(4741) <= a and b;
    layer2_outputs(4742) <= a and not b;
    layer2_outputs(4743) <= '0';
    layer2_outputs(4744) <= a;
    layer2_outputs(4745) <= not b or a;
    layer2_outputs(4746) <= a;
    layer2_outputs(4747) <= a and b;
    layer2_outputs(4748) <= not b or a;
    layer2_outputs(4749) <= a;
    layer2_outputs(4750) <= not (a or b);
    layer2_outputs(4751) <= a;
    layer2_outputs(4752) <= not (a xor b);
    layer2_outputs(4753) <= a and b;
    layer2_outputs(4754) <= a or b;
    layer2_outputs(4755) <= b;
    layer2_outputs(4756) <= a and not b;
    layer2_outputs(4757) <= b;
    layer2_outputs(4758) <= b;
    layer2_outputs(4759) <= not (a or b);
    layer2_outputs(4760) <= not b;
    layer2_outputs(4761) <= '0';
    layer2_outputs(4762) <= a and b;
    layer2_outputs(4763) <= not b or a;
    layer2_outputs(4764) <= a or b;
    layer2_outputs(4765) <= a xor b;
    layer2_outputs(4766) <= b;
    layer2_outputs(4767) <= a;
    layer2_outputs(4768) <= '0';
    layer2_outputs(4769) <= a and not b;
    layer2_outputs(4770) <= not b or a;
    layer2_outputs(4771) <= not b;
    layer2_outputs(4772) <= not (a or b);
    layer2_outputs(4773) <= '1';
    layer2_outputs(4774) <= '0';
    layer2_outputs(4775) <= not a or b;
    layer2_outputs(4776) <= not (a or b);
    layer2_outputs(4777) <= '1';
    layer2_outputs(4778) <= not (a xor b);
    layer2_outputs(4779) <= not (a and b);
    layer2_outputs(4780) <= not (a and b);
    layer2_outputs(4781) <= a and b;
    layer2_outputs(4782) <= a and not b;
    layer2_outputs(4783) <= not (a xor b);
    layer2_outputs(4784) <= not b;
    layer2_outputs(4785) <= not a;
    layer2_outputs(4786) <= a;
    layer2_outputs(4787) <= not a or b;
    layer2_outputs(4788) <= a xor b;
    layer2_outputs(4789) <= a and b;
    layer2_outputs(4790) <= a;
    layer2_outputs(4791) <= not (a xor b);
    layer2_outputs(4792) <= a and b;
    layer2_outputs(4793) <= not a;
    layer2_outputs(4794) <= b and not a;
    layer2_outputs(4795) <= '0';
    layer2_outputs(4796) <= b;
    layer2_outputs(4797) <= not (a and b);
    layer2_outputs(4798) <= not (a or b);
    layer2_outputs(4799) <= b;
    layer2_outputs(4800) <= b;
    layer2_outputs(4801) <= not b or a;
    layer2_outputs(4802) <= not (a or b);
    layer2_outputs(4803) <= a;
    layer2_outputs(4804) <= a or b;
    layer2_outputs(4805) <= a and not b;
    layer2_outputs(4806) <= a;
    layer2_outputs(4807) <= b and not a;
    layer2_outputs(4808) <= not a;
    layer2_outputs(4809) <= b;
    layer2_outputs(4810) <= b;
    layer2_outputs(4811) <= '1';
    layer2_outputs(4812) <= not (a and b);
    layer2_outputs(4813) <= b;
    layer2_outputs(4814) <= not b or a;
    layer2_outputs(4815) <= not b;
    layer2_outputs(4816) <= a;
    layer2_outputs(4817) <= not (a or b);
    layer2_outputs(4818) <= b;
    layer2_outputs(4819) <= '1';
    layer2_outputs(4820) <= not (a or b);
    layer2_outputs(4821) <= b;
    layer2_outputs(4822) <= not b or a;
    layer2_outputs(4823) <= not b or a;
    layer2_outputs(4824) <= '0';
    layer2_outputs(4825) <= a;
    layer2_outputs(4826) <= not (a and b);
    layer2_outputs(4827) <= a;
    layer2_outputs(4828) <= b;
    layer2_outputs(4829) <= not (a or b);
    layer2_outputs(4830) <= a or b;
    layer2_outputs(4831) <= not a;
    layer2_outputs(4832) <= b;
    layer2_outputs(4833) <= '0';
    layer2_outputs(4834) <= not a or b;
    layer2_outputs(4835) <= a or b;
    layer2_outputs(4836) <= not b;
    layer2_outputs(4837) <= a;
    layer2_outputs(4838) <= a and b;
    layer2_outputs(4839) <= a or b;
    layer2_outputs(4840) <= not a;
    layer2_outputs(4841) <= not b;
    layer2_outputs(4842) <= a xor b;
    layer2_outputs(4843) <= a;
    layer2_outputs(4844) <= '1';
    layer2_outputs(4845) <= not b or a;
    layer2_outputs(4846) <= not a;
    layer2_outputs(4847) <= '0';
    layer2_outputs(4848) <= b;
    layer2_outputs(4849) <= a or b;
    layer2_outputs(4850) <= '0';
    layer2_outputs(4851) <= a and not b;
    layer2_outputs(4852) <= '1';
    layer2_outputs(4853) <= '1';
    layer2_outputs(4854) <= not (a and b);
    layer2_outputs(4855) <= a and not b;
    layer2_outputs(4856) <= not b;
    layer2_outputs(4857) <= b;
    layer2_outputs(4858) <= b;
    layer2_outputs(4859) <= b;
    layer2_outputs(4860) <= '1';
    layer2_outputs(4861) <= not (a xor b);
    layer2_outputs(4862) <= a;
    layer2_outputs(4863) <= b and not a;
    layer2_outputs(4864) <= a;
    layer2_outputs(4865) <= not b or a;
    layer2_outputs(4866) <= '1';
    layer2_outputs(4867) <= a or b;
    layer2_outputs(4868) <= b;
    layer2_outputs(4869) <= not (a or b);
    layer2_outputs(4870) <= b and not a;
    layer2_outputs(4871) <= a and not b;
    layer2_outputs(4872) <= not (a and b);
    layer2_outputs(4873) <= '0';
    layer2_outputs(4874) <= not b;
    layer2_outputs(4875) <= a and b;
    layer2_outputs(4876) <= a and not b;
    layer2_outputs(4877) <= not a;
    layer2_outputs(4878) <= not (a or b);
    layer2_outputs(4879) <= not a or b;
    layer2_outputs(4880) <= a and b;
    layer2_outputs(4881) <= a and not b;
    layer2_outputs(4882) <= not (a and b);
    layer2_outputs(4883) <= not b;
    layer2_outputs(4884) <= not a or b;
    layer2_outputs(4885) <= b;
    layer2_outputs(4886) <= not b or a;
    layer2_outputs(4887) <= a;
    layer2_outputs(4888) <= not a;
    layer2_outputs(4889) <= a and b;
    layer2_outputs(4890) <= a or b;
    layer2_outputs(4891) <= not a;
    layer2_outputs(4892) <= not a;
    layer2_outputs(4893) <= not b or a;
    layer2_outputs(4894) <= b and not a;
    layer2_outputs(4895) <= a and not b;
    layer2_outputs(4896) <= not a;
    layer2_outputs(4897) <= '1';
    layer2_outputs(4898) <= not (a or b);
    layer2_outputs(4899) <= not a or b;
    layer2_outputs(4900) <= '1';
    layer2_outputs(4901) <= not (a and b);
    layer2_outputs(4902) <= a and not b;
    layer2_outputs(4903) <= not a;
    layer2_outputs(4904) <= a;
    layer2_outputs(4905) <= b and not a;
    layer2_outputs(4906) <= a or b;
    layer2_outputs(4907) <= not b;
    layer2_outputs(4908) <= '1';
    layer2_outputs(4909) <= b and not a;
    layer2_outputs(4910) <= not b or a;
    layer2_outputs(4911) <= a and b;
    layer2_outputs(4912) <= not (a xor b);
    layer2_outputs(4913) <= not a;
    layer2_outputs(4914) <= not a;
    layer2_outputs(4915) <= b;
    layer2_outputs(4916) <= not b or a;
    layer2_outputs(4917) <= b and not a;
    layer2_outputs(4918) <= a and not b;
    layer2_outputs(4919) <= a and not b;
    layer2_outputs(4920) <= not a;
    layer2_outputs(4921) <= not a;
    layer2_outputs(4922) <= a and b;
    layer2_outputs(4923) <= a and not b;
    layer2_outputs(4924) <= not (a or b);
    layer2_outputs(4925) <= not (a and b);
    layer2_outputs(4926) <= b;
    layer2_outputs(4927) <= a or b;
    layer2_outputs(4928) <= '0';
    layer2_outputs(4929) <= '0';
    layer2_outputs(4930) <= a;
    layer2_outputs(4931) <= b;
    layer2_outputs(4932) <= not a;
    layer2_outputs(4933) <= not (a xor b);
    layer2_outputs(4934) <= a and b;
    layer2_outputs(4935) <= a and b;
    layer2_outputs(4936) <= not (a and b);
    layer2_outputs(4937) <= not a;
    layer2_outputs(4938) <= a and b;
    layer2_outputs(4939) <= not (a xor b);
    layer2_outputs(4940) <= not a;
    layer2_outputs(4941) <= not a or b;
    layer2_outputs(4942) <= a xor b;
    layer2_outputs(4943) <= a and not b;
    layer2_outputs(4944) <= not a or b;
    layer2_outputs(4945) <= b and not a;
    layer2_outputs(4946) <= a;
    layer2_outputs(4947) <= b;
    layer2_outputs(4948) <= b;
    layer2_outputs(4949) <= b;
    layer2_outputs(4950) <= not (a and b);
    layer2_outputs(4951) <= a or b;
    layer2_outputs(4952) <= a and b;
    layer2_outputs(4953) <= a;
    layer2_outputs(4954) <= a and not b;
    layer2_outputs(4955) <= b;
    layer2_outputs(4956) <= not (a or b);
    layer2_outputs(4957) <= not a or b;
    layer2_outputs(4958) <= b;
    layer2_outputs(4959) <= b;
    layer2_outputs(4960) <= '1';
    layer2_outputs(4961) <= b;
    layer2_outputs(4962) <= not (a and b);
    layer2_outputs(4963) <= not a or b;
    layer2_outputs(4964) <= not b or a;
    layer2_outputs(4965) <= a;
    layer2_outputs(4966) <= '0';
    layer2_outputs(4967) <= not (a or b);
    layer2_outputs(4968) <= not a or b;
    layer2_outputs(4969) <= a xor b;
    layer2_outputs(4970) <= a and not b;
    layer2_outputs(4971) <= '1';
    layer2_outputs(4972) <= b;
    layer2_outputs(4973) <= a and b;
    layer2_outputs(4974) <= a and not b;
    layer2_outputs(4975) <= b and not a;
    layer2_outputs(4976) <= not (a or b);
    layer2_outputs(4977) <= not b;
    layer2_outputs(4978) <= a;
    layer2_outputs(4979) <= a and not b;
    layer2_outputs(4980) <= not b or a;
    layer2_outputs(4981) <= not a or b;
    layer2_outputs(4982) <= b;
    layer2_outputs(4983) <= a and b;
    layer2_outputs(4984) <= not (a or b);
    layer2_outputs(4985) <= not b or a;
    layer2_outputs(4986) <= not (a or b);
    layer2_outputs(4987) <= not b or a;
    layer2_outputs(4988) <= not (a or b);
    layer2_outputs(4989) <= not a;
    layer2_outputs(4990) <= not b;
    layer2_outputs(4991) <= not (a or b);
    layer2_outputs(4992) <= b;
    layer2_outputs(4993) <= not a;
    layer2_outputs(4994) <= a and b;
    layer2_outputs(4995) <= not a;
    layer2_outputs(4996) <= not b;
    layer2_outputs(4997) <= '1';
    layer2_outputs(4998) <= not a or b;
    layer2_outputs(4999) <= a and b;
    layer2_outputs(5000) <= not (a and b);
    layer2_outputs(5001) <= not (a and b);
    layer2_outputs(5002) <= b;
    layer2_outputs(5003) <= not b or a;
    layer2_outputs(5004) <= a and not b;
    layer2_outputs(5005) <= a and not b;
    layer2_outputs(5006) <= not b;
    layer2_outputs(5007) <= '0';
    layer2_outputs(5008) <= a and not b;
    layer2_outputs(5009) <= b;
    layer2_outputs(5010) <= a or b;
    layer2_outputs(5011) <= a and not b;
    layer2_outputs(5012) <= a xor b;
    layer2_outputs(5013) <= a;
    layer2_outputs(5014) <= a and b;
    layer2_outputs(5015) <= not (a xor b);
    layer2_outputs(5016) <= b;
    layer2_outputs(5017) <= a or b;
    layer2_outputs(5018) <= a and b;
    layer2_outputs(5019) <= b and not a;
    layer2_outputs(5020) <= not (a and b);
    layer2_outputs(5021) <= not (a xor b);
    layer2_outputs(5022) <= b;
    layer2_outputs(5023) <= not a;
    layer2_outputs(5024) <= a and not b;
    layer2_outputs(5025) <= not a or b;
    layer2_outputs(5026) <= not (a and b);
    layer2_outputs(5027) <= not a;
    layer2_outputs(5028) <= a or b;
    layer2_outputs(5029) <= not b or a;
    layer2_outputs(5030) <= a or b;
    layer2_outputs(5031) <= not a;
    layer2_outputs(5032) <= a;
    layer2_outputs(5033) <= not a or b;
    layer2_outputs(5034) <= a and b;
    layer2_outputs(5035) <= a and not b;
    layer2_outputs(5036) <= not b;
    layer2_outputs(5037) <= a and not b;
    layer2_outputs(5038) <= not a;
    layer2_outputs(5039) <= not b;
    layer2_outputs(5040) <= not b;
    layer2_outputs(5041) <= not b;
    layer2_outputs(5042) <= '0';
    layer2_outputs(5043) <= a xor b;
    layer2_outputs(5044) <= not (a or b);
    layer2_outputs(5045) <= not a;
    layer2_outputs(5046) <= a or b;
    layer2_outputs(5047) <= not a;
    layer2_outputs(5048) <= not a or b;
    layer2_outputs(5049) <= not a;
    layer2_outputs(5050) <= not (a or b);
    layer2_outputs(5051) <= a and not b;
    layer2_outputs(5052) <= not a;
    layer2_outputs(5053) <= a and b;
    layer2_outputs(5054) <= '0';
    layer2_outputs(5055) <= '1';
    layer2_outputs(5056) <= a xor b;
    layer2_outputs(5057) <= a or b;
    layer2_outputs(5058) <= not b or a;
    layer2_outputs(5059) <= '0';
    layer2_outputs(5060) <= b;
    layer2_outputs(5061) <= a and b;
    layer2_outputs(5062) <= not b;
    layer2_outputs(5063) <= not b;
    layer2_outputs(5064) <= not (a or b);
    layer2_outputs(5065) <= not b;
    layer2_outputs(5066) <= a or b;
    layer2_outputs(5067) <= a or b;
    layer2_outputs(5068) <= a and not b;
    layer2_outputs(5069) <= not b;
    layer2_outputs(5070) <= b and not a;
    layer2_outputs(5071) <= not a;
    layer2_outputs(5072) <= b;
    layer2_outputs(5073) <= not (a or b);
    layer2_outputs(5074) <= not b;
    layer2_outputs(5075) <= a and not b;
    layer2_outputs(5076) <= b;
    layer2_outputs(5077) <= b and not a;
    layer2_outputs(5078) <= not (a and b);
    layer2_outputs(5079) <= a and not b;
    layer2_outputs(5080) <= b;
    layer2_outputs(5081) <= b and not a;
    layer2_outputs(5082) <= '0';
    layer2_outputs(5083) <= not b;
    layer2_outputs(5084) <= not a or b;
    layer2_outputs(5085) <= a and b;
    layer2_outputs(5086) <= b and not a;
    layer2_outputs(5087) <= a xor b;
    layer2_outputs(5088) <= b;
    layer2_outputs(5089) <= a;
    layer2_outputs(5090) <= not b;
    layer2_outputs(5091) <= a;
    layer2_outputs(5092) <= not a;
    layer2_outputs(5093) <= '1';
    layer2_outputs(5094) <= a or b;
    layer2_outputs(5095) <= not a;
    layer2_outputs(5096) <= not a;
    layer2_outputs(5097) <= not (a or b);
    layer2_outputs(5098) <= not (a xor b);
    layer2_outputs(5099) <= a and b;
    layer2_outputs(5100) <= a and b;
    layer2_outputs(5101) <= not (a or b);
    layer2_outputs(5102) <= not b or a;
    layer2_outputs(5103) <= a and b;
    layer2_outputs(5104) <= b and not a;
    layer2_outputs(5105) <= not (a and b);
    layer2_outputs(5106) <= not (a xor b);
    layer2_outputs(5107) <= a or b;
    layer2_outputs(5108) <= not b;
    layer2_outputs(5109) <= not (a and b);
    layer2_outputs(5110) <= not (a or b);
    layer2_outputs(5111) <= not (a and b);
    layer2_outputs(5112) <= a and not b;
    layer2_outputs(5113) <= b and not a;
    layer2_outputs(5114) <= a and not b;
    layer2_outputs(5115) <= a;
    layer2_outputs(5116) <= b;
    layer2_outputs(5117) <= not b;
    layer2_outputs(5118) <= a xor b;
    layer2_outputs(5119) <= a and b;
    layer2_outputs(5120) <= a and not b;
    layer2_outputs(5121) <= a and b;
    layer2_outputs(5122) <= a and not b;
    layer2_outputs(5123) <= a;
    layer2_outputs(5124) <= not b or a;
    layer2_outputs(5125) <= not b or a;
    layer2_outputs(5126) <= not a or b;
    layer2_outputs(5127) <= not b;
    layer2_outputs(5128) <= not a;
    layer2_outputs(5129) <= not a or b;
    layer2_outputs(5130) <= not b;
    layer2_outputs(5131) <= not (a or b);
    layer2_outputs(5132) <= a xor b;
    layer2_outputs(5133) <= a or b;
    layer2_outputs(5134) <= not b;
    layer2_outputs(5135) <= not a or b;
    layer2_outputs(5136) <= not b or a;
    layer2_outputs(5137) <= not a;
    layer2_outputs(5138) <= not b;
    layer2_outputs(5139) <= not a or b;
    layer2_outputs(5140) <= not (a xor b);
    layer2_outputs(5141) <= not (a or b);
    layer2_outputs(5142) <= '0';
    layer2_outputs(5143) <= not a or b;
    layer2_outputs(5144) <= '1';
    layer2_outputs(5145) <= not a or b;
    layer2_outputs(5146) <= b;
    layer2_outputs(5147) <= '1';
    layer2_outputs(5148) <= not (a or b);
    layer2_outputs(5149) <= not (a or b);
    layer2_outputs(5150) <= b;
    layer2_outputs(5151) <= b;
    layer2_outputs(5152) <= not a;
    layer2_outputs(5153) <= not a;
    layer2_outputs(5154) <= '0';
    layer2_outputs(5155) <= not b or a;
    layer2_outputs(5156) <= b;
    layer2_outputs(5157) <= a or b;
    layer2_outputs(5158) <= not b;
    layer2_outputs(5159) <= not a or b;
    layer2_outputs(5160) <= not (a or b);
    layer2_outputs(5161) <= b;
    layer2_outputs(5162) <= b and not a;
    layer2_outputs(5163) <= not (a or b);
    layer2_outputs(5164) <= a;
    layer2_outputs(5165) <= not (a and b);
    layer2_outputs(5166) <= a and not b;
    layer2_outputs(5167) <= a;
    layer2_outputs(5168) <= not b;
    layer2_outputs(5169) <= a and b;
    layer2_outputs(5170) <= a;
    layer2_outputs(5171) <= not a or b;
    layer2_outputs(5172) <= b and not a;
    layer2_outputs(5173) <= b;
    layer2_outputs(5174) <= not a or b;
    layer2_outputs(5175) <= b and not a;
    layer2_outputs(5176) <= not (a and b);
    layer2_outputs(5177) <= not b or a;
    layer2_outputs(5178) <= not (a and b);
    layer2_outputs(5179) <= not b or a;
    layer2_outputs(5180) <= b;
    layer2_outputs(5181) <= not b;
    layer2_outputs(5182) <= a;
    layer2_outputs(5183) <= not a;
    layer2_outputs(5184) <= not a;
    layer2_outputs(5185) <= a and not b;
    layer2_outputs(5186) <= not a;
    layer2_outputs(5187) <= '1';
    layer2_outputs(5188) <= b;
    layer2_outputs(5189) <= '0';
    layer2_outputs(5190) <= not (a and b);
    layer2_outputs(5191) <= b;
    layer2_outputs(5192) <= not (a and b);
    layer2_outputs(5193) <= not (a or b);
    layer2_outputs(5194) <= not b;
    layer2_outputs(5195) <= not (a or b);
    layer2_outputs(5196) <= not (a and b);
    layer2_outputs(5197) <= b;
    layer2_outputs(5198) <= not b;
    layer2_outputs(5199) <= b;
    layer2_outputs(5200) <= a;
    layer2_outputs(5201) <= '1';
    layer2_outputs(5202) <= not b or a;
    layer2_outputs(5203) <= a or b;
    layer2_outputs(5204) <= a and b;
    layer2_outputs(5205) <= b and not a;
    layer2_outputs(5206) <= not (a xor b);
    layer2_outputs(5207) <= a or b;
    layer2_outputs(5208) <= '1';
    layer2_outputs(5209) <= not a or b;
    layer2_outputs(5210) <= not a or b;
    layer2_outputs(5211) <= b;
    layer2_outputs(5212) <= not (a and b);
    layer2_outputs(5213) <= a;
    layer2_outputs(5214) <= not a;
    layer2_outputs(5215) <= b;
    layer2_outputs(5216) <= '1';
    layer2_outputs(5217) <= not a or b;
    layer2_outputs(5218) <= b;
    layer2_outputs(5219) <= not (a or b);
    layer2_outputs(5220) <= not a or b;
    layer2_outputs(5221) <= a and b;
    layer2_outputs(5222) <= '1';
    layer2_outputs(5223) <= a;
    layer2_outputs(5224) <= not a or b;
    layer2_outputs(5225) <= a or b;
    layer2_outputs(5226) <= not a or b;
    layer2_outputs(5227) <= not (a xor b);
    layer2_outputs(5228) <= not b;
    layer2_outputs(5229) <= '1';
    layer2_outputs(5230) <= not b;
    layer2_outputs(5231) <= not a;
    layer2_outputs(5232) <= b;
    layer2_outputs(5233) <= a;
    layer2_outputs(5234) <= b;
    layer2_outputs(5235) <= not b;
    layer2_outputs(5236) <= not (a or b);
    layer2_outputs(5237) <= not (a and b);
    layer2_outputs(5238) <= a or b;
    layer2_outputs(5239) <= b and not a;
    layer2_outputs(5240) <= a;
    layer2_outputs(5241) <= not a or b;
    layer2_outputs(5242) <= b and not a;
    layer2_outputs(5243) <= not (a and b);
    layer2_outputs(5244) <= b and not a;
    layer2_outputs(5245) <= not b;
    layer2_outputs(5246) <= not b or a;
    layer2_outputs(5247) <= '1';
    layer2_outputs(5248) <= '0';
    layer2_outputs(5249) <= a;
    layer2_outputs(5250) <= not (a and b);
    layer2_outputs(5251) <= not b or a;
    layer2_outputs(5252) <= b;
    layer2_outputs(5253) <= '1';
    layer2_outputs(5254) <= a;
    layer2_outputs(5255) <= not b;
    layer2_outputs(5256) <= not a or b;
    layer2_outputs(5257) <= b and not a;
    layer2_outputs(5258) <= not (a and b);
    layer2_outputs(5259) <= b and not a;
    layer2_outputs(5260) <= a and b;
    layer2_outputs(5261) <= a;
    layer2_outputs(5262) <= b and not a;
    layer2_outputs(5263) <= a;
    layer2_outputs(5264) <= not b or a;
    layer2_outputs(5265) <= a or b;
    layer2_outputs(5266) <= a and not b;
    layer2_outputs(5267) <= a and not b;
    layer2_outputs(5268) <= b;
    layer2_outputs(5269) <= not b or a;
    layer2_outputs(5270) <= not a;
    layer2_outputs(5271) <= not a or b;
    layer2_outputs(5272) <= a or b;
    layer2_outputs(5273) <= not a or b;
    layer2_outputs(5274) <= a or b;
    layer2_outputs(5275) <= a or b;
    layer2_outputs(5276) <= not (a or b);
    layer2_outputs(5277) <= '1';
    layer2_outputs(5278) <= '1';
    layer2_outputs(5279) <= not a or b;
    layer2_outputs(5280) <= '1';
    layer2_outputs(5281) <= not a or b;
    layer2_outputs(5282) <= not (a or b);
    layer2_outputs(5283) <= not (a xor b);
    layer2_outputs(5284) <= b;
    layer2_outputs(5285) <= a and not b;
    layer2_outputs(5286) <= a;
    layer2_outputs(5287) <= '0';
    layer2_outputs(5288) <= a and not b;
    layer2_outputs(5289) <= not a or b;
    layer2_outputs(5290) <= not (a and b);
    layer2_outputs(5291) <= a and not b;
    layer2_outputs(5292) <= not b;
    layer2_outputs(5293) <= not (a and b);
    layer2_outputs(5294) <= '1';
    layer2_outputs(5295) <= not (a and b);
    layer2_outputs(5296) <= not a or b;
    layer2_outputs(5297) <= b and not a;
    layer2_outputs(5298) <= a and not b;
    layer2_outputs(5299) <= a;
    layer2_outputs(5300) <= a;
    layer2_outputs(5301) <= not (a or b);
    layer2_outputs(5302) <= not b or a;
    layer2_outputs(5303) <= not (a and b);
    layer2_outputs(5304) <= not a or b;
    layer2_outputs(5305) <= a and b;
    layer2_outputs(5306) <= not (a or b);
    layer2_outputs(5307) <= a;
    layer2_outputs(5308) <= not a;
    layer2_outputs(5309) <= not b;
    layer2_outputs(5310) <= not a or b;
    layer2_outputs(5311) <= '0';
    layer2_outputs(5312) <= not a;
    layer2_outputs(5313) <= '1';
    layer2_outputs(5314) <= not (a and b);
    layer2_outputs(5315) <= not b or a;
    layer2_outputs(5316) <= not (a and b);
    layer2_outputs(5317) <= not (a and b);
    layer2_outputs(5318) <= '1';
    layer2_outputs(5319) <= not a or b;
    layer2_outputs(5320) <= a or b;
    layer2_outputs(5321) <= b and not a;
    layer2_outputs(5322) <= a and b;
    layer2_outputs(5323) <= not b;
    layer2_outputs(5324) <= '0';
    layer2_outputs(5325) <= b;
    layer2_outputs(5326) <= a and not b;
    layer2_outputs(5327) <= b and not a;
    layer2_outputs(5328) <= not a or b;
    layer2_outputs(5329) <= b;
    layer2_outputs(5330) <= not a;
    layer2_outputs(5331) <= b and not a;
    layer2_outputs(5332) <= not (a or b);
    layer2_outputs(5333) <= not (a xor b);
    layer2_outputs(5334) <= not a or b;
    layer2_outputs(5335) <= b and not a;
    layer2_outputs(5336) <= not (a and b);
    layer2_outputs(5337) <= not (a and b);
    layer2_outputs(5338) <= not b or a;
    layer2_outputs(5339) <= not (a xor b);
    layer2_outputs(5340) <= a;
    layer2_outputs(5341) <= '0';
    layer2_outputs(5342) <= a;
    layer2_outputs(5343) <= a;
    layer2_outputs(5344) <= a and not b;
    layer2_outputs(5345) <= not (a and b);
    layer2_outputs(5346) <= not a or b;
    layer2_outputs(5347) <= a and b;
    layer2_outputs(5348) <= a and b;
    layer2_outputs(5349) <= not (a or b);
    layer2_outputs(5350) <= a;
    layer2_outputs(5351) <= '1';
    layer2_outputs(5352) <= a;
    layer2_outputs(5353) <= '1';
    layer2_outputs(5354) <= '1';
    layer2_outputs(5355) <= not a;
    layer2_outputs(5356) <= b;
    layer2_outputs(5357) <= a and not b;
    layer2_outputs(5358) <= b;
    layer2_outputs(5359) <= not a;
    layer2_outputs(5360) <= not a;
    layer2_outputs(5361) <= b;
    layer2_outputs(5362) <= a and b;
    layer2_outputs(5363) <= a;
    layer2_outputs(5364) <= a and not b;
    layer2_outputs(5365) <= not a;
    layer2_outputs(5366) <= not b or a;
    layer2_outputs(5367) <= '0';
    layer2_outputs(5368) <= not a;
    layer2_outputs(5369) <= a or b;
    layer2_outputs(5370) <= b and not a;
    layer2_outputs(5371) <= a and b;
    layer2_outputs(5372) <= not a or b;
    layer2_outputs(5373) <= '0';
    layer2_outputs(5374) <= a;
    layer2_outputs(5375) <= not (a and b);
    layer2_outputs(5376) <= b and not a;
    layer2_outputs(5377) <= not (a or b);
    layer2_outputs(5378) <= not (a and b);
    layer2_outputs(5379) <= a or b;
    layer2_outputs(5380) <= a;
    layer2_outputs(5381) <= a and not b;
    layer2_outputs(5382) <= a or b;
    layer2_outputs(5383) <= not b or a;
    layer2_outputs(5384) <= a;
    layer2_outputs(5385) <= not (a and b);
    layer2_outputs(5386) <= not b;
    layer2_outputs(5387) <= not (a or b);
    layer2_outputs(5388) <= not b or a;
    layer2_outputs(5389) <= '1';
    layer2_outputs(5390) <= not b or a;
    layer2_outputs(5391) <= b;
    layer2_outputs(5392) <= b;
    layer2_outputs(5393) <= a or b;
    layer2_outputs(5394) <= a or b;
    layer2_outputs(5395) <= '1';
    layer2_outputs(5396) <= not a;
    layer2_outputs(5397) <= a;
    layer2_outputs(5398) <= a;
    layer2_outputs(5399) <= a and not b;
    layer2_outputs(5400) <= '1';
    layer2_outputs(5401) <= a and b;
    layer2_outputs(5402) <= a xor b;
    layer2_outputs(5403) <= not b or a;
    layer2_outputs(5404) <= not a;
    layer2_outputs(5405) <= a or b;
    layer2_outputs(5406) <= not a;
    layer2_outputs(5407) <= not a;
    layer2_outputs(5408) <= not a;
    layer2_outputs(5409) <= not (a or b);
    layer2_outputs(5410) <= not a;
    layer2_outputs(5411) <= b;
    layer2_outputs(5412) <= a xor b;
    layer2_outputs(5413) <= '0';
    layer2_outputs(5414) <= a and b;
    layer2_outputs(5415) <= a or b;
    layer2_outputs(5416) <= a and b;
    layer2_outputs(5417) <= not (a and b);
    layer2_outputs(5418) <= not b;
    layer2_outputs(5419) <= not b;
    layer2_outputs(5420) <= not a or b;
    layer2_outputs(5421) <= not (a or b);
    layer2_outputs(5422) <= not (a or b);
    layer2_outputs(5423) <= a;
    layer2_outputs(5424) <= a and not b;
    layer2_outputs(5425) <= b and not a;
    layer2_outputs(5426) <= b and not a;
    layer2_outputs(5427) <= not (a or b);
    layer2_outputs(5428) <= '1';
    layer2_outputs(5429) <= not a;
    layer2_outputs(5430) <= a xor b;
    layer2_outputs(5431) <= a xor b;
    layer2_outputs(5432) <= b;
    layer2_outputs(5433) <= b;
    layer2_outputs(5434) <= not a or b;
    layer2_outputs(5435) <= a and not b;
    layer2_outputs(5436) <= a and b;
    layer2_outputs(5437) <= not (a xor b);
    layer2_outputs(5438) <= '1';
    layer2_outputs(5439) <= a and not b;
    layer2_outputs(5440) <= a or b;
    layer2_outputs(5441) <= '1';
    layer2_outputs(5442) <= not (a and b);
    layer2_outputs(5443) <= a;
    layer2_outputs(5444) <= not a or b;
    layer2_outputs(5445) <= a and not b;
    layer2_outputs(5446) <= not (a xor b);
    layer2_outputs(5447) <= a;
    layer2_outputs(5448) <= not a;
    layer2_outputs(5449) <= not b;
    layer2_outputs(5450) <= b and not a;
    layer2_outputs(5451) <= '1';
    layer2_outputs(5452) <= '1';
    layer2_outputs(5453) <= b and not a;
    layer2_outputs(5454) <= a;
    layer2_outputs(5455) <= a and not b;
    layer2_outputs(5456) <= not a;
    layer2_outputs(5457) <= b;
    layer2_outputs(5458) <= not b or a;
    layer2_outputs(5459) <= not a or b;
    layer2_outputs(5460) <= a and not b;
    layer2_outputs(5461) <= a and not b;
    layer2_outputs(5462) <= a and b;
    layer2_outputs(5463) <= not b;
    layer2_outputs(5464) <= b;
    layer2_outputs(5465) <= a and b;
    layer2_outputs(5466) <= b;
    layer2_outputs(5467) <= not (a or b);
    layer2_outputs(5468) <= not b;
    layer2_outputs(5469) <= a or b;
    layer2_outputs(5470) <= b;
    layer2_outputs(5471) <= not b or a;
    layer2_outputs(5472) <= a and b;
    layer2_outputs(5473) <= '1';
    layer2_outputs(5474) <= a;
    layer2_outputs(5475) <= a and b;
    layer2_outputs(5476) <= a and b;
    layer2_outputs(5477) <= not (a and b);
    layer2_outputs(5478) <= a and b;
    layer2_outputs(5479) <= b and not a;
    layer2_outputs(5480) <= not a;
    layer2_outputs(5481) <= not (a and b);
    layer2_outputs(5482) <= b;
    layer2_outputs(5483) <= a or b;
    layer2_outputs(5484) <= a and not b;
    layer2_outputs(5485) <= not a or b;
    layer2_outputs(5486) <= a and b;
    layer2_outputs(5487) <= not b;
    layer2_outputs(5488) <= not (a or b);
    layer2_outputs(5489) <= a xor b;
    layer2_outputs(5490) <= a and not b;
    layer2_outputs(5491) <= not (a and b);
    layer2_outputs(5492) <= not (a xor b);
    layer2_outputs(5493) <= b and not a;
    layer2_outputs(5494) <= not (a xor b);
    layer2_outputs(5495) <= not b;
    layer2_outputs(5496) <= a and not b;
    layer2_outputs(5497) <= b and not a;
    layer2_outputs(5498) <= not b or a;
    layer2_outputs(5499) <= b;
    layer2_outputs(5500) <= not a;
    layer2_outputs(5501) <= not a;
    layer2_outputs(5502) <= a;
    layer2_outputs(5503) <= not (a and b);
    layer2_outputs(5504) <= not b;
    layer2_outputs(5505) <= not b;
    layer2_outputs(5506) <= not a or b;
    layer2_outputs(5507) <= not b or a;
    layer2_outputs(5508) <= not a or b;
    layer2_outputs(5509) <= a or b;
    layer2_outputs(5510) <= not (a and b);
    layer2_outputs(5511) <= not (a xor b);
    layer2_outputs(5512) <= a and not b;
    layer2_outputs(5513) <= not a;
    layer2_outputs(5514) <= not (a or b);
    layer2_outputs(5515) <= not (a xor b);
    layer2_outputs(5516) <= a and not b;
    layer2_outputs(5517) <= a;
    layer2_outputs(5518) <= not a;
    layer2_outputs(5519) <= '1';
    layer2_outputs(5520) <= a and not b;
    layer2_outputs(5521) <= b;
    layer2_outputs(5522) <= b and not a;
    layer2_outputs(5523) <= '1';
    layer2_outputs(5524) <= '1';
    layer2_outputs(5525) <= not (a or b);
    layer2_outputs(5526) <= not (a and b);
    layer2_outputs(5527) <= not (a and b);
    layer2_outputs(5528) <= b;
    layer2_outputs(5529) <= not a;
    layer2_outputs(5530) <= '0';
    layer2_outputs(5531) <= not b or a;
    layer2_outputs(5532) <= '1';
    layer2_outputs(5533) <= a and not b;
    layer2_outputs(5534) <= a xor b;
    layer2_outputs(5535) <= '1';
    layer2_outputs(5536) <= not b or a;
    layer2_outputs(5537) <= not (a or b);
    layer2_outputs(5538) <= '0';
    layer2_outputs(5539) <= a or b;
    layer2_outputs(5540) <= b and not a;
    layer2_outputs(5541) <= '1';
    layer2_outputs(5542) <= a and b;
    layer2_outputs(5543) <= not b;
    layer2_outputs(5544) <= a and b;
    layer2_outputs(5545) <= not (a or b);
    layer2_outputs(5546) <= b;
    layer2_outputs(5547) <= a and not b;
    layer2_outputs(5548) <= a;
    layer2_outputs(5549) <= not (a xor b);
    layer2_outputs(5550) <= not a or b;
    layer2_outputs(5551) <= a and b;
    layer2_outputs(5552) <= '1';
    layer2_outputs(5553) <= a;
    layer2_outputs(5554) <= a or b;
    layer2_outputs(5555) <= not b or a;
    layer2_outputs(5556) <= not a or b;
    layer2_outputs(5557) <= not a;
    layer2_outputs(5558) <= not a;
    layer2_outputs(5559) <= b and not a;
    layer2_outputs(5560) <= not b;
    layer2_outputs(5561) <= not (a or b);
    layer2_outputs(5562) <= b;
    layer2_outputs(5563) <= a or b;
    layer2_outputs(5564) <= not a or b;
    layer2_outputs(5565) <= not (a or b);
    layer2_outputs(5566) <= not b;
    layer2_outputs(5567) <= '1';
    layer2_outputs(5568) <= not b;
    layer2_outputs(5569) <= not (a or b);
    layer2_outputs(5570) <= not a or b;
    layer2_outputs(5571) <= not (a and b);
    layer2_outputs(5572) <= b;
    layer2_outputs(5573) <= b and not a;
    layer2_outputs(5574) <= a;
    layer2_outputs(5575) <= '1';
    layer2_outputs(5576) <= b;
    layer2_outputs(5577) <= a and b;
    layer2_outputs(5578) <= a;
    layer2_outputs(5579) <= b;
    layer2_outputs(5580) <= a and b;
    layer2_outputs(5581) <= not (a or b);
    layer2_outputs(5582) <= not a;
    layer2_outputs(5583) <= a and b;
    layer2_outputs(5584) <= not b;
    layer2_outputs(5585) <= not (a and b);
    layer2_outputs(5586) <= a;
    layer2_outputs(5587) <= a or b;
    layer2_outputs(5588) <= a and b;
    layer2_outputs(5589) <= a;
    layer2_outputs(5590) <= not (a and b);
    layer2_outputs(5591) <= b and not a;
    layer2_outputs(5592) <= a and not b;
    layer2_outputs(5593) <= not (a xor b);
    layer2_outputs(5594) <= a;
    layer2_outputs(5595) <= not b;
    layer2_outputs(5596) <= not (a xor b);
    layer2_outputs(5597) <= not (a and b);
    layer2_outputs(5598) <= '1';
    layer2_outputs(5599) <= not a or b;
    layer2_outputs(5600) <= a and not b;
    layer2_outputs(5601) <= not a;
    layer2_outputs(5602) <= a or b;
    layer2_outputs(5603) <= b;
    layer2_outputs(5604) <= not a or b;
    layer2_outputs(5605) <= a xor b;
    layer2_outputs(5606) <= not b;
    layer2_outputs(5607) <= a and b;
    layer2_outputs(5608) <= not a or b;
    layer2_outputs(5609) <= not a;
    layer2_outputs(5610) <= not a or b;
    layer2_outputs(5611) <= not a or b;
    layer2_outputs(5612) <= '1';
    layer2_outputs(5613) <= a xor b;
    layer2_outputs(5614) <= a;
    layer2_outputs(5615) <= a and not b;
    layer2_outputs(5616) <= not b;
    layer2_outputs(5617) <= b;
    layer2_outputs(5618) <= a or b;
    layer2_outputs(5619) <= a and b;
    layer2_outputs(5620) <= not (a or b);
    layer2_outputs(5621) <= '0';
    layer2_outputs(5622) <= not b;
    layer2_outputs(5623) <= b;
    layer2_outputs(5624) <= a;
    layer2_outputs(5625) <= not (a xor b);
    layer2_outputs(5626) <= b and not a;
    layer2_outputs(5627) <= '0';
    layer2_outputs(5628) <= not b or a;
    layer2_outputs(5629) <= not a;
    layer2_outputs(5630) <= not b or a;
    layer2_outputs(5631) <= a xor b;
    layer2_outputs(5632) <= '1';
    layer2_outputs(5633) <= a and not b;
    layer2_outputs(5634) <= a and not b;
    layer2_outputs(5635) <= '0';
    layer2_outputs(5636) <= not (a and b);
    layer2_outputs(5637) <= a and not b;
    layer2_outputs(5638) <= a;
    layer2_outputs(5639) <= not b;
    layer2_outputs(5640) <= not a or b;
    layer2_outputs(5641) <= a or b;
    layer2_outputs(5642) <= not b;
    layer2_outputs(5643) <= b;
    layer2_outputs(5644) <= b and not a;
    layer2_outputs(5645) <= a;
    layer2_outputs(5646) <= a xor b;
    layer2_outputs(5647) <= not (a and b);
    layer2_outputs(5648) <= not a;
    layer2_outputs(5649) <= a and not b;
    layer2_outputs(5650) <= not b;
    layer2_outputs(5651) <= '0';
    layer2_outputs(5652) <= not a or b;
    layer2_outputs(5653) <= a and not b;
    layer2_outputs(5654) <= not a;
    layer2_outputs(5655) <= not b;
    layer2_outputs(5656) <= '0';
    layer2_outputs(5657) <= b;
    layer2_outputs(5658) <= not a;
    layer2_outputs(5659) <= a and b;
    layer2_outputs(5660) <= b;
    layer2_outputs(5661) <= not (a or b);
    layer2_outputs(5662) <= not a or b;
    layer2_outputs(5663) <= not b or a;
    layer2_outputs(5664) <= not b or a;
    layer2_outputs(5665) <= not (a or b);
    layer2_outputs(5666) <= not (a or b);
    layer2_outputs(5667) <= not a;
    layer2_outputs(5668) <= a and not b;
    layer2_outputs(5669) <= not a;
    layer2_outputs(5670) <= a and b;
    layer2_outputs(5671) <= not (a or b);
    layer2_outputs(5672) <= a and b;
    layer2_outputs(5673) <= a or b;
    layer2_outputs(5674) <= not a or b;
    layer2_outputs(5675) <= not a;
    layer2_outputs(5676) <= a or b;
    layer2_outputs(5677) <= b;
    layer2_outputs(5678) <= a or b;
    layer2_outputs(5679) <= '0';
    layer2_outputs(5680) <= not (a xor b);
    layer2_outputs(5681) <= not (a or b);
    layer2_outputs(5682) <= a;
    layer2_outputs(5683) <= not a;
    layer2_outputs(5684) <= not a;
    layer2_outputs(5685) <= '0';
    layer2_outputs(5686) <= b and not a;
    layer2_outputs(5687) <= a or b;
    layer2_outputs(5688) <= not b;
    layer2_outputs(5689) <= a and b;
    layer2_outputs(5690) <= '0';
    layer2_outputs(5691) <= a and not b;
    layer2_outputs(5692) <= a;
    layer2_outputs(5693) <= a and not b;
    layer2_outputs(5694) <= '0';
    layer2_outputs(5695) <= not a;
    layer2_outputs(5696) <= not b;
    layer2_outputs(5697) <= not b;
    layer2_outputs(5698) <= a and not b;
    layer2_outputs(5699) <= a xor b;
    layer2_outputs(5700) <= not b;
    layer2_outputs(5701) <= a and b;
    layer2_outputs(5702) <= not (a or b);
    layer2_outputs(5703) <= a and not b;
    layer2_outputs(5704) <= not (a and b);
    layer2_outputs(5705) <= '0';
    layer2_outputs(5706) <= a and b;
    layer2_outputs(5707) <= not b or a;
    layer2_outputs(5708) <= '1';
    layer2_outputs(5709) <= a xor b;
    layer2_outputs(5710) <= not a or b;
    layer2_outputs(5711) <= a or b;
    layer2_outputs(5712) <= a;
    layer2_outputs(5713) <= b and not a;
    layer2_outputs(5714) <= not b;
    layer2_outputs(5715) <= b;
    layer2_outputs(5716) <= b;
    layer2_outputs(5717) <= b;
    layer2_outputs(5718) <= b;
    layer2_outputs(5719) <= not b or a;
    layer2_outputs(5720) <= not a or b;
    layer2_outputs(5721) <= not b;
    layer2_outputs(5722) <= b and not a;
    layer2_outputs(5723) <= not a;
    layer2_outputs(5724) <= a xor b;
    layer2_outputs(5725) <= not a or b;
    layer2_outputs(5726) <= '0';
    layer2_outputs(5727) <= not b;
    layer2_outputs(5728) <= not a;
    layer2_outputs(5729) <= '1';
    layer2_outputs(5730) <= not b;
    layer2_outputs(5731) <= '1';
    layer2_outputs(5732) <= not b or a;
    layer2_outputs(5733) <= a and not b;
    layer2_outputs(5734) <= a or b;
    layer2_outputs(5735) <= a xor b;
    layer2_outputs(5736) <= not b or a;
    layer2_outputs(5737) <= not (a or b);
    layer2_outputs(5738) <= b;
    layer2_outputs(5739) <= b and not a;
    layer2_outputs(5740) <= b;
    layer2_outputs(5741) <= a and b;
    layer2_outputs(5742) <= not (a or b);
    layer2_outputs(5743) <= not a;
    layer2_outputs(5744) <= not (a and b);
    layer2_outputs(5745) <= not b;
    layer2_outputs(5746) <= not b or a;
    layer2_outputs(5747) <= not (a or b);
    layer2_outputs(5748) <= b and not a;
    layer2_outputs(5749) <= a and b;
    layer2_outputs(5750) <= not b;
    layer2_outputs(5751) <= '0';
    layer2_outputs(5752) <= not (a or b);
    layer2_outputs(5753) <= a and not b;
    layer2_outputs(5754) <= not a;
    layer2_outputs(5755) <= a;
    layer2_outputs(5756) <= a and not b;
    layer2_outputs(5757) <= a and not b;
    layer2_outputs(5758) <= not (a or b);
    layer2_outputs(5759) <= not (a and b);
    layer2_outputs(5760) <= not (a xor b);
    layer2_outputs(5761) <= not (a or b);
    layer2_outputs(5762) <= a and not b;
    layer2_outputs(5763) <= b;
    layer2_outputs(5764) <= a and not b;
    layer2_outputs(5765) <= not a;
    layer2_outputs(5766) <= '1';
    layer2_outputs(5767) <= a;
    layer2_outputs(5768) <= b;
    layer2_outputs(5769) <= not (a and b);
    layer2_outputs(5770) <= b;
    layer2_outputs(5771) <= not b;
    layer2_outputs(5772) <= not (a or b);
    layer2_outputs(5773) <= '0';
    layer2_outputs(5774) <= not a;
    layer2_outputs(5775) <= not (a or b);
    layer2_outputs(5776) <= a xor b;
    layer2_outputs(5777) <= not a;
    layer2_outputs(5778) <= '1';
    layer2_outputs(5779) <= not (a or b);
    layer2_outputs(5780) <= not (a and b);
    layer2_outputs(5781) <= not (a or b);
    layer2_outputs(5782) <= not a or b;
    layer2_outputs(5783) <= not a or b;
    layer2_outputs(5784) <= a;
    layer2_outputs(5785) <= not b or a;
    layer2_outputs(5786) <= a and b;
    layer2_outputs(5787) <= not (a and b);
    layer2_outputs(5788) <= a and not b;
    layer2_outputs(5789) <= not (a xor b);
    layer2_outputs(5790) <= not b;
    layer2_outputs(5791) <= a or b;
    layer2_outputs(5792) <= not a;
    layer2_outputs(5793) <= '0';
    layer2_outputs(5794) <= b;
    layer2_outputs(5795) <= b and not a;
    layer2_outputs(5796) <= '1';
    layer2_outputs(5797) <= not b or a;
    layer2_outputs(5798) <= not a;
    layer2_outputs(5799) <= b and not a;
    layer2_outputs(5800) <= not b or a;
    layer2_outputs(5801) <= not (a or b);
    layer2_outputs(5802) <= not (a xor b);
    layer2_outputs(5803) <= a xor b;
    layer2_outputs(5804) <= b and not a;
    layer2_outputs(5805) <= '1';
    layer2_outputs(5806) <= b and not a;
    layer2_outputs(5807) <= a;
    layer2_outputs(5808) <= a or b;
    layer2_outputs(5809) <= not a or b;
    layer2_outputs(5810) <= b;
    layer2_outputs(5811) <= a or b;
    layer2_outputs(5812) <= not (a xor b);
    layer2_outputs(5813) <= not a;
    layer2_outputs(5814) <= not b;
    layer2_outputs(5815) <= not a or b;
    layer2_outputs(5816) <= '0';
    layer2_outputs(5817) <= not a;
    layer2_outputs(5818) <= not (a xor b);
    layer2_outputs(5819) <= a or b;
    layer2_outputs(5820) <= not b;
    layer2_outputs(5821) <= a and b;
    layer2_outputs(5822) <= not b;
    layer2_outputs(5823) <= not b or a;
    layer2_outputs(5824) <= not (a or b);
    layer2_outputs(5825) <= a xor b;
    layer2_outputs(5826) <= not a;
    layer2_outputs(5827) <= not (a and b);
    layer2_outputs(5828) <= not b or a;
    layer2_outputs(5829) <= a;
    layer2_outputs(5830) <= a and not b;
    layer2_outputs(5831) <= not a;
    layer2_outputs(5832) <= not (a or b);
    layer2_outputs(5833) <= not (a xor b);
    layer2_outputs(5834) <= a or b;
    layer2_outputs(5835) <= not a;
    layer2_outputs(5836) <= not (a or b);
    layer2_outputs(5837) <= not b;
    layer2_outputs(5838) <= not (a and b);
    layer2_outputs(5839) <= not (a or b);
    layer2_outputs(5840) <= a or b;
    layer2_outputs(5841) <= not (a xor b);
    layer2_outputs(5842) <= b;
    layer2_outputs(5843) <= b;
    layer2_outputs(5844) <= not (a xor b);
    layer2_outputs(5845) <= a;
    layer2_outputs(5846) <= not a;
    layer2_outputs(5847) <= a and not b;
    layer2_outputs(5848) <= not (a and b);
    layer2_outputs(5849) <= not (a and b);
    layer2_outputs(5850) <= b;
    layer2_outputs(5851) <= not b;
    layer2_outputs(5852) <= b and not a;
    layer2_outputs(5853) <= b;
    layer2_outputs(5854) <= b;
    layer2_outputs(5855) <= a or b;
    layer2_outputs(5856) <= a and b;
    layer2_outputs(5857) <= not a;
    layer2_outputs(5858) <= not b;
    layer2_outputs(5859) <= not (a and b);
    layer2_outputs(5860) <= '1';
    layer2_outputs(5861) <= a;
    layer2_outputs(5862) <= not b or a;
    layer2_outputs(5863) <= a or b;
    layer2_outputs(5864) <= a or b;
    layer2_outputs(5865) <= '0';
    layer2_outputs(5866) <= not a or b;
    layer2_outputs(5867) <= not (a or b);
    layer2_outputs(5868) <= not a;
    layer2_outputs(5869) <= not a or b;
    layer2_outputs(5870) <= a and b;
    layer2_outputs(5871) <= a;
    layer2_outputs(5872) <= a and not b;
    layer2_outputs(5873) <= not a;
    layer2_outputs(5874) <= not b or a;
    layer2_outputs(5875) <= a and not b;
    layer2_outputs(5876) <= not a or b;
    layer2_outputs(5877) <= b;
    layer2_outputs(5878) <= b and not a;
    layer2_outputs(5879) <= a and not b;
    layer2_outputs(5880) <= not b or a;
    layer2_outputs(5881) <= not b or a;
    layer2_outputs(5882) <= a or b;
    layer2_outputs(5883) <= a;
    layer2_outputs(5884) <= a and not b;
    layer2_outputs(5885) <= not (a or b);
    layer2_outputs(5886) <= b;
    layer2_outputs(5887) <= a and b;
    layer2_outputs(5888) <= not b;
    layer2_outputs(5889) <= b and not a;
    layer2_outputs(5890) <= not b;
    layer2_outputs(5891) <= a and b;
    layer2_outputs(5892) <= a xor b;
    layer2_outputs(5893) <= not b or a;
    layer2_outputs(5894) <= not a;
    layer2_outputs(5895) <= not a;
    layer2_outputs(5896) <= not a;
    layer2_outputs(5897) <= '0';
    layer2_outputs(5898) <= a and not b;
    layer2_outputs(5899) <= '1';
    layer2_outputs(5900) <= not a;
    layer2_outputs(5901) <= a xor b;
    layer2_outputs(5902) <= a and not b;
    layer2_outputs(5903) <= not b or a;
    layer2_outputs(5904) <= not (a xor b);
    layer2_outputs(5905) <= '1';
    layer2_outputs(5906) <= b;
    layer2_outputs(5907) <= not b;
    layer2_outputs(5908) <= '1';
    layer2_outputs(5909) <= b;
    layer2_outputs(5910) <= b;
    layer2_outputs(5911) <= a xor b;
    layer2_outputs(5912) <= not (a xor b);
    layer2_outputs(5913) <= not a;
    layer2_outputs(5914) <= not a;
    layer2_outputs(5915) <= b;
    layer2_outputs(5916) <= '0';
    layer2_outputs(5917) <= a;
    layer2_outputs(5918) <= not (a and b);
    layer2_outputs(5919) <= not (a and b);
    layer2_outputs(5920) <= not (a xor b);
    layer2_outputs(5921) <= a xor b;
    layer2_outputs(5922) <= not a or b;
    layer2_outputs(5923) <= b and not a;
    layer2_outputs(5924) <= a;
    layer2_outputs(5925) <= not b;
    layer2_outputs(5926) <= b;
    layer2_outputs(5927) <= not (a and b);
    layer2_outputs(5928) <= not a;
    layer2_outputs(5929) <= not b;
    layer2_outputs(5930) <= not (a and b);
    layer2_outputs(5931) <= '0';
    layer2_outputs(5932) <= not (a and b);
    layer2_outputs(5933) <= not (a and b);
    layer2_outputs(5934) <= b and not a;
    layer2_outputs(5935) <= not (a xor b);
    layer2_outputs(5936) <= not (a and b);
    layer2_outputs(5937) <= a;
    layer2_outputs(5938) <= a and b;
    layer2_outputs(5939) <= '0';
    layer2_outputs(5940) <= not b;
    layer2_outputs(5941) <= a xor b;
    layer2_outputs(5942) <= not a;
    layer2_outputs(5943) <= not a;
    layer2_outputs(5944) <= not a or b;
    layer2_outputs(5945) <= a and not b;
    layer2_outputs(5946) <= a or b;
    layer2_outputs(5947) <= not a or b;
    layer2_outputs(5948) <= '1';
    layer2_outputs(5949) <= b and not a;
    layer2_outputs(5950) <= a and not b;
    layer2_outputs(5951) <= not (a or b);
    layer2_outputs(5952) <= b;
    layer2_outputs(5953) <= '1';
    layer2_outputs(5954) <= '1';
    layer2_outputs(5955) <= not b or a;
    layer2_outputs(5956) <= a and not b;
    layer2_outputs(5957) <= a and not b;
    layer2_outputs(5958) <= '1';
    layer2_outputs(5959) <= not b;
    layer2_outputs(5960) <= not b;
    layer2_outputs(5961) <= not a;
    layer2_outputs(5962) <= not (a or b);
    layer2_outputs(5963) <= '0';
    layer2_outputs(5964) <= a;
    layer2_outputs(5965) <= b;
    layer2_outputs(5966) <= not b;
    layer2_outputs(5967) <= a;
    layer2_outputs(5968) <= a;
    layer2_outputs(5969) <= a and b;
    layer2_outputs(5970) <= not b;
    layer2_outputs(5971) <= b;
    layer2_outputs(5972) <= a or b;
    layer2_outputs(5973) <= not a;
    layer2_outputs(5974) <= not (a and b);
    layer2_outputs(5975) <= '1';
    layer2_outputs(5976) <= a;
    layer2_outputs(5977) <= '0';
    layer2_outputs(5978) <= a or b;
    layer2_outputs(5979) <= '0';
    layer2_outputs(5980) <= '0';
    layer2_outputs(5981) <= not a;
    layer2_outputs(5982) <= not (a and b);
    layer2_outputs(5983) <= not b;
    layer2_outputs(5984) <= not (a or b);
    layer2_outputs(5985) <= a and not b;
    layer2_outputs(5986) <= a and not b;
    layer2_outputs(5987) <= a and b;
    layer2_outputs(5988) <= not a or b;
    layer2_outputs(5989) <= a and b;
    layer2_outputs(5990) <= not (a xor b);
    layer2_outputs(5991) <= a or b;
    layer2_outputs(5992) <= a and b;
    layer2_outputs(5993) <= a;
    layer2_outputs(5994) <= b;
    layer2_outputs(5995) <= not b;
    layer2_outputs(5996) <= b;
    layer2_outputs(5997) <= b;
    layer2_outputs(5998) <= a;
    layer2_outputs(5999) <= not (a and b);
    layer2_outputs(6000) <= b and not a;
    layer2_outputs(6001) <= not a;
    layer2_outputs(6002) <= a or b;
    layer2_outputs(6003) <= a and b;
    layer2_outputs(6004) <= not (a and b);
    layer2_outputs(6005) <= not a or b;
    layer2_outputs(6006) <= b;
    layer2_outputs(6007) <= b;
    layer2_outputs(6008) <= not (a and b);
    layer2_outputs(6009) <= b;
    layer2_outputs(6010) <= not a or b;
    layer2_outputs(6011) <= a;
    layer2_outputs(6012) <= not (a or b);
    layer2_outputs(6013) <= '0';
    layer2_outputs(6014) <= b;
    layer2_outputs(6015) <= b;
    layer2_outputs(6016) <= b;
    layer2_outputs(6017) <= not (a or b);
    layer2_outputs(6018) <= not b;
    layer2_outputs(6019) <= a and b;
    layer2_outputs(6020) <= not b;
    layer2_outputs(6021) <= not (a and b);
    layer2_outputs(6022) <= a and b;
    layer2_outputs(6023) <= a;
    layer2_outputs(6024) <= b and not a;
    layer2_outputs(6025) <= not b or a;
    layer2_outputs(6026) <= a and b;
    layer2_outputs(6027) <= '0';
    layer2_outputs(6028) <= not a;
    layer2_outputs(6029) <= b;
    layer2_outputs(6030) <= not b;
    layer2_outputs(6031) <= '0';
    layer2_outputs(6032) <= '0';
    layer2_outputs(6033) <= not b;
    layer2_outputs(6034) <= a and b;
    layer2_outputs(6035) <= b;
    layer2_outputs(6036) <= not (a and b);
    layer2_outputs(6037) <= b;
    layer2_outputs(6038) <= a and not b;
    layer2_outputs(6039) <= not (a xor b);
    layer2_outputs(6040) <= not a;
    layer2_outputs(6041) <= not a;
    layer2_outputs(6042) <= a and not b;
    layer2_outputs(6043) <= not b;
    layer2_outputs(6044) <= not a or b;
    layer2_outputs(6045) <= not b;
    layer2_outputs(6046) <= '0';
    layer2_outputs(6047) <= a and not b;
    layer2_outputs(6048) <= a or b;
    layer2_outputs(6049) <= not b;
    layer2_outputs(6050) <= not a;
    layer2_outputs(6051) <= not (a or b);
    layer2_outputs(6052) <= '0';
    layer2_outputs(6053) <= not a or b;
    layer2_outputs(6054) <= a and b;
    layer2_outputs(6055) <= b;
    layer2_outputs(6056) <= b;
    layer2_outputs(6057) <= '0';
    layer2_outputs(6058) <= not (a and b);
    layer2_outputs(6059) <= not b;
    layer2_outputs(6060) <= a xor b;
    layer2_outputs(6061) <= not (a or b);
    layer2_outputs(6062) <= not b;
    layer2_outputs(6063) <= not a;
    layer2_outputs(6064) <= '1';
    layer2_outputs(6065) <= not b;
    layer2_outputs(6066) <= '0';
    layer2_outputs(6067) <= '0';
    layer2_outputs(6068) <= not a;
    layer2_outputs(6069) <= a or b;
    layer2_outputs(6070) <= not a;
    layer2_outputs(6071) <= b;
    layer2_outputs(6072) <= a;
    layer2_outputs(6073) <= not a or b;
    layer2_outputs(6074) <= not b;
    layer2_outputs(6075) <= not (a or b);
    layer2_outputs(6076) <= '0';
    layer2_outputs(6077) <= a;
    layer2_outputs(6078) <= '1';
    layer2_outputs(6079) <= a;
    layer2_outputs(6080) <= '1';
    layer2_outputs(6081) <= a and b;
    layer2_outputs(6082) <= '0';
    layer2_outputs(6083) <= not b or a;
    layer2_outputs(6084) <= '1';
    layer2_outputs(6085) <= '1';
    layer2_outputs(6086) <= not (a or b);
    layer2_outputs(6087) <= not a;
    layer2_outputs(6088) <= b and not a;
    layer2_outputs(6089) <= not b;
    layer2_outputs(6090) <= not b;
    layer2_outputs(6091) <= b and not a;
    layer2_outputs(6092) <= not (a and b);
    layer2_outputs(6093) <= a;
    layer2_outputs(6094) <= b;
    layer2_outputs(6095) <= a and b;
    layer2_outputs(6096) <= b;
    layer2_outputs(6097) <= not a;
    layer2_outputs(6098) <= not (a or b);
    layer2_outputs(6099) <= not a;
    layer2_outputs(6100) <= b;
    layer2_outputs(6101) <= a and b;
    layer2_outputs(6102) <= not b or a;
    layer2_outputs(6103) <= a and b;
    layer2_outputs(6104) <= b and not a;
    layer2_outputs(6105) <= not b or a;
    layer2_outputs(6106) <= not (a or b);
    layer2_outputs(6107) <= a or b;
    layer2_outputs(6108) <= not (a or b);
    layer2_outputs(6109) <= a or b;
    layer2_outputs(6110) <= not (a or b);
    layer2_outputs(6111) <= a xor b;
    layer2_outputs(6112) <= not (a or b);
    layer2_outputs(6113) <= a or b;
    layer2_outputs(6114) <= a;
    layer2_outputs(6115) <= a;
    layer2_outputs(6116) <= not (a xor b);
    layer2_outputs(6117) <= a;
    layer2_outputs(6118) <= b and not a;
    layer2_outputs(6119) <= a and not b;
    layer2_outputs(6120) <= not a or b;
    layer2_outputs(6121) <= a;
    layer2_outputs(6122) <= not b;
    layer2_outputs(6123) <= b;
    layer2_outputs(6124) <= '0';
    layer2_outputs(6125) <= b and not a;
    layer2_outputs(6126) <= not a;
    layer2_outputs(6127) <= '1';
    layer2_outputs(6128) <= '1';
    layer2_outputs(6129) <= not b or a;
    layer2_outputs(6130) <= not b or a;
    layer2_outputs(6131) <= b and not a;
    layer2_outputs(6132) <= not a or b;
    layer2_outputs(6133) <= not (a xor b);
    layer2_outputs(6134) <= '0';
    layer2_outputs(6135) <= a xor b;
    layer2_outputs(6136) <= b;
    layer2_outputs(6137) <= not a;
    layer2_outputs(6138) <= not a or b;
    layer2_outputs(6139) <= b;
    layer2_outputs(6140) <= a xor b;
    layer2_outputs(6141) <= a or b;
    layer2_outputs(6142) <= a and b;
    layer2_outputs(6143) <= not a;
    layer2_outputs(6144) <= '0';
    layer2_outputs(6145) <= a and not b;
    layer2_outputs(6146) <= '1';
    layer2_outputs(6147) <= a or b;
    layer2_outputs(6148) <= not a;
    layer2_outputs(6149) <= not (a xor b);
    layer2_outputs(6150) <= a or b;
    layer2_outputs(6151) <= not (a and b);
    layer2_outputs(6152) <= not a or b;
    layer2_outputs(6153) <= not b;
    layer2_outputs(6154) <= not a;
    layer2_outputs(6155) <= '0';
    layer2_outputs(6156) <= a and b;
    layer2_outputs(6157) <= not a or b;
    layer2_outputs(6158) <= not a or b;
    layer2_outputs(6159) <= a or b;
    layer2_outputs(6160) <= not b;
    layer2_outputs(6161) <= '0';
    layer2_outputs(6162) <= a and b;
    layer2_outputs(6163) <= a and not b;
    layer2_outputs(6164) <= '0';
    layer2_outputs(6165) <= b;
    layer2_outputs(6166) <= not b;
    layer2_outputs(6167) <= b;
    layer2_outputs(6168) <= '1';
    layer2_outputs(6169) <= a and not b;
    layer2_outputs(6170) <= b and not a;
    layer2_outputs(6171) <= a or b;
    layer2_outputs(6172) <= not (a and b);
    layer2_outputs(6173) <= a or b;
    layer2_outputs(6174) <= a or b;
    layer2_outputs(6175) <= not a;
    layer2_outputs(6176) <= a xor b;
    layer2_outputs(6177) <= not a;
    layer2_outputs(6178) <= '0';
    layer2_outputs(6179) <= a and not b;
    layer2_outputs(6180) <= a and b;
    layer2_outputs(6181) <= b;
    layer2_outputs(6182) <= a;
    layer2_outputs(6183) <= not (a and b);
    layer2_outputs(6184) <= a and b;
    layer2_outputs(6185) <= b;
    layer2_outputs(6186) <= b;
    layer2_outputs(6187) <= a or b;
    layer2_outputs(6188) <= b;
    layer2_outputs(6189) <= a xor b;
    layer2_outputs(6190) <= b;
    layer2_outputs(6191) <= not (a and b);
    layer2_outputs(6192) <= a;
    layer2_outputs(6193) <= not b;
    layer2_outputs(6194) <= a and b;
    layer2_outputs(6195) <= not (a and b);
    layer2_outputs(6196) <= not b or a;
    layer2_outputs(6197) <= not a;
    layer2_outputs(6198) <= not (a xor b);
    layer2_outputs(6199) <= not (a and b);
    layer2_outputs(6200) <= '1';
    layer2_outputs(6201) <= not b or a;
    layer2_outputs(6202) <= not a or b;
    layer2_outputs(6203) <= b and not a;
    layer2_outputs(6204) <= '0';
    layer2_outputs(6205) <= b and not a;
    layer2_outputs(6206) <= not a or b;
    layer2_outputs(6207) <= a and not b;
    layer2_outputs(6208) <= b and not a;
    layer2_outputs(6209) <= a and not b;
    layer2_outputs(6210) <= a or b;
    layer2_outputs(6211) <= not (a or b);
    layer2_outputs(6212) <= b;
    layer2_outputs(6213) <= not (a xor b);
    layer2_outputs(6214) <= a xor b;
    layer2_outputs(6215) <= not a;
    layer2_outputs(6216) <= a and b;
    layer2_outputs(6217) <= not b;
    layer2_outputs(6218) <= '0';
    layer2_outputs(6219) <= a;
    layer2_outputs(6220) <= not b;
    layer2_outputs(6221) <= b and not a;
    layer2_outputs(6222) <= not (a and b);
    layer2_outputs(6223) <= not b;
    layer2_outputs(6224) <= not a or b;
    layer2_outputs(6225) <= a and b;
    layer2_outputs(6226) <= b and not a;
    layer2_outputs(6227) <= a;
    layer2_outputs(6228) <= b and not a;
    layer2_outputs(6229) <= '0';
    layer2_outputs(6230) <= b;
    layer2_outputs(6231) <= a;
    layer2_outputs(6232) <= not (a or b);
    layer2_outputs(6233) <= a and b;
    layer2_outputs(6234) <= a;
    layer2_outputs(6235) <= not (a and b);
    layer2_outputs(6236) <= a;
    layer2_outputs(6237) <= not b or a;
    layer2_outputs(6238) <= not (a or b);
    layer2_outputs(6239) <= not b;
    layer2_outputs(6240) <= a and b;
    layer2_outputs(6241) <= not b;
    layer2_outputs(6242) <= not b;
    layer2_outputs(6243) <= a;
    layer2_outputs(6244) <= a and not b;
    layer2_outputs(6245) <= '1';
    layer2_outputs(6246) <= not a or b;
    layer2_outputs(6247) <= not (a xor b);
    layer2_outputs(6248) <= not (a and b);
    layer2_outputs(6249) <= a xor b;
    layer2_outputs(6250) <= not (a and b);
    layer2_outputs(6251) <= a or b;
    layer2_outputs(6252) <= a;
    layer2_outputs(6253) <= '1';
    layer2_outputs(6254) <= b and not a;
    layer2_outputs(6255) <= '0';
    layer2_outputs(6256) <= a;
    layer2_outputs(6257) <= not b or a;
    layer2_outputs(6258) <= a or b;
    layer2_outputs(6259) <= a xor b;
    layer2_outputs(6260) <= not b;
    layer2_outputs(6261) <= b;
    layer2_outputs(6262) <= a;
    layer2_outputs(6263) <= b and not a;
    layer2_outputs(6264) <= a and not b;
    layer2_outputs(6265) <= not (a or b);
    layer2_outputs(6266) <= not b;
    layer2_outputs(6267) <= not a;
    layer2_outputs(6268) <= a xor b;
    layer2_outputs(6269) <= not b;
    layer2_outputs(6270) <= a;
    layer2_outputs(6271) <= '1';
    layer2_outputs(6272) <= not b;
    layer2_outputs(6273) <= b and not a;
    layer2_outputs(6274) <= not a or b;
    layer2_outputs(6275) <= not a;
    layer2_outputs(6276) <= '1';
    layer2_outputs(6277) <= a;
    layer2_outputs(6278) <= b;
    layer2_outputs(6279) <= not a;
    layer2_outputs(6280) <= '0';
    layer2_outputs(6281) <= not b or a;
    layer2_outputs(6282) <= not (a and b);
    layer2_outputs(6283) <= a and b;
    layer2_outputs(6284) <= not (a and b);
    layer2_outputs(6285) <= a;
    layer2_outputs(6286) <= not (a and b);
    layer2_outputs(6287) <= a or b;
    layer2_outputs(6288) <= not a;
    layer2_outputs(6289) <= not b or a;
    layer2_outputs(6290) <= a and b;
    layer2_outputs(6291) <= not b or a;
    layer2_outputs(6292) <= '1';
    layer2_outputs(6293) <= '1';
    layer2_outputs(6294) <= not a or b;
    layer2_outputs(6295) <= '0';
    layer2_outputs(6296) <= b;
    layer2_outputs(6297) <= '1';
    layer2_outputs(6298) <= not b or a;
    layer2_outputs(6299) <= not (a and b);
    layer2_outputs(6300) <= not (a and b);
    layer2_outputs(6301) <= not a or b;
    layer2_outputs(6302) <= not b or a;
    layer2_outputs(6303) <= not b;
    layer2_outputs(6304) <= not a;
    layer2_outputs(6305) <= b;
    layer2_outputs(6306) <= b and not a;
    layer2_outputs(6307) <= a;
    layer2_outputs(6308) <= a and not b;
    layer2_outputs(6309) <= a;
    layer2_outputs(6310) <= not (a and b);
    layer2_outputs(6311) <= '1';
    layer2_outputs(6312) <= a and b;
    layer2_outputs(6313) <= a and b;
    layer2_outputs(6314) <= not a or b;
    layer2_outputs(6315) <= not a;
    layer2_outputs(6316) <= b;
    layer2_outputs(6317) <= b;
    layer2_outputs(6318) <= a and b;
    layer2_outputs(6319) <= not b or a;
    layer2_outputs(6320) <= a or b;
    layer2_outputs(6321) <= b and not a;
    layer2_outputs(6322) <= not b or a;
    layer2_outputs(6323) <= a;
    layer2_outputs(6324) <= b and not a;
    layer2_outputs(6325) <= not a or b;
    layer2_outputs(6326) <= a and b;
    layer2_outputs(6327) <= b and not a;
    layer2_outputs(6328) <= not (a and b);
    layer2_outputs(6329) <= a;
    layer2_outputs(6330) <= b;
    layer2_outputs(6331) <= '0';
    layer2_outputs(6332) <= b;
    layer2_outputs(6333) <= not (a xor b);
    layer2_outputs(6334) <= not a;
    layer2_outputs(6335) <= a and b;
    layer2_outputs(6336) <= not a or b;
    layer2_outputs(6337) <= a;
    layer2_outputs(6338) <= not a;
    layer2_outputs(6339) <= a and not b;
    layer2_outputs(6340) <= not a;
    layer2_outputs(6341) <= not b or a;
    layer2_outputs(6342) <= b;
    layer2_outputs(6343) <= b and not a;
    layer2_outputs(6344) <= not a or b;
    layer2_outputs(6345) <= not b;
    layer2_outputs(6346) <= '1';
    layer2_outputs(6347) <= b;
    layer2_outputs(6348) <= a and b;
    layer2_outputs(6349) <= a and b;
    layer2_outputs(6350) <= not b;
    layer2_outputs(6351) <= b;
    layer2_outputs(6352) <= a;
    layer2_outputs(6353) <= not a or b;
    layer2_outputs(6354) <= '1';
    layer2_outputs(6355) <= not b or a;
    layer2_outputs(6356) <= a or b;
    layer2_outputs(6357) <= a;
    layer2_outputs(6358) <= not b;
    layer2_outputs(6359) <= not a or b;
    layer2_outputs(6360) <= not b;
    layer2_outputs(6361) <= b and not a;
    layer2_outputs(6362) <= a;
    layer2_outputs(6363) <= not b or a;
    layer2_outputs(6364) <= a and b;
    layer2_outputs(6365) <= a or b;
    layer2_outputs(6366) <= a and b;
    layer2_outputs(6367) <= b and not a;
    layer2_outputs(6368) <= '1';
    layer2_outputs(6369) <= not a;
    layer2_outputs(6370) <= '1';
    layer2_outputs(6371) <= not (a xor b);
    layer2_outputs(6372) <= not a;
    layer2_outputs(6373) <= not (a xor b);
    layer2_outputs(6374) <= not a or b;
    layer2_outputs(6375) <= not (a and b);
    layer2_outputs(6376) <= a or b;
    layer2_outputs(6377) <= a and b;
    layer2_outputs(6378) <= b and not a;
    layer2_outputs(6379) <= not a;
    layer2_outputs(6380) <= a xor b;
    layer2_outputs(6381) <= '1';
    layer2_outputs(6382) <= not (a and b);
    layer2_outputs(6383) <= not a;
    layer2_outputs(6384) <= not b;
    layer2_outputs(6385) <= not (a or b);
    layer2_outputs(6386) <= a and b;
    layer2_outputs(6387) <= a and b;
    layer2_outputs(6388) <= a and not b;
    layer2_outputs(6389) <= not b;
    layer2_outputs(6390) <= a;
    layer2_outputs(6391) <= '0';
    layer2_outputs(6392) <= not (a xor b);
    layer2_outputs(6393) <= not b;
    layer2_outputs(6394) <= '0';
    layer2_outputs(6395) <= a or b;
    layer2_outputs(6396) <= not a;
    layer2_outputs(6397) <= not (a xor b);
    layer2_outputs(6398) <= not b or a;
    layer2_outputs(6399) <= a or b;
    layer2_outputs(6400) <= not b or a;
    layer2_outputs(6401) <= a and b;
    layer2_outputs(6402) <= b and not a;
    layer2_outputs(6403) <= not a;
    layer2_outputs(6404) <= not (a and b);
    layer2_outputs(6405) <= a or b;
    layer2_outputs(6406) <= a and not b;
    layer2_outputs(6407) <= b and not a;
    layer2_outputs(6408) <= b;
    layer2_outputs(6409) <= not (a or b);
    layer2_outputs(6410) <= not (a and b);
    layer2_outputs(6411) <= a xor b;
    layer2_outputs(6412) <= not b or a;
    layer2_outputs(6413) <= b;
    layer2_outputs(6414) <= b and not a;
    layer2_outputs(6415) <= not (a or b);
    layer2_outputs(6416) <= not (a or b);
    layer2_outputs(6417) <= not b;
    layer2_outputs(6418) <= not (a and b);
    layer2_outputs(6419) <= a or b;
    layer2_outputs(6420) <= '0';
    layer2_outputs(6421) <= b and not a;
    layer2_outputs(6422) <= not b;
    layer2_outputs(6423) <= not b;
    layer2_outputs(6424) <= not (a xor b);
    layer2_outputs(6425) <= a or b;
    layer2_outputs(6426) <= not (a xor b);
    layer2_outputs(6427) <= not (a and b);
    layer2_outputs(6428) <= not b;
    layer2_outputs(6429) <= b;
    layer2_outputs(6430) <= not (a and b);
    layer2_outputs(6431) <= b;
    layer2_outputs(6432) <= b;
    layer2_outputs(6433) <= not a;
    layer2_outputs(6434) <= not b or a;
    layer2_outputs(6435) <= b;
    layer2_outputs(6436) <= a and b;
    layer2_outputs(6437) <= not b or a;
    layer2_outputs(6438) <= not b;
    layer2_outputs(6439) <= a and b;
    layer2_outputs(6440) <= not (a or b);
    layer2_outputs(6441) <= a;
    layer2_outputs(6442) <= not b or a;
    layer2_outputs(6443) <= a and not b;
    layer2_outputs(6444) <= b;
    layer2_outputs(6445) <= not (a or b);
    layer2_outputs(6446) <= a and not b;
    layer2_outputs(6447) <= a and b;
    layer2_outputs(6448) <= b;
    layer2_outputs(6449) <= not (a and b);
    layer2_outputs(6450) <= not b;
    layer2_outputs(6451) <= '1';
    layer2_outputs(6452) <= not (a or b);
    layer2_outputs(6453) <= not (a or b);
    layer2_outputs(6454) <= a and not b;
    layer2_outputs(6455) <= not a or b;
    layer2_outputs(6456) <= not b;
    layer2_outputs(6457) <= a xor b;
    layer2_outputs(6458) <= a xor b;
    layer2_outputs(6459) <= a and not b;
    layer2_outputs(6460) <= not (a and b);
    layer2_outputs(6461) <= b;
    layer2_outputs(6462) <= not a;
    layer2_outputs(6463) <= not b;
    layer2_outputs(6464) <= b and not a;
    layer2_outputs(6465) <= not a or b;
    layer2_outputs(6466) <= not b or a;
    layer2_outputs(6467) <= a and b;
    layer2_outputs(6468) <= a xor b;
    layer2_outputs(6469) <= not (a or b);
    layer2_outputs(6470) <= '1';
    layer2_outputs(6471) <= a and b;
    layer2_outputs(6472) <= b;
    layer2_outputs(6473) <= not b or a;
    layer2_outputs(6474) <= not b or a;
    layer2_outputs(6475) <= a or b;
    layer2_outputs(6476) <= not (a or b);
    layer2_outputs(6477) <= not b;
    layer2_outputs(6478) <= a or b;
    layer2_outputs(6479) <= '1';
    layer2_outputs(6480) <= b;
    layer2_outputs(6481) <= b;
    layer2_outputs(6482) <= a and b;
    layer2_outputs(6483) <= not (a or b);
    layer2_outputs(6484) <= not a or b;
    layer2_outputs(6485) <= b;
    layer2_outputs(6486) <= b;
    layer2_outputs(6487) <= not (a and b);
    layer2_outputs(6488) <= a and not b;
    layer2_outputs(6489) <= a or b;
    layer2_outputs(6490) <= a and b;
    layer2_outputs(6491) <= not b;
    layer2_outputs(6492) <= a or b;
    layer2_outputs(6493) <= a and b;
    layer2_outputs(6494) <= not (a or b);
    layer2_outputs(6495) <= a or b;
    layer2_outputs(6496) <= not (a or b);
    layer2_outputs(6497) <= b;
    layer2_outputs(6498) <= '0';
    layer2_outputs(6499) <= '1';
    layer2_outputs(6500) <= not a;
    layer2_outputs(6501) <= b and not a;
    layer2_outputs(6502) <= not (a or b);
    layer2_outputs(6503) <= a or b;
    layer2_outputs(6504) <= '1';
    layer2_outputs(6505) <= not b;
    layer2_outputs(6506) <= b and not a;
    layer2_outputs(6507) <= not (a and b);
    layer2_outputs(6508) <= not b or a;
    layer2_outputs(6509) <= a and b;
    layer2_outputs(6510) <= not a;
    layer2_outputs(6511) <= not (a or b);
    layer2_outputs(6512) <= '1';
    layer2_outputs(6513) <= not (a xor b);
    layer2_outputs(6514) <= a or b;
    layer2_outputs(6515) <= not a;
    layer2_outputs(6516) <= not a or b;
    layer2_outputs(6517) <= not (a or b);
    layer2_outputs(6518) <= not (a or b);
    layer2_outputs(6519) <= not a;
    layer2_outputs(6520) <= not b;
    layer2_outputs(6521) <= a and not b;
    layer2_outputs(6522) <= a or b;
    layer2_outputs(6523) <= '0';
    layer2_outputs(6524) <= b;
    layer2_outputs(6525) <= not a or b;
    layer2_outputs(6526) <= b;
    layer2_outputs(6527) <= a;
    layer2_outputs(6528) <= not b or a;
    layer2_outputs(6529) <= b and not a;
    layer2_outputs(6530) <= not b or a;
    layer2_outputs(6531) <= not (a and b);
    layer2_outputs(6532) <= '0';
    layer2_outputs(6533) <= a and not b;
    layer2_outputs(6534) <= not (a and b);
    layer2_outputs(6535) <= b;
    layer2_outputs(6536) <= a;
    layer2_outputs(6537) <= not a;
    layer2_outputs(6538) <= '0';
    layer2_outputs(6539) <= b and not a;
    layer2_outputs(6540) <= b and not a;
    layer2_outputs(6541) <= b;
    layer2_outputs(6542) <= not (a or b);
    layer2_outputs(6543) <= a or b;
    layer2_outputs(6544) <= not b;
    layer2_outputs(6545) <= b;
    layer2_outputs(6546) <= b;
    layer2_outputs(6547) <= a or b;
    layer2_outputs(6548) <= not b;
    layer2_outputs(6549) <= not (a and b);
    layer2_outputs(6550) <= not b or a;
    layer2_outputs(6551) <= a;
    layer2_outputs(6552) <= b and not a;
    layer2_outputs(6553) <= b;
    layer2_outputs(6554) <= not a;
    layer2_outputs(6555) <= a and b;
    layer2_outputs(6556) <= b;
    layer2_outputs(6557) <= not b;
    layer2_outputs(6558) <= not b;
    layer2_outputs(6559) <= a or b;
    layer2_outputs(6560) <= not b;
    layer2_outputs(6561) <= b and not a;
    layer2_outputs(6562) <= a and b;
    layer2_outputs(6563) <= a and not b;
    layer2_outputs(6564) <= not b;
    layer2_outputs(6565) <= '0';
    layer2_outputs(6566) <= a and b;
    layer2_outputs(6567) <= a and b;
    layer2_outputs(6568) <= not b;
    layer2_outputs(6569) <= a;
    layer2_outputs(6570) <= a or b;
    layer2_outputs(6571) <= not a;
    layer2_outputs(6572) <= a and b;
    layer2_outputs(6573) <= not a or b;
    layer2_outputs(6574) <= a and not b;
    layer2_outputs(6575) <= not (a xor b);
    layer2_outputs(6576) <= b;
    layer2_outputs(6577) <= a;
    layer2_outputs(6578) <= not (a or b);
    layer2_outputs(6579) <= not a or b;
    layer2_outputs(6580) <= not a or b;
    layer2_outputs(6581) <= not a;
    layer2_outputs(6582) <= a or b;
    layer2_outputs(6583) <= b;
    layer2_outputs(6584) <= not b;
    layer2_outputs(6585) <= not (a xor b);
    layer2_outputs(6586) <= a and not b;
    layer2_outputs(6587) <= not a or b;
    layer2_outputs(6588) <= not (a or b);
    layer2_outputs(6589) <= b;
    layer2_outputs(6590) <= a and b;
    layer2_outputs(6591) <= not a or b;
    layer2_outputs(6592) <= '0';
    layer2_outputs(6593) <= '1';
    layer2_outputs(6594) <= b and not a;
    layer2_outputs(6595) <= not b;
    layer2_outputs(6596) <= '0';
    layer2_outputs(6597) <= a xor b;
    layer2_outputs(6598) <= not b or a;
    layer2_outputs(6599) <= not a;
    layer2_outputs(6600) <= a and b;
    layer2_outputs(6601) <= b;
    layer2_outputs(6602) <= a and b;
    layer2_outputs(6603) <= not b;
    layer2_outputs(6604) <= not b or a;
    layer2_outputs(6605) <= not (a and b);
    layer2_outputs(6606) <= not (a xor b);
    layer2_outputs(6607) <= not (a or b);
    layer2_outputs(6608) <= a xor b;
    layer2_outputs(6609) <= a and not b;
    layer2_outputs(6610) <= not (a and b);
    layer2_outputs(6611) <= a;
    layer2_outputs(6612) <= not (a or b);
    layer2_outputs(6613) <= b and not a;
    layer2_outputs(6614) <= a or b;
    layer2_outputs(6615) <= not b or a;
    layer2_outputs(6616) <= not b;
    layer2_outputs(6617) <= not b or a;
    layer2_outputs(6618) <= a;
    layer2_outputs(6619) <= not a;
    layer2_outputs(6620) <= a and not b;
    layer2_outputs(6621) <= not b or a;
    layer2_outputs(6622) <= '1';
    layer2_outputs(6623) <= '1';
    layer2_outputs(6624) <= not (a or b);
    layer2_outputs(6625) <= not (a and b);
    layer2_outputs(6626) <= '0';
    layer2_outputs(6627) <= not (a and b);
    layer2_outputs(6628) <= a or b;
    layer2_outputs(6629) <= not a;
    layer2_outputs(6630) <= not (a or b);
    layer2_outputs(6631) <= b and not a;
    layer2_outputs(6632) <= not b or a;
    layer2_outputs(6633) <= a;
    layer2_outputs(6634) <= not (a and b);
    layer2_outputs(6635) <= a and b;
    layer2_outputs(6636) <= b;
    layer2_outputs(6637) <= '1';
    layer2_outputs(6638) <= a and not b;
    layer2_outputs(6639) <= b and not a;
    layer2_outputs(6640) <= not a;
    layer2_outputs(6641) <= a;
    layer2_outputs(6642) <= a and not b;
    layer2_outputs(6643) <= not b;
    layer2_outputs(6644) <= '1';
    layer2_outputs(6645) <= a xor b;
    layer2_outputs(6646) <= b and not a;
    layer2_outputs(6647) <= a xor b;
    layer2_outputs(6648) <= a xor b;
    layer2_outputs(6649) <= not b;
    layer2_outputs(6650) <= '0';
    layer2_outputs(6651) <= a or b;
    layer2_outputs(6652) <= not (a or b);
    layer2_outputs(6653) <= not (a xor b);
    layer2_outputs(6654) <= a and b;
    layer2_outputs(6655) <= not b;
    layer2_outputs(6656) <= a and not b;
    layer2_outputs(6657) <= not b;
    layer2_outputs(6658) <= '1';
    layer2_outputs(6659) <= a and b;
    layer2_outputs(6660) <= not (a or b);
    layer2_outputs(6661) <= not (a or b);
    layer2_outputs(6662) <= a;
    layer2_outputs(6663) <= a;
    layer2_outputs(6664) <= not (a and b);
    layer2_outputs(6665) <= b;
    layer2_outputs(6666) <= not (a and b);
    layer2_outputs(6667) <= b and not a;
    layer2_outputs(6668) <= a or b;
    layer2_outputs(6669) <= not a;
    layer2_outputs(6670) <= a and not b;
    layer2_outputs(6671) <= not a;
    layer2_outputs(6672) <= not b or a;
    layer2_outputs(6673) <= '1';
    layer2_outputs(6674) <= a or b;
    layer2_outputs(6675) <= a and not b;
    layer2_outputs(6676) <= b and not a;
    layer2_outputs(6677) <= not b;
    layer2_outputs(6678) <= not (a and b);
    layer2_outputs(6679) <= b;
    layer2_outputs(6680) <= not (a or b);
    layer2_outputs(6681) <= not b;
    layer2_outputs(6682) <= a xor b;
    layer2_outputs(6683) <= not b;
    layer2_outputs(6684) <= b and not a;
    layer2_outputs(6685) <= a and not b;
    layer2_outputs(6686) <= a and b;
    layer2_outputs(6687) <= not b;
    layer2_outputs(6688) <= not b;
    layer2_outputs(6689) <= not a;
    layer2_outputs(6690) <= not b;
    layer2_outputs(6691) <= b and not a;
    layer2_outputs(6692) <= a;
    layer2_outputs(6693) <= b;
    layer2_outputs(6694) <= a and b;
    layer2_outputs(6695) <= not b or a;
    layer2_outputs(6696) <= not b;
    layer2_outputs(6697) <= a or b;
    layer2_outputs(6698) <= b;
    layer2_outputs(6699) <= b;
    layer2_outputs(6700) <= '1';
    layer2_outputs(6701) <= not a;
    layer2_outputs(6702) <= not (a or b);
    layer2_outputs(6703) <= not a or b;
    layer2_outputs(6704) <= a and b;
    layer2_outputs(6705) <= a;
    layer2_outputs(6706) <= a xor b;
    layer2_outputs(6707) <= b and not a;
    layer2_outputs(6708) <= not a;
    layer2_outputs(6709) <= not a;
    layer2_outputs(6710) <= not b or a;
    layer2_outputs(6711) <= a or b;
    layer2_outputs(6712) <= b;
    layer2_outputs(6713) <= not b;
    layer2_outputs(6714) <= a and not b;
    layer2_outputs(6715) <= not a or b;
    layer2_outputs(6716) <= not a or b;
    layer2_outputs(6717) <= not b or a;
    layer2_outputs(6718) <= not (a and b);
    layer2_outputs(6719) <= not (a and b);
    layer2_outputs(6720) <= not b or a;
    layer2_outputs(6721) <= b and not a;
    layer2_outputs(6722) <= not a or b;
    layer2_outputs(6723) <= a xor b;
    layer2_outputs(6724) <= a and not b;
    layer2_outputs(6725) <= a and not b;
    layer2_outputs(6726) <= not (a or b);
    layer2_outputs(6727) <= a;
    layer2_outputs(6728) <= not (a xor b);
    layer2_outputs(6729) <= not a;
    layer2_outputs(6730) <= a xor b;
    layer2_outputs(6731) <= not a or b;
    layer2_outputs(6732) <= '0';
    layer2_outputs(6733) <= a and b;
    layer2_outputs(6734) <= a and not b;
    layer2_outputs(6735) <= a and not b;
    layer2_outputs(6736) <= not b or a;
    layer2_outputs(6737) <= a and b;
    layer2_outputs(6738) <= not (a or b);
    layer2_outputs(6739) <= not b or a;
    layer2_outputs(6740) <= a and b;
    layer2_outputs(6741) <= a;
    layer2_outputs(6742) <= not b or a;
    layer2_outputs(6743) <= not (a and b);
    layer2_outputs(6744) <= a and b;
    layer2_outputs(6745) <= not b or a;
    layer2_outputs(6746) <= a;
    layer2_outputs(6747) <= a and not b;
    layer2_outputs(6748) <= a;
    layer2_outputs(6749) <= b and not a;
    layer2_outputs(6750) <= not a;
    layer2_outputs(6751) <= a or b;
    layer2_outputs(6752) <= a or b;
    layer2_outputs(6753) <= not a;
    layer2_outputs(6754) <= a;
    layer2_outputs(6755) <= not a;
    layer2_outputs(6756) <= not b;
    layer2_outputs(6757) <= a or b;
    layer2_outputs(6758) <= not b;
    layer2_outputs(6759) <= not (a or b);
    layer2_outputs(6760) <= not (a or b);
    layer2_outputs(6761) <= '0';
    layer2_outputs(6762) <= not b;
    layer2_outputs(6763) <= b and not a;
    layer2_outputs(6764) <= not (a and b);
    layer2_outputs(6765) <= not a or b;
    layer2_outputs(6766) <= not (a or b);
    layer2_outputs(6767) <= a or b;
    layer2_outputs(6768) <= a;
    layer2_outputs(6769) <= not a or b;
    layer2_outputs(6770) <= '1';
    layer2_outputs(6771) <= b;
    layer2_outputs(6772) <= '1';
    layer2_outputs(6773) <= a xor b;
    layer2_outputs(6774) <= a and b;
    layer2_outputs(6775) <= not (a and b);
    layer2_outputs(6776) <= a or b;
    layer2_outputs(6777) <= a;
    layer2_outputs(6778) <= a;
    layer2_outputs(6779) <= b and not a;
    layer2_outputs(6780) <= a;
    layer2_outputs(6781) <= a and b;
    layer2_outputs(6782) <= b;
    layer2_outputs(6783) <= a;
    layer2_outputs(6784) <= b;
    layer2_outputs(6785) <= not a;
    layer2_outputs(6786) <= a xor b;
    layer2_outputs(6787) <= not (a or b);
    layer2_outputs(6788) <= a or b;
    layer2_outputs(6789) <= b;
    layer2_outputs(6790) <= a or b;
    layer2_outputs(6791) <= b;
    layer2_outputs(6792) <= not (a or b);
    layer2_outputs(6793) <= not b;
    layer2_outputs(6794) <= b;
    layer2_outputs(6795) <= not (a or b);
    layer2_outputs(6796) <= not (a or b);
    layer2_outputs(6797) <= b and not a;
    layer2_outputs(6798) <= not a or b;
    layer2_outputs(6799) <= not b or a;
    layer2_outputs(6800) <= not a;
    layer2_outputs(6801) <= b;
    layer2_outputs(6802) <= a and b;
    layer2_outputs(6803) <= not (a and b);
    layer2_outputs(6804) <= b;
    layer2_outputs(6805) <= a and b;
    layer2_outputs(6806) <= a and b;
    layer2_outputs(6807) <= b;
    layer2_outputs(6808) <= not (a xor b);
    layer2_outputs(6809) <= a xor b;
    layer2_outputs(6810) <= not b;
    layer2_outputs(6811) <= b;
    layer2_outputs(6812) <= not a;
    layer2_outputs(6813) <= not a;
    layer2_outputs(6814) <= not (a or b);
    layer2_outputs(6815) <= a and not b;
    layer2_outputs(6816) <= not (a xor b);
    layer2_outputs(6817) <= '1';
    layer2_outputs(6818) <= a;
    layer2_outputs(6819) <= a or b;
    layer2_outputs(6820) <= b;
    layer2_outputs(6821) <= b and not a;
    layer2_outputs(6822) <= not (a and b);
    layer2_outputs(6823) <= a or b;
    layer2_outputs(6824) <= not (a and b);
    layer2_outputs(6825) <= a or b;
    layer2_outputs(6826) <= a or b;
    layer2_outputs(6827) <= '1';
    layer2_outputs(6828) <= not b;
    layer2_outputs(6829) <= '0';
    layer2_outputs(6830) <= not a;
    layer2_outputs(6831) <= not (a xor b);
    layer2_outputs(6832) <= a;
    layer2_outputs(6833) <= a;
    layer2_outputs(6834) <= not a;
    layer2_outputs(6835) <= a and not b;
    layer2_outputs(6836) <= a;
    layer2_outputs(6837) <= not (a or b);
    layer2_outputs(6838) <= '1';
    layer2_outputs(6839) <= not (a or b);
    layer2_outputs(6840) <= not b or a;
    layer2_outputs(6841) <= a;
    layer2_outputs(6842) <= not a or b;
    layer2_outputs(6843) <= a;
    layer2_outputs(6844) <= a;
    layer2_outputs(6845) <= not b or a;
    layer2_outputs(6846) <= not a or b;
    layer2_outputs(6847) <= a and b;
    layer2_outputs(6848) <= '1';
    layer2_outputs(6849) <= not b or a;
    layer2_outputs(6850) <= a or b;
    layer2_outputs(6851) <= a and not b;
    layer2_outputs(6852) <= not b;
    layer2_outputs(6853) <= '1';
    layer2_outputs(6854) <= not b or a;
    layer2_outputs(6855) <= b;
    layer2_outputs(6856) <= not a or b;
    layer2_outputs(6857) <= not a or b;
    layer2_outputs(6858) <= b and not a;
    layer2_outputs(6859) <= not a;
    layer2_outputs(6860) <= not b or a;
    layer2_outputs(6861) <= a;
    layer2_outputs(6862) <= a or b;
    layer2_outputs(6863) <= not (a and b);
    layer2_outputs(6864) <= '0';
    layer2_outputs(6865) <= '1';
    layer2_outputs(6866) <= '0';
    layer2_outputs(6867) <= not b;
    layer2_outputs(6868) <= a;
    layer2_outputs(6869) <= not (a and b);
    layer2_outputs(6870) <= a or b;
    layer2_outputs(6871) <= a;
    layer2_outputs(6872) <= '1';
    layer2_outputs(6873) <= not (a and b);
    layer2_outputs(6874) <= a and b;
    layer2_outputs(6875) <= not a or b;
    layer2_outputs(6876) <= not b or a;
    layer2_outputs(6877) <= a;
    layer2_outputs(6878) <= b;
    layer2_outputs(6879) <= not b;
    layer2_outputs(6880) <= not b;
    layer2_outputs(6881) <= not b or a;
    layer2_outputs(6882) <= b and not a;
    layer2_outputs(6883) <= not a or b;
    layer2_outputs(6884) <= '1';
    layer2_outputs(6885) <= b;
    layer2_outputs(6886) <= a or b;
    layer2_outputs(6887) <= not (a and b);
    layer2_outputs(6888) <= not b;
    layer2_outputs(6889) <= b and not a;
    layer2_outputs(6890) <= b;
    layer2_outputs(6891) <= '0';
    layer2_outputs(6892) <= b;
    layer2_outputs(6893) <= a;
    layer2_outputs(6894) <= '0';
    layer2_outputs(6895) <= a;
    layer2_outputs(6896) <= a or b;
    layer2_outputs(6897) <= '1';
    layer2_outputs(6898) <= a xor b;
    layer2_outputs(6899) <= a and b;
    layer2_outputs(6900) <= '1';
    layer2_outputs(6901) <= a or b;
    layer2_outputs(6902) <= a or b;
    layer2_outputs(6903) <= b and not a;
    layer2_outputs(6904) <= not (a xor b);
    layer2_outputs(6905) <= not (a xor b);
    layer2_outputs(6906) <= a and not b;
    layer2_outputs(6907) <= not (a or b);
    layer2_outputs(6908) <= b;
    layer2_outputs(6909) <= not (a xor b);
    layer2_outputs(6910) <= a or b;
    layer2_outputs(6911) <= b and not a;
    layer2_outputs(6912) <= not b;
    layer2_outputs(6913) <= b;
    layer2_outputs(6914) <= '0';
    layer2_outputs(6915) <= not b;
    layer2_outputs(6916) <= b;
    layer2_outputs(6917) <= not (a or b);
    layer2_outputs(6918) <= not a or b;
    layer2_outputs(6919) <= not (a xor b);
    layer2_outputs(6920) <= a and not b;
    layer2_outputs(6921) <= not b or a;
    layer2_outputs(6922) <= a or b;
    layer2_outputs(6923) <= a and not b;
    layer2_outputs(6924) <= a;
    layer2_outputs(6925) <= not (a or b);
    layer2_outputs(6926) <= b;
    layer2_outputs(6927) <= not b;
    layer2_outputs(6928) <= b;
    layer2_outputs(6929) <= a and not b;
    layer2_outputs(6930) <= a xor b;
    layer2_outputs(6931) <= not b;
    layer2_outputs(6932) <= a or b;
    layer2_outputs(6933) <= b;
    layer2_outputs(6934) <= not (a or b);
    layer2_outputs(6935) <= b and not a;
    layer2_outputs(6936) <= a and b;
    layer2_outputs(6937) <= not (a xor b);
    layer2_outputs(6938) <= not b or a;
    layer2_outputs(6939) <= b and not a;
    layer2_outputs(6940) <= not a or b;
    layer2_outputs(6941) <= not a;
    layer2_outputs(6942) <= '0';
    layer2_outputs(6943) <= b;
    layer2_outputs(6944) <= not a;
    layer2_outputs(6945) <= b;
    layer2_outputs(6946) <= b;
    layer2_outputs(6947) <= a and b;
    layer2_outputs(6948) <= a xor b;
    layer2_outputs(6949) <= not a;
    layer2_outputs(6950) <= b and not a;
    layer2_outputs(6951) <= '0';
    layer2_outputs(6952) <= not b;
    layer2_outputs(6953) <= b and not a;
    layer2_outputs(6954) <= a and not b;
    layer2_outputs(6955) <= b;
    layer2_outputs(6956) <= a xor b;
    layer2_outputs(6957) <= a and not b;
    layer2_outputs(6958) <= a;
    layer2_outputs(6959) <= not a or b;
    layer2_outputs(6960) <= b and not a;
    layer2_outputs(6961) <= a;
    layer2_outputs(6962) <= a;
    layer2_outputs(6963) <= b and not a;
    layer2_outputs(6964) <= a;
    layer2_outputs(6965) <= a or b;
    layer2_outputs(6966) <= not b;
    layer2_outputs(6967) <= not a or b;
    layer2_outputs(6968) <= not (a or b);
    layer2_outputs(6969) <= '0';
    layer2_outputs(6970) <= a;
    layer2_outputs(6971) <= not a or b;
    layer2_outputs(6972) <= not a or b;
    layer2_outputs(6973) <= a or b;
    layer2_outputs(6974) <= not b;
    layer2_outputs(6975) <= not (a or b);
    layer2_outputs(6976) <= '0';
    layer2_outputs(6977) <= not b or a;
    layer2_outputs(6978) <= b;
    layer2_outputs(6979) <= a xor b;
    layer2_outputs(6980) <= not (a or b);
    layer2_outputs(6981) <= not a;
    layer2_outputs(6982) <= a and b;
    layer2_outputs(6983) <= b and not a;
    layer2_outputs(6984) <= '1';
    layer2_outputs(6985) <= b and not a;
    layer2_outputs(6986) <= '1';
    layer2_outputs(6987) <= not (a and b);
    layer2_outputs(6988) <= a or b;
    layer2_outputs(6989) <= '0';
    layer2_outputs(6990) <= a or b;
    layer2_outputs(6991) <= not a;
    layer2_outputs(6992) <= not (a or b);
    layer2_outputs(6993) <= a or b;
    layer2_outputs(6994) <= a and b;
    layer2_outputs(6995) <= a and b;
    layer2_outputs(6996) <= not b or a;
    layer2_outputs(6997) <= '0';
    layer2_outputs(6998) <= not a or b;
    layer2_outputs(6999) <= not (a or b);
    layer2_outputs(7000) <= a and b;
    layer2_outputs(7001) <= not b;
    layer2_outputs(7002) <= a xor b;
    layer2_outputs(7003) <= not b;
    layer2_outputs(7004) <= not a;
    layer2_outputs(7005) <= not b;
    layer2_outputs(7006) <= '1';
    layer2_outputs(7007) <= b;
    layer2_outputs(7008) <= a and b;
    layer2_outputs(7009) <= a;
    layer2_outputs(7010) <= b and not a;
    layer2_outputs(7011) <= not b;
    layer2_outputs(7012) <= not b;
    layer2_outputs(7013) <= a xor b;
    layer2_outputs(7014) <= not a;
    layer2_outputs(7015) <= not (a and b);
    layer2_outputs(7016) <= b and not a;
    layer2_outputs(7017) <= a or b;
    layer2_outputs(7018) <= not b;
    layer2_outputs(7019) <= a and not b;
    layer2_outputs(7020) <= a and not b;
    layer2_outputs(7021) <= not a;
    layer2_outputs(7022) <= a and b;
    layer2_outputs(7023) <= '0';
    layer2_outputs(7024) <= not b or a;
    layer2_outputs(7025) <= a and b;
    layer2_outputs(7026) <= not (a or b);
    layer2_outputs(7027) <= b and not a;
    layer2_outputs(7028) <= not (a xor b);
    layer2_outputs(7029) <= not (a and b);
    layer2_outputs(7030) <= not b or a;
    layer2_outputs(7031) <= not a;
    layer2_outputs(7032) <= not b or a;
    layer2_outputs(7033) <= a and not b;
    layer2_outputs(7034) <= not (a and b);
    layer2_outputs(7035) <= '1';
    layer2_outputs(7036) <= not a;
    layer2_outputs(7037) <= b;
    layer2_outputs(7038) <= '0';
    layer2_outputs(7039) <= b and not a;
    layer2_outputs(7040) <= not (a or b);
    layer2_outputs(7041) <= a or b;
    layer2_outputs(7042) <= not b;
    layer2_outputs(7043) <= a;
    layer2_outputs(7044) <= '0';
    layer2_outputs(7045) <= not b;
    layer2_outputs(7046) <= b and not a;
    layer2_outputs(7047) <= a xor b;
    layer2_outputs(7048) <= not b;
    layer2_outputs(7049) <= not a;
    layer2_outputs(7050) <= a and b;
    layer2_outputs(7051) <= a and not b;
    layer2_outputs(7052) <= a;
    layer2_outputs(7053) <= a or b;
    layer2_outputs(7054) <= b and not a;
    layer2_outputs(7055) <= not b;
    layer2_outputs(7056) <= a xor b;
    layer2_outputs(7057) <= a and not b;
    layer2_outputs(7058) <= a and not b;
    layer2_outputs(7059) <= not (a or b);
    layer2_outputs(7060) <= a and not b;
    layer2_outputs(7061) <= a or b;
    layer2_outputs(7062) <= b;
    layer2_outputs(7063) <= a;
    layer2_outputs(7064) <= not b;
    layer2_outputs(7065) <= not a;
    layer2_outputs(7066) <= not b or a;
    layer2_outputs(7067) <= not b or a;
    layer2_outputs(7068) <= a and not b;
    layer2_outputs(7069) <= not b or a;
    layer2_outputs(7070) <= not (a or b);
    layer2_outputs(7071) <= a or b;
    layer2_outputs(7072) <= not a;
    layer2_outputs(7073) <= a and not b;
    layer2_outputs(7074) <= not (a or b);
    layer2_outputs(7075) <= a and b;
    layer2_outputs(7076) <= not a or b;
    layer2_outputs(7077) <= a xor b;
    layer2_outputs(7078) <= not b or a;
    layer2_outputs(7079) <= a xor b;
    layer2_outputs(7080) <= not a;
    layer2_outputs(7081) <= a and not b;
    layer2_outputs(7082) <= not (a and b);
    layer2_outputs(7083) <= '0';
    layer2_outputs(7084) <= not a;
    layer2_outputs(7085) <= not a;
    layer2_outputs(7086) <= b;
    layer2_outputs(7087) <= not (a and b);
    layer2_outputs(7088) <= a or b;
    layer2_outputs(7089) <= not b or a;
    layer2_outputs(7090) <= a;
    layer2_outputs(7091) <= not (a and b);
    layer2_outputs(7092) <= not b;
    layer2_outputs(7093) <= not a;
    layer2_outputs(7094) <= a and not b;
    layer2_outputs(7095) <= not b;
    layer2_outputs(7096) <= a;
    layer2_outputs(7097) <= a and b;
    layer2_outputs(7098) <= not (a and b);
    layer2_outputs(7099) <= b;
    layer2_outputs(7100) <= a and not b;
    layer2_outputs(7101) <= not (a or b);
    layer2_outputs(7102) <= not (a and b);
    layer2_outputs(7103) <= not (a and b);
    layer2_outputs(7104) <= a or b;
    layer2_outputs(7105) <= not (a or b);
    layer2_outputs(7106) <= not a or b;
    layer2_outputs(7107) <= a;
    layer2_outputs(7108) <= not (a and b);
    layer2_outputs(7109) <= not (a or b);
    layer2_outputs(7110) <= not b or a;
    layer2_outputs(7111) <= not (a xor b);
    layer2_outputs(7112) <= not b;
    layer2_outputs(7113) <= a and b;
    layer2_outputs(7114) <= not a;
    layer2_outputs(7115) <= not a;
    layer2_outputs(7116) <= not (a and b);
    layer2_outputs(7117) <= not b;
    layer2_outputs(7118) <= not a;
    layer2_outputs(7119) <= not b;
    layer2_outputs(7120) <= b;
    layer2_outputs(7121) <= a;
    layer2_outputs(7122) <= not (a xor b);
    layer2_outputs(7123) <= not a or b;
    layer2_outputs(7124) <= a xor b;
    layer2_outputs(7125) <= not a;
    layer2_outputs(7126) <= a and not b;
    layer2_outputs(7127) <= b;
    layer2_outputs(7128) <= not b or a;
    layer2_outputs(7129) <= not a;
    layer2_outputs(7130) <= b;
    layer2_outputs(7131) <= not b;
    layer2_outputs(7132) <= not (a and b);
    layer2_outputs(7133) <= not (a and b);
    layer2_outputs(7134) <= not a or b;
    layer2_outputs(7135) <= not b;
    layer2_outputs(7136) <= not b or a;
    layer2_outputs(7137) <= a and b;
    layer2_outputs(7138) <= a or b;
    layer2_outputs(7139) <= a;
    layer2_outputs(7140) <= not b or a;
    layer2_outputs(7141) <= not a;
    layer2_outputs(7142) <= not a or b;
    layer2_outputs(7143) <= b and not a;
    layer2_outputs(7144) <= a and b;
    layer2_outputs(7145) <= '0';
    layer2_outputs(7146) <= a and b;
    layer2_outputs(7147) <= a;
    layer2_outputs(7148) <= '0';
    layer2_outputs(7149) <= not a or b;
    layer2_outputs(7150) <= not (a xor b);
    layer2_outputs(7151) <= b;
    layer2_outputs(7152) <= a or b;
    layer2_outputs(7153) <= not a or b;
    layer2_outputs(7154) <= not b or a;
    layer2_outputs(7155) <= a;
    layer2_outputs(7156) <= b and not a;
    layer2_outputs(7157) <= '0';
    layer2_outputs(7158) <= not (a and b);
    layer2_outputs(7159) <= a or b;
    layer2_outputs(7160) <= a;
    layer2_outputs(7161) <= a and not b;
    layer2_outputs(7162) <= b and not a;
    layer2_outputs(7163) <= b and not a;
    layer2_outputs(7164) <= not a or b;
    layer2_outputs(7165) <= not b or a;
    layer2_outputs(7166) <= a xor b;
    layer2_outputs(7167) <= not a or b;
    layer2_outputs(7168) <= not (a and b);
    layer2_outputs(7169) <= b;
    layer2_outputs(7170) <= a and b;
    layer2_outputs(7171) <= not a;
    layer2_outputs(7172) <= not (a or b);
    layer2_outputs(7173) <= a and b;
    layer2_outputs(7174) <= b and not a;
    layer2_outputs(7175) <= not a or b;
    layer2_outputs(7176) <= b;
    layer2_outputs(7177) <= a;
    layer2_outputs(7178) <= b and not a;
    layer2_outputs(7179) <= not b;
    layer2_outputs(7180) <= not (a and b);
    layer2_outputs(7181) <= not b;
    layer2_outputs(7182) <= not a;
    layer2_outputs(7183) <= not (a and b);
    layer2_outputs(7184) <= a;
    layer2_outputs(7185) <= '0';
    layer2_outputs(7186) <= not (a and b);
    layer2_outputs(7187) <= a and not b;
    layer2_outputs(7188) <= '0';
    layer2_outputs(7189) <= '1';
    layer2_outputs(7190) <= not (a xor b);
    layer2_outputs(7191) <= a;
    layer2_outputs(7192) <= b and not a;
    layer2_outputs(7193) <= not a;
    layer2_outputs(7194) <= not (a or b);
    layer2_outputs(7195) <= a;
    layer2_outputs(7196) <= b;
    layer2_outputs(7197) <= not a;
    layer2_outputs(7198) <= not (a and b);
    layer2_outputs(7199) <= b;
    layer2_outputs(7200) <= '1';
    layer2_outputs(7201) <= not b;
    layer2_outputs(7202) <= not a;
    layer2_outputs(7203) <= a or b;
    layer2_outputs(7204) <= not b;
    layer2_outputs(7205) <= b;
    layer2_outputs(7206) <= a or b;
    layer2_outputs(7207) <= a;
    layer2_outputs(7208) <= not b;
    layer2_outputs(7209) <= not (a or b);
    layer2_outputs(7210) <= b and not a;
    layer2_outputs(7211) <= a and not b;
    layer2_outputs(7212) <= a;
    layer2_outputs(7213) <= not (a and b);
    layer2_outputs(7214) <= a and b;
    layer2_outputs(7215) <= b;
    layer2_outputs(7216) <= not b;
    layer2_outputs(7217) <= not a;
    layer2_outputs(7218) <= '0';
    layer2_outputs(7219) <= not b;
    layer2_outputs(7220) <= not b;
    layer2_outputs(7221) <= b;
    layer2_outputs(7222) <= not b;
    layer2_outputs(7223) <= not b or a;
    layer2_outputs(7224) <= a and not b;
    layer2_outputs(7225) <= not b;
    layer2_outputs(7226) <= not (a and b);
    layer2_outputs(7227) <= a;
    layer2_outputs(7228) <= '0';
    layer2_outputs(7229) <= '0';
    layer2_outputs(7230) <= not a or b;
    layer2_outputs(7231) <= a and not b;
    layer2_outputs(7232) <= a;
    layer2_outputs(7233) <= not b;
    layer2_outputs(7234) <= not b or a;
    layer2_outputs(7235) <= not b or a;
    layer2_outputs(7236) <= not (a xor b);
    layer2_outputs(7237) <= '1';
    layer2_outputs(7238) <= b and not a;
    layer2_outputs(7239) <= a;
    layer2_outputs(7240) <= '1';
    layer2_outputs(7241) <= not b or a;
    layer2_outputs(7242) <= not (a and b);
    layer2_outputs(7243) <= '0';
    layer2_outputs(7244) <= not b;
    layer2_outputs(7245) <= not b;
    layer2_outputs(7246) <= a;
    layer2_outputs(7247) <= not a;
    layer2_outputs(7248) <= not (a or b);
    layer2_outputs(7249) <= a or b;
    layer2_outputs(7250) <= '0';
    layer2_outputs(7251) <= a and b;
    layer2_outputs(7252) <= b;
    layer2_outputs(7253) <= b;
    layer2_outputs(7254) <= b and not a;
    layer2_outputs(7255) <= not a or b;
    layer2_outputs(7256) <= b and not a;
    layer2_outputs(7257) <= a and not b;
    layer2_outputs(7258) <= a and b;
    layer2_outputs(7259) <= not (a or b);
    layer2_outputs(7260) <= '0';
    layer2_outputs(7261) <= not (a and b);
    layer2_outputs(7262) <= not a;
    layer2_outputs(7263) <= not a;
    layer2_outputs(7264) <= not b or a;
    layer2_outputs(7265) <= a and b;
    layer2_outputs(7266) <= not (a and b);
    layer2_outputs(7267) <= '0';
    layer2_outputs(7268) <= '0';
    layer2_outputs(7269) <= a and b;
    layer2_outputs(7270) <= b and not a;
    layer2_outputs(7271) <= not b or a;
    layer2_outputs(7272) <= not a or b;
    layer2_outputs(7273) <= not b;
    layer2_outputs(7274) <= not (a or b);
    layer2_outputs(7275) <= not a or b;
    layer2_outputs(7276) <= not b;
    layer2_outputs(7277) <= a;
    layer2_outputs(7278) <= not a;
    layer2_outputs(7279) <= not a or b;
    layer2_outputs(7280) <= not (a or b);
    layer2_outputs(7281) <= b and not a;
    layer2_outputs(7282) <= '1';
    layer2_outputs(7283) <= a or b;
    layer2_outputs(7284) <= not a or b;
    layer2_outputs(7285) <= '1';
    layer2_outputs(7286) <= not b;
    layer2_outputs(7287) <= not b or a;
    layer2_outputs(7288) <= not a or b;
    layer2_outputs(7289) <= a;
    layer2_outputs(7290) <= '1';
    layer2_outputs(7291) <= b and not a;
    layer2_outputs(7292) <= b;
    layer2_outputs(7293) <= not (a or b);
    layer2_outputs(7294) <= a and not b;
    layer2_outputs(7295) <= not a or b;
    layer2_outputs(7296) <= a and not b;
    layer2_outputs(7297) <= not b or a;
    layer2_outputs(7298) <= a and b;
    layer2_outputs(7299) <= not a;
    layer2_outputs(7300) <= a and b;
    layer2_outputs(7301) <= not a or b;
    layer2_outputs(7302) <= a;
    layer2_outputs(7303) <= not b or a;
    layer2_outputs(7304) <= a and b;
    layer2_outputs(7305) <= b and not a;
    layer2_outputs(7306) <= not (a xor b);
    layer2_outputs(7307) <= not b or a;
    layer2_outputs(7308) <= not (a xor b);
    layer2_outputs(7309) <= not (a or b);
    layer2_outputs(7310) <= not a;
    layer2_outputs(7311) <= not a;
    layer2_outputs(7312) <= a and not b;
    layer2_outputs(7313) <= a xor b;
    layer2_outputs(7314) <= not b;
    layer2_outputs(7315) <= not b;
    layer2_outputs(7316) <= a;
    layer2_outputs(7317) <= b;
    layer2_outputs(7318) <= not (a or b);
    layer2_outputs(7319) <= not a;
    layer2_outputs(7320) <= '0';
    layer2_outputs(7321) <= '0';
    layer2_outputs(7322) <= not (a xor b);
    layer2_outputs(7323) <= a;
    layer2_outputs(7324) <= not a;
    layer2_outputs(7325) <= not b;
    layer2_outputs(7326) <= a and not b;
    layer2_outputs(7327) <= a and not b;
    layer2_outputs(7328) <= not a or b;
    layer2_outputs(7329) <= not a or b;
    layer2_outputs(7330) <= not a;
    layer2_outputs(7331) <= '0';
    layer2_outputs(7332) <= b and not a;
    layer2_outputs(7333) <= a;
    layer2_outputs(7334) <= a and b;
    layer2_outputs(7335) <= '1';
    layer2_outputs(7336) <= b;
    layer2_outputs(7337) <= b and not a;
    layer2_outputs(7338) <= a and not b;
    layer2_outputs(7339) <= a;
    layer2_outputs(7340) <= not (a or b);
    layer2_outputs(7341) <= b and not a;
    layer2_outputs(7342) <= not b;
    layer2_outputs(7343) <= a;
    layer2_outputs(7344) <= not (a xor b);
    layer2_outputs(7345) <= a and not b;
    layer2_outputs(7346) <= not b;
    layer2_outputs(7347) <= b;
    layer2_outputs(7348) <= not (a and b);
    layer2_outputs(7349) <= not (a and b);
    layer2_outputs(7350) <= a xor b;
    layer2_outputs(7351) <= '1';
    layer2_outputs(7352) <= not (a xor b);
    layer2_outputs(7353) <= a and not b;
    layer2_outputs(7354) <= not a or b;
    layer2_outputs(7355) <= not a or b;
    layer2_outputs(7356) <= a;
    layer2_outputs(7357) <= a xor b;
    layer2_outputs(7358) <= not (a xor b);
    layer2_outputs(7359) <= b;
    layer2_outputs(7360) <= not a or b;
    layer2_outputs(7361) <= a;
    layer2_outputs(7362) <= not a;
    layer2_outputs(7363) <= not a or b;
    layer2_outputs(7364) <= not a or b;
    layer2_outputs(7365) <= '0';
    layer2_outputs(7366) <= not a;
    layer2_outputs(7367) <= a and b;
    layer2_outputs(7368) <= a xor b;
    layer2_outputs(7369) <= '1';
    layer2_outputs(7370) <= '0';
    layer2_outputs(7371) <= a and not b;
    layer2_outputs(7372) <= '1';
    layer2_outputs(7373) <= a xor b;
    layer2_outputs(7374) <= not b or a;
    layer2_outputs(7375) <= not a;
    layer2_outputs(7376) <= b;
    layer2_outputs(7377) <= a;
    layer2_outputs(7378) <= a and b;
    layer2_outputs(7379) <= a;
    layer2_outputs(7380) <= '1';
    layer2_outputs(7381) <= a or b;
    layer2_outputs(7382) <= not a;
    layer2_outputs(7383) <= '1';
    layer2_outputs(7384) <= '0';
    layer2_outputs(7385) <= a and b;
    layer2_outputs(7386) <= not a;
    layer2_outputs(7387) <= '0';
    layer2_outputs(7388) <= b;
    layer2_outputs(7389) <= b and not a;
    layer2_outputs(7390) <= not b;
    layer2_outputs(7391) <= '0';
    layer2_outputs(7392) <= not (a or b);
    layer2_outputs(7393) <= not (a or b);
    layer2_outputs(7394) <= a or b;
    layer2_outputs(7395) <= b;
    layer2_outputs(7396) <= a or b;
    layer2_outputs(7397) <= '1';
    layer2_outputs(7398) <= not (a and b);
    layer2_outputs(7399) <= not (a xor b);
    layer2_outputs(7400) <= a and b;
    layer2_outputs(7401) <= not a or b;
    layer2_outputs(7402) <= a or b;
    layer2_outputs(7403) <= '1';
    layer2_outputs(7404) <= a and not b;
    layer2_outputs(7405) <= not b;
    layer2_outputs(7406) <= a and not b;
    layer2_outputs(7407) <= not a;
    layer2_outputs(7408) <= not b or a;
    layer2_outputs(7409) <= not a;
    layer2_outputs(7410) <= a or b;
    layer2_outputs(7411) <= not b;
    layer2_outputs(7412) <= a and b;
    layer2_outputs(7413) <= not (a or b);
    layer2_outputs(7414) <= a and b;
    layer2_outputs(7415) <= a xor b;
    layer2_outputs(7416) <= '0';
    layer2_outputs(7417) <= not (a or b);
    layer2_outputs(7418) <= a;
    layer2_outputs(7419) <= not b;
    layer2_outputs(7420) <= a xor b;
    layer2_outputs(7421) <= b and not a;
    layer2_outputs(7422) <= b;
    layer2_outputs(7423) <= not b;
    layer2_outputs(7424) <= a and not b;
    layer2_outputs(7425) <= not a;
    layer2_outputs(7426) <= '1';
    layer2_outputs(7427) <= not (a xor b);
    layer2_outputs(7428) <= not (a or b);
    layer2_outputs(7429) <= not (a and b);
    layer2_outputs(7430) <= b and not a;
    layer2_outputs(7431) <= a and not b;
    layer2_outputs(7432) <= b;
    layer2_outputs(7433) <= b and not a;
    layer2_outputs(7434) <= not a or b;
    layer2_outputs(7435) <= a and b;
    layer2_outputs(7436) <= not a or b;
    layer2_outputs(7437) <= not (a and b);
    layer2_outputs(7438) <= not (a and b);
    layer2_outputs(7439) <= not a or b;
    layer2_outputs(7440) <= not a;
    layer2_outputs(7441) <= a or b;
    layer2_outputs(7442) <= '0';
    layer2_outputs(7443) <= b and not a;
    layer2_outputs(7444) <= not b;
    layer2_outputs(7445) <= '1';
    layer2_outputs(7446) <= not b or a;
    layer2_outputs(7447) <= not a;
    layer2_outputs(7448) <= b and not a;
    layer2_outputs(7449) <= b;
    layer2_outputs(7450) <= not a;
    layer2_outputs(7451) <= a and not b;
    layer2_outputs(7452) <= not b;
    layer2_outputs(7453) <= a and b;
    layer2_outputs(7454) <= not b or a;
    layer2_outputs(7455) <= not b or a;
    layer2_outputs(7456) <= not a or b;
    layer2_outputs(7457) <= a;
    layer2_outputs(7458) <= not (a or b);
    layer2_outputs(7459) <= b;
    layer2_outputs(7460) <= not a;
    layer2_outputs(7461) <= not (a and b);
    layer2_outputs(7462) <= not b or a;
    layer2_outputs(7463) <= not (a and b);
    layer2_outputs(7464) <= a and not b;
    layer2_outputs(7465) <= a;
    layer2_outputs(7466) <= not a or b;
    layer2_outputs(7467) <= not a or b;
    layer2_outputs(7468) <= '1';
    layer2_outputs(7469) <= not b;
    layer2_outputs(7470) <= not b or a;
    layer2_outputs(7471) <= '0';
    layer2_outputs(7472) <= not a or b;
    layer2_outputs(7473) <= a or b;
    layer2_outputs(7474) <= not a;
    layer2_outputs(7475) <= a and not b;
    layer2_outputs(7476) <= not b;
    layer2_outputs(7477) <= not a;
    layer2_outputs(7478) <= not a or b;
    layer2_outputs(7479) <= '1';
    layer2_outputs(7480) <= a;
    layer2_outputs(7481) <= a and not b;
    layer2_outputs(7482) <= b and not a;
    layer2_outputs(7483) <= not b;
    layer2_outputs(7484) <= b;
    layer2_outputs(7485) <= a;
    layer2_outputs(7486) <= b;
    layer2_outputs(7487) <= a and not b;
    layer2_outputs(7488) <= a and b;
    layer2_outputs(7489) <= '1';
    layer2_outputs(7490) <= not a;
    layer2_outputs(7491) <= not a;
    layer2_outputs(7492) <= '0';
    layer2_outputs(7493) <= not (a and b);
    layer2_outputs(7494) <= not (a or b);
    layer2_outputs(7495) <= not a or b;
    layer2_outputs(7496) <= a;
    layer2_outputs(7497) <= not b or a;
    layer2_outputs(7498) <= '1';
    layer2_outputs(7499) <= '1';
    layer2_outputs(7500) <= a or b;
    layer2_outputs(7501) <= not b;
    layer2_outputs(7502) <= not (a xor b);
    layer2_outputs(7503) <= a or b;
    layer2_outputs(7504) <= b and not a;
    layer2_outputs(7505) <= not (a or b);
    layer2_outputs(7506) <= a and not b;
    layer2_outputs(7507) <= not (a xor b);
    layer2_outputs(7508) <= a;
    layer2_outputs(7509) <= not a or b;
    layer2_outputs(7510) <= b;
    layer2_outputs(7511) <= not (a or b);
    layer2_outputs(7512) <= a and not b;
    layer2_outputs(7513) <= not a or b;
    layer2_outputs(7514) <= '1';
    layer2_outputs(7515) <= not (a and b);
    layer2_outputs(7516) <= b;
    layer2_outputs(7517) <= not a;
    layer2_outputs(7518) <= a and b;
    layer2_outputs(7519) <= not (a xor b);
    layer2_outputs(7520) <= a and not b;
    layer2_outputs(7521) <= b;
    layer2_outputs(7522) <= '1';
    layer2_outputs(7523) <= '1';
    layer2_outputs(7524) <= a and not b;
    layer2_outputs(7525) <= a and not b;
    layer2_outputs(7526) <= not (a xor b);
    layer2_outputs(7527) <= a and not b;
    layer2_outputs(7528) <= not b;
    layer2_outputs(7529) <= a and not b;
    layer2_outputs(7530) <= not b or a;
    layer2_outputs(7531) <= a and not b;
    layer2_outputs(7532) <= a or b;
    layer2_outputs(7533) <= a and not b;
    layer2_outputs(7534) <= '0';
    layer2_outputs(7535) <= not b or a;
    layer2_outputs(7536) <= '1';
    layer2_outputs(7537) <= not a;
    layer2_outputs(7538) <= b;
    layer2_outputs(7539) <= not a or b;
    layer2_outputs(7540) <= b;
    layer2_outputs(7541) <= a xor b;
    layer2_outputs(7542) <= not (a and b);
    layer2_outputs(7543) <= not a;
    layer2_outputs(7544) <= a and not b;
    layer2_outputs(7545) <= not b;
    layer2_outputs(7546) <= '1';
    layer2_outputs(7547) <= not (a and b);
    layer2_outputs(7548) <= not (a and b);
    layer2_outputs(7549) <= not a;
    layer2_outputs(7550) <= b;
    layer2_outputs(7551) <= a and b;
    layer2_outputs(7552) <= a and not b;
    layer2_outputs(7553) <= not a;
    layer2_outputs(7554) <= b;
    layer2_outputs(7555) <= not a or b;
    layer2_outputs(7556) <= b;
    layer2_outputs(7557) <= not (a and b);
    layer2_outputs(7558) <= b and not a;
    layer2_outputs(7559) <= not a or b;
    layer2_outputs(7560) <= a and not b;
    layer2_outputs(7561) <= a;
    layer2_outputs(7562) <= not (a and b);
    layer2_outputs(7563) <= not a or b;
    layer2_outputs(7564) <= a or b;
    layer2_outputs(7565) <= not (a and b);
    layer2_outputs(7566) <= a and not b;
    layer2_outputs(7567) <= not b;
    layer2_outputs(7568) <= b;
    layer2_outputs(7569) <= a and not b;
    layer2_outputs(7570) <= '0';
    layer2_outputs(7571) <= a and not b;
    layer2_outputs(7572) <= a and not b;
    layer2_outputs(7573) <= b and not a;
    layer2_outputs(7574) <= a or b;
    layer2_outputs(7575) <= not b or a;
    layer2_outputs(7576) <= not a or b;
    layer2_outputs(7577) <= a or b;
    layer2_outputs(7578) <= not a;
    layer2_outputs(7579) <= '0';
    layer2_outputs(7580) <= not a;
    layer2_outputs(7581) <= b;
    layer2_outputs(7582) <= a;
    layer2_outputs(7583) <= not b;
    layer2_outputs(7584) <= '1';
    layer2_outputs(7585) <= a or b;
    layer2_outputs(7586) <= not (a and b);
    layer2_outputs(7587) <= not (a or b);
    layer2_outputs(7588) <= a and not b;
    layer2_outputs(7589) <= b and not a;
    layer2_outputs(7590) <= b;
    layer2_outputs(7591) <= not (a or b);
    layer2_outputs(7592) <= not a or b;
    layer2_outputs(7593) <= not b;
    layer2_outputs(7594) <= not (a or b);
    layer2_outputs(7595) <= a or b;
    layer2_outputs(7596) <= not (a xor b);
    layer2_outputs(7597) <= b and not a;
    layer2_outputs(7598) <= not a;
    layer2_outputs(7599) <= a;
    layer2_outputs(7600) <= a and b;
    layer2_outputs(7601) <= a;
    layer2_outputs(7602) <= a and not b;
    layer2_outputs(7603) <= a and b;
    layer2_outputs(7604) <= not a;
    layer2_outputs(7605) <= not a or b;
    layer2_outputs(7606) <= b and not a;
    layer2_outputs(7607) <= '1';
    layer2_outputs(7608) <= not (a or b);
    layer2_outputs(7609) <= '0';
    layer2_outputs(7610) <= not (a and b);
    layer2_outputs(7611) <= not b;
    layer2_outputs(7612) <= a or b;
    layer2_outputs(7613) <= not a or b;
    layer2_outputs(7614) <= not b or a;
    layer2_outputs(7615) <= a;
    layer2_outputs(7616) <= a or b;
    layer2_outputs(7617) <= not a;
    layer2_outputs(7618) <= '0';
    layer2_outputs(7619) <= '1';
    layer2_outputs(7620) <= a and not b;
    layer2_outputs(7621) <= not b;
    layer2_outputs(7622) <= not b;
    layer2_outputs(7623) <= not (a or b);
    layer2_outputs(7624) <= b and not a;
    layer2_outputs(7625) <= a xor b;
    layer2_outputs(7626) <= not b or a;
    layer2_outputs(7627) <= '0';
    layer2_outputs(7628) <= not b;
    layer2_outputs(7629) <= '0';
    layer2_outputs(7630) <= not b;
    layer2_outputs(7631) <= not a or b;
    layer2_outputs(7632) <= a and not b;
    layer2_outputs(7633) <= not (a or b);
    layer2_outputs(7634) <= not b or a;
    layer2_outputs(7635) <= a and b;
    layer2_outputs(7636) <= not a or b;
    layer2_outputs(7637) <= a;
    layer2_outputs(7638) <= not (a xor b);
    layer2_outputs(7639) <= not b or a;
    layer2_outputs(7640) <= '0';
    layer2_outputs(7641) <= a and b;
    layer2_outputs(7642) <= a;
    layer2_outputs(7643) <= not b or a;
    layer2_outputs(7644) <= not (a or b);
    layer2_outputs(7645) <= a;
    layer2_outputs(7646) <= b;
    layer2_outputs(7647) <= not b;
    layer2_outputs(7648) <= not a or b;
    layer2_outputs(7649) <= a;
    layer2_outputs(7650) <= not (a or b);
    layer2_outputs(7651) <= a xor b;
    layer2_outputs(7652) <= '1';
    layer2_outputs(7653) <= not a or b;
    layer2_outputs(7654) <= not b;
    layer2_outputs(7655) <= '1';
    layer2_outputs(7656) <= a;
    layer2_outputs(7657) <= a xor b;
    layer2_outputs(7658) <= not a or b;
    layer2_outputs(7659) <= not a or b;
    layer2_outputs(7660) <= not b;
    layer2_outputs(7661) <= a and not b;
    layer2_outputs(7662) <= b;
    layer2_outputs(7663) <= a and b;
    layer2_outputs(7664) <= '1';
    layer2_outputs(7665) <= a and not b;
    layer2_outputs(7666) <= not a;
    layer2_outputs(7667) <= a and not b;
    layer2_outputs(7668) <= b;
    layer2_outputs(7669) <= a and b;
    layer2_outputs(7670) <= not b;
    layer2_outputs(7671) <= a or b;
    layer2_outputs(7672) <= '1';
    layer2_outputs(7673) <= not (a and b);
    layer2_outputs(7674) <= not a;
    layer2_outputs(7675) <= '0';
    layer2_outputs(7676) <= not a;
    layer2_outputs(7677) <= a and b;
    layer2_outputs(7678) <= not a;
    layer2_outputs(7679) <= '1';
    layer2_outputs(7680) <= b;
    layer2_outputs(7681) <= not b;
    layer2_outputs(7682) <= a and not b;
    layer2_outputs(7683) <= not b or a;
    layer2_outputs(7684) <= not b or a;
    layer2_outputs(7685) <= a and b;
    layer2_outputs(7686) <= b;
    layer2_outputs(7687) <= not (a and b);
    layer2_outputs(7688) <= not b or a;
    layer2_outputs(7689) <= not a;
    layer2_outputs(7690) <= not b;
    layer2_outputs(7691) <= not a;
    layer2_outputs(7692) <= not b;
    layer2_outputs(7693) <= '0';
    layer2_outputs(7694) <= b and not a;
    layer2_outputs(7695) <= '1';
    layer2_outputs(7696) <= a and b;
    layer2_outputs(7697) <= a and b;
    layer2_outputs(7698) <= a and b;
    layer2_outputs(7699) <= a and b;
    layer2_outputs(7700) <= a;
    layer2_outputs(7701) <= a or b;
    layer2_outputs(7702) <= b and not a;
    layer2_outputs(7703) <= '0';
    layer2_outputs(7704) <= not a or b;
    layer2_outputs(7705) <= a;
    layer2_outputs(7706) <= '1';
    layer2_outputs(7707) <= '1';
    layer2_outputs(7708) <= a and not b;
    layer2_outputs(7709) <= '0';
    layer2_outputs(7710) <= a and b;
    layer2_outputs(7711) <= a;
    layer2_outputs(7712) <= a and b;
    layer2_outputs(7713) <= not b;
    layer2_outputs(7714) <= b and not a;
    layer2_outputs(7715) <= a;
    layer2_outputs(7716) <= not b or a;
    layer2_outputs(7717) <= a or b;
    layer2_outputs(7718) <= not a;
    layer2_outputs(7719) <= a or b;
    layer2_outputs(7720) <= a and b;
    layer2_outputs(7721) <= not b or a;
    layer2_outputs(7722) <= not a or b;
    layer2_outputs(7723) <= b;
    layer2_outputs(7724) <= a;
    layer2_outputs(7725) <= b;
    layer2_outputs(7726) <= b;
    layer2_outputs(7727) <= not b;
    layer2_outputs(7728) <= not (a and b);
    layer2_outputs(7729) <= b and not a;
    layer2_outputs(7730) <= not (a or b);
    layer2_outputs(7731) <= b and not a;
    layer2_outputs(7732) <= '1';
    layer2_outputs(7733) <= not a;
    layer2_outputs(7734) <= a and not b;
    layer2_outputs(7735) <= not a or b;
    layer2_outputs(7736) <= not (a xor b);
    layer2_outputs(7737) <= b and not a;
    layer2_outputs(7738) <= b and not a;
    layer2_outputs(7739) <= not b;
    layer2_outputs(7740) <= not (a or b);
    layer2_outputs(7741) <= a and not b;
    layer2_outputs(7742) <= not b;
    layer2_outputs(7743) <= b and not a;
    layer2_outputs(7744) <= not b or a;
    layer2_outputs(7745) <= '1';
    layer2_outputs(7746) <= not b or a;
    layer2_outputs(7747) <= not a;
    layer2_outputs(7748) <= not a or b;
    layer2_outputs(7749) <= not b or a;
    layer2_outputs(7750) <= a or b;
    layer2_outputs(7751) <= b;
    layer2_outputs(7752) <= '1';
    layer2_outputs(7753) <= a and b;
    layer2_outputs(7754) <= not b;
    layer2_outputs(7755) <= '0';
    layer2_outputs(7756) <= not a;
    layer2_outputs(7757) <= a;
    layer2_outputs(7758) <= a;
    layer2_outputs(7759) <= not a;
    layer2_outputs(7760) <= not b;
    layer2_outputs(7761) <= a;
    layer2_outputs(7762) <= not a;
    layer2_outputs(7763) <= not a or b;
    layer2_outputs(7764) <= not a or b;
    layer2_outputs(7765) <= '1';
    layer2_outputs(7766) <= a and b;
    layer2_outputs(7767) <= b and not a;
    layer2_outputs(7768) <= not b or a;
    layer2_outputs(7769) <= not b;
    layer2_outputs(7770) <= a or b;
    layer2_outputs(7771) <= not (a or b);
    layer2_outputs(7772) <= b and not a;
    layer2_outputs(7773) <= not a;
    layer2_outputs(7774) <= b;
    layer2_outputs(7775) <= a xor b;
    layer2_outputs(7776) <= a;
    layer2_outputs(7777) <= a and not b;
    layer2_outputs(7778) <= not (a or b);
    layer2_outputs(7779) <= not b;
    layer2_outputs(7780) <= a and b;
    layer2_outputs(7781) <= not b or a;
    layer2_outputs(7782) <= not (a or b);
    layer2_outputs(7783) <= not b;
    layer2_outputs(7784) <= not b;
    layer2_outputs(7785) <= b and not a;
    layer2_outputs(7786) <= b and not a;
    layer2_outputs(7787) <= '1';
    layer2_outputs(7788) <= a;
    layer2_outputs(7789) <= not (a or b);
    layer2_outputs(7790) <= not b or a;
    layer2_outputs(7791) <= b;
    layer2_outputs(7792) <= not a;
    layer2_outputs(7793) <= b;
    layer2_outputs(7794) <= b;
    layer2_outputs(7795) <= not b or a;
    layer2_outputs(7796) <= not b or a;
    layer2_outputs(7797) <= a;
    layer2_outputs(7798) <= not (a or b);
    layer2_outputs(7799) <= not a or b;
    layer2_outputs(7800) <= b and not a;
    layer2_outputs(7801) <= not b;
    layer2_outputs(7802) <= not (a or b);
    layer2_outputs(7803) <= not a or b;
    layer2_outputs(7804) <= b and not a;
    layer2_outputs(7805) <= '0';
    layer2_outputs(7806) <= not a;
    layer2_outputs(7807) <= not b;
    layer2_outputs(7808) <= '1';
    layer2_outputs(7809) <= a;
    layer2_outputs(7810) <= a;
    layer2_outputs(7811) <= a and not b;
    layer2_outputs(7812) <= a;
    layer2_outputs(7813) <= not b;
    layer2_outputs(7814) <= not b;
    layer2_outputs(7815) <= b;
    layer2_outputs(7816) <= not b or a;
    layer2_outputs(7817) <= a or b;
    layer2_outputs(7818) <= not b;
    layer2_outputs(7819) <= a and not b;
    layer2_outputs(7820) <= a;
    layer2_outputs(7821) <= not b;
    layer2_outputs(7822) <= not b;
    layer2_outputs(7823) <= a and b;
    layer2_outputs(7824) <= not b;
    layer2_outputs(7825) <= a or b;
    layer2_outputs(7826) <= not b;
    layer2_outputs(7827) <= not a or b;
    layer2_outputs(7828) <= '0';
    layer2_outputs(7829) <= '1';
    layer2_outputs(7830) <= not (a or b);
    layer2_outputs(7831) <= b;
    layer2_outputs(7832) <= not b or a;
    layer2_outputs(7833) <= not (a and b);
    layer2_outputs(7834) <= not (a or b);
    layer2_outputs(7835) <= '1';
    layer2_outputs(7836) <= not (a and b);
    layer2_outputs(7837) <= not (a or b);
    layer2_outputs(7838) <= not (a xor b);
    layer2_outputs(7839) <= a;
    layer2_outputs(7840) <= b and not a;
    layer2_outputs(7841) <= not (a xor b);
    layer2_outputs(7842) <= not (a and b);
    layer2_outputs(7843) <= '0';
    layer2_outputs(7844) <= b and not a;
    layer2_outputs(7845) <= b;
    layer2_outputs(7846) <= not a or b;
    layer2_outputs(7847) <= b;
    layer2_outputs(7848) <= b;
    layer2_outputs(7849) <= not b or a;
    layer2_outputs(7850) <= a;
    layer2_outputs(7851) <= a;
    layer2_outputs(7852) <= not (a xor b);
    layer2_outputs(7853) <= not b;
    layer2_outputs(7854) <= not a;
    layer2_outputs(7855) <= not a or b;
    layer2_outputs(7856) <= a and not b;
    layer2_outputs(7857) <= '1';
    layer2_outputs(7858) <= not b;
    layer2_outputs(7859) <= not (a and b);
    layer2_outputs(7860) <= a or b;
    layer2_outputs(7861) <= b and not a;
    layer2_outputs(7862) <= b;
    layer2_outputs(7863) <= a or b;
    layer2_outputs(7864) <= a or b;
    layer2_outputs(7865) <= b and not a;
    layer2_outputs(7866) <= a;
    layer2_outputs(7867) <= not (a xor b);
    layer2_outputs(7868) <= not a;
    layer2_outputs(7869) <= not b or a;
    layer2_outputs(7870) <= not (a or b);
    layer2_outputs(7871) <= a and b;
    layer2_outputs(7872) <= not b;
    layer2_outputs(7873) <= not a;
    layer2_outputs(7874) <= '1';
    layer2_outputs(7875) <= a;
    layer2_outputs(7876) <= a or b;
    layer2_outputs(7877) <= a and b;
    layer2_outputs(7878) <= not a;
    layer2_outputs(7879) <= a and not b;
    layer2_outputs(7880) <= b and not a;
    layer2_outputs(7881) <= '0';
    layer2_outputs(7882) <= not a or b;
    layer2_outputs(7883) <= not b;
    layer2_outputs(7884) <= not a or b;
    layer2_outputs(7885) <= b;
    layer2_outputs(7886) <= a or b;
    layer2_outputs(7887) <= not (a or b);
    layer2_outputs(7888) <= a or b;
    layer2_outputs(7889) <= not (a xor b);
    layer2_outputs(7890) <= a and not b;
    layer2_outputs(7891) <= '0';
    layer2_outputs(7892) <= not (a and b);
    layer2_outputs(7893) <= not b;
    layer2_outputs(7894) <= not b or a;
    layer2_outputs(7895) <= not b;
    layer2_outputs(7896) <= a or b;
    layer2_outputs(7897) <= b and not a;
    layer2_outputs(7898) <= not a;
    layer2_outputs(7899) <= a or b;
    layer2_outputs(7900) <= not b or a;
    layer2_outputs(7901) <= a;
    layer2_outputs(7902) <= '1';
    layer2_outputs(7903) <= b;
    layer2_outputs(7904) <= not (a and b);
    layer2_outputs(7905) <= '0';
    layer2_outputs(7906) <= a and not b;
    layer2_outputs(7907) <= b;
    layer2_outputs(7908) <= not a;
    layer2_outputs(7909) <= '1';
    layer2_outputs(7910) <= a and not b;
    layer2_outputs(7911) <= b and not a;
    layer2_outputs(7912) <= b and not a;
    layer2_outputs(7913) <= not a or b;
    layer2_outputs(7914) <= not (a and b);
    layer2_outputs(7915) <= b;
    layer2_outputs(7916) <= a;
    layer2_outputs(7917) <= not (a and b);
    layer2_outputs(7918) <= not a;
    layer2_outputs(7919) <= not b or a;
    layer2_outputs(7920) <= a or b;
    layer2_outputs(7921) <= not a or b;
    layer2_outputs(7922) <= '0';
    layer2_outputs(7923) <= '1';
    layer2_outputs(7924) <= b;
    layer2_outputs(7925) <= a and not b;
    layer2_outputs(7926) <= '1';
    layer2_outputs(7927) <= not (a xor b);
    layer2_outputs(7928) <= not (a and b);
    layer2_outputs(7929) <= a;
    layer2_outputs(7930) <= not a;
    layer2_outputs(7931) <= not a or b;
    layer2_outputs(7932) <= not (a and b);
    layer2_outputs(7933) <= not a;
    layer2_outputs(7934) <= not (a and b);
    layer2_outputs(7935) <= not a;
    layer2_outputs(7936) <= a or b;
    layer2_outputs(7937) <= not (a and b);
    layer2_outputs(7938) <= a;
    layer2_outputs(7939) <= not b;
    layer2_outputs(7940) <= b and not a;
    layer2_outputs(7941) <= a and b;
    layer2_outputs(7942) <= not a;
    layer2_outputs(7943) <= b and not a;
    layer2_outputs(7944) <= not a;
    layer2_outputs(7945) <= a;
    layer2_outputs(7946) <= not (a or b);
    layer2_outputs(7947) <= b;
    layer2_outputs(7948) <= a or b;
    layer2_outputs(7949) <= not (a and b);
    layer2_outputs(7950) <= not b or a;
    layer2_outputs(7951) <= a or b;
    layer2_outputs(7952) <= not b;
    layer2_outputs(7953) <= a and b;
    layer2_outputs(7954) <= not (a xor b);
    layer2_outputs(7955) <= not b;
    layer2_outputs(7956) <= a and not b;
    layer2_outputs(7957) <= a xor b;
    layer2_outputs(7958) <= '0';
    layer2_outputs(7959) <= a or b;
    layer2_outputs(7960) <= a and b;
    layer2_outputs(7961) <= '1';
    layer2_outputs(7962) <= not a;
    layer2_outputs(7963) <= '0';
    layer2_outputs(7964) <= not b or a;
    layer2_outputs(7965) <= a or b;
    layer2_outputs(7966) <= not (a or b);
    layer2_outputs(7967) <= a;
    layer2_outputs(7968) <= a xor b;
    layer2_outputs(7969) <= not a;
    layer2_outputs(7970) <= not (a or b);
    layer2_outputs(7971) <= '1';
    layer2_outputs(7972) <= not b;
    layer2_outputs(7973) <= not (a and b);
    layer2_outputs(7974) <= not a;
    layer2_outputs(7975) <= '0';
    layer2_outputs(7976) <= not (a and b);
    layer2_outputs(7977) <= a;
    layer2_outputs(7978) <= a;
    layer2_outputs(7979) <= b;
    layer2_outputs(7980) <= not (a xor b);
    layer2_outputs(7981) <= b;
    layer2_outputs(7982) <= not b;
    layer2_outputs(7983) <= not (a or b);
    layer2_outputs(7984) <= a;
    layer2_outputs(7985) <= b;
    layer2_outputs(7986) <= a or b;
    layer2_outputs(7987) <= a and b;
    layer2_outputs(7988) <= not b;
    layer2_outputs(7989) <= '0';
    layer2_outputs(7990) <= a and b;
    layer2_outputs(7991) <= b and not a;
    layer2_outputs(7992) <= not (a and b);
    layer2_outputs(7993) <= a and b;
    layer2_outputs(7994) <= not a or b;
    layer2_outputs(7995) <= '0';
    layer2_outputs(7996) <= a;
    layer2_outputs(7997) <= b;
    layer2_outputs(7998) <= a and not b;
    layer2_outputs(7999) <= a and b;
    layer2_outputs(8000) <= a;
    layer2_outputs(8001) <= not b or a;
    layer2_outputs(8002) <= b;
    layer2_outputs(8003) <= a or b;
    layer2_outputs(8004) <= a and b;
    layer2_outputs(8005) <= '1';
    layer2_outputs(8006) <= b;
    layer2_outputs(8007) <= '0';
    layer2_outputs(8008) <= not (a and b);
    layer2_outputs(8009) <= '0';
    layer2_outputs(8010) <= '1';
    layer2_outputs(8011) <= a and b;
    layer2_outputs(8012) <= not (a or b);
    layer2_outputs(8013) <= not b or a;
    layer2_outputs(8014) <= a;
    layer2_outputs(8015) <= not (a or b);
    layer2_outputs(8016) <= '0';
    layer2_outputs(8017) <= b and not a;
    layer2_outputs(8018) <= a and b;
    layer2_outputs(8019) <= a xor b;
    layer2_outputs(8020) <= not (a and b);
    layer2_outputs(8021) <= b and not a;
    layer2_outputs(8022) <= a or b;
    layer2_outputs(8023) <= not b;
    layer2_outputs(8024) <= a;
    layer2_outputs(8025) <= a and not b;
    layer2_outputs(8026) <= not (a and b);
    layer2_outputs(8027) <= not (a or b);
    layer2_outputs(8028) <= a and not b;
    layer2_outputs(8029) <= a and not b;
    layer2_outputs(8030) <= not a;
    layer2_outputs(8031) <= not a or b;
    layer2_outputs(8032) <= not b;
    layer2_outputs(8033) <= b and not a;
    layer2_outputs(8034) <= not b;
    layer2_outputs(8035) <= b;
    layer2_outputs(8036) <= b;
    layer2_outputs(8037) <= a;
    layer2_outputs(8038) <= a or b;
    layer2_outputs(8039) <= '1';
    layer2_outputs(8040) <= not (a and b);
    layer2_outputs(8041) <= a or b;
    layer2_outputs(8042) <= a;
    layer2_outputs(8043) <= a;
    layer2_outputs(8044) <= not b or a;
    layer2_outputs(8045) <= a and not b;
    layer2_outputs(8046) <= not b;
    layer2_outputs(8047) <= a and not b;
    layer2_outputs(8048) <= a and b;
    layer2_outputs(8049) <= not (a xor b);
    layer2_outputs(8050) <= not b;
    layer2_outputs(8051) <= a and b;
    layer2_outputs(8052) <= b;
    layer2_outputs(8053) <= not a;
    layer2_outputs(8054) <= '0';
    layer2_outputs(8055) <= not b or a;
    layer2_outputs(8056) <= not a;
    layer2_outputs(8057) <= '1';
    layer2_outputs(8058) <= b;
    layer2_outputs(8059) <= not b;
    layer2_outputs(8060) <= '1';
    layer2_outputs(8061) <= not b;
    layer2_outputs(8062) <= a and b;
    layer2_outputs(8063) <= b and not a;
    layer2_outputs(8064) <= b and not a;
    layer2_outputs(8065) <= b and not a;
    layer2_outputs(8066) <= not (a and b);
    layer2_outputs(8067) <= a and b;
    layer2_outputs(8068) <= not b;
    layer2_outputs(8069) <= not (a or b);
    layer2_outputs(8070) <= not b;
    layer2_outputs(8071) <= not b;
    layer2_outputs(8072) <= not b or a;
    layer2_outputs(8073) <= a and not b;
    layer2_outputs(8074) <= not a;
    layer2_outputs(8075) <= b;
    layer2_outputs(8076) <= a;
    layer2_outputs(8077) <= b;
    layer2_outputs(8078) <= not b;
    layer2_outputs(8079) <= b and not a;
    layer2_outputs(8080) <= '0';
    layer2_outputs(8081) <= a;
    layer2_outputs(8082) <= a or b;
    layer2_outputs(8083) <= not a;
    layer2_outputs(8084) <= '1';
    layer2_outputs(8085) <= a;
    layer2_outputs(8086) <= not b;
    layer2_outputs(8087) <= a;
    layer2_outputs(8088) <= not a;
    layer2_outputs(8089) <= not (a and b);
    layer2_outputs(8090) <= not (a xor b);
    layer2_outputs(8091) <= a;
    layer2_outputs(8092) <= not b or a;
    layer2_outputs(8093) <= a or b;
    layer2_outputs(8094) <= '0';
    layer2_outputs(8095) <= not (a xor b);
    layer2_outputs(8096) <= b;
    layer2_outputs(8097) <= a and b;
    layer2_outputs(8098) <= not a;
    layer2_outputs(8099) <= not (a and b);
    layer2_outputs(8100) <= a or b;
    layer2_outputs(8101) <= not (a xor b);
    layer2_outputs(8102) <= not a;
    layer2_outputs(8103) <= '1';
    layer2_outputs(8104) <= a or b;
    layer2_outputs(8105) <= not a;
    layer2_outputs(8106) <= a and b;
    layer2_outputs(8107) <= a and b;
    layer2_outputs(8108) <= not (a and b);
    layer2_outputs(8109) <= a;
    layer2_outputs(8110) <= not a;
    layer2_outputs(8111) <= not b;
    layer2_outputs(8112) <= b and not a;
    layer2_outputs(8113) <= not a;
    layer2_outputs(8114) <= b;
    layer2_outputs(8115) <= not b or a;
    layer2_outputs(8116) <= not a or b;
    layer2_outputs(8117) <= not (a or b);
    layer2_outputs(8118) <= not (a and b);
    layer2_outputs(8119) <= a and not b;
    layer2_outputs(8120) <= '1';
    layer2_outputs(8121) <= '1';
    layer2_outputs(8122) <= a or b;
    layer2_outputs(8123) <= a or b;
    layer2_outputs(8124) <= b;
    layer2_outputs(8125) <= '0';
    layer2_outputs(8126) <= a;
    layer2_outputs(8127) <= not (a and b);
    layer2_outputs(8128) <= a and not b;
    layer2_outputs(8129) <= '0';
    layer2_outputs(8130) <= not a or b;
    layer2_outputs(8131) <= a or b;
    layer2_outputs(8132) <= a;
    layer2_outputs(8133) <= '0';
    layer2_outputs(8134) <= a and not b;
    layer2_outputs(8135) <= not (a and b);
    layer2_outputs(8136) <= not b or a;
    layer2_outputs(8137) <= a or b;
    layer2_outputs(8138) <= b;
    layer2_outputs(8139) <= not b or a;
    layer2_outputs(8140) <= not (a or b);
    layer2_outputs(8141) <= b;
    layer2_outputs(8142) <= not (a xor b);
    layer2_outputs(8143) <= b;
    layer2_outputs(8144) <= b;
    layer2_outputs(8145) <= not a;
    layer2_outputs(8146) <= not (a or b);
    layer2_outputs(8147) <= b;
    layer2_outputs(8148) <= b and not a;
    layer2_outputs(8149) <= not b;
    layer2_outputs(8150) <= a;
    layer2_outputs(8151) <= not a or b;
    layer2_outputs(8152) <= a and b;
    layer2_outputs(8153) <= not (a xor b);
    layer2_outputs(8154) <= '1';
    layer2_outputs(8155) <= not (a or b);
    layer2_outputs(8156) <= a and not b;
    layer2_outputs(8157) <= a;
    layer2_outputs(8158) <= b;
    layer2_outputs(8159) <= a and not b;
    layer2_outputs(8160) <= not a;
    layer2_outputs(8161) <= not a or b;
    layer2_outputs(8162) <= not a;
    layer2_outputs(8163) <= not (a or b);
    layer2_outputs(8164) <= b;
    layer2_outputs(8165) <= b and not a;
    layer2_outputs(8166) <= a xor b;
    layer2_outputs(8167) <= a;
    layer2_outputs(8168) <= a and b;
    layer2_outputs(8169) <= not a;
    layer2_outputs(8170) <= not a or b;
    layer2_outputs(8171) <= a;
    layer2_outputs(8172) <= not a or b;
    layer2_outputs(8173) <= not b;
    layer2_outputs(8174) <= a or b;
    layer2_outputs(8175) <= a and b;
    layer2_outputs(8176) <= a;
    layer2_outputs(8177) <= a;
    layer2_outputs(8178) <= '0';
    layer2_outputs(8179) <= a and b;
    layer2_outputs(8180) <= not (a and b);
    layer2_outputs(8181) <= a or b;
    layer2_outputs(8182) <= not (a and b);
    layer2_outputs(8183) <= a;
    layer2_outputs(8184) <= a;
    layer2_outputs(8185) <= not a or b;
    layer2_outputs(8186) <= a or b;
    layer2_outputs(8187) <= a;
    layer2_outputs(8188) <= not (a or b);
    layer2_outputs(8189) <= a;
    layer2_outputs(8190) <= a and b;
    layer2_outputs(8191) <= not a;
    layer2_outputs(8192) <= b;
    layer2_outputs(8193) <= a and b;
    layer2_outputs(8194) <= a or b;
    layer2_outputs(8195) <= a and b;
    layer2_outputs(8196) <= not (a xor b);
    layer2_outputs(8197) <= not (a or b);
    layer2_outputs(8198) <= '1';
    layer2_outputs(8199) <= a or b;
    layer2_outputs(8200) <= a or b;
    layer2_outputs(8201) <= '0';
    layer2_outputs(8202) <= a;
    layer2_outputs(8203) <= not (a and b);
    layer2_outputs(8204) <= a or b;
    layer2_outputs(8205) <= a;
    layer2_outputs(8206) <= a;
    layer2_outputs(8207) <= b;
    layer2_outputs(8208) <= b and not a;
    layer2_outputs(8209) <= a and b;
    layer2_outputs(8210) <= a and b;
    layer2_outputs(8211) <= '1';
    layer2_outputs(8212) <= '0';
    layer2_outputs(8213) <= a;
    layer2_outputs(8214) <= not b;
    layer2_outputs(8215) <= not b;
    layer2_outputs(8216) <= b;
    layer2_outputs(8217) <= a and b;
    layer2_outputs(8218) <= not (a or b);
    layer2_outputs(8219) <= not (a or b);
    layer2_outputs(8220) <= not a;
    layer2_outputs(8221) <= not b or a;
    layer2_outputs(8222) <= b;
    layer2_outputs(8223) <= b and not a;
    layer2_outputs(8224) <= b;
    layer2_outputs(8225) <= '1';
    layer2_outputs(8226) <= not a or b;
    layer2_outputs(8227) <= not a or b;
    layer2_outputs(8228) <= b;
    layer2_outputs(8229) <= not b;
    layer2_outputs(8230) <= not (a and b);
    layer2_outputs(8231) <= a;
    layer2_outputs(8232) <= a;
    layer2_outputs(8233) <= not b;
    layer2_outputs(8234) <= a;
    layer2_outputs(8235) <= a and b;
    layer2_outputs(8236) <= '1';
    layer2_outputs(8237) <= not a or b;
    layer2_outputs(8238) <= a or b;
    layer2_outputs(8239) <= a or b;
    layer2_outputs(8240) <= a;
    layer2_outputs(8241) <= not (a and b);
    layer2_outputs(8242) <= not b or a;
    layer2_outputs(8243) <= '0';
    layer2_outputs(8244) <= '1';
    layer2_outputs(8245) <= a;
    layer2_outputs(8246) <= b and not a;
    layer2_outputs(8247) <= b and not a;
    layer2_outputs(8248) <= b;
    layer2_outputs(8249) <= a;
    layer2_outputs(8250) <= not (a or b);
    layer2_outputs(8251) <= b and not a;
    layer2_outputs(8252) <= a and b;
    layer2_outputs(8253) <= not b or a;
    layer2_outputs(8254) <= a and not b;
    layer2_outputs(8255) <= not (a or b);
    layer2_outputs(8256) <= a or b;
    layer2_outputs(8257) <= not a;
    layer2_outputs(8258) <= b;
    layer2_outputs(8259) <= a xor b;
    layer2_outputs(8260) <= a or b;
    layer2_outputs(8261) <= not a;
    layer2_outputs(8262) <= not a or b;
    layer2_outputs(8263) <= a and b;
    layer2_outputs(8264) <= not (a xor b);
    layer2_outputs(8265) <= not a;
    layer2_outputs(8266) <= b and not a;
    layer2_outputs(8267) <= a xor b;
    layer2_outputs(8268) <= b;
    layer2_outputs(8269) <= a or b;
    layer2_outputs(8270) <= not a or b;
    layer2_outputs(8271) <= a;
    layer2_outputs(8272) <= not a;
    layer2_outputs(8273) <= not b or a;
    layer2_outputs(8274) <= a and not b;
    layer2_outputs(8275) <= not b or a;
    layer2_outputs(8276) <= not a or b;
    layer2_outputs(8277) <= b and not a;
    layer2_outputs(8278) <= not (a or b);
    layer2_outputs(8279) <= '1';
    layer2_outputs(8280) <= not (a and b);
    layer2_outputs(8281) <= not b;
    layer2_outputs(8282) <= not b or a;
    layer2_outputs(8283) <= b;
    layer2_outputs(8284) <= a;
    layer2_outputs(8285) <= not b;
    layer2_outputs(8286) <= not (a xor b);
    layer2_outputs(8287) <= b and not a;
    layer2_outputs(8288) <= a;
    layer2_outputs(8289) <= not a or b;
    layer2_outputs(8290) <= not a;
    layer2_outputs(8291) <= not (a and b);
    layer2_outputs(8292) <= b and not a;
    layer2_outputs(8293) <= a;
    layer2_outputs(8294) <= not (a and b);
    layer2_outputs(8295) <= a and b;
    layer2_outputs(8296) <= not b;
    layer2_outputs(8297) <= not b or a;
    layer2_outputs(8298) <= b;
    layer2_outputs(8299) <= a or b;
    layer2_outputs(8300) <= a and b;
    layer2_outputs(8301) <= a and b;
    layer2_outputs(8302) <= not (a or b);
    layer2_outputs(8303) <= '0';
    layer2_outputs(8304) <= b and not a;
    layer2_outputs(8305) <= a and b;
    layer2_outputs(8306) <= not a or b;
    layer2_outputs(8307) <= b;
    layer2_outputs(8308) <= a;
    layer2_outputs(8309) <= a;
    layer2_outputs(8310) <= a;
    layer2_outputs(8311) <= a xor b;
    layer2_outputs(8312) <= not (a or b);
    layer2_outputs(8313) <= not (a or b);
    layer2_outputs(8314) <= not a;
    layer2_outputs(8315) <= not a;
    layer2_outputs(8316) <= not (a or b);
    layer2_outputs(8317) <= a and not b;
    layer2_outputs(8318) <= a and not b;
    layer2_outputs(8319) <= not a;
    layer2_outputs(8320) <= not (a or b);
    layer2_outputs(8321) <= a and not b;
    layer2_outputs(8322) <= a xor b;
    layer2_outputs(8323) <= a and b;
    layer2_outputs(8324) <= b and not a;
    layer2_outputs(8325) <= a and not b;
    layer2_outputs(8326) <= not b or a;
    layer2_outputs(8327) <= a and b;
    layer2_outputs(8328) <= b and not a;
    layer2_outputs(8329) <= not a or b;
    layer2_outputs(8330) <= a or b;
    layer2_outputs(8331) <= a;
    layer2_outputs(8332) <= not b;
    layer2_outputs(8333) <= a and b;
    layer2_outputs(8334) <= '1';
    layer2_outputs(8335) <= a or b;
    layer2_outputs(8336) <= not (a or b);
    layer2_outputs(8337) <= not a;
    layer2_outputs(8338) <= not a or b;
    layer2_outputs(8339) <= a;
    layer2_outputs(8340) <= not a;
    layer2_outputs(8341) <= a or b;
    layer2_outputs(8342) <= a and b;
    layer2_outputs(8343) <= a and not b;
    layer2_outputs(8344) <= a;
    layer2_outputs(8345) <= not (a or b);
    layer2_outputs(8346) <= a and not b;
    layer2_outputs(8347) <= not b or a;
    layer2_outputs(8348) <= not (a or b);
    layer2_outputs(8349) <= b;
    layer2_outputs(8350) <= a;
    layer2_outputs(8351) <= not a or b;
    layer2_outputs(8352) <= not b;
    layer2_outputs(8353) <= not a;
    layer2_outputs(8354) <= '0';
    layer2_outputs(8355) <= not (a and b);
    layer2_outputs(8356) <= '0';
    layer2_outputs(8357) <= not (a or b);
    layer2_outputs(8358) <= a or b;
    layer2_outputs(8359) <= a or b;
    layer2_outputs(8360) <= '0';
    layer2_outputs(8361) <= not (a and b);
    layer2_outputs(8362) <= not a;
    layer2_outputs(8363) <= a and b;
    layer2_outputs(8364) <= a;
    layer2_outputs(8365) <= a xor b;
    layer2_outputs(8366) <= not a or b;
    layer2_outputs(8367) <= a or b;
    layer2_outputs(8368) <= a;
    layer2_outputs(8369) <= not a or b;
    layer2_outputs(8370) <= a and b;
    layer2_outputs(8371) <= a xor b;
    layer2_outputs(8372) <= not a or b;
    layer2_outputs(8373) <= not (a and b);
    layer2_outputs(8374) <= a or b;
    layer2_outputs(8375) <= not b;
    layer2_outputs(8376) <= a;
    layer2_outputs(8377) <= a and b;
    layer2_outputs(8378) <= not b or a;
    layer2_outputs(8379) <= not b or a;
    layer2_outputs(8380) <= '0';
    layer2_outputs(8381) <= b and not a;
    layer2_outputs(8382) <= not (a and b);
    layer2_outputs(8383) <= a and b;
    layer2_outputs(8384) <= '1';
    layer2_outputs(8385) <= not (a and b);
    layer2_outputs(8386) <= not a or b;
    layer2_outputs(8387) <= not a;
    layer2_outputs(8388) <= not (a and b);
    layer2_outputs(8389) <= not a or b;
    layer2_outputs(8390) <= a and not b;
    layer2_outputs(8391) <= '1';
    layer2_outputs(8392) <= not b or a;
    layer2_outputs(8393) <= a and b;
    layer2_outputs(8394) <= not (a or b);
    layer2_outputs(8395) <= '0';
    layer2_outputs(8396) <= a and b;
    layer2_outputs(8397) <= '0';
    layer2_outputs(8398) <= a or b;
    layer2_outputs(8399) <= b and not a;
    layer2_outputs(8400) <= b;
    layer2_outputs(8401) <= a or b;
    layer2_outputs(8402) <= a and b;
    layer2_outputs(8403) <= a;
    layer2_outputs(8404) <= not (a and b);
    layer2_outputs(8405) <= not (a or b);
    layer2_outputs(8406) <= b;
    layer2_outputs(8407) <= '1';
    layer2_outputs(8408) <= not b or a;
    layer2_outputs(8409) <= a or b;
    layer2_outputs(8410) <= not (a or b);
    layer2_outputs(8411) <= not (a and b);
    layer2_outputs(8412) <= not b or a;
    layer2_outputs(8413) <= '1';
    layer2_outputs(8414) <= '0';
    layer2_outputs(8415) <= '1';
    layer2_outputs(8416) <= not (a xor b);
    layer2_outputs(8417) <= b and not a;
    layer2_outputs(8418) <= not (a or b);
    layer2_outputs(8419) <= '1';
    layer2_outputs(8420) <= b and not a;
    layer2_outputs(8421) <= not b;
    layer2_outputs(8422) <= b and not a;
    layer2_outputs(8423) <= not a or b;
    layer2_outputs(8424) <= b;
    layer2_outputs(8425) <= a;
    layer2_outputs(8426) <= not b or a;
    layer2_outputs(8427) <= not a or b;
    layer2_outputs(8428) <= not a or b;
    layer2_outputs(8429) <= a xor b;
    layer2_outputs(8430) <= not b or a;
    layer2_outputs(8431) <= a;
    layer2_outputs(8432) <= a;
    layer2_outputs(8433) <= a and b;
    layer2_outputs(8434) <= not b or a;
    layer2_outputs(8435) <= a and not b;
    layer2_outputs(8436) <= '1';
    layer2_outputs(8437) <= b;
    layer2_outputs(8438) <= a;
    layer2_outputs(8439) <= a and not b;
    layer2_outputs(8440) <= not b or a;
    layer2_outputs(8441) <= not (a and b);
    layer2_outputs(8442) <= not (a and b);
    layer2_outputs(8443) <= not a or b;
    layer2_outputs(8444) <= not b or a;
    layer2_outputs(8445) <= not b;
    layer2_outputs(8446) <= a;
    layer2_outputs(8447) <= not a;
    layer2_outputs(8448) <= a or b;
    layer2_outputs(8449) <= a or b;
    layer2_outputs(8450) <= not b;
    layer2_outputs(8451) <= not (a and b);
    layer2_outputs(8452) <= a;
    layer2_outputs(8453) <= not a;
    layer2_outputs(8454) <= not (a and b);
    layer2_outputs(8455) <= not (a xor b);
    layer2_outputs(8456) <= not b;
    layer2_outputs(8457) <= a and b;
    layer2_outputs(8458) <= not (a and b);
    layer2_outputs(8459) <= a and not b;
    layer2_outputs(8460) <= a or b;
    layer2_outputs(8461) <= '1';
    layer2_outputs(8462) <= not a or b;
    layer2_outputs(8463) <= not b;
    layer2_outputs(8464) <= not (a or b);
    layer2_outputs(8465) <= not b;
    layer2_outputs(8466) <= a and not b;
    layer2_outputs(8467) <= b;
    layer2_outputs(8468) <= b and not a;
    layer2_outputs(8469) <= b;
    layer2_outputs(8470) <= not a;
    layer2_outputs(8471) <= b;
    layer2_outputs(8472) <= a and not b;
    layer2_outputs(8473) <= a xor b;
    layer2_outputs(8474) <= a and not b;
    layer2_outputs(8475) <= a and not b;
    layer2_outputs(8476) <= a and not b;
    layer2_outputs(8477) <= not b;
    layer2_outputs(8478) <= a and not b;
    layer2_outputs(8479) <= a and b;
    layer2_outputs(8480) <= a or b;
    layer2_outputs(8481) <= '1';
    layer2_outputs(8482) <= a;
    layer2_outputs(8483) <= a and b;
    layer2_outputs(8484) <= not a;
    layer2_outputs(8485) <= not a;
    layer2_outputs(8486) <= '0';
    layer2_outputs(8487) <= a or b;
    layer2_outputs(8488) <= not b;
    layer2_outputs(8489) <= a and not b;
    layer2_outputs(8490) <= b;
    layer2_outputs(8491) <= a and b;
    layer2_outputs(8492) <= not a or b;
    layer2_outputs(8493) <= not (a or b);
    layer2_outputs(8494) <= not b or a;
    layer2_outputs(8495) <= a or b;
    layer2_outputs(8496) <= b and not a;
    layer2_outputs(8497) <= a or b;
    layer2_outputs(8498) <= not b;
    layer2_outputs(8499) <= not (a and b);
    layer2_outputs(8500) <= not b or a;
    layer2_outputs(8501) <= not a;
    layer2_outputs(8502) <= a and not b;
    layer2_outputs(8503) <= a xor b;
    layer2_outputs(8504) <= a and not b;
    layer2_outputs(8505) <= not a;
    layer2_outputs(8506) <= a;
    layer2_outputs(8507) <= a;
    layer2_outputs(8508) <= b;
    layer2_outputs(8509) <= a and not b;
    layer2_outputs(8510) <= not b or a;
    layer2_outputs(8511) <= a;
    layer2_outputs(8512) <= a;
    layer2_outputs(8513) <= a;
    layer2_outputs(8514) <= not b;
    layer2_outputs(8515) <= not b or a;
    layer2_outputs(8516) <= not (a and b);
    layer2_outputs(8517) <= a;
    layer2_outputs(8518) <= not a or b;
    layer2_outputs(8519) <= a and b;
    layer2_outputs(8520) <= not b;
    layer2_outputs(8521) <= not a;
    layer2_outputs(8522) <= '0';
    layer2_outputs(8523) <= a;
    layer2_outputs(8524) <= not b or a;
    layer2_outputs(8525) <= not a or b;
    layer2_outputs(8526) <= b;
    layer2_outputs(8527) <= a and b;
    layer2_outputs(8528) <= '0';
    layer2_outputs(8529) <= a;
    layer2_outputs(8530) <= not a;
    layer2_outputs(8531) <= a and b;
    layer2_outputs(8532) <= a and not b;
    layer2_outputs(8533) <= '1';
    layer2_outputs(8534) <= not (a and b);
    layer2_outputs(8535) <= a xor b;
    layer2_outputs(8536) <= '0';
    layer2_outputs(8537) <= not b;
    layer2_outputs(8538) <= not b;
    layer2_outputs(8539) <= not b or a;
    layer2_outputs(8540) <= b;
    layer2_outputs(8541) <= not (a and b);
    layer2_outputs(8542) <= '1';
    layer2_outputs(8543) <= '1';
    layer2_outputs(8544) <= not a;
    layer2_outputs(8545) <= '1';
    layer2_outputs(8546) <= not b or a;
    layer2_outputs(8547) <= a;
    layer2_outputs(8548) <= not b;
    layer2_outputs(8549) <= not a;
    layer2_outputs(8550) <= b;
    layer2_outputs(8551) <= a;
    layer2_outputs(8552) <= not (a and b);
    layer2_outputs(8553) <= not a or b;
    layer2_outputs(8554) <= '0';
    layer2_outputs(8555) <= a;
    layer2_outputs(8556) <= a and b;
    layer2_outputs(8557) <= not b;
    layer2_outputs(8558) <= not b or a;
    layer2_outputs(8559) <= not (a and b);
    layer2_outputs(8560) <= b;
    layer2_outputs(8561) <= b and not a;
    layer2_outputs(8562) <= a and not b;
    layer2_outputs(8563) <= not b or a;
    layer2_outputs(8564) <= '1';
    layer2_outputs(8565) <= not a or b;
    layer2_outputs(8566) <= '1';
    layer2_outputs(8567) <= a;
    layer2_outputs(8568) <= b;
    layer2_outputs(8569) <= not a or b;
    layer2_outputs(8570) <= a and b;
    layer2_outputs(8571) <= b;
    layer2_outputs(8572) <= b;
    layer2_outputs(8573) <= b;
    layer2_outputs(8574) <= '1';
    layer2_outputs(8575) <= not a;
    layer2_outputs(8576) <= '0';
    layer2_outputs(8577) <= not b;
    layer2_outputs(8578) <= b;
    layer2_outputs(8579) <= a and b;
    layer2_outputs(8580) <= not b;
    layer2_outputs(8581) <= not b;
    layer2_outputs(8582) <= not a;
    layer2_outputs(8583) <= b;
    layer2_outputs(8584) <= '1';
    layer2_outputs(8585) <= not a;
    layer2_outputs(8586) <= b;
    layer2_outputs(8587) <= a and b;
    layer2_outputs(8588) <= '1';
    layer2_outputs(8589) <= b;
    layer2_outputs(8590) <= not (a xor b);
    layer2_outputs(8591) <= not a or b;
    layer2_outputs(8592) <= not a;
    layer2_outputs(8593) <= a and b;
    layer2_outputs(8594) <= b and not a;
    layer2_outputs(8595) <= not (a xor b);
    layer2_outputs(8596) <= b and not a;
    layer2_outputs(8597) <= '0';
    layer2_outputs(8598) <= not a;
    layer2_outputs(8599) <= not b;
    layer2_outputs(8600) <= not b or a;
    layer2_outputs(8601) <= a or b;
    layer2_outputs(8602) <= not a;
    layer2_outputs(8603) <= not b;
    layer2_outputs(8604) <= not a;
    layer2_outputs(8605) <= not (a and b);
    layer2_outputs(8606) <= a xor b;
    layer2_outputs(8607) <= b;
    layer2_outputs(8608) <= not b;
    layer2_outputs(8609) <= '0';
    layer2_outputs(8610) <= a or b;
    layer2_outputs(8611) <= not b or a;
    layer2_outputs(8612) <= not b or a;
    layer2_outputs(8613) <= not b or a;
    layer2_outputs(8614) <= '1';
    layer2_outputs(8615) <= a;
    layer2_outputs(8616) <= not b or a;
    layer2_outputs(8617) <= b and not a;
    layer2_outputs(8618) <= not b or a;
    layer2_outputs(8619) <= a or b;
    layer2_outputs(8620) <= a;
    layer2_outputs(8621) <= a or b;
    layer2_outputs(8622) <= a and b;
    layer2_outputs(8623) <= not (a xor b);
    layer2_outputs(8624) <= '1';
    layer2_outputs(8625) <= not (a xor b);
    layer2_outputs(8626) <= not (a and b);
    layer2_outputs(8627) <= not b or a;
    layer2_outputs(8628) <= a and not b;
    layer2_outputs(8629) <= not a;
    layer2_outputs(8630) <= not a;
    layer2_outputs(8631) <= a;
    layer2_outputs(8632) <= not b or a;
    layer2_outputs(8633) <= not (a xor b);
    layer2_outputs(8634) <= a;
    layer2_outputs(8635) <= not (a xor b);
    layer2_outputs(8636) <= b;
    layer2_outputs(8637) <= not b or a;
    layer2_outputs(8638) <= not b or a;
    layer2_outputs(8639) <= not b or a;
    layer2_outputs(8640) <= b and not a;
    layer2_outputs(8641) <= b;
    layer2_outputs(8642) <= not b or a;
    layer2_outputs(8643) <= not b;
    layer2_outputs(8644) <= not a or b;
    layer2_outputs(8645) <= a and not b;
    layer2_outputs(8646) <= not (a xor b);
    layer2_outputs(8647) <= not (a xor b);
    layer2_outputs(8648) <= a or b;
    layer2_outputs(8649) <= a and b;
    layer2_outputs(8650) <= a and not b;
    layer2_outputs(8651) <= not b or a;
    layer2_outputs(8652) <= not a;
    layer2_outputs(8653) <= a and b;
    layer2_outputs(8654) <= not b or a;
    layer2_outputs(8655) <= a or b;
    layer2_outputs(8656) <= not b or a;
    layer2_outputs(8657) <= b;
    layer2_outputs(8658) <= not (a or b);
    layer2_outputs(8659) <= a and b;
    layer2_outputs(8660) <= a;
    layer2_outputs(8661) <= a or b;
    layer2_outputs(8662) <= not (a and b);
    layer2_outputs(8663) <= b;
    layer2_outputs(8664) <= not (a xor b);
    layer2_outputs(8665) <= not b or a;
    layer2_outputs(8666) <= a;
    layer2_outputs(8667) <= a and not b;
    layer2_outputs(8668) <= '0';
    layer2_outputs(8669) <= not (a and b);
    layer2_outputs(8670) <= b and not a;
    layer2_outputs(8671) <= a and not b;
    layer2_outputs(8672) <= not a;
    layer2_outputs(8673) <= a and b;
    layer2_outputs(8674) <= b;
    layer2_outputs(8675) <= a;
    layer2_outputs(8676) <= b;
    layer2_outputs(8677) <= '0';
    layer2_outputs(8678) <= a and b;
    layer2_outputs(8679) <= a or b;
    layer2_outputs(8680) <= a;
    layer2_outputs(8681) <= not b;
    layer2_outputs(8682) <= a xor b;
    layer2_outputs(8683) <= not b;
    layer2_outputs(8684) <= b and not a;
    layer2_outputs(8685) <= not b or a;
    layer2_outputs(8686) <= not (a or b);
    layer2_outputs(8687) <= '1';
    layer2_outputs(8688) <= a and not b;
    layer2_outputs(8689) <= not b;
    layer2_outputs(8690) <= not a or b;
    layer2_outputs(8691) <= not (a or b);
    layer2_outputs(8692) <= b and not a;
    layer2_outputs(8693) <= not (a and b);
    layer2_outputs(8694) <= '1';
    layer2_outputs(8695) <= not (a or b);
    layer2_outputs(8696) <= not b;
    layer2_outputs(8697) <= a and b;
    layer2_outputs(8698) <= '0';
    layer2_outputs(8699) <= not a or b;
    layer2_outputs(8700) <= b;
    layer2_outputs(8701) <= b;
    layer2_outputs(8702) <= a xor b;
    layer2_outputs(8703) <= b;
    layer2_outputs(8704) <= not (a xor b);
    layer2_outputs(8705) <= not b or a;
    layer2_outputs(8706) <= b and not a;
    layer2_outputs(8707) <= a and b;
    layer2_outputs(8708) <= b;
    layer2_outputs(8709) <= not a or b;
    layer2_outputs(8710) <= a and not b;
    layer2_outputs(8711) <= a and not b;
    layer2_outputs(8712) <= a and not b;
    layer2_outputs(8713) <= not (a or b);
    layer2_outputs(8714) <= not (a and b);
    layer2_outputs(8715) <= not (a and b);
    layer2_outputs(8716) <= a;
    layer2_outputs(8717) <= a or b;
    layer2_outputs(8718) <= not a;
    layer2_outputs(8719) <= not a;
    layer2_outputs(8720) <= not (a xor b);
    layer2_outputs(8721) <= not (a or b);
    layer2_outputs(8722) <= b and not a;
    layer2_outputs(8723) <= not a;
    layer2_outputs(8724) <= a and b;
    layer2_outputs(8725) <= not (a xor b);
    layer2_outputs(8726) <= b;
    layer2_outputs(8727) <= not b or a;
    layer2_outputs(8728) <= not a;
    layer2_outputs(8729) <= not (a and b);
    layer2_outputs(8730) <= not a or b;
    layer2_outputs(8731) <= not b;
    layer2_outputs(8732) <= b and not a;
    layer2_outputs(8733) <= '0';
    layer2_outputs(8734) <= not a or b;
    layer2_outputs(8735) <= b;
    layer2_outputs(8736) <= '0';
    layer2_outputs(8737) <= not b;
    layer2_outputs(8738) <= not (a or b);
    layer2_outputs(8739) <= a and not b;
    layer2_outputs(8740) <= '1';
    layer2_outputs(8741) <= not a;
    layer2_outputs(8742) <= not (a xor b);
    layer2_outputs(8743) <= b and not a;
    layer2_outputs(8744) <= a and b;
    layer2_outputs(8745) <= b;
    layer2_outputs(8746) <= a and not b;
    layer2_outputs(8747) <= not a;
    layer2_outputs(8748) <= a and not b;
    layer2_outputs(8749) <= not a;
    layer2_outputs(8750) <= not a;
    layer2_outputs(8751) <= a and b;
    layer2_outputs(8752) <= not (a xor b);
    layer2_outputs(8753) <= not a;
    layer2_outputs(8754) <= b;
    layer2_outputs(8755) <= not b;
    layer2_outputs(8756) <= a and b;
    layer2_outputs(8757) <= a xor b;
    layer2_outputs(8758) <= b and not a;
    layer2_outputs(8759) <= not b;
    layer2_outputs(8760) <= not (a or b);
    layer2_outputs(8761) <= a and not b;
    layer2_outputs(8762) <= not (a and b);
    layer2_outputs(8763) <= a;
    layer2_outputs(8764) <= not (a and b);
    layer2_outputs(8765) <= not a or b;
    layer2_outputs(8766) <= not (a xor b);
    layer2_outputs(8767) <= '0';
    layer2_outputs(8768) <= not a or b;
    layer2_outputs(8769) <= not (a xor b);
    layer2_outputs(8770) <= a and not b;
    layer2_outputs(8771) <= not b or a;
    layer2_outputs(8772) <= '0';
    layer2_outputs(8773) <= not b;
    layer2_outputs(8774) <= not a or b;
    layer2_outputs(8775) <= not a or b;
    layer2_outputs(8776) <= not a;
    layer2_outputs(8777) <= not b;
    layer2_outputs(8778) <= a and not b;
    layer2_outputs(8779) <= b and not a;
    layer2_outputs(8780) <= '1';
    layer2_outputs(8781) <= '0';
    layer2_outputs(8782) <= not a;
    layer2_outputs(8783) <= a;
    layer2_outputs(8784) <= not b or a;
    layer2_outputs(8785) <= not (a or b);
    layer2_outputs(8786) <= b;
    layer2_outputs(8787) <= not a or b;
    layer2_outputs(8788) <= not (a or b);
    layer2_outputs(8789) <= not a;
    layer2_outputs(8790) <= a or b;
    layer2_outputs(8791) <= a;
    layer2_outputs(8792) <= a and b;
    layer2_outputs(8793) <= not a;
    layer2_outputs(8794) <= b;
    layer2_outputs(8795) <= not (a or b);
    layer2_outputs(8796) <= b and not a;
    layer2_outputs(8797) <= b and not a;
    layer2_outputs(8798) <= not (a or b);
    layer2_outputs(8799) <= not a or b;
    layer2_outputs(8800) <= not a;
    layer2_outputs(8801) <= not (a or b);
    layer2_outputs(8802) <= not a or b;
    layer2_outputs(8803) <= not (a xor b);
    layer2_outputs(8804) <= '0';
    layer2_outputs(8805) <= '1';
    layer2_outputs(8806) <= a;
    layer2_outputs(8807) <= not (a and b);
    layer2_outputs(8808) <= a xor b;
    layer2_outputs(8809) <= a;
    layer2_outputs(8810) <= not b;
    layer2_outputs(8811) <= a or b;
    layer2_outputs(8812) <= not b;
    layer2_outputs(8813) <= a or b;
    layer2_outputs(8814) <= a and b;
    layer2_outputs(8815) <= not a;
    layer2_outputs(8816) <= a and b;
    layer2_outputs(8817) <= not a or b;
    layer2_outputs(8818) <= not a;
    layer2_outputs(8819) <= b and not a;
    layer2_outputs(8820) <= not b;
    layer2_outputs(8821) <= '0';
    layer2_outputs(8822) <= not a;
    layer2_outputs(8823) <= a;
    layer2_outputs(8824) <= b and not a;
    layer2_outputs(8825) <= b and not a;
    layer2_outputs(8826) <= a xor b;
    layer2_outputs(8827) <= b and not a;
    layer2_outputs(8828) <= b and not a;
    layer2_outputs(8829) <= a or b;
    layer2_outputs(8830) <= a;
    layer2_outputs(8831) <= b;
    layer2_outputs(8832) <= b;
    layer2_outputs(8833) <= b;
    layer2_outputs(8834) <= a;
    layer2_outputs(8835) <= not (a or b);
    layer2_outputs(8836) <= not (a and b);
    layer2_outputs(8837) <= not a;
    layer2_outputs(8838) <= not a or b;
    layer2_outputs(8839) <= not a or b;
    layer2_outputs(8840) <= '0';
    layer2_outputs(8841) <= a xor b;
    layer2_outputs(8842) <= a and not b;
    layer2_outputs(8843) <= a xor b;
    layer2_outputs(8844) <= b;
    layer2_outputs(8845) <= '1';
    layer2_outputs(8846) <= '0';
    layer2_outputs(8847) <= not b or a;
    layer2_outputs(8848) <= not b or a;
    layer2_outputs(8849) <= not (a or b);
    layer2_outputs(8850) <= not b or a;
    layer2_outputs(8851) <= not b;
    layer2_outputs(8852) <= not b;
    layer2_outputs(8853) <= not (a and b);
    layer2_outputs(8854) <= b and not a;
    layer2_outputs(8855) <= a and b;
    layer2_outputs(8856) <= not (a xor b);
    layer2_outputs(8857) <= not a;
    layer2_outputs(8858) <= '1';
    layer2_outputs(8859) <= not a;
    layer2_outputs(8860) <= '0';
    layer2_outputs(8861) <= not (a or b);
    layer2_outputs(8862) <= not a;
    layer2_outputs(8863) <= a;
    layer2_outputs(8864) <= b;
    layer2_outputs(8865) <= a xor b;
    layer2_outputs(8866) <= not a or b;
    layer2_outputs(8867) <= not (a and b);
    layer2_outputs(8868) <= a and not b;
    layer2_outputs(8869) <= a;
    layer2_outputs(8870) <= a and b;
    layer2_outputs(8871) <= not b or a;
    layer2_outputs(8872) <= not (a xor b);
    layer2_outputs(8873) <= '0';
    layer2_outputs(8874) <= a and b;
    layer2_outputs(8875) <= not b;
    layer2_outputs(8876) <= a;
    layer2_outputs(8877) <= not a;
    layer2_outputs(8878) <= not a;
    layer2_outputs(8879) <= b and not a;
    layer2_outputs(8880) <= b and not a;
    layer2_outputs(8881) <= a;
    layer2_outputs(8882) <= not b or a;
    layer2_outputs(8883) <= not a or b;
    layer2_outputs(8884) <= not b or a;
    layer2_outputs(8885) <= a and not b;
    layer2_outputs(8886) <= '0';
    layer2_outputs(8887) <= a;
    layer2_outputs(8888) <= b;
    layer2_outputs(8889) <= not (a and b);
    layer2_outputs(8890) <= a and not b;
    layer2_outputs(8891) <= not (a xor b);
    layer2_outputs(8892) <= not (a and b);
    layer2_outputs(8893) <= not a;
    layer2_outputs(8894) <= not b or a;
    layer2_outputs(8895) <= '0';
    layer2_outputs(8896) <= b and not a;
    layer2_outputs(8897) <= '0';
    layer2_outputs(8898) <= not b or a;
    layer2_outputs(8899) <= not a or b;
    layer2_outputs(8900) <= a;
    layer2_outputs(8901) <= '0';
    layer2_outputs(8902) <= not b;
    layer2_outputs(8903) <= not b or a;
    layer2_outputs(8904) <= not a;
    layer2_outputs(8905) <= not b or a;
    layer2_outputs(8906) <= b and not a;
    layer2_outputs(8907) <= a and b;
    layer2_outputs(8908) <= not a or b;
    layer2_outputs(8909) <= b and not a;
    layer2_outputs(8910) <= a and b;
    layer2_outputs(8911) <= not b;
    layer2_outputs(8912) <= not b;
    layer2_outputs(8913) <= '1';
    layer2_outputs(8914) <= not b;
    layer2_outputs(8915) <= not (a or b);
    layer2_outputs(8916) <= a;
    layer2_outputs(8917) <= '1';
    layer2_outputs(8918) <= '1';
    layer2_outputs(8919) <= a and b;
    layer2_outputs(8920) <= not (a and b);
    layer2_outputs(8921) <= not b or a;
    layer2_outputs(8922) <= not b or a;
    layer2_outputs(8923) <= '0';
    layer2_outputs(8924) <= not a;
    layer2_outputs(8925) <= not b;
    layer2_outputs(8926) <= '1';
    layer2_outputs(8927) <= not (a and b);
    layer2_outputs(8928) <= not a or b;
    layer2_outputs(8929) <= a xor b;
    layer2_outputs(8930) <= not (a and b);
    layer2_outputs(8931) <= a;
    layer2_outputs(8932) <= '0';
    layer2_outputs(8933) <= a or b;
    layer2_outputs(8934) <= not b;
    layer2_outputs(8935) <= a and b;
    layer2_outputs(8936) <= b;
    layer2_outputs(8937) <= not a;
    layer2_outputs(8938) <= not b;
    layer2_outputs(8939) <= b;
    layer2_outputs(8940) <= b;
    layer2_outputs(8941) <= not a;
    layer2_outputs(8942) <= a and not b;
    layer2_outputs(8943) <= not (a and b);
    layer2_outputs(8944) <= '1';
    layer2_outputs(8945) <= not b or a;
    layer2_outputs(8946) <= not b or a;
    layer2_outputs(8947) <= a xor b;
    layer2_outputs(8948) <= b and not a;
    layer2_outputs(8949) <= '1';
    layer2_outputs(8950) <= a or b;
    layer2_outputs(8951) <= '0';
    layer2_outputs(8952) <= a and not b;
    layer2_outputs(8953) <= not (a and b);
    layer2_outputs(8954) <= a and not b;
    layer2_outputs(8955) <= b and not a;
    layer2_outputs(8956) <= a;
    layer2_outputs(8957) <= b and not a;
    layer2_outputs(8958) <= not (a or b);
    layer2_outputs(8959) <= a and not b;
    layer2_outputs(8960) <= a or b;
    layer2_outputs(8961) <= not b;
    layer2_outputs(8962) <= b;
    layer2_outputs(8963) <= not (a and b);
    layer2_outputs(8964) <= '1';
    layer2_outputs(8965) <= not (a and b);
    layer2_outputs(8966) <= not (a and b);
    layer2_outputs(8967) <= b and not a;
    layer2_outputs(8968) <= '0';
    layer2_outputs(8969) <= not b or a;
    layer2_outputs(8970) <= b and not a;
    layer2_outputs(8971) <= not b;
    layer2_outputs(8972) <= '1';
    layer2_outputs(8973) <= not b or a;
    layer2_outputs(8974) <= not b;
    layer2_outputs(8975) <= not (a and b);
    layer2_outputs(8976) <= a;
    layer2_outputs(8977) <= b and not a;
    layer2_outputs(8978) <= a xor b;
    layer2_outputs(8979) <= not a or b;
    layer2_outputs(8980) <= b;
    layer2_outputs(8981) <= a and not b;
    layer2_outputs(8982) <= b;
    layer2_outputs(8983) <= not a;
    layer2_outputs(8984) <= a and not b;
    layer2_outputs(8985) <= not (a or b);
    layer2_outputs(8986) <= a xor b;
    layer2_outputs(8987) <= a;
    layer2_outputs(8988) <= a;
    layer2_outputs(8989) <= a and b;
    layer2_outputs(8990) <= b and not a;
    layer2_outputs(8991) <= not (a or b);
    layer2_outputs(8992) <= a;
    layer2_outputs(8993) <= a and b;
    layer2_outputs(8994) <= a;
    layer2_outputs(8995) <= not (a and b);
    layer2_outputs(8996) <= b;
    layer2_outputs(8997) <= not b;
    layer2_outputs(8998) <= b;
    layer2_outputs(8999) <= not (a and b);
    layer2_outputs(9000) <= a and b;
    layer2_outputs(9001) <= b;
    layer2_outputs(9002) <= '0';
    layer2_outputs(9003) <= a;
    layer2_outputs(9004) <= '1';
    layer2_outputs(9005) <= not b or a;
    layer2_outputs(9006) <= not b or a;
    layer2_outputs(9007) <= a xor b;
    layer2_outputs(9008) <= not b;
    layer2_outputs(9009) <= b;
    layer2_outputs(9010) <= not a or b;
    layer2_outputs(9011) <= b;
    layer2_outputs(9012) <= b;
    layer2_outputs(9013) <= not a or b;
    layer2_outputs(9014) <= not (a or b);
    layer2_outputs(9015) <= a and not b;
    layer2_outputs(9016) <= not b or a;
    layer2_outputs(9017) <= '1';
    layer2_outputs(9018) <= b;
    layer2_outputs(9019) <= a;
    layer2_outputs(9020) <= a xor b;
    layer2_outputs(9021) <= a;
    layer2_outputs(9022) <= a and not b;
    layer2_outputs(9023) <= not (a xor b);
    layer2_outputs(9024) <= not a or b;
    layer2_outputs(9025) <= b and not a;
    layer2_outputs(9026) <= not (a or b);
    layer2_outputs(9027) <= '1';
    layer2_outputs(9028) <= not (a or b);
    layer2_outputs(9029) <= a xor b;
    layer2_outputs(9030) <= a;
    layer2_outputs(9031) <= not b or a;
    layer2_outputs(9032) <= not (a or b);
    layer2_outputs(9033) <= not (a or b);
    layer2_outputs(9034) <= a and b;
    layer2_outputs(9035) <= a and b;
    layer2_outputs(9036) <= a or b;
    layer2_outputs(9037) <= a;
    layer2_outputs(9038) <= '0';
    layer2_outputs(9039) <= not (a xor b);
    layer2_outputs(9040) <= not (a or b);
    layer2_outputs(9041) <= b and not a;
    layer2_outputs(9042) <= not b;
    layer2_outputs(9043) <= not (a or b);
    layer2_outputs(9044) <= b;
    layer2_outputs(9045) <= not a;
    layer2_outputs(9046) <= not (a and b);
    layer2_outputs(9047) <= not a;
    layer2_outputs(9048) <= b and not a;
    layer2_outputs(9049) <= not b;
    layer2_outputs(9050) <= not (a or b);
    layer2_outputs(9051) <= not a;
    layer2_outputs(9052) <= not a or b;
    layer2_outputs(9053) <= not (a or b);
    layer2_outputs(9054) <= not a;
    layer2_outputs(9055) <= not b;
    layer2_outputs(9056) <= a and b;
    layer2_outputs(9057) <= a and not b;
    layer2_outputs(9058) <= a xor b;
    layer2_outputs(9059) <= not b;
    layer2_outputs(9060) <= a and b;
    layer2_outputs(9061) <= a xor b;
    layer2_outputs(9062) <= '0';
    layer2_outputs(9063) <= a and not b;
    layer2_outputs(9064) <= not a or b;
    layer2_outputs(9065) <= '1';
    layer2_outputs(9066) <= not b;
    layer2_outputs(9067) <= b and not a;
    layer2_outputs(9068) <= not a or b;
    layer2_outputs(9069) <= not b;
    layer2_outputs(9070) <= b and not a;
    layer2_outputs(9071) <= not b or a;
    layer2_outputs(9072) <= a;
    layer2_outputs(9073) <= a and not b;
    layer2_outputs(9074) <= a or b;
    layer2_outputs(9075) <= not b or a;
    layer2_outputs(9076) <= not b;
    layer2_outputs(9077) <= not b;
    layer2_outputs(9078) <= b and not a;
    layer2_outputs(9079) <= not a or b;
    layer2_outputs(9080) <= b;
    layer2_outputs(9081) <= a xor b;
    layer2_outputs(9082) <= b;
    layer2_outputs(9083) <= '0';
    layer2_outputs(9084) <= b;
    layer2_outputs(9085) <= not a;
    layer2_outputs(9086) <= '0';
    layer2_outputs(9087) <= not (a or b);
    layer2_outputs(9088) <= b and not a;
    layer2_outputs(9089) <= not (a and b);
    layer2_outputs(9090) <= '0';
    layer2_outputs(9091) <= not b;
    layer2_outputs(9092) <= not (a and b);
    layer2_outputs(9093) <= b;
    layer2_outputs(9094) <= not a or b;
    layer2_outputs(9095) <= not (a or b);
    layer2_outputs(9096) <= a;
    layer2_outputs(9097) <= a and not b;
    layer2_outputs(9098) <= b and not a;
    layer2_outputs(9099) <= '1';
    layer2_outputs(9100) <= '1';
    layer2_outputs(9101) <= not b;
    layer2_outputs(9102) <= a and not b;
    layer2_outputs(9103) <= not a;
    layer2_outputs(9104) <= not a;
    layer2_outputs(9105) <= not b;
    layer2_outputs(9106) <= a and b;
    layer2_outputs(9107) <= not b or a;
    layer2_outputs(9108) <= '0';
    layer2_outputs(9109) <= not (a and b);
    layer2_outputs(9110) <= a and b;
    layer2_outputs(9111) <= b and not a;
    layer2_outputs(9112) <= b;
    layer2_outputs(9113) <= a and not b;
    layer2_outputs(9114) <= '0';
    layer2_outputs(9115) <= b;
    layer2_outputs(9116) <= '0';
    layer2_outputs(9117) <= b and not a;
    layer2_outputs(9118) <= a xor b;
    layer2_outputs(9119) <= a;
    layer2_outputs(9120) <= not b or a;
    layer2_outputs(9121) <= '1';
    layer2_outputs(9122) <= b and not a;
    layer2_outputs(9123) <= a;
    layer2_outputs(9124) <= b;
    layer2_outputs(9125) <= not b;
    layer2_outputs(9126) <= a;
    layer2_outputs(9127) <= a xor b;
    layer2_outputs(9128) <= not a or b;
    layer2_outputs(9129) <= b;
    layer2_outputs(9130) <= a or b;
    layer2_outputs(9131) <= not (a or b);
    layer2_outputs(9132) <= '1';
    layer2_outputs(9133) <= not b;
    layer2_outputs(9134) <= a and b;
    layer2_outputs(9135) <= not b or a;
    layer2_outputs(9136) <= '0';
    layer2_outputs(9137) <= not (a or b);
    layer2_outputs(9138) <= a and b;
    layer2_outputs(9139) <= b and not a;
    layer2_outputs(9140) <= not b;
    layer2_outputs(9141) <= b;
    layer2_outputs(9142) <= not (a or b);
    layer2_outputs(9143) <= not (a or b);
    layer2_outputs(9144) <= not b;
    layer2_outputs(9145) <= '1';
    layer2_outputs(9146) <= not a;
    layer2_outputs(9147) <= b and not a;
    layer2_outputs(9148) <= not (a and b);
    layer2_outputs(9149) <= not (a or b);
    layer2_outputs(9150) <= not a;
    layer2_outputs(9151) <= '1';
    layer2_outputs(9152) <= b and not a;
    layer2_outputs(9153) <= '0';
    layer2_outputs(9154) <= a or b;
    layer2_outputs(9155) <= not (a and b);
    layer2_outputs(9156) <= not (a and b);
    layer2_outputs(9157) <= not a or b;
    layer2_outputs(9158) <= not (a xor b);
    layer2_outputs(9159) <= not a;
    layer2_outputs(9160) <= a and not b;
    layer2_outputs(9161) <= a;
    layer2_outputs(9162) <= not b;
    layer2_outputs(9163) <= a xor b;
    layer2_outputs(9164) <= b;
    layer2_outputs(9165) <= not a;
    layer2_outputs(9166) <= not b or a;
    layer2_outputs(9167) <= b;
    layer2_outputs(9168) <= a or b;
    layer2_outputs(9169) <= a and not b;
    layer2_outputs(9170) <= a or b;
    layer2_outputs(9171) <= not b or a;
    layer2_outputs(9172) <= not b or a;
    layer2_outputs(9173) <= a;
    layer2_outputs(9174) <= a or b;
    layer2_outputs(9175) <= a or b;
    layer2_outputs(9176) <= a and not b;
    layer2_outputs(9177) <= not (a and b);
    layer2_outputs(9178) <= a;
    layer2_outputs(9179) <= a xor b;
    layer2_outputs(9180) <= b;
    layer2_outputs(9181) <= a;
    layer2_outputs(9182) <= not (a or b);
    layer2_outputs(9183) <= b;
    layer2_outputs(9184) <= not b;
    layer2_outputs(9185) <= a and b;
    layer2_outputs(9186) <= not a or b;
    layer2_outputs(9187) <= b;
    layer2_outputs(9188) <= a and b;
    layer2_outputs(9189) <= a xor b;
    layer2_outputs(9190) <= not (a or b);
    layer2_outputs(9191) <= a and b;
    layer2_outputs(9192) <= '1';
    layer2_outputs(9193) <= not a or b;
    layer2_outputs(9194) <= not (a or b);
    layer2_outputs(9195) <= '1';
    layer2_outputs(9196) <= not (a and b);
    layer2_outputs(9197) <= b and not a;
    layer2_outputs(9198) <= not b;
    layer2_outputs(9199) <= b;
    layer2_outputs(9200) <= a;
    layer2_outputs(9201) <= not (a and b);
    layer2_outputs(9202) <= b;
    layer2_outputs(9203) <= not (a or b);
    layer2_outputs(9204) <= not b or a;
    layer2_outputs(9205) <= a and b;
    layer2_outputs(9206) <= not (a and b);
    layer2_outputs(9207) <= a and not b;
    layer2_outputs(9208) <= '0';
    layer2_outputs(9209) <= not b or a;
    layer2_outputs(9210) <= not (a xor b);
    layer2_outputs(9211) <= '1';
    layer2_outputs(9212) <= a and b;
    layer2_outputs(9213) <= b;
    layer2_outputs(9214) <= '1';
    layer2_outputs(9215) <= a or b;
    layer2_outputs(9216) <= b and not a;
    layer2_outputs(9217) <= a and not b;
    layer2_outputs(9218) <= not a;
    layer2_outputs(9219) <= not (a or b);
    layer2_outputs(9220) <= not a;
    layer2_outputs(9221) <= '1';
    layer2_outputs(9222) <= not (a and b);
    layer2_outputs(9223) <= a;
    layer2_outputs(9224) <= a or b;
    layer2_outputs(9225) <= a and not b;
    layer2_outputs(9226) <= not (a and b);
    layer2_outputs(9227) <= not a or b;
    layer2_outputs(9228) <= not b;
    layer2_outputs(9229) <= b and not a;
    layer2_outputs(9230) <= a xor b;
    layer2_outputs(9231) <= a or b;
    layer2_outputs(9232) <= b;
    layer2_outputs(9233) <= a xor b;
    layer2_outputs(9234) <= b;
    layer2_outputs(9235) <= not b;
    layer2_outputs(9236) <= not (a or b);
    layer2_outputs(9237) <= a;
    layer2_outputs(9238) <= not b or a;
    layer2_outputs(9239) <= b and not a;
    layer2_outputs(9240) <= a or b;
    layer2_outputs(9241) <= a;
    layer2_outputs(9242) <= a;
    layer2_outputs(9243) <= not b or a;
    layer2_outputs(9244) <= b;
    layer2_outputs(9245) <= '0';
    layer2_outputs(9246) <= b;
    layer2_outputs(9247) <= not a or b;
    layer2_outputs(9248) <= a or b;
    layer2_outputs(9249) <= a and not b;
    layer2_outputs(9250) <= not b;
    layer2_outputs(9251) <= a;
    layer2_outputs(9252) <= a and b;
    layer2_outputs(9253) <= not (a or b);
    layer2_outputs(9254) <= a;
    layer2_outputs(9255) <= not b;
    layer2_outputs(9256) <= not (a xor b);
    layer2_outputs(9257) <= b and not a;
    layer2_outputs(9258) <= a;
    layer2_outputs(9259) <= not (a and b);
    layer2_outputs(9260) <= not b or a;
    layer2_outputs(9261) <= a and b;
    layer2_outputs(9262) <= a or b;
    layer2_outputs(9263) <= a or b;
    layer2_outputs(9264) <= a or b;
    layer2_outputs(9265) <= not a;
    layer2_outputs(9266) <= a and b;
    layer2_outputs(9267) <= '1';
    layer2_outputs(9268) <= not (a and b);
    layer2_outputs(9269) <= '1';
    layer2_outputs(9270) <= not (a and b);
    layer2_outputs(9271) <= a;
    layer2_outputs(9272) <= not a or b;
    layer2_outputs(9273) <= not a;
    layer2_outputs(9274) <= not b or a;
    layer2_outputs(9275) <= a and b;
    layer2_outputs(9276) <= b;
    layer2_outputs(9277) <= a;
    layer2_outputs(9278) <= a;
    layer2_outputs(9279) <= '1';
    layer2_outputs(9280) <= not a or b;
    layer2_outputs(9281) <= a or b;
    layer2_outputs(9282) <= '1';
    layer2_outputs(9283) <= not a;
    layer2_outputs(9284) <= not b;
    layer2_outputs(9285) <= a;
    layer2_outputs(9286) <= not (a xor b);
    layer2_outputs(9287) <= not a or b;
    layer2_outputs(9288) <= not (a xor b);
    layer2_outputs(9289) <= not a;
    layer2_outputs(9290) <= not (a or b);
    layer2_outputs(9291) <= not a or b;
    layer2_outputs(9292) <= not (a or b);
    layer2_outputs(9293) <= not b or a;
    layer2_outputs(9294) <= a and b;
    layer2_outputs(9295) <= not (a or b);
    layer2_outputs(9296) <= b;
    layer2_outputs(9297) <= a;
    layer2_outputs(9298) <= not b;
    layer2_outputs(9299) <= not (a and b);
    layer2_outputs(9300) <= a and not b;
    layer2_outputs(9301) <= a xor b;
    layer2_outputs(9302) <= not b or a;
    layer2_outputs(9303) <= not (a and b);
    layer2_outputs(9304) <= a xor b;
    layer2_outputs(9305) <= b;
    layer2_outputs(9306) <= a and not b;
    layer2_outputs(9307) <= '0';
    layer2_outputs(9308) <= not (a or b);
    layer2_outputs(9309) <= not b;
    layer2_outputs(9310) <= b and not a;
    layer2_outputs(9311) <= b;
    layer2_outputs(9312) <= b;
    layer2_outputs(9313) <= not (a xor b);
    layer2_outputs(9314) <= a or b;
    layer2_outputs(9315) <= not a or b;
    layer2_outputs(9316) <= '0';
    layer2_outputs(9317) <= a;
    layer2_outputs(9318) <= not b or a;
    layer2_outputs(9319) <= not (a and b);
    layer2_outputs(9320) <= not b;
    layer2_outputs(9321) <= b and not a;
    layer2_outputs(9322) <= '0';
    layer2_outputs(9323) <= not a;
    layer2_outputs(9324) <= not b;
    layer2_outputs(9325) <= not (a and b);
    layer2_outputs(9326) <= not b or a;
    layer2_outputs(9327) <= not a;
    layer2_outputs(9328) <= a or b;
    layer2_outputs(9329) <= not a;
    layer2_outputs(9330) <= b and not a;
    layer2_outputs(9331) <= a or b;
    layer2_outputs(9332) <= not a;
    layer2_outputs(9333) <= not (a and b);
    layer2_outputs(9334) <= a;
    layer2_outputs(9335) <= '0';
    layer2_outputs(9336) <= not b or a;
    layer2_outputs(9337) <= a or b;
    layer2_outputs(9338) <= not a;
    layer2_outputs(9339) <= a xor b;
    layer2_outputs(9340) <= b;
    layer2_outputs(9341) <= '1';
    layer2_outputs(9342) <= '0';
    layer2_outputs(9343) <= b and not a;
    layer2_outputs(9344) <= not (a or b);
    layer2_outputs(9345) <= a and not b;
    layer2_outputs(9346) <= a and not b;
    layer2_outputs(9347) <= b;
    layer2_outputs(9348) <= not (a or b);
    layer2_outputs(9349) <= not (a or b);
    layer2_outputs(9350) <= '1';
    layer2_outputs(9351) <= '1';
    layer2_outputs(9352) <= b and not a;
    layer2_outputs(9353) <= not (a or b);
    layer2_outputs(9354) <= not b;
    layer2_outputs(9355) <= not b;
    layer2_outputs(9356) <= b;
    layer2_outputs(9357) <= a;
    layer2_outputs(9358) <= not a;
    layer2_outputs(9359) <= b;
    layer2_outputs(9360) <= not (a or b);
    layer2_outputs(9361) <= a;
    layer2_outputs(9362) <= not b;
    layer2_outputs(9363) <= a;
    layer2_outputs(9364) <= a and not b;
    layer2_outputs(9365) <= b and not a;
    layer2_outputs(9366) <= not a or b;
    layer2_outputs(9367) <= b and not a;
    layer2_outputs(9368) <= not b;
    layer2_outputs(9369) <= not b or a;
    layer2_outputs(9370) <= not b or a;
    layer2_outputs(9371) <= not (a and b);
    layer2_outputs(9372) <= a;
    layer2_outputs(9373) <= not (a xor b);
    layer2_outputs(9374) <= '0';
    layer2_outputs(9375) <= not b or a;
    layer2_outputs(9376) <= a;
    layer2_outputs(9377) <= a;
    layer2_outputs(9378) <= not a;
    layer2_outputs(9379) <= b and not a;
    layer2_outputs(9380) <= a;
    layer2_outputs(9381) <= a xor b;
    layer2_outputs(9382) <= a;
    layer2_outputs(9383) <= a;
    layer2_outputs(9384) <= not (a or b);
    layer2_outputs(9385) <= not (a or b);
    layer2_outputs(9386) <= not b or a;
    layer2_outputs(9387) <= b and not a;
    layer2_outputs(9388) <= b;
    layer2_outputs(9389) <= a;
    layer2_outputs(9390) <= a or b;
    layer2_outputs(9391) <= a;
    layer2_outputs(9392) <= '0';
    layer2_outputs(9393) <= not (a or b);
    layer2_outputs(9394) <= not b or a;
    layer2_outputs(9395) <= '0';
    layer2_outputs(9396) <= not b;
    layer2_outputs(9397) <= a and b;
    layer2_outputs(9398) <= b;
    layer2_outputs(9399) <= not b or a;
    layer2_outputs(9400) <= b and not a;
    layer2_outputs(9401) <= not a;
    layer2_outputs(9402) <= not b;
    layer2_outputs(9403) <= '0';
    layer2_outputs(9404) <= '1';
    layer2_outputs(9405) <= b;
    layer2_outputs(9406) <= b;
    layer2_outputs(9407) <= a and not b;
    layer2_outputs(9408) <= '0';
    layer2_outputs(9409) <= not b;
    layer2_outputs(9410) <= a or b;
    layer2_outputs(9411) <= a and not b;
    layer2_outputs(9412) <= a and b;
    layer2_outputs(9413) <= not (a xor b);
    layer2_outputs(9414) <= '1';
    layer2_outputs(9415) <= b and not a;
    layer2_outputs(9416) <= a or b;
    layer2_outputs(9417) <= a;
    layer2_outputs(9418) <= a and not b;
    layer2_outputs(9419) <= b and not a;
    layer2_outputs(9420) <= a;
    layer2_outputs(9421) <= not a;
    layer2_outputs(9422) <= not (a or b);
    layer2_outputs(9423) <= not b or a;
    layer2_outputs(9424) <= b and not a;
    layer2_outputs(9425) <= a and b;
    layer2_outputs(9426) <= b;
    layer2_outputs(9427) <= not a or b;
    layer2_outputs(9428) <= not a or b;
    layer2_outputs(9429) <= a;
    layer2_outputs(9430) <= a;
    layer2_outputs(9431) <= b and not a;
    layer2_outputs(9432) <= a and b;
    layer2_outputs(9433) <= not b;
    layer2_outputs(9434) <= not b;
    layer2_outputs(9435) <= b;
    layer2_outputs(9436) <= a and b;
    layer2_outputs(9437) <= b;
    layer2_outputs(9438) <= a and b;
    layer2_outputs(9439) <= a xor b;
    layer2_outputs(9440) <= not a or b;
    layer2_outputs(9441) <= not (a xor b);
    layer2_outputs(9442) <= not (a or b);
    layer2_outputs(9443) <= '0';
    layer2_outputs(9444) <= b and not a;
    layer2_outputs(9445) <= a and b;
    layer2_outputs(9446) <= a and b;
    layer2_outputs(9447) <= b;
    layer2_outputs(9448) <= '0';
    layer2_outputs(9449) <= not a or b;
    layer2_outputs(9450) <= a;
    layer2_outputs(9451) <= not a;
    layer2_outputs(9452) <= not (a or b);
    layer2_outputs(9453) <= not b;
    layer2_outputs(9454) <= b;
    layer2_outputs(9455) <= not (a or b);
    layer2_outputs(9456) <= not b;
    layer2_outputs(9457) <= a and b;
    layer2_outputs(9458) <= not (a or b);
    layer2_outputs(9459) <= not (a and b);
    layer2_outputs(9460) <= '1';
    layer2_outputs(9461) <= '0';
    layer2_outputs(9462) <= a;
    layer2_outputs(9463) <= not b;
    layer2_outputs(9464) <= not (a or b);
    layer2_outputs(9465) <= not b or a;
    layer2_outputs(9466) <= not b or a;
    layer2_outputs(9467) <= a;
    layer2_outputs(9468) <= b;
    layer2_outputs(9469) <= not a;
    layer2_outputs(9470) <= '1';
    layer2_outputs(9471) <= b and not a;
    layer2_outputs(9472) <= not b;
    layer2_outputs(9473) <= not a;
    layer2_outputs(9474) <= b;
    layer2_outputs(9475) <= not b;
    layer2_outputs(9476) <= '1';
    layer2_outputs(9477) <= not (a or b);
    layer2_outputs(9478) <= not b or a;
    layer2_outputs(9479) <= not b;
    layer2_outputs(9480) <= '1';
    layer2_outputs(9481) <= not a or b;
    layer2_outputs(9482) <= '1';
    layer2_outputs(9483) <= a and b;
    layer2_outputs(9484) <= not b or a;
    layer2_outputs(9485) <= a or b;
    layer2_outputs(9486) <= a or b;
    layer2_outputs(9487) <= b and not a;
    layer2_outputs(9488) <= not b or a;
    layer2_outputs(9489) <= b;
    layer2_outputs(9490) <= b;
    layer2_outputs(9491) <= not (a or b);
    layer2_outputs(9492) <= not (a or b);
    layer2_outputs(9493) <= not a;
    layer2_outputs(9494) <= not (a xor b);
    layer2_outputs(9495) <= b and not a;
    layer2_outputs(9496) <= not (a and b);
    layer2_outputs(9497) <= not b;
    layer2_outputs(9498) <= b and not a;
    layer2_outputs(9499) <= not a;
    layer2_outputs(9500) <= not b;
    layer2_outputs(9501) <= not a or b;
    layer2_outputs(9502) <= a and not b;
    layer2_outputs(9503) <= '0';
    layer2_outputs(9504) <= not a;
    layer2_outputs(9505) <= a or b;
    layer2_outputs(9506) <= a and not b;
    layer2_outputs(9507) <= not (a or b);
    layer2_outputs(9508) <= not b or a;
    layer2_outputs(9509) <= '0';
    layer2_outputs(9510) <= a or b;
    layer2_outputs(9511) <= b;
    layer2_outputs(9512) <= b;
    layer2_outputs(9513) <= not b;
    layer2_outputs(9514) <= not a or b;
    layer2_outputs(9515) <= not a;
    layer2_outputs(9516) <= not b;
    layer2_outputs(9517) <= a and b;
    layer2_outputs(9518) <= '1';
    layer2_outputs(9519) <= '0';
    layer2_outputs(9520) <= b;
    layer2_outputs(9521) <= b;
    layer2_outputs(9522) <= '1';
    layer2_outputs(9523) <= a and not b;
    layer2_outputs(9524) <= not (a xor b);
    layer2_outputs(9525) <= b;
    layer2_outputs(9526) <= not (a or b);
    layer2_outputs(9527) <= a;
    layer2_outputs(9528) <= not a or b;
    layer2_outputs(9529) <= not (a or b);
    layer2_outputs(9530) <= '1';
    layer2_outputs(9531) <= not a;
    layer2_outputs(9532) <= not (a or b);
    layer2_outputs(9533) <= a or b;
    layer2_outputs(9534) <= a xor b;
    layer2_outputs(9535) <= '0';
    layer2_outputs(9536) <= not b or a;
    layer2_outputs(9537) <= b;
    layer2_outputs(9538) <= not (a or b);
    layer2_outputs(9539) <= a and not b;
    layer2_outputs(9540) <= not b;
    layer2_outputs(9541) <= not (a or b);
    layer2_outputs(9542) <= b;
    layer2_outputs(9543) <= not b or a;
    layer2_outputs(9544) <= a or b;
    layer2_outputs(9545) <= not (a or b);
    layer2_outputs(9546) <= '1';
    layer2_outputs(9547) <= not a or b;
    layer2_outputs(9548) <= a and not b;
    layer2_outputs(9549) <= not a;
    layer2_outputs(9550) <= a;
    layer2_outputs(9551) <= b and not a;
    layer2_outputs(9552) <= b and not a;
    layer2_outputs(9553) <= not (a or b);
    layer2_outputs(9554) <= a xor b;
    layer2_outputs(9555) <= '1';
    layer2_outputs(9556) <= b and not a;
    layer2_outputs(9557) <= not (a and b);
    layer2_outputs(9558) <= '1';
    layer2_outputs(9559) <= not a;
    layer2_outputs(9560) <= b and not a;
    layer2_outputs(9561) <= a;
    layer2_outputs(9562) <= '1';
    layer2_outputs(9563) <= not b or a;
    layer2_outputs(9564) <= not (a and b);
    layer2_outputs(9565) <= a and b;
    layer2_outputs(9566) <= not b or a;
    layer2_outputs(9567) <= '0';
    layer2_outputs(9568) <= not a or b;
    layer2_outputs(9569) <= '0';
    layer2_outputs(9570) <= not b or a;
    layer2_outputs(9571) <= not (a xor b);
    layer2_outputs(9572) <= a and b;
    layer2_outputs(9573) <= b;
    layer2_outputs(9574) <= a and not b;
    layer2_outputs(9575) <= not a or b;
    layer2_outputs(9576) <= b and not a;
    layer2_outputs(9577) <= a;
    layer2_outputs(9578) <= not b;
    layer2_outputs(9579) <= not a;
    layer2_outputs(9580) <= b;
    layer2_outputs(9581) <= b and not a;
    layer2_outputs(9582) <= a and b;
    layer2_outputs(9583) <= not a or b;
    layer2_outputs(9584) <= a or b;
    layer2_outputs(9585) <= not b;
    layer2_outputs(9586) <= b;
    layer2_outputs(9587) <= not b;
    layer2_outputs(9588) <= not (a xor b);
    layer2_outputs(9589) <= not a;
    layer2_outputs(9590) <= not b or a;
    layer2_outputs(9591) <= a;
    layer2_outputs(9592) <= a;
    layer2_outputs(9593) <= '0';
    layer2_outputs(9594) <= not a;
    layer2_outputs(9595) <= a;
    layer2_outputs(9596) <= b;
    layer2_outputs(9597) <= not a or b;
    layer2_outputs(9598) <= a xor b;
    layer2_outputs(9599) <= not a;
    layer2_outputs(9600) <= not (a xor b);
    layer2_outputs(9601) <= not a or b;
    layer2_outputs(9602) <= a and b;
    layer2_outputs(9603) <= not a;
    layer2_outputs(9604) <= '1';
    layer2_outputs(9605) <= a and not b;
    layer2_outputs(9606) <= b and not a;
    layer2_outputs(9607) <= b;
    layer2_outputs(9608) <= not (a or b);
    layer2_outputs(9609) <= a xor b;
    layer2_outputs(9610) <= not (a and b);
    layer2_outputs(9611) <= not b;
    layer2_outputs(9612) <= b;
    layer2_outputs(9613) <= not (a and b);
    layer2_outputs(9614) <= b and not a;
    layer2_outputs(9615) <= b;
    layer2_outputs(9616) <= a and not b;
    layer2_outputs(9617) <= not (a and b);
    layer2_outputs(9618) <= b;
    layer2_outputs(9619) <= not b or a;
    layer2_outputs(9620) <= b;
    layer2_outputs(9621) <= b;
    layer2_outputs(9622) <= not (a or b);
    layer2_outputs(9623) <= not a;
    layer2_outputs(9624) <= '1';
    layer2_outputs(9625) <= b and not a;
    layer2_outputs(9626) <= '0';
    layer2_outputs(9627) <= not (a and b);
    layer2_outputs(9628) <= not a;
    layer2_outputs(9629) <= a and b;
    layer2_outputs(9630) <= b;
    layer2_outputs(9631) <= a and not b;
    layer2_outputs(9632) <= b;
    layer2_outputs(9633) <= '0';
    layer2_outputs(9634) <= not a;
    layer2_outputs(9635) <= '1';
    layer2_outputs(9636) <= '0';
    layer2_outputs(9637) <= a and b;
    layer2_outputs(9638) <= not a or b;
    layer2_outputs(9639) <= not b or a;
    layer2_outputs(9640) <= a;
    layer2_outputs(9641) <= '1';
    layer2_outputs(9642) <= a xor b;
    layer2_outputs(9643) <= not a;
    layer2_outputs(9644) <= not (a or b);
    layer2_outputs(9645) <= '1';
    layer2_outputs(9646) <= a and not b;
    layer2_outputs(9647) <= '1';
    layer2_outputs(9648) <= b and not a;
    layer2_outputs(9649) <= not b or a;
    layer2_outputs(9650) <= not a;
    layer2_outputs(9651) <= b and not a;
    layer2_outputs(9652) <= not b;
    layer2_outputs(9653) <= not b;
    layer2_outputs(9654) <= a;
    layer2_outputs(9655) <= not b or a;
    layer2_outputs(9656) <= a;
    layer2_outputs(9657) <= not (a and b);
    layer2_outputs(9658) <= b and not a;
    layer2_outputs(9659) <= not a or b;
    layer2_outputs(9660) <= a xor b;
    layer2_outputs(9661) <= '1';
    layer2_outputs(9662) <= '0';
    layer2_outputs(9663) <= not a or b;
    layer2_outputs(9664) <= not b;
    layer2_outputs(9665) <= not (a or b);
    layer2_outputs(9666) <= not a;
    layer2_outputs(9667) <= a or b;
    layer2_outputs(9668) <= b;
    layer2_outputs(9669) <= '1';
    layer2_outputs(9670) <= not b or a;
    layer2_outputs(9671) <= a or b;
    layer2_outputs(9672) <= b;
    layer2_outputs(9673) <= not a or b;
    layer2_outputs(9674) <= not a;
    layer2_outputs(9675) <= a xor b;
    layer2_outputs(9676) <= a or b;
    layer2_outputs(9677) <= a and not b;
    layer2_outputs(9678) <= not (a xor b);
    layer2_outputs(9679) <= a and not b;
    layer2_outputs(9680) <= not b;
    layer2_outputs(9681) <= not b or a;
    layer2_outputs(9682) <= a;
    layer2_outputs(9683) <= a and b;
    layer2_outputs(9684) <= not (a and b);
    layer2_outputs(9685) <= not (a and b);
    layer2_outputs(9686) <= not b;
    layer2_outputs(9687) <= not b or a;
    layer2_outputs(9688) <= not b;
    layer2_outputs(9689) <= not b;
    layer2_outputs(9690) <= not (a and b);
    layer2_outputs(9691) <= a;
    layer2_outputs(9692) <= '0';
    layer2_outputs(9693) <= not (a xor b);
    layer2_outputs(9694) <= not b;
    layer2_outputs(9695) <= not (a or b);
    layer2_outputs(9696) <= not a;
    layer2_outputs(9697) <= b and not a;
    layer2_outputs(9698) <= not b;
    layer2_outputs(9699) <= not a;
    layer2_outputs(9700) <= not b or a;
    layer2_outputs(9701) <= not b;
    layer2_outputs(9702) <= not a;
    layer2_outputs(9703) <= not (a and b);
    layer2_outputs(9704) <= b;
    layer2_outputs(9705) <= a or b;
    layer2_outputs(9706) <= not b;
    layer2_outputs(9707) <= not a;
    layer2_outputs(9708) <= b;
    layer2_outputs(9709) <= b and not a;
    layer2_outputs(9710) <= a and not b;
    layer2_outputs(9711) <= a;
    layer2_outputs(9712) <= '1';
    layer2_outputs(9713) <= b and not a;
    layer2_outputs(9714) <= not (a or b);
    layer2_outputs(9715) <= '1';
    layer2_outputs(9716) <= not (a or b);
    layer2_outputs(9717) <= a and not b;
    layer2_outputs(9718) <= a;
    layer2_outputs(9719) <= a or b;
    layer2_outputs(9720) <= not a or b;
    layer2_outputs(9721) <= b;
    layer2_outputs(9722) <= '1';
    layer2_outputs(9723) <= not b;
    layer2_outputs(9724) <= not b;
    layer2_outputs(9725) <= not (a xor b);
    layer2_outputs(9726) <= b and not a;
    layer2_outputs(9727) <= not a;
    layer2_outputs(9728) <= not a;
    layer2_outputs(9729) <= not b;
    layer2_outputs(9730) <= a and b;
    layer2_outputs(9731) <= a and b;
    layer2_outputs(9732) <= a or b;
    layer2_outputs(9733) <= b;
    layer2_outputs(9734) <= not (a and b);
    layer2_outputs(9735) <= b;
    layer2_outputs(9736) <= not b;
    layer2_outputs(9737) <= not (a and b);
    layer2_outputs(9738) <= a or b;
    layer2_outputs(9739) <= not (a and b);
    layer2_outputs(9740) <= not b;
    layer2_outputs(9741) <= not a;
    layer2_outputs(9742) <= b and not a;
    layer2_outputs(9743) <= b;
    layer2_outputs(9744) <= '1';
    layer2_outputs(9745) <= '0';
    layer2_outputs(9746) <= a;
    layer2_outputs(9747) <= not (a and b);
    layer2_outputs(9748) <= not a or b;
    layer2_outputs(9749) <= b;
    layer2_outputs(9750) <= not a;
    layer2_outputs(9751) <= a xor b;
    layer2_outputs(9752) <= not b or a;
    layer2_outputs(9753) <= not b;
    layer2_outputs(9754) <= a and not b;
    layer2_outputs(9755) <= '0';
    layer2_outputs(9756) <= a and b;
    layer2_outputs(9757) <= not a;
    layer2_outputs(9758) <= not b;
    layer2_outputs(9759) <= not a;
    layer2_outputs(9760) <= a;
    layer2_outputs(9761) <= '0';
    layer2_outputs(9762) <= not (a or b);
    layer2_outputs(9763) <= a or b;
    layer2_outputs(9764) <= a and not b;
    layer2_outputs(9765) <= a and not b;
    layer2_outputs(9766) <= not (a and b);
    layer2_outputs(9767) <= a;
    layer2_outputs(9768) <= a and not b;
    layer2_outputs(9769) <= not (a and b);
    layer2_outputs(9770) <= not (a and b);
    layer2_outputs(9771) <= not (a xor b);
    layer2_outputs(9772) <= not a;
    layer2_outputs(9773) <= not b or a;
    layer2_outputs(9774) <= b;
    layer2_outputs(9775) <= a;
    layer2_outputs(9776) <= b;
    layer2_outputs(9777) <= not (a and b);
    layer2_outputs(9778) <= not b or a;
    layer2_outputs(9779) <= b;
    layer2_outputs(9780) <= not a or b;
    layer2_outputs(9781) <= not a;
    layer2_outputs(9782) <= b and not a;
    layer2_outputs(9783) <= not (a and b);
    layer2_outputs(9784) <= b and not a;
    layer2_outputs(9785) <= a;
    layer2_outputs(9786) <= not b or a;
    layer2_outputs(9787) <= not b or a;
    layer2_outputs(9788) <= a and b;
    layer2_outputs(9789) <= b and not a;
    layer2_outputs(9790) <= '0';
    layer2_outputs(9791) <= a;
    layer2_outputs(9792) <= b and not a;
    layer2_outputs(9793) <= a and not b;
    layer2_outputs(9794) <= not a;
    layer2_outputs(9795) <= '1';
    layer2_outputs(9796) <= a xor b;
    layer2_outputs(9797) <= b;
    layer2_outputs(9798) <= not b or a;
    layer2_outputs(9799) <= not a;
    layer2_outputs(9800) <= '1';
    layer2_outputs(9801) <= not (a or b);
    layer2_outputs(9802) <= a;
    layer2_outputs(9803) <= b;
    layer2_outputs(9804) <= a and b;
    layer2_outputs(9805) <= a or b;
    layer2_outputs(9806) <= '0';
    layer2_outputs(9807) <= a;
    layer2_outputs(9808) <= not a;
    layer2_outputs(9809) <= not b or a;
    layer2_outputs(9810) <= not (a or b);
    layer2_outputs(9811) <= not (a or b);
    layer2_outputs(9812) <= not a;
    layer2_outputs(9813) <= '1';
    layer2_outputs(9814) <= not b;
    layer2_outputs(9815) <= not b or a;
    layer2_outputs(9816) <= not a or b;
    layer2_outputs(9817) <= not b or a;
    layer2_outputs(9818) <= b and not a;
    layer2_outputs(9819) <= not a;
    layer2_outputs(9820) <= not b;
    layer2_outputs(9821) <= b;
    layer2_outputs(9822) <= not (a xor b);
    layer2_outputs(9823) <= not b;
    layer2_outputs(9824) <= a and not b;
    layer2_outputs(9825) <= a or b;
    layer2_outputs(9826) <= a and b;
    layer2_outputs(9827) <= not b;
    layer2_outputs(9828) <= a;
    layer2_outputs(9829) <= b and not a;
    layer2_outputs(9830) <= b;
    layer2_outputs(9831) <= a or b;
    layer2_outputs(9832) <= a;
    layer2_outputs(9833) <= a and b;
    layer2_outputs(9834) <= not (a and b);
    layer2_outputs(9835) <= not a or b;
    layer2_outputs(9836) <= not (a xor b);
    layer2_outputs(9837) <= not b or a;
    layer2_outputs(9838) <= not (a and b);
    layer2_outputs(9839) <= not (a xor b);
    layer2_outputs(9840) <= not b or a;
    layer2_outputs(9841) <= a and not b;
    layer2_outputs(9842) <= not (a or b);
    layer2_outputs(9843) <= not (a or b);
    layer2_outputs(9844) <= b;
    layer2_outputs(9845) <= '1';
    layer2_outputs(9846) <= a;
    layer2_outputs(9847) <= a;
    layer2_outputs(9848) <= not (a and b);
    layer2_outputs(9849) <= not b;
    layer2_outputs(9850) <= '1';
    layer2_outputs(9851) <= not a;
    layer2_outputs(9852) <= a;
    layer2_outputs(9853) <= not a or b;
    layer2_outputs(9854) <= a and b;
    layer2_outputs(9855) <= a xor b;
    layer2_outputs(9856) <= not b or a;
    layer2_outputs(9857) <= a;
    layer2_outputs(9858) <= b;
    layer2_outputs(9859) <= '1';
    layer2_outputs(9860) <= a;
    layer2_outputs(9861) <= b;
    layer2_outputs(9862) <= not b or a;
    layer2_outputs(9863) <= not b or a;
    layer2_outputs(9864) <= '0';
    layer2_outputs(9865) <= not a or b;
    layer2_outputs(9866) <= a and not b;
    layer2_outputs(9867) <= '1';
    layer2_outputs(9868) <= a and not b;
    layer2_outputs(9869) <= not a or b;
    layer2_outputs(9870) <= a and not b;
    layer2_outputs(9871) <= not (a or b);
    layer2_outputs(9872) <= '0';
    layer2_outputs(9873) <= a or b;
    layer2_outputs(9874) <= b;
    layer2_outputs(9875) <= b;
    layer2_outputs(9876) <= not (a xor b);
    layer2_outputs(9877) <= a and b;
    layer2_outputs(9878) <= a xor b;
    layer2_outputs(9879) <= '1';
    layer2_outputs(9880) <= not b or a;
    layer2_outputs(9881) <= not (a and b);
    layer2_outputs(9882) <= '1';
    layer2_outputs(9883) <= '1';
    layer2_outputs(9884) <= not b;
    layer2_outputs(9885) <= not (a and b);
    layer2_outputs(9886) <= a or b;
    layer2_outputs(9887) <= b;
    layer2_outputs(9888) <= a or b;
    layer2_outputs(9889) <= a or b;
    layer2_outputs(9890) <= a;
    layer2_outputs(9891) <= not a or b;
    layer2_outputs(9892) <= not a;
    layer2_outputs(9893) <= not (a or b);
    layer2_outputs(9894) <= b;
    layer2_outputs(9895) <= not a;
    layer2_outputs(9896) <= not b or a;
    layer2_outputs(9897) <= not b;
    layer2_outputs(9898) <= not a;
    layer2_outputs(9899) <= '0';
    layer2_outputs(9900) <= a;
    layer2_outputs(9901) <= not a;
    layer2_outputs(9902) <= a and b;
    layer2_outputs(9903) <= not (a xor b);
    layer2_outputs(9904) <= a and b;
    layer2_outputs(9905) <= b and not a;
    layer2_outputs(9906) <= not a;
    layer2_outputs(9907) <= a;
    layer2_outputs(9908) <= '1';
    layer2_outputs(9909) <= not a;
    layer2_outputs(9910) <= not b or a;
    layer2_outputs(9911) <= not (a xor b);
    layer2_outputs(9912) <= a xor b;
    layer2_outputs(9913) <= not (a xor b);
    layer2_outputs(9914) <= '1';
    layer2_outputs(9915) <= a or b;
    layer2_outputs(9916) <= a;
    layer2_outputs(9917) <= b;
    layer2_outputs(9918) <= not a;
    layer2_outputs(9919) <= not a;
    layer2_outputs(9920) <= b;
    layer2_outputs(9921) <= a or b;
    layer2_outputs(9922) <= not (a xor b);
    layer2_outputs(9923) <= not b or a;
    layer2_outputs(9924) <= not (a and b);
    layer2_outputs(9925) <= a and b;
    layer2_outputs(9926) <= a or b;
    layer2_outputs(9927) <= a and not b;
    layer2_outputs(9928) <= not (a xor b);
    layer2_outputs(9929) <= not b or a;
    layer2_outputs(9930) <= not (a or b);
    layer2_outputs(9931) <= b;
    layer2_outputs(9932) <= a;
    layer2_outputs(9933) <= not b;
    layer2_outputs(9934) <= not (a and b);
    layer2_outputs(9935) <= b and not a;
    layer2_outputs(9936) <= a or b;
    layer2_outputs(9937) <= b;
    layer2_outputs(9938) <= not a;
    layer2_outputs(9939) <= a or b;
    layer2_outputs(9940) <= b;
    layer2_outputs(9941) <= b;
    layer2_outputs(9942) <= not (a xor b);
    layer2_outputs(9943) <= a and not b;
    layer2_outputs(9944) <= b and not a;
    layer2_outputs(9945) <= not b or a;
    layer2_outputs(9946) <= b and not a;
    layer2_outputs(9947) <= a and b;
    layer2_outputs(9948) <= not b;
    layer2_outputs(9949) <= not a or b;
    layer2_outputs(9950) <= not b;
    layer2_outputs(9951) <= not a or b;
    layer2_outputs(9952) <= b and not a;
    layer2_outputs(9953) <= a and b;
    layer2_outputs(9954) <= not a or b;
    layer2_outputs(9955) <= not a;
    layer2_outputs(9956) <= a or b;
    layer2_outputs(9957) <= a;
    layer2_outputs(9958) <= '0';
    layer2_outputs(9959) <= b;
    layer2_outputs(9960) <= not a or b;
    layer2_outputs(9961) <= '0';
    layer2_outputs(9962) <= a and b;
    layer2_outputs(9963) <= a;
    layer2_outputs(9964) <= a;
    layer2_outputs(9965) <= a and not b;
    layer2_outputs(9966) <= a and b;
    layer2_outputs(9967) <= not (a xor b);
    layer2_outputs(9968) <= a and b;
    layer2_outputs(9969) <= b and not a;
    layer2_outputs(9970) <= not (a and b);
    layer2_outputs(9971) <= b;
    layer2_outputs(9972) <= not a;
    layer2_outputs(9973) <= not a;
    layer2_outputs(9974) <= '1';
    layer2_outputs(9975) <= '0';
    layer2_outputs(9976) <= not a;
    layer2_outputs(9977) <= a and not b;
    layer2_outputs(9978) <= not (a or b);
    layer2_outputs(9979) <= not a;
    layer2_outputs(9980) <= a and b;
    layer2_outputs(9981) <= a or b;
    layer2_outputs(9982) <= not a or b;
    layer2_outputs(9983) <= a;
    layer2_outputs(9984) <= not b;
    layer2_outputs(9985) <= not (a and b);
    layer2_outputs(9986) <= not b or a;
    layer2_outputs(9987) <= not a;
    layer2_outputs(9988) <= not (a or b);
    layer2_outputs(9989) <= '0';
    layer2_outputs(9990) <= a;
    layer2_outputs(9991) <= not a;
    layer2_outputs(9992) <= not a or b;
    layer2_outputs(9993) <= b and not a;
    layer2_outputs(9994) <= a and not b;
    layer2_outputs(9995) <= b and not a;
    layer2_outputs(9996) <= not b;
    layer2_outputs(9997) <= b;
    layer2_outputs(9998) <= a or b;
    layer2_outputs(9999) <= a xor b;
    layer2_outputs(10000) <= a and b;
    layer2_outputs(10001) <= '1';
    layer2_outputs(10002) <= '1';
    layer2_outputs(10003) <= not b or a;
    layer2_outputs(10004) <= a or b;
    layer2_outputs(10005) <= a and b;
    layer2_outputs(10006) <= a;
    layer2_outputs(10007) <= b;
    layer2_outputs(10008) <= not b;
    layer2_outputs(10009) <= not a;
    layer2_outputs(10010) <= a and not b;
    layer2_outputs(10011) <= not a or b;
    layer2_outputs(10012) <= not a;
    layer2_outputs(10013) <= not (a and b);
    layer2_outputs(10014) <= a and b;
    layer2_outputs(10015) <= not a;
    layer2_outputs(10016) <= a and not b;
    layer2_outputs(10017) <= a xor b;
    layer2_outputs(10018) <= '1';
    layer2_outputs(10019) <= '0';
    layer2_outputs(10020) <= not a or b;
    layer2_outputs(10021) <= not (a and b);
    layer2_outputs(10022) <= b;
    layer2_outputs(10023) <= not a or b;
    layer2_outputs(10024) <= not a;
    layer2_outputs(10025) <= b and not a;
    layer2_outputs(10026) <= a;
    layer2_outputs(10027) <= a xor b;
    layer2_outputs(10028) <= b and not a;
    layer2_outputs(10029) <= a and not b;
    layer2_outputs(10030) <= not b;
    layer2_outputs(10031) <= not b;
    layer2_outputs(10032) <= not a;
    layer2_outputs(10033) <= not b;
    layer2_outputs(10034) <= b;
    layer2_outputs(10035) <= a or b;
    layer2_outputs(10036) <= '1';
    layer2_outputs(10037) <= a xor b;
    layer2_outputs(10038) <= not b;
    layer2_outputs(10039) <= '0';
    layer2_outputs(10040) <= not a;
    layer2_outputs(10041) <= not (a xor b);
    layer2_outputs(10042) <= not (a or b);
    layer2_outputs(10043) <= not a or b;
    layer2_outputs(10044) <= not b or a;
    layer2_outputs(10045) <= a;
    layer2_outputs(10046) <= not (a or b);
    layer2_outputs(10047) <= b;
    layer2_outputs(10048) <= not a or b;
    layer2_outputs(10049) <= not b;
    layer2_outputs(10050) <= not (a and b);
    layer2_outputs(10051) <= not (a and b);
    layer2_outputs(10052) <= a or b;
    layer2_outputs(10053) <= not (a and b);
    layer2_outputs(10054) <= b and not a;
    layer2_outputs(10055) <= not (a xor b);
    layer2_outputs(10056) <= not (a xor b);
    layer2_outputs(10057) <= a and b;
    layer2_outputs(10058) <= not a;
    layer2_outputs(10059) <= a and b;
    layer2_outputs(10060) <= a and b;
    layer2_outputs(10061) <= a or b;
    layer2_outputs(10062) <= a and not b;
    layer2_outputs(10063) <= a and not b;
    layer2_outputs(10064) <= '0';
    layer2_outputs(10065) <= not b;
    layer2_outputs(10066) <= not a or b;
    layer2_outputs(10067) <= a and not b;
    layer2_outputs(10068) <= '0';
    layer2_outputs(10069) <= a and not b;
    layer2_outputs(10070) <= a and b;
    layer2_outputs(10071) <= a and not b;
    layer2_outputs(10072) <= a;
    layer2_outputs(10073) <= a and not b;
    layer2_outputs(10074) <= a and not b;
    layer2_outputs(10075) <= not (a xor b);
    layer2_outputs(10076) <= not b;
    layer2_outputs(10077) <= b;
    layer2_outputs(10078) <= not (a or b);
    layer2_outputs(10079) <= not (a or b);
    layer2_outputs(10080) <= a and not b;
    layer2_outputs(10081) <= not (a or b);
    layer2_outputs(10082) <= not b;
    layer2_outputs(10083) <= a or b;
    layer2_outputs(10084) <= a;
    layer2_outputs(10085) <= not (a or b);
    layer2_outputs(10086) <= a and b;
    layer2_outputs(10087) <= a and b;
    layer2_outputs(10088) <= not a or b;
    layer2_outputs(10089) <= a and b;
    layer2_outputs(10090) <= not (a and b);
    layer2_outputs(10091) <= b and not a;
    layer2_outputs(10092) <= a and not b;
    layer2_outputs(10093) <= '0';
    layer2_outputs(10094) <= not b;
    layer2_outputs(10095) <= a;
    layer2_outputs(10096) <= a and b;
    layer2_outputs(10097) <= a or b;
    layer2_outputs(10098) <= '1';
    layer2_outputs(10099) <= '0';
    layer2_outputs(10100) <= a;
    layer2_outputs(10101) <= not (a and b);
    layer2_outputs(10102) <= not b or a;
    layer2_outputs(10103) <= not b;
    layer2_outputs(10104) <= b and not a;
    layer2_outputs(10105) <= not b or a;
    layer2_outputs(10106) <= a and not b;
    layer2_outputs(10107) <= not (a or b);
    layer2_outputs(10108) <= b and not a;
    layer2_outputs(10109) <= a;
    layer2_outputs(10110) <= b and not a;
    layer2_outputs(10111) <= not a or b;
    layer2_outputs(10112) <= '1';
    layer2_outputs(10113) <= '1';
    layer2_outputs(10114) <= not a or b;
    layer2_outputs(10115) <= b;
    layer2_outputs(10116) <= not (a xor b);
    layer2_outputs(10117) <= a and not b;
    layer2_outputs(10118) <= a and b;
    layer2_outputs(10119) <= '0';
    layer2_outputs(10120) <= not (a or b);
    layer2_outputs(10121) <= not (a and b);
    layer2_outputs(10122) <= a;
    layer2_outputs(10123) <= not b;
    layer2_outputs(10124) <= '1';
    layer2_outputs(10125) <= a and b;
    layer2_outputs(10126) <= not a;
    layer2_outputs(10127) <= '1';
    layer2_outputs(10128) <= '1';
    layer2_outputs(10129) <= a or b;
    layer2_outputs(10130) <= not (a xor b);
    layer2_outputs(10131) <= not b;
    layer2_outputs(10132) <= not a;
    layer2_outputs(10133) <= '1';
    layer2_outputs(10134) <= b and not a;
    layer2_outputs(10135) <= b and not a;
    layer2_outputs(10136) <= not b or a;
    layer2_outputs(10137) <= a;
    layer2_outputs(10138) <= '0';
    layer2_outputs(10139) <= b and not a;
    layer2_outputs(10140) <= b;
    layer2_outputs(10141) <= '0';
    layer2_outputs(10142) <= a and not b;
    layer2_outputs(10143) <= b and not a;
    layer2_outputs(10144) <= a xor b;
    layer2_outputs(10145) <= not (a or b);
    layer2_outputs(10146) <= a and not b;
    layer2_outputs(10147) <= a and b;
    layer2_outputs(10148) <= not a;
    layer2_outputs(10149) <= a and not b;
    layer2_outputs(10150) <= not (a and b);
    layer2_outputs(10151) <= a;
    layer2_outputs(10152) <= not a or b;
    layer2_outputs(10153) <= '0';
    layer2_outputs(10154) <= not b or a;
    layer2_outputs(10155) <= '1';
    layer2_outputs(10156) <= not b or a;
    layer2_outputs(10157) <= '0';
    layer2_outputs(10158) <= not (a xor b);
    layer2_outputs(10159) <= not (a and b);
    layer2_outputs(10160) <= not a or b;
    layer2_outputs(10161) <= b;
    layer2_outputs(10162) <= not a;
    layer2_outputs(10163) <= a and b;
    layer2_outputs(10164) <= a;
    layer2_outputs(10165) <= b;
    layer2_outputs(10166) <= not b;
    layer2_outputs(10167) <= a;
    layer2_outputs(10168) <= a and not b;
    layer2_outputs(10169) <= a and b;
    layer2_outputs(10170) <= a or b;
    layer2_outputs(10171) <= not a or b;
    layer2_outputs(10172) <= '0';
    layer2_outputs(10173) <= '1';
    layer2_outputs(10174) <= a or b;
    layer2_outputs(10175) <= '1';
    layer2_outputs(10176) <= not b or a;
    layer2_outputs(10177) <= not b or a;
    layer2_outputs(10178) <= b and not a;
    layer2_outputs(10179) <= not b or a;
    layer2_outputs(10180) <= not b;
    layer2_outputs(10181) <= a or b;
    layer2_outputs(10182) <= b;
    layer2_outputs(10183) <= b;
    layer2_outputs(10184) <= a or b;
    layer2_outputs(10185) <= not b;
    layer2_outputs(10186) <= b and not a;
    layer2_outputs(10187) <= not b;
    layer2_outputs(10188) <= '0';
    layer2_outputs(10189) <= a;
    layer2_outputs(10190) <= not (a and b);
    layer2_outputs(10191) <= b;
    layer2_outputs(10192) <= b;
    layer2_outputs(10193) <= a xor b;
    layer2_outputs(10194) <= '0';
    layer2_outputs(10195) <= a or b;
    layer2_outputs(10196) <= b;
    layer2_outputs(10197) <= b;
    layer2_outputs(10198) <= not b or a;
    layer2_outputs(10199) <= not a or b;
    layer2_outputs(10200) <= a and not b;
    layer2_outputs(10201) <= not (a and b);
    layer2_outputs(10202) <= a;
    layer2_outputs(10203) <= not a or b;
    layer2_outputs(10204) <= a or b;
    layer2_outputs(10205) <= not a;
    layer2_outputs(10206) <= not (a or b);
    layer2_outputs(10207) <= a;
    layer2_outputs(10208) <= b and not a;
    layer2_outputs(10209) <= b;
    layer2_outputs(10210) <= not (a and b);
    layer2_outputs(10211) <= b;
    layer2_outputs(10212) <= a xor b;
    layer2_outputs(10213) <= not a;
    layer2_outputs(10214) <= not b;
    layer2_outputs(10215) <= not (a and b);
    layer2_outputs(10216) <= a and not b;
    layer2_outputs(10217) <= a and b;
    layer2_outputs(10218) <= a or b;
    layer2_outputs(10219) <= b;
    layer2_outputs(10220) <= not (a or b);
    layer2_outputs(10221) <= '0';
    layer2_outputs(10222) <= a and b;
    layer2_outputs(10223) <= b and not a;
    layer2_outputs(10224) <= not a;
    layer2_outputs(10225) <= a;
    layer2_outputs(10226) <= not (a and b);
    layer2_outputs(10227) <= not (a and b);
    layer2_outputs(10228) <= not (a or b);
    layer2_outputs(10229) <= a xor b;
    layer2_outputs(10230) <= a and not b;
    layer2_outputs(10231) <= not a;
    layer2_outputs(10232) <= not (a or b);
    layer2_outputs(10233) <= not b or a;
    layer2_outputs(10234) <= a;
    layer2_outputs(10235) <= not a;
    layer2_outputs(10236) <= not b or a;
    layer2_outputs(10237) <= not b;
    layer2_outputs(10238) <= a and not b;
    layer2_outputs(10239) <= not (a and b);
    layer3_outputs(0) <= a;
    layer3_outputs(1) <= b;
    layer3_outputs(2) <= a and b;
    layer3_outputs(3) <= b;
    layer3_outputs(4) <= not (a xor b);
    layer3_outputs(5) <= b;
    layer3_outputs(6) <= not (a or b);
    layer3_outputs(7) <= not (a xor b);
    layer3_outputs(8) <= not b;
    layer3_outputs(9) <= not a;
    layer3_outputs(10) <= a;
    layer3_outputs(11) <= a xor b;
    layer3_outputs(12) <= a or b;
    layer3_outputs(13) <= not b or a;
    layer3_outputs(14) <= a or b;
    layer3_outputs(15) <= not a;
    layer3_outputs(16) <= a and not b;
    layer3_outputs(17) <= not b;
    layer3_outputs(18) <= a and b;
    layer3_outputs(19) <= not (a xor b);
    layer3_outputs(20) <= a or b;
    layer3_outputs(21) <= '0';
    layer3_outputs(22) <= not (a or b);
    layer3_outputs(23) <= not a;
    layer3_outputs(24) <= not b;
    layer3_outputs(25) <= not a;
    layer3_outputs(26) <= a and b;
    layer3_outputs(27) <= '1';
    layer3_outputs(28) <= not b;
    layer3_outputs(29) <= b;
    layer3_outputs(30) <= '1';
    layer3_outputs(31) <= a xor b;
    layer3_outputs(32) <= not a;
    layer3_outputs(33) <= not a;
    layer3_outputs(34) <= b;
    layer3_outputs(35) <= not b or a;
    layer3_outputs(36) <= not (a or b);
    layer3_outputs(37) <= '1';
    layer3_outputs(38) <= a;
    layer3_outputs(39) <= '0';
    layer3_outputs(40) <= b;
    layer3_outputs(41) <= not (a xor b);
    layer3_outputs(42) <= '1';
    layer3_outputs(43) <= a;
    layer3_outputs(44) <= a and not b;
    layer3_outputs(45) <= not a or b;
    layer3_outputs(46) <= not a;
    layer3_outputs(47) <= not a;
    layer3_outputs(48) <= b;
    layer3_outputs(49) <= '1';
    layer3_outputs(50) <= not (a and b);
    layer3_outputs(51) <= a and b;
    layer3_outputs(52) <= not (a or b);
    layer3_outputs(53) <= a;
    layer3_outputs(54) <= not b or a;
    layer3_outputs(55) <= '1';
    layer3_outputs(56) <= a;
    layer3_outputs(57) <= b;
    layer3_outputs(58) <= not a;
    layer3_outputs(59) <= not (a xor b);
    layer3_outputs(60) <= a;
    layer3_outputs(61) <= not (a or b);
    layer3_outputs(62) <= a;
    layer3_outputs(63) <= not b or a;
    layer3_outputs(64) <= not a or b;
    layer3_outputs(65) <= a xor b;
    layer3_outputs(66) <= not b;
    layer3_outputs(67) <= not b or a;
    layer3_outputs(68) <= not (a xor b);
    layer3_outputs(69) <= not a or b;
    layer3_outputs(70) <= not (a or b);
    layer3_outputs(71) <= a xor b;
    layer3_outputs(72) <= b and not a;
    layer3_outputs(73) <= a;
    layer3_outputs(74) <= a;
    layer3_outputs(75) <= a or b;
    layer3_outputs(76) <= a;
    layer3_outputs(77) <= b;
    layer3_outputs(78) <= a;
    layer3_outputs(79) <= a and b;
    layer3_outputs(80) <= not (a and b);
    layer3_outputs(81) <= b;
    layer3_outputs(82) <= not (a and b);
    layer3_outputs(83) <= not a or b;
    layer3_outputs(84) <= a and b;
    layer3_outputs(85) <= a or b;
    layer3_outputs(86) <= a;
    layer3_outputs(87) <= a or b;
    layer3_outputs(88) <= b and not a;
    layer3_outputs(89) <= a;
    layer3_outputs(90) <= a and not b;
    layer3_outputs(91) <= a or b;
    layer3_outputs(92) <= b;
    layer3_outputs(93) <= not b;
    layer3_outputs(94) <= a;
    layer3_outputs(95) <= a;
    layer3_outputs(96) <= not b or a;
    layer3_outputs(97) <= a;
    layer3_outputs(98) <= not (a and b);
    layer3_outputs(99) <= not (a and b);
    layer3_outputs(100) <= b;
    layer3_outputs(101) <= not a or b;
    layer3_outputs(102) <= b;
    layer3_outputs(103) <= a xor b;
    layer3_outputs(104) <= not a;
    layer3_outputs(105) <= b and not a;
    layer3_outputs(106) <= a;
    layer3_outputs(107) <= a and b;
    layer3_outputs(108) <= not (a or b);
    layer3_outputs(109) <= not (a and b);
    layer3_outputs(110) <= not a or b;
    layer3_outputs(111) <= not b;
    layer3_outputs(112) <= b;
    layer3_outputs(113) <= not a;
    layer3_outputs(114) <= a;
    layer3_outputs(115) <= not (a or b);
    layer3_outputs(116) <= not a;
    layer3_outputs(117) <= not (a and b);
    layer3_outputs(118) <= not a;
    layer3_outputs(119) <= not (a and b);
    layer3_outputs(120) <= not a;
    layer3_outputs(121) <= b;
    layer3_outputs(122) <= not a;
    layer3_outputs(123) <= not a;
    layer3_outputs(124) <= not (a or b);
    layer3_outputs(125) <= a;
    layer3_outputs(126) <= not a;
    layer3_outputs(127) <= not b;
    layer3_outputs(128) <= not (a and b);
    layer3_outputs(129) <= not b;
    layer3_outputs(130) <= not (a and b);
    layer3_outputs(131) <= a or b;
    layer3_outputs(132) <= '1';
    layer3_outputs(133) <= b;
    layer3_outputs(134) <= a or b;
    layer3_outputs(135) <= not a;
    layer3_outputs(136) <= not b;
    layer3_outputs(137) <= a or b;
    layer3_outputs(138) <= not (a and b);
    layer3_outputs(139) <= a;
    layer3_outputs(140) <= '0';
    layer3_outputs(141) <= a or b;
    layer3_outputs(142) <= a;
    layer3_outputs(143) <= a and b;
    layer3_outputs(144) <= not a or b;
    layer3_outputs(145) <= b;
    layer3_outputs(146) <= b and not a;
    layer3_outputs(147) <= '0';
    layer3_outputs(148) <= a or b;
    layer3_outputs(149) <= b and not a;
    layer3_outputs(150) <= b and not a;
    layer3_outputs(151) <= not (a and b);
    layer3_outputs(152) <= b;
    layer3_outputs(153) <= a and not b;
    layer3_outputs(154) <= not a;
    layer3_outputs(155) <= '1';
    layer3_outputs(156) <= not a or b;
    layer3_outputs(157) <= a and not b;
    layer3_outputs(158) <= not b;
    layer3_outputs(159) <= not b;
    layer3_outputs(160) <= not b;
    layer3_outputs(161) <= a and not b;
    layer3_outputs(162) <= not (a and b);
    layer3_outputs(163) <= a;
    layer3_outputs(164) <= '0';
    layer3_outputs(165) <= not a or b;
    layer3_outputs(166) <= a or b;
    layer3_outputs(167) <= a and b;
    layer3_outputs(168) <= not b or a;
    layer3_outputs(169) <= not b;
    layer3_outputs(170) <= not a or b;
    layer3_outputs(171) <= a and b;
    layer3_outputs(172) <= '0';
    layer3_outputs(173) <= b;
    layer3_outputs(174) <= '1';
    layer3_outputs(175) <= b;
    layer3_outputs(176) <= a and b;
    layer3_outputs(177) <= not (a xor b);
    layer3_outputs(178) <= not b or a;
    layer3_outputs(179) <= not (a and b);
    layer3_outputs(180) <= a and b;
    layer3_outputs(181) <= b and not a;
    layer3_outputs(182) <= not b;
    layer3_outputs(183) <= b and not a;
    layer3_outputs(184) <= '1';
    layer3_outputs(185) <= not (a xor b);
    layer3_outputs(186) <= '1';
    layer3_outputs(187) <= b;
    layer3_outputs(188) <= not (a and b);
    layer3_outputs(189) <= not a;
    layer3_outputs(190) <= b and not a;
    layer3_outputs(191) <= a or b;
    layer3_outputs(192) <= a;
    layer3_outputs(193) <= '0';
    layer3_outputs(194) <= a and b;
    layer3_outputs(195) <= a;
    layer3_outputs(196) <= not b;
    layer3_outputs(197) <= a;
    layer3_outputs(198) <= b;
    layer3_outputs(199) <= a;
    layer3_outputs(200) <= a or b;
    layer3_outputs(201) <= not a;
    layer3_outputs(202) <= a and not b;
    layer3_outputs(203) <= a and b;
    layer3_outputs(204) <= a or b;
    layer3_outputs(205) <= a and b;
    layer3_outputs(206) <= not b;
    layer3_outputs(207) <= not a;
    layer3_outputs(208) <= not a;
    layer3_outputs(209) <= a xor b;
    layer3_outputs(210) <= not a;
    layer3_outputs(211) <= not a or b;
    layer3_outputs(212) <= b and not a;
    layer3_outputs(213) <= b and not a;
    layer3_outputs(214) <= b and not a;
    layer3_outputs(215) <= '1';
    layer3_outputs(216) <= not a;
    layer3_outputs(217) <= a and not b;
    layer3_outputs(218) <= b and not a;
    layer3_outputs(219) <= b;
    layer3_outputs(220) <= a xor b;
    layer3_outputs(221) <= a xor b;
    layer3_outputs(222) <= not b;
    layer3_outputs(223) <= not b;
    layer3_outputs(224) <= not a or b;
    layer3_outputs(225) <= b and not a;
    layer3_outputs(226) <= '0';
    layer3_outputs(227) <= b;
    layer3_outputs(228) <= a and not b;
    layer3_outputs(229) <= a;
    layer3_outputs(230) <= not b;
    layer3_outputs(231) <= not (a or b);
    layer3_outputs(232) <= a xor b;
    layer3_outputs(233) <= a and not b;
    layer3_outputs(234) <= not b;
    layer3_outputs(235) <= not (a and b);
    layer3_outputs(236) <= not a or b;
    layer3_outputs(237) <= not a;
    layer3_outputs(238) <= not a;
    layer3_outputs(239) <= a or b;
    layer3_outputs(240) <= a and b;
    layer3_outputs(241) <= a;
    layer3_outputs(242) <= not a or b;
    layer3_outputs(243) <= a and b;
    layer3_outputs(244) <= not (a or b);
    layer3_outputs(245) <= not b;
    layer3_outputs(246) <= '0';
    layer3_outputs(247) <= not (a and b);
    layer3_outputs(248) <= not (a or b);
    layer3_outputs(249) <= a xor b;
    layer3_outputs(250) <= b;
    layer3_outputs(251) <= not (a or b);
    layer3_outputs(252) <= not b or a;
    layer3_outputs(253) <= a;
    layer3_outputs(254) <= b and not a;
    layer3_outputs(255) <= not b;
    layer3_outputs(256) <= a;
    layer3_outputs(257) <= a and b;
    layer3_outputs(258) <= not b;
    layer3_outputs(259) <= not a or b;
    layer3_outputs(260) <= a or b;
    layer3_outputs(261) <= a;
    layer3_outputs(262) <= not a;
    layer3_outputs(263) <= b and not a;
    layer3_outputs(264) <= a and not b;
    layer3_outputs(265) <= not a;
    layer3_outputs(266) <= not (a and b);
    layer3_outputs(267) <= a xor b;
    layer3_outputs(268) <= not (a and b);
    layer3_outputs(269) <= b;
    layer3_outputs(270) <= not a or b;
    layer3_outputs(271) <= a and b;
    layer3_outputs(272) <= '0';
    layer3_outputs(273) <= not (a or b);
    layer3_outputs(274) <= a;
    layer3_outputs(275) <= not (a and b);
    layer3_outputs(276) <= a and b;
    layer3_outputs(277) <= not b;
    layer3_outputs(278) <= a and not b;
    layer3_outputs(279) <= a;
    layer3_outputs(280) <= '0';
    layer3_outputs(281) <= not a or b;
    layer3_outputs(282) <= a;
    layer3_outputs(283) <= not a;
    layer3_outputs(284) <= not a;
    layer3_outputs(285) <= a xor b;
    layer3_outputs(286) <= a or b;
    layer3_outputs(287) <= not (a xor b);
    layer3_outputs(288) <= not a or b;
    layer3_outputs(289) <= not a;
    layer3_outputs(290) <= b and not a;
    layer3_outputs(291) <= a and not b;
    layer3_outputs(292) <= not b;
    layer3_outputs(293) <= a xor b;
    layer3_outputs(294) <= a;
    layer3_outputs(295) <= b;
    layer3_outputs(296) <= not a;
    layer3_outputs(297) <= b and not a;
    layer3_outputs(298) <= '1';
    layer3_outputs(299) <= a;
    layer3_outputs(300) <= a and not b;
    layer3_outputs(301) <= a or b;
    layer3_outputs(302) <= not a;
    layer3_outputs(303) <= not b;
    layer3_outputs(304) <= not (a and b);
    layer3_outputs(305) <= not b;
    layer3_outputs(306) <= not (a or b);
    layer3_outputs(307) <= a or b;
    layer3_outputs(308) <= not (a or b);
    layer3_outputs(309) <= '1';
    layer3_outputs(310) <= b and not a;
    layer3_outputs(311) <= b;
    layer3_outputs(312) <= b and not a;
    layer3_outputs(313) <= a;
    layer3_outputs(314) <= a;
    layer3_outputs(315) <= not a;
    layer3_outputs(316) <= not b;
    layer3_outputs(317) <= b;
    layer3_outputs(318) <= a and not b;
    layer3_outputs(319) <= not a or b;
    layer3_outputs(320) <= b;
    layer3_outputs(321) <= not a;
    layer3_outputs(322) <= b;
    layer3_outputs(323) <= b;
    layer3_outputs(324) <= a and not b;
    layer3_outputs(325) <= a;
    layer3_outputs(326) <= not b;
    layer3_outputs(327) <= not (a and b);
    layer3_outputs(328) <= not a;
    layer3_outputs(329) <= b and not a;
    layer3_outputs(330) <= not b;
    layer3_outputs(331) <= a and b;
    layer3_outputs(332) <= a;
    layer3_outputs(333) <= a and not b;
    layer3_outputs(334) <= not a;
    layer3_outputs(335) <= a;
    layer3_outputs(336) <= not (a and b);
    layer3_outputs(337) <= a;
    layer3_outputs(338) <= a and b;
    layer3_outputs(339) <= not b or a;
    layer3_outputs(340) <= not a;
    layer3_outputs(341) <= '1';
    layer3_outputs(342) <= a or b;
    layer3_outputs(343) <= a and not b;
    layer3_outputs(344) <= '0';
    layer3_outputs(345) <= a xor b;
    layer3_outputs(346) <= '1';
    layer3_outputs(347) <= not (a or b);
    layer3_outputs(348) <= a xor b;
    layer3_outputs(349) <= a and not b;
    layer3_outputs(350) <= a xor b;
    layer3_outputs(351) <= b;
    layer3_outputs(352) <= not a or b;
    layer3_outputs(353) <= not a;
    layer3_outputs(354) <= '1';
    layer3_outputs(355) <= not (a or b);
    layer3_outputs(356) <= not (a and b);
    layer3_outputs(357) <= a and not b;
    layer3_outputs(358) <= a xor b;
    layer3_outputs(359) <= not b or a;
    layer3_outputs(360) <= b;
    layer3_outputs(361) <= not b;
    layer3_outputs(362) <= a or b;
    layer3_outputs(363) <= not b or a;
    layer3_outputs(364) <= a and not b;
    layer3_outputs(365) <= b and not a;
    layer3_outputs(366) <= a or b;
    layer3_outputs(367) <= not b;
    layer3_outputs(368) <= b;
    layer3_outputs(369) <= not b;
    layer3_outputs(370) <= not (a or b);
    layer3_outputs(371) <= not a or b;
    layer3_outputs(372) <= a and not b;
    layer3_outputs(373) <= a or b;
    layer3_outputs(374) <= not a;
    layer3_outputs(375) <= not a or b;
    layer3_outputs(376) <= '1';
    layer3_outputs(377) <= b;
    layer3_outputs(378) <= b;
    layer3_outputs(379) <= '1';
    layer3_outputs(380) <= not b or a;
    layer3_outputs(381) <= a and not b;
    layer3_outputs(382) <= not b;
    layer3_outputs(383) <= not a;
    layer3_outputs(384) <= not a;
    layer3_outputs(385) <= b;
    layer3_outputs(386) <= not b;
    layer3_outputs(387) <= '0';
    layer3_outputs(388) <= not a or b;
    layer3_outputs(389) <= not b or a;
    layer3_outputs(390) <= a;
    layer3_outputs(391) <= a;
    layer3_outputs(392) <= not b;
    layer3_outputs(393) <= '1';
    layer3_outputs(394) <= '0';
    layer3_outputs(395) <= not (a and b);
    layer3_outputs(396) <= not (a and b);
    layer3_outputs(397) <= not (a xor b);
    layer3_outputs(398) <= b;
    layer3_outputs(399) <= b;
    layer3_outputs(400) <= not a or b;
    layer3_outputs(401) <= not b;
    layer3_outputs(402) <= not b;
    layer3_outputs(403) <= not b or a;
    layer3_outputs(404) <= not b or a;
    layer3_outputs(405) <= not a or b;
    layer3_outputs(406) <= not a;
    layer3_outputs(407) <= not b or a;
    layer3_outputs(408) <= not b or a;
    layer3_outputs(409) <= not b;
    layer3_outputs(410) <= not a;
    layer3_outputs(411) <= a and not b;
    layer3_outputs(412) <= not a or b;
    layer3_outputs(413) <= a and not b;
    layer3_outputs(414) <= a and b;
    layer3_outputs(415) <= b;
    layer3_outputs(416) <= a and b;
    layer3_outputs(417) <= not b or a;
    layer3_outputs(418) <= not (a and b);
    layer3_outputs(419) <= not (a and b);
    layer3_outputs(420) <= not (a or b);
    layer3_outputs(421) <= b;
    layer3_outputs(422) <= not a;
    layer3_outputs(423) <= not a;
    layer3_outputs(424) <= not (a xor b);
    layer3_outputs(425) <= a or b;
    layer3_outputs(426) <= a or b;
    layer3_outputs(427) <= '1';
    layer3_outputs(428) <= '1';
    layer3_outputs(429) <= '1';
    layer3_outputs(430) <= not a or b;
    layer3_outputs(431) <= a and not b;
    layer3_outputs(432) <= not (a and b);
    layer3_outputs(433) <= not a;
    layer3_outputs(434) <= not b or a;
    layer3_outputs(435) <= b;
    layer3_outputs(436) <= b and not a;
    layer3_outputs(437) <= not b;
    layer3_outputs(438) <= a and b;
    layer3_outputs(439) <= a and not b;
    layer3_outputs(440) <= not b;
    layer3_outputs(441) <= not b or a;
    layer3_outputs(442) <= not (a or b);
    layer3_outputs(443) <= a xor b;
    layer3_outputs(444) <= '1';
    layer3_outputs(445) <= a and not b;
    layer3_outputs(446) <= not (a and b);
    layer3_outputs(447) <= not a;
    layer3_outputs(448) <= a and not b;
    layer3_outputs(449) <= b;
    layer3_outputs(450) <= not (a and b);
    layer3_outputs(451) <= b;
    layer3_outputs(452) <= a;
    layer3_outputs(453) <= '1';
    layer3_outputs(454) <= not (a or b);
    layer3_outputs(455) <= b;
    layer3_outputs(456) <= a;
    layer3_outputs(457) <= not (a xor b);
    layer3_outputs(458) <= not (a or b);
    layer3_outputs(459) <= b and not a;
    layer3_outputs(460) <= not (a or b);
    layer3_outputs(461) <= not (a or b);
    layer3_outputs(462) <= '1';
    layer3_outputs(463) <= not (a xor b);
    layer3_outputs(464) <= a or b;
    layer3_outputs(465) <= not a;
    layer3_outputs(466) <= not b or a;
    layer3_outputs(467) <= a and b;
    layer3_outputs(468) <= a and b;
    layer3_outputs(469) <= not a or b;
    layer3_outputs(470) <= not a;
    layer3_outputs(471) <= b;
    layer3_outputs(472) <= not b;
    layer3_outputs(473) <= b and not a;
    layer3_outputs(474) <= a;
    layer3_outputs(475) <= a or b;
    layer3_outputs(476) <= a;
    layer3_outputs(477) <= b;
    layer3_outputs(478) <= a;
    layer3_outputs(479) <= not a;
    layer3_outputs(480) <= a and b;
    layer3_outputs(481) <= a xor b;
    layer3_outputs(482) <= not a;
    layer3_outputs(483) <= not (a and b);
    layer3_outputs(484) <= b;
    layer3_outputs(485) <= b;
    layer3_outputs(486) <= b;
    layer3_outputs(487) <= a and not b;
    layer3_outputs(488) <= a;
    layer3_outputs(489) <= a xor b;
    layer3_outputs(490) <= b;
    layer3_outputs(491) <= '0';
    layer3_outputs(492) <= a or b;
    layer3_outputs(493) <= not b;
    layer3_outputs(494) <= a or b;
    layer3_outputs(495) <= b and not a;
    layer3_outputs(496) <= a and not b;
    layer3_outputs(497) <= a or b;
    layer3_outputs(498) <= a and b;
    layer3_outputs(499) <= not a or b;
    layer3_outputs(500) <= not a;
    layer3_outputs(501) <= '1';
    layer3_outputs(502) <= a and b;
    layer3_outputs(503) <= a and b;
    layer3_outputs(504) <= a or b;
    layer3_outputs(505) <= '0';
    layer3_outputs(506) <= '1';
    layer3_outputs(507) <= not b or a;
    layer3_outputs(508) <= not (a or b);
    layer3_outputs(509) <= not (a and b);
    layer3_outputs(510) <= not b;
    layer3_outputs(511) <= not (a xor b);
    layer3_outputs(512) <= '0';
    layer3_outputs(513) <= not b or a;
    layer3_outputs(514) <= not b or a;
    layer3_outputs(515) <= not b or a;
    layer3_outputs(516) <= a;
    layer3_outputs(517) <= not a;
    layer3_outputs(518) <= not (a or b);
    layer3_outputs(519) <= '0';
    layer3_outputs(520) <= not (a and b);
    layer3_outputs(521) <= not a or b;
    layer3_outputs(522) <= not a or b;
    layer3_outputs(523) <= not b;
    layer3_outputs(524) <= b;
    layer3_outputs(525) <= not a;
    layer3_outputs(526) <= b;
    layer3_outputs(527) <= not b or a;
    layer3_outputs(528) <= a and b;
    layer3_outputs(529) <= a;
    layer3_outputs(530) <= b and not a;
    layer3_outputs(531) <= not a;
    layer3_outputs(532) <= not (a or b);
    layer3_outputs(533) <= not a or b;
    layer3_outputs(534) <= '1';
    layer3_outputs(535) <= not a;
    layer3_outputs(536) <= a and b;
    layer3_outputs(537) <= a and not b;
    layer3_outputs(538) <= not b;
    layer3_outputs(539) <= a and b;
    layer3_outputs(540) <= b;
    layer3_outputs(541) <= '1';
    layer3_outputs(542) <= '0';
    layer3_outputs(543) <= '0';
    layer3_outputs(544) <= not b or a;
    layer3_outputs(545) <= a;
    layer3_outputs(546) <= not b;
    layer3_outputs(547) <= b and not a;
    layer3_outputs(548) <= not a or b;
    layer3_outputs(549) <= not a or b;
    layer3_outputs(550) <= a;
    layer3_outputs(551) <= not (a and b);
    layer3_outputs(552) <= not b or a;
    layer3_outputs(553) <= a or b;
    layer3_outputs(554) <= not b;
    layer3_outputs(555) <= not b or a;
    layer3_outputs(556) <= not (a or b);
    layer3_outputs(557) <= not b or a;
    layer3_outputs(558) <= not (a or b);
    layer3_outputs(559) <= b;
    layer3_outputs(560) <= not b or a;
    layer3_outputs(561) <= not a;
    layer3_outputs(562) <= b;
    layer3_outputs(563) <= '0';
    layer3_outputs(564) <= '0';
    layer3_outputs(565) <= not (a and b);
    layer3_outputs(566) <= b;
    layer3_outputs(567) <= not a or b;
    layer3_outputs(568) <= not (a and b);
    layer3_outputs(569) <= not b;
    layer3_outputs(570) <= not (a or b);
    layer3_outputs(571) <= a;
    layer3_outputs(572) <= b;
    layer3_outputs(573) <= not (a xor b);
    layer3_outputs(574) <= b;
    layer3_outputs(575) <= b;
    layer3_outputs(576) <= not b or a;
    layer3_outputs(577) <= '1';
    layer3_outputs(578) <= not b or a;
    layer3_outputs(579) <= '0';
    layer3_outputs(580) <= not a;
    layer3_outputs(581) <= not a;
    layer3_outputs(582) <= not a or b;
    layer3_outputs(583) <= b;
    layer3_outputs(584) <= '0';
    layer3_outputs(585) <= '1';
    layer3_outputs(586) <= not (a or b);
    layer3_outputs(587) <= b;
    layer3_outputs(588) <= a or b;
    layer3_outputs(589) <= not a;
    layer3_outputs(590) <= not (a or b);
    layer3_outputs(591) <= not b;
    layer3_outputs(592) <= not a or b;
    layer3_outputs(593) <= not (a and b);
    layer3_outputs(594) <= not b or a;
    layer3_outputs(595) <= not (a and b);
    layer3_outputs(596) <= not b or a;
    layer3_outputs(597) <= a or b;
    layer3_outputs(598) <= '1';
    layer3_outputs(599) <= a;
    layer3_outputs(600) <= not (a and b);
    layer3_outputs(601) <= not (a xor b);
    layer3_outputs(602) <= a and b;
    layer3_outputs(603) <= not b;
    layer3_outputs(604) <= not b or a;
    layer3_outputs(605) <= a and b;
    layer3_outputs(606) <= a or b;
    layer3_outputs(607) <= not a;
    layer3_outputs(608) <= a or b;
    layer3_outputs(609) <= a and not b;
    layer3_outputs(610) <= a and not b;
    layer3_outputs(611) <= not b;
    layer3_outputs(612) <= '0';
    layer3_outputs(613) <= not (a and b);
    layer3_outputs(614) <= a and b;
    layer3_outputs(615) <= not a or b;
    layer3_outputs(616) <= '0';
    layer3_outputs(617) <= not (a and b);
    layer3_outputs(618) <= not a or b;
    layer3_outputs(619) <= not (a or b);
    layer3_outputs(620) <= b;
    layer3_outputs(621) <= not a or b;
    layer3_outputs(622) <= a and b;
    layer3_outputs(623) <= a;
    layer3_outputs(624) <= a;
    layer3_outputs(625) <= a and b;
    layer3_outputs(626) <= a xor b;
    layer3_outputs(627) <= not a;
    layer3_outputs(628) <= not b;
    layer3_outputs(629) <= '0';
    layer3_outputs(630) <= b and not a;
    layer3_outputs(631) <= not (a and b);
    layer3_outputs(632) <= a;
    layer3_outputs(633) <= a and b;
    layer3_outputs(634) <= not (a xor b);
    layer3_outputs(635) <= '0';
    layer3_outputs(636) <= '1';
    layer3_outputs(637) <= b and not a;
    layer3_outputs(638) <= a or b;
    layer3_outputs(639) <= not b;
    layer3_outputs(640) <= not (a xor b);
    layer3_outputs(641) <= not a or b;
    layer3_outputs(642) <= a;
    layer3_outputs(643) <= not (a and b);
    layer3_outputs(644) <= not (a and b);
    layer3_outputs(645) <= b;
    layer3_outputs(646) <= a or b;
    layer3_outputs(647) <= not (a and b);
    layer3_outputs(648) <= b;
    layer3_outputs(649) <= a xor b;
    layer3_outputs(650) <= not (a and b);
    layer3_outputs(651) <= not a;
    layer3_outputs(652) <= a;
    layer3_outputs(653) <= not b;
    layer3_outputs(654) <= a;
    layer3_outputs(655) <= a and b;
    layer3_outputs(656) <= a and not b;
    layer3_outputs(657) <= not (a or b);
    layer3_outputs(658) <= not (a and b);
    layer3_outputs(659) <= b;
    layer3_outputs(660) <= not a;
    layer3_outputs(661) <= not a or b;
    layer3_outputs(662) <= not b or a;
    layer3_outputs(663) <= a and not b;
    layer3_outputs(664) <= a;
    layer3_outputs(665) <= b and not a;
    layer3_outputs(666) <= not (a xor b);
    layer3_outputs(667) <= not b;
    layer3_outputs(668) <= not a or b;
    layer3_outputs(669) <= b and not a;
    layer3_outputs(670) <= a;
    layer3_outputs(671) <= not a;
    layer3_outputs(672) <= not a;
    layer3_outputs(673) <= a and not b;
    layer3_outputs(674) <= not (a and b);
    layer3_outputs(675) <= a xor b;
    layer3_outputs(676) <= not b or a;
    layer3_outputs(677) <= a or b;
    layer3_outputs(678) <= '0';
    layer3_outputs(679) <= a and not b;
    layer3_outputs(680) <= b and not a;
    layer3_outputs(681) <= a;
    layer3_outputs(682) <= not (a or b);
    layer3_outputs(683) <= '0';
    layer3_outputs(684) <= not b or a;
    layer3_outputs(685) <= '0';
    layer3_outputs(686) <= a xor b;
    layer3_outputs(687) <= a and not b;
    layer3_outputs(688) <= not (a xor b);
    layer3_outputs(689) <= a and b;
    layer3_outputs(690) <= '0';
    layer3_outputs(691) <= a xor b;
    layer3_outputs(692) <= a and b;
    layer3_outputs(693) <= not a;
    layer3_outputs(694) <= not a or b;
    layer3_outputs(695) <= b and not a;
    layer3_outputs(696) <= not b;
    layer3_outputs(697) <= not (a or b);
    layer3_outputs(698) <= a xor b;
    layer3_outputs(699) <= not b or a;
    layer3_outputs(700) <= not a or b;
    layer3_outputs(701) <= not a or b;
    layer3_outputs(702) <= b and not a;
    layer3_outputs(703) <= b;
    layer3_outputs(704) <= a or b;
    layer3_outputs(705) <= a or b;
    layer3_outputs(706) <= a or b;
    layer3_outputs(707) <= a and b;
    layer3_outputs(708) <= not b or a;
    layer3_outputs(709) <= not (a or b);
    layer3_outputs(710) <= not b;
    layer3_outputs(711) <= not (a or b);
    layer3_outputs(712) <= a and b;
    layer3_outputs(713) <= not (a and b);
    layer3_outputs(714) <= b;
    layer3_outputs(715) <= '1';
    layer3_outputs(716) <= not (a or b);
    layer3_outputs(717) <= b;
    layer3_outputs(718) <= a xor b;
    layer3_outputs(719) <= not a or b;
    layer3_outputs(720) <= a and b;
    layer3_outputs(721) <= not (a or b);
    layer3_outputs(722) <= not b;
    layer3_outputs(723) <= a or b;
    layer3_outputs(724) <= not a or b;
    layer3_outputs(725) <= not (a or b);
    layer3_outputs(726) <= not b;
    layer3_outputs(727) <= not (a and b);
    layer3_outputs(728) <= b;
    layer3_outputs(729) <= not b;
    layer3_outputs(730) <= a;
    layer3_outputs(731) <= a and b;
    layer3_outputs(732) <= a and not b;
    layer3_outputs(733) <= not a or b;
    layer3_outputs(734) <= not a;
    layer3_outputs(735) <= not (a and b);
    layer3_outputs(736) <= a and not b;
    layer3_outputs(737) <= a;
    layer3_outputs(738) <= a;
    layer3_outputs(739) <= a;
    layer3_outputs(740) <= b and not a;
    layer3_outputs(741) <= b;
    layer3_outputs(742) <= not b;
    layer3_outputs(743) <= not b or a;
    layer3_outputs(744) <= a;
    layer3_outputs(745) <= b and not a;
    layer3_outputs(746) <= '1';
    layer3_outputs(747) <= not (a and b);
    layer3_outputs(748) <= not (a or b);
    layer3_outputs(749) <= not b or a;
    layer3_outputs(750) <= a and not b;
    layer3_outputs(751) <= not (a xor b);
    layer3_outputs(752) <= a;
    layer3_outputs(753) <= not (a xor b);
    layer3_outputs(754) <= b and not a;
    layer3_outputs(755) <= not a;
    layer3_outputs(756) <= not a;
    layer3_outputs(757) <= a or b;
    layer3_outputs(758) <= a and not b;
    layer3_outputs(759) <= b and not a;
    layer3_outputs(760) <= '0';
    layer3_outputs(761) <= not b;
    layer3_outputs(762) <= '0';
    layer3_outputs(763) <= not b;
    layer3_outputs(764) <= not b;
    layer3_outputs(765) <= not a or b;
    layer3_outputs(766) <= not b or a;
    layer3_outputs(767) <= a and b;
    layer3_outputs(768) <= not (a and b);
    layer3_outputs(769) <= not a;
    layer3_outputs(770) <= not (a xor b);
    layer3_outputs(771) <= '1';
    layer3_outputs(772) <= b and not a;
    layer3_outputs(773) <= b;
    layer3_outputs(774) <= b;
    layer3_outputs(775) <= not (a and b);
    layer3_outputs(776) <= '0';
    layer3_outputs(777) <= a and not b;
    layer3_outputs(778) <= not a or b;
    layer3_outputs(779) <= not b;
    layer3_outputs(780) <= not (a or b);
    layer3_outputs(781) <= not a;
    layer3_outputs(782) <= not (a and b);
    layer3_outputs(783) <= not a or b;
    layer3_outputs(784) <= not (a xor b);
    layer3_outputs(785) <= a and b;
    layer3_outputs(786) <= not b;
    layer3_outputs(787) <= a;
    layer3_outputs(788) <= not (a or b);
    layer3_outputs(789) <= a;
    layer3_outputs(790) <= b and not a;
    layer3_outputs(791) <= not (a xor b);
    layer3_outputs(792) <= a or b;
    layer3_outputs(793) <= not a or b;
    layer3_outputs(794) <= not (a and b);
    layer3_outputs(795) <= not a or b;
    layer3_outputs(796) <= a;
    layer3_outputs(797) <= a or b;
    layer3_outputs(798) <= b and not a;
    layer3_outputs(799) <= b and not a;
    layer3_outputs(800) <= a and b;
    layer3_outputs(801) <= not b or a;
    layer3_outputs(802) <= not (a or b);
    layer3_outputs(803) <= not (a and b);
    layer3_outputs(804) <= b and not a;
    layer3_outputs(805) <= a and not b;
    layer3_outputs(806) <= a and b;
    layer3_outputs(807) <= a or b;
    layer3_outputs(808) <= a and b;
    layer3_outputs(809) <= not b or a;
    layer3_outputs(810) <= a and not b;
    layer3_outputs(811) <= a or b;
    layer3_outputs(812) <= not (a and b);
    layer3_outputs(813) <= '0';
    layer3_outputs(814) <= not b or a;
    layer3_outputs(815) <= b;
    layer3_outputs(816) <= not b;
    layer3_outputs(817) <= a and not b;
    layer3_outputs(818) <= a and b;
    layer3_outputs(819) <= '1';
    layer3_outputs(820) <= not a;
    layer3_outputs(821) <= not a or b;
    layer3_outputs(822) <= not a;
    layer3_outputs(823) <= b;
    layer3_outputs(824) <= not a;
    layer3_outputs(825) <= not (a and b);
    layer3_outputs(826) <= b;
    layer3_outputs(827) <= b;
    layer3_outputs(828) <= not b or a;
    layer3_outputs(829) <= not (a and b);
    layer3_outputs(830) <= not a;
    layer3_outputs(831) <= b;
    layer3_outputs(832) <= b;
    layer3_outputs(833) <= not (a and b);
    layer3_outputs(834) <= b;
    layer3_outputs(835) <= not (a and b);
    layer3_outputs(836) <= a;
    layer3_outputs(837) <= a or b;
    layer3_outputs(838) <= a or b;
    layer3_outputs(839) <= b and not a;
    layer3_outputs(840) <= not b;
    layer3_outputs(841) <= not b;
    layer3_outputs(842) <= a and b;
    layer3_outputs(843) <= not a;
    layer3_outputs(844) <= a and b;
    layer3_outputs(845) <= '0';
    layer3_outputs(846) <= a;
    layer3_outputs(847) <= not (a xor b);
    layer3_outputs(848) <= not a;
    layer3_outputs(849) <= not (a and b);
    layer3_outputs(850) <= a;
    layer3_outputs(851) <= a and b;
    layer3_outputs(852) <= not b;
    layer3_outputs(853) <= a or b;
    layer3_outputs(854) <= a xor b;
    layer3_outputs(855) <= b and not a;
    layer3_outputs(856) <= '1';
    layer3_outputs(857) <= a xor b;
    layer3_outputs(858) <= not a or b;
    layer3_outputs(859) <= a;
    layer3_outputs(860) <= a xor b;
    layer3_outputs(861) <= a;
    layer3_outputs(862) <= not b or a;
    layer3_outputs(863) <= a;
    layer3_outputs(864) <= a and not b;
    layer3_outputs(865) <= a;
    layer3_outputs(866) <= '0';
    layer3_outputs(867) <= not a;
    layer3_outputs(868) <= a and not b;
    layer3_outputs(869) <= a and not b;
    layer3_outputs(870) <= b and not a;
    layer3_outputs(871) <= not a or b;
    layer3_outputs(872) <= not a or b;
    layer3_outputs(873) <= not a;
    layer3_outputs(874) <= not b;
    layer3_outputs(875) <= a and not b;
    layer3_outputs(876) <= a xor b;
    layer3_outputs(877) <= not a or b;
    layer3_outputs(878) <= a;
    layer3_outputs(879) <= not (a or b);
    layer3_outputs(880) <= not (a xor b);
    layer3_outputs(881) <= not (a and b);
    layer3_outputs(882) <= a or b;
    layer3_outputs(883) <= not a;
    layer3_outputs(884) <= a xor b;
    layer3_outputs(885) <= not (a or b);
    layer3_outputs(886) <= b;
    layer3_outputs(887) <= not b;
    layer3_outputs(888) <= not b;
    layer3_outputs(889) <= '0';
    layer3_outputs(890) <= not a;
    layer3_outputs(891) <= not b or a;
    layer3_outputs(892) <= a or b;
    layer3_outputs(893) <= '0';
    layer3_outputs(894) <= b and not a;
    layer3_outputs(895) <= '0';
    layer3_outputs(896) <= not a;
    layer3_outputs(897) <= not a;
    layer3_outputs(898) <= a;
    layer3_outputs(899) <= a xor b;
    layer3_outputs(900) <= not (a and b);
    layer3_outputs(901) <= a;
    layer3_outputs(902) <= not a;
    layer3_outputs(903) <= not b;
    layer3_outputs(904) <= '1';
    layer3_outputs(905) <= not (a xor b);
    layer3_outputs(906) <= b and not a;
    layer3_outputs(907) <= b;
    layer3_outputs(908) <= a;
    layer3_outputs(909) <= b and not a;
    layer3_outputs(910) <= a or b;
    layer3_outputs(911) <= not b;
    layer3_outputs(912) <= not b;
    layer3_outputs(913) <= a or b;
    layer3_outputs(914) <= not (a xor b);
    layer3_outputs(915) <= not a or b;
    layer3_outputs(916) <= b and not a;
    layer3_outputs(917) <= a or b;
    layer3_outputs(918) <= not (a or b);
    layer3_outputs(919) <= not (a or b);
    layer3_outputs(920) <= a or b;
    layer3_outputs(921) <= a or b;
    layer3_outputs(922) <= not (a and b);
    layer3_outputs(923) <= '0';
    layer3_outputs(924) <= b and not a;
    layer3_outputs(925) <= a;
    layer3_outputs(926) <= not b;
    layer3_outputs(927) <= not b;
    layer3_outputs(928) <= not b;
    layer3_outputs(929) <= a;
    layer3_outputs(930) <= a xor b;
    layer3_outputs(931) <= a xor b;
    layer3_outputs(932) <= not b;
    layer3_outputs(933) <= not a or b;
    layer3_outputs(934) <= not (a xor b);
    layer3_outputs(935) <= a or b;
    layer3_outputs(936) <= not a;
    layer3_outputs(937) <= a xor b;
    layer3_outputs(938) <= a and not b;
    layer3_outputs(939) <= b and not a;
    layer3_outputs(940) <= not (a and b);
    layer3_outputs(941) <= b;
    layer3_outputs(942) <= not a;
    layer3_outputs(943) <= a;
    layer3_outputs(944) <= a xor b;
    layer3_outputs(945) <= b and not a;
    layer3_outputs(946) <= not (a and b);
    layer3_outputs(947) <= '0';
    layer3_outputs(948) <= not a or b;
    layer3_outputs(949) <= b;
    layer3_outputs(950) <= not b or a;
    layer3_outputs(951) <= not (a and b);
    layer3_outputs(952) <= not a;
    layer3_outputs(953) <= not b or a;
    layer3_outputs(954) <= not b or a;
    layer3_outputs(955) <= a or b;
    layer3_outputs(956) <= not (a and b);
    layer3_outputs(957) <= b and not a;
    layer3_outputs(958) <= not a;
    layer3_outputs(959) <= not (a or b);
    layer3_outputs(960) <= not b;
    layer3_outputs(961) <= not b or a;
    layer3_outputs(962) <= not a;
    layer3_outputs(963) <= not a;
    layer3_outputs(964) <= a or b;
    layer3_outputs(965) <= b and not a;
    layer3_outputs(966) <= a and not b;
    layer3_outputs(967) <= a;
    layer3_outputs(968) <= b and not a;
    layer3_outputs(969) <= not (a or b);
    layer3_outputs(970) <= a or b;
    layer3_outputs(971) <= b and not a;
    layer3_outputs(972) <= a and b;
    layer3_outputs(973) <= not (a and b);
    layer3_outputs(974) <= not a or b;
    layer3_outputs(975) <= not (a or b);
    layer3_outputs(976) <= '0';
    layer3_outputs(977) <= a;
    layer3_outputs(978) <= not a or b;
    layer3_outputs(979) <= '1';
    layer3_outputs(980) <= a or b;
    layer3_outputs(981) <= not a;
    layer3_outputs(982) <= b;
    layer3_outputs(983) <= a;
    layer3_outputs(984) <= not a;
    layer3_outputs(985) <= b;
    layer3_outputs(986) <= not b or a;
    layer3_outputs(987) <= not a or b;
    layer3_outputs(988) <= '1';
    layer3_outputs(989) <= not a;
    layer3_outputs(990) <= '1';
    layer3_outputs(991) <= b;
    layer3_outputs(992) <= not b;
    layer3_outputs(993) <= not b;
    layer3_outputs(994) <= a;
    layer3_outputs(995) <= a xor b;
    layer3_outputs(996) <= not (a or b);
    layer3_outputs(997) <= a;
    layer3_outputs(998) <= b;
    layer3_outputs(999) <= not a or b;
    layer3_outputs(1000) <= a and not b;
    layer3_outputs(1001) <= not (a or b);
    layer3_outputs(1002) <= b and not a;
    layer3_outputs(1003) <= a xor b;
    layer3_outputs(1004) <= not b;
    layer3_outputs(1005) <= a or b;
    layer3_outputs(1006) <= not a or b;
    layer3_outputs(1007) <= a;
    layer3_outputs(1008) <= a and not b;
    layer3_outputs(1009) <= a;
    layer3_outputs(1010) <= not (a xor b);
    layer3_outputs(1011) <= not b;
    layer3_outputs(1012) <= a;
    layer3_outputs(1013) <= b and not a;
    layer3_outputs(1014) <= a;
    layer3_outputs(1015) <= '1';
    layer3_outputs(1016) <= a and not b;
    layer3_outputs(1017) <= b and not a;
    layer3_outputs(1018) <= a and b;
    layer3_outputs(1019) <= a and not b;
    layer3_outputs(1020) <= not b or a;
    layer3_outputs(1021) <= a and not b;
    layer3_outputs(1022) <= b;
    layer3_outputs(1023) <= a;
    layer3_outputs(1024) <= not b or a;
    layer3_outputs(1025) <= a;
    layer3_outputs(1026) <= not b or a;
    layer3_outputs(1027) <= a or b;
    layer3_outputs(1028) <= not (a and b);
    layer3_outputs(1029) <= '0';
    layer3_outputs(1030) <= not (a or b);
    layer3_outputs(1031) <= a xor b;
    layer3_outputs(1032) <= a xor b;
    layer3_outputs(1033) <= not (a or b);
    layer3_outputs(1034) <= a and b;
    layer3_outputs(1035) <= not (a or b);
    layer3_outputs(1036) <= not a or b;
    layer3_outputs(1037) <= '1';
    layer3_outputs(1038) <= a and b;
    layer3_outputs(1039) <= a or b;
    layer3_outputs(1040) <= not (a or b);
    layer3_outputs(1041) <= not a or b;
    layer3_outputs(1042) <= '0';
    layer3_outputs(1043) <= not (a and b);
    layer3_outputs(1044) <= not b or a;
    layer3_outputs(1045) <= a xor b;
    layer3_outputs(1046) <= b;
    layer3_outputs(1047) <= not b;
    layer3_outputs(1048) <= b and not a;
    layer3_outputs(1049) <= not b;
    layer3_outputs(1050) <= a or b;
    layer3_outputs(1051) <= not a;
    layer3_outputs(1052) <= not a or b;
    layer3_outputs(1053) <= a and not b;
    layer3_outputs(1054) <= not a;
    layer3_outputs(1055) <= a xor b;
    layer3_outputs(1056) <= a or b;
    layer3_outputs(1057) <= not a;
    layer3_outputs(1058) <= not a;
    layer3_outputs(1059) <= b;
    layer3_outputs(1060) <= not b;
    layer3_outputs(1061) <= not a or b;
    layer3_outputs(1062) <= not (a and b);
    layer3_outputs(1063) <= b;
    layer3_outputs(1064) <= not (a and b);
    layer3_outputs(1065) <= not b or a;
    layer3_outputs(1066) <= not a;
    layer3_outputs(1067) <= b;
    layer3_outputs(1068) <= not (a xor b);
    layer3_outputs(1069) <= a or b;
    layer3_outputs(1070) <= not (a and b);
    layer3_outputs(1071) <= not b or a;
    layer3_outputs(1072) <= b;
    layer3_outputs(1073) <= not a;
    layer3_outputs(1074) <= a;
    layer3_outputs(1075) <= not a;
    layer3_outputs(1076) <= a and b;
    layer3_outputs(1077) <= not a or b;
    layer3_outputs(1078) <= b and not a;
    layer3_outputs(1079) <= a and b;
    layer3_outputs(1080) <= '0';
    layer3_outputs(1081) <= a and b;
    layer3_outputs(1082) <= b;
    layer3_outputs(1083) <= a and not b;
    layer3_outputs(1084) <= '1';
    layer3_outputs(1085) <= '0';
    layer3_outputs(1086) <= a and b;
    layer3_outputs(1087) <= a;
    layer3_outputs(1088) <= '0';
    layer3_outputs(1089) <= b;
    layer3_outputs(1090) <= not b;
    layer3_outputs(1091) <= a xor b;
    layer3_outputs(1092) <= '1';
    layer3_outputs(1093) <= not b or a;
    layer3_outputs(1094) <= not b or a;
    layer3_outputs(1095) <= not a;
    layer3_outputs(1096) <= b;
    layer3_outputs(1097) <= not (a xor b);
    layer3_outputs(1098) <= not a;
    layer3_outputs(1099) <= not (a xor b);
    layer3_outputs(1100) <= b;
    layer3_outputs(1101) <= not b;
    layer3_outputs(1102) <= b and not a;
    layer3_outputs(1103) <= not (a or b);
    layer3_outputs(1104) <= not a or b;
    layer3_outputs(1105) <= not a;
    layer3_outputs(1106) <= '0';
    layer3_outputs(1107) <= not (a or b);
    layer3_outputs(1108) <= a or b;
    layer3_outputs(1109) <= not (a or b);
    layer3_outputs(1110) <= a;
    layer3_outputs(1111) <= not b;
    layer3_outputs(1112) <= a or b;
    layer3_outputs(1113) <= not a or b;
    layer3_outputs(1114) <= not a or b;
    layer3_outputs(1115) <= not a;
    layer3_outputs(1116) <= a and not b;
    layer3_outputs(1117) <= b and not a;
    layer3_outputs(1118) <= a and b;
    layer3_outputs(1119) <= a and b;
    layer3_outputs(1120) <= not (a and b);
    layer3_outputs(1121) <= b and not a;
    layer3_outputs(1122) <= a;
    layer3_outputs(1123) <= b;
    layer3_outputs(1124) <= a;
    layer3_outputs(1125) <= not b or a;
    layer3_outputs(1126) <= not a;
    layer3_outputs(1127) <= a and not b;
    layer3_outputs(1128) <= a;
    layer3_outputs(1129) <= not (a and b);
    layer3_outputs(1130) <= not a or b;
    layer3_outputs(1131) <= not (a or b);
    layer3_outputs(1132) <= a or b;
    layer3_outputs(1133) <= not b;
    layer3_outputs(1134) <= a and not b;
    layer3_outputs(1135) <= not a or b;
    layer3_outputs(1136) <= b and not a;
    layer3_outputs(1137) <= not (a or b);
    layer3_outputs(1138) <= b and not a;
    layer3_outputs(1139) <= a and not b;
    layer3_outputs(1140) <= not (a xor b);
    layer3_outputs(1141) <= not (a and b);
    layer3_outputs(1142) <= b;
    layer3_outputs(1143) <= a;
    layer3_outputs(1144) <= a;
    layer3_outputs(1145) <= a;
    layer3_outputs(1146) <= not (a and b);
    layer3_outputs(1147) <= b;
    layer3_outputs(1148) <= not (a and b);
    layer3_outputs(1149) <= a;
    layer3_outputs(1150) <= not a;
    layer3_outputs(1151) <= not a;
    layer3_outputs(1152) <= b;
    layer3_outputs(1153) <= not b;
    layer3_outputs(1154) <= a xor b;
    layer3_outputs(1155) <= not (a and b);
    layer3_outputs(1156) <= a xor b;
    layer3_outputs(1157) <= not b or a;
    layer3_outputs(1158) <= not b;
    layer3_outputs(1159) <= not b or a;
    layer3_outputs(1160) <= not (a or b);
    layer3_outputs(1161) <= not (a and b);
    layer3_outputs(1162) <= b and not a;
    layer3_outputs(1163) <= not b;
    layer3_outputs(1164) <= '0';
    layer3_outputs(1165) <= a;
    layer3_outputs(1166) <= not b or a;
    layer3_outputs(1167) <= not (a and b);
    layer3_outputs(1168) <= not b;
    layer3_outputs(1169) <= a and b;
    layer3_outputs(1170) <= not a;
    layer3_outputs(1171) <= b and not a;
    layer3_outputs(1172) <= b and not a;
    layer3_outputs(1173) <= not b;
    layer3_outputs(1174) <= not b;
    layer3_outputs(1175) <= a and b;
    layer3_outputs(1176) <= not b;
    layer3_outputs(1177) <= b;
    layer3_outputs(1178) <= not a or b;
    layer3_outputs(1179) <= a and b;
    layer3_outputs(1180) <= not b or a;
    layer3_outputs(1181) <= a and b;
    layer3_outputs(1182) <= a and not b;
    layer3_outputs(1183) <= not a;
    layer3_outputs(1184) <= not a;
    layer3_outputs(1185) <= a xor b;
    layer3_outputs(1186) <= not a;
    layer3_outputs(1187) <= not b;
    layer3_outputs(1188) <= not b or a;
    layer3_outputs(1189) <= a and not b;
    layer3_outputs(1190) <= not a;
    layer3_outputs(1191) <= a or b;
    layer3_outputs(1192) <= a and b;
    layer3_outputs(1193) <= not (a xor b);
    layer3_outputs(1194) <= b;
    layer3_outputs(1195) <= a;
    layer3_outputs(1196) <= a and not b;
    layer3_outputs(1197) <= not (a and b);
    layer3_outputs(1198) <= a or b;
    layer3_outputs(1199) <= not (a or b);
    layer3_outputs(1200) <= b and not a;
    layer3_outputs(1201) <= a xor b;
    layer3_outputs(1202) <= not (a or b);
    layer3_outputs(1203) <= not a;
    layer3_outputs(1204) <= not a;
    layer3_outputs(1205) <= not (a xor b);
    layer3_outputs(1206) <= not a;
    layer3_outputs(1207) <= not a or b;
    layer3_outputs(1208) <= '1';
    layer3_outputs(1209) <= a or b;
    layer3_outputs(1210) <= not (a or b);
    layer3_outputs(1211) <= not (a or b);
    layer3_outputs(1212) <= a and b;
    layer3_outputs(1213) <= not a or b;
    layer3_outputs(1214) <= a or b;
    layer3_outputs(1215) <= not a or b;
    layer3_outputs(1216) <= a;
    layer3_outputs(1217) <= not a or b;
    layer3_outputs(1218) <= a;
    layer3_outputs(1219) <= a or b;
    layer3_outputs(1220) <= b and not a;
    layer3_outputs(1221) <= not (a xor b);
    layer3_outputs(1222) <= not a or b;
    layer3_outputs(1223) <= a and not b;
    layer3_outputs(1224) <= a and b;
    layer3_outputs(1225) <= b;
    layer3_outputs(1226) <= b and not a;
    layer3_outputs(1227) <= not b or a;
    layer3_outputs(1228) <= not a;
    layer3_outputs(1229) <= a and b;
    layer3_outputs(1230) <= '1';
    layer3_outputs(1231) <= not b or a;
    layer3_outputs(1232) <= a;
    layer3_outputs(1233) <= '0';
    layer3_outputs(1234) <= not b or a;
    layer3_outputs(1235) <= not (a or b);
    layer3_outputs(1236) <= a and b;
    layer3_outputs(1237) <= not b or a;
    layer3_outputs(1238) <= not b or a;
    layer3_outputs(1239) <= not a;
    layer3_outputs(1240) <= a xor b;
    layer3_outputs(1241) <= b and not a;
    layer3_outputs(1242) <= b and not a;
    layer3_outputs(1243) <= not a;
    layer3_outputs(1244) <= b and not a;
    layer3_outputs(1245) <= not (a or b);
    layer3_outputs(1246) <= '0';
    layer3_outputs(1247) <= not a;
    layer3_outputs(1248) <= not (a or b);
    layer3_outputs(1249) <= a or b;
    layer3_outputs(1250) <= a;
    layer3_outputs(1251) <= not b or a;
    layer3_outputs(1252) <= '1';
    layer3_outputs(1253) <= not b;
    layer3_outputs(1254) <= a and b;
    layer3_outputs(1255) <= a and b;
    layer3_outputs(1256) <= a and not b;
    layer3_outputs(1257) <= not b;
    layer3_outputs(1258) <= a;
    layer3_outputs(1259) <= b;
    layer3_outputs(1260) <= a xor b;
    layer3_outputs(1261) <= not a or b;
    layer3_outputs(1262) <= b and not a;
    layer3_outputs(1263) <= not b;
    layer3_outputs(1264) <= b and not a;
    layer3_outputs(1265) <= b;
    layer3_outputs(1266) <= not a;
    layer3_outputs(1267) <= not b or a;
    layer3_outputs(1268) <= b and not a;
    layer3_outputs(1269) <= not b;
    layer3_outputs(1270) <= a and b;
    layer3_outputs(1271) <= not a;
    layer3_outputs(1272) <= b;
    layer3_outputs(1273) <= a or b;
    layer3_outputs(1274) <= not b;
    layer3_outputs(1275) <= not b or a;
    layer3_outputs(1276) <= a and b;
    layer3_outputs(1277) <= a or b;
    layer3_outputs(1278) <= b;
    layer3_outputs(1279) <= not a;
    layer3_outputs(1280) <= b;
    layer3_outputs(1281) <= a and not b;
    layer3_outputs(1282) <= b;
    layer3_outputs(1283) <= b and not a;
    layer3_outputs(1284) <= not (a and b);
    layer3_outputs(1285) <= not a or b;
    layer3_outputs(1286) <= a and not b;
    layer3_outputs(1287) <= not a or b;
    layer3_outputs(1288) <= b and not a;
    layer3_outputs(1289) <= not b;
    layer3_outputs(1290) <= a and not b;
    layer3_outputs(1291) <= not a;
    layer3_outputs(1292) <= '1';
    layer3_outputs(1293) <= b and not a;
    layer3_outputs(1294) <= a and not b;
    layer3_outputs(1295) <= not b;
    layer3_outputs(1296) <= not b;
    layer3_outputs(1297) <= '1';
    layer3_outputs(1298) <= not a;
    layer3_outputs(1299) <= a or b;
    layer3_outputs(1300) <= not (a xor b);
    layer3_outputs(1301) <= '0';
    layer3_outputs(1302) <= b and not a;
    layer3_outputs(1303) <= b;
    layer3_outputs(1304) <= not a;
    layer3_outputs(1305) <= not a;
    layer3_outputs(1306) <= b;
    layer3_outputs(1307) <= not a or b;
    layer3_outputs(1308) <= not a;
    layer3_outputs(1309) <= a and not b;
    layer3_outputs(1310) <= a xor b;
    layer3_outputs(1311) <= a;
    layer3_outputs(1312) <= b;
    layer3_outputs(1313) <= not (a or b);
    layer3_outputs(1314) <= not (a or b);
    layer3_outputs(1315) <= not (a and b);
    layer3_outputs(1316) <= not a;
    layer3_outputs(1317) <= a or b;
    layer3_outputs(1318) <= b;
    layer3_outputs(1319) <= a;
    layer3_outputs(1320) <= not b;
    layer3_outputs(1321) <= not (a and b);
    layer3_outputs(1322) <= not (a xor b);
    layer3_outputs(1323) <= a xor b;
    layer3_outputs(1324) <= not (a xor b);
    layer3_outputs(1325) <= a and not b;
    layer3_outputs(1326) <= not (a or b);
    layer3_outputs(1327) <= not (a or b);
    layer3_outputs(1328) <= not (a or b);
    layer3_outputs(1329) <= a and not b;
    layer3_outputs(1330) <= a and not b;
    layer3_outputs(1331) <= not (a xor b);
    layer3_outputs(1332) <= not a;
    layer3_outputs(1333) <= b;
    layer3_outputs(1334) <= not (a or b);
    layer3_outputs(1335) <= not (a and b);
    layer3_outputs(1336) <= a and not b;
    layer3_outputs(1337) <= b and not a;
    layer3_outputs(1338) <= a or b;
    layer3_outputs(1339) <= b;
    layer3_outputs(1340) <= a and not b;
    layer3_outputs(1341) <= b;
    layer3_outputs(1342) <= not b;
    layer3_outputs(1343) <= b;
    layer3_outputs(1344) <= not (a or b);
    layer3_outputs(1345) <= a;
    layer3_outputs(1346) <= not b or a;
    layer3_outputs(1347) <= a;
    layer3_outputs(1348) <= not (a xor b);
    layer3_outputs(1349) <= not a or b;
    layer3_outputs(1350) <= b;
    layer3_outputs(1351) <= a;
    layer3_outputs(1352) <= not a or b;
    layer3_outputs(1353) <= not a;
    layer3_outputs(1354) <= not (a xor b);
    layer3_outputs(1355) <= not a;
    layer3_outputs(1356) <= a and not b;
    layer3_outputs(1357) <= a and not b;
    layer3_outputs(1358) <= b and not a;
    layer3_outputs(1359) <= not b;
    layer3_outputs(1360) <= a and b;
    layer3_outputs(1361) <= not (a or b);
    layer3_outputs(1362) <= not (a and b);
    layer3_outputs(1363) <= a;
    layer3_outputs(1364) <= not a or b;
    layer3_outputs(1365) <= not (a or b);
    layer3_outputs(1366) <= a and b;
    layer3_outputs(1367) <= not a;
    layer3_outputs(1368) <= b and not a;
    layer3_outputs(1369) <= not (a and b);
    layer3_outputs(1370) <= a or b;
    layer3_outputs(1371) <= a or b;
    layer3_outputs(1372) <= not a;
    layer3_outputs(1373) <= not b;
    layer3_outputs(1374) <= not b;
    layer3_outputs(1375) <= not b;
    layer3_outputs(1376) <= b;
    layer3_outputs(1377) <= a;
    layer3_outputs(1378) <= a;
    layer3_outputs(1379) <= not a;
    layer3_outputs(1380) <= not b;
    layer3_outputs(1381) <= not (a or b);
    layer3_outputs(1382) <= not a or b;
    layer3_outputs(1383) <= a;
    layer3_outputs(1384) <= not b;
    layer3_outputs(1385) <= a or b;
    layer3_outputs(1386) <= a or b;
    layer3_outputs(1387) <= a;
    layer3_outputs(1388) <= a xor b;
    layer3_outputs(1389) <= not (a or b);
    layer3_outputs(1390) <= a xor b;
    layer3_outputs(1391) <= not a;
    layer3_outputs(1392) <= not b or a;
    layer3_outputs(1393) <= a xor b;
    layer3_outputs(1394) <= a;
    layer3_outputs(1395) <= '1';
    layer3_outputs(1396) <= not a;
    layer3_outputs(1397) <= b and not a;
    layer3_outputs(1398) <= not b;
    layer3_outputs(1399) <= not a;
    layer3_outputs(1400) <= b;
    layer3_outputs(1401) <= a;
    layer3_outputs(1402) <= not b or a;
    layer3_outputs(1403) <= not a;
    layer3_outputs(1404) <= a or b;
    layer3_outputs(1405) <= a or b;
    layer3_outputs(1406) <= a and b;
    layer3_outputs(1407) <= not (a xor b);
    layer3_outputs(1408) <= a and not b;
    layer3_outputs(1409) <= not a;
    layer3_outputs(1410) <= not a or b;
    layer3_outputs(1411) <= not a or b;
    layer3_outputs(1412) <= a or b;
    layer3_outputs(1413) <= not (a and b);
    layer3_outputs(1414) <= a or b;
    layer3_outputs(1415) <= b and not a;
    layer3_outputs(1416) <= '0';
    layer3_outputs(1417) <= not b or a;
    layer3_outputs(1418) <= '0';
    layer3_outputs(1419) <= '0';
    layer3_outputs(1420) <= a and b;
    layer3_outputs(1421) <= a or b;
    layer3_outputs(1422) <= b and not a;
    layer3_outputs(1423) <= a;
    layer3_outputs(1424) <= not b or a;
    layer3_outputs(1425) <= not (a or b);
    layer3_outputs(1426) <= not (a xor b);
    layer3_outputs(1427) <= a or b;
    layer3_outputs(1428) <= not b;
    layer3_outputs(1429) <= not b;
    layer3_outputs(1430) <= not b;
    layer3_outputs(1431) <= not a;
    layer3_outputs(1432) <= not b or a;
    layer3_outputs(1433) <= not b;
    layer3_outputs(1434) <= not a;
    layer3_outputs(1435) <= not b or a;
    layer3_outputs(1436) <= not (a or b);
    layer3_outputs(1437) <= a and not b;
    layer3_outputs(1438) <= not (a and b);
    layer3_outputs(1439) <= not (a and b);
    layer3_outputs(1440) <= a;
    layer3_outputs(1441) <= not a;
    layer3_outputs(1442) <= not a;
    layer3_outputs(1443) <= b;
    layer3_outputs(1444) <= not b or a;
    layer3_outputs(1445) <= a and not b;
    layer3_outputs(1446) <= b;
    layer3_outputs(1447) <= a or b;
    layer3_outputs(1448) <= not (a and b);
    layer3_outputs(1449) <= b;
    layer3_outputs(1450) <= not (a xor b);
    layer3_outputs(1451) <= not a;
    layer3_outputs(1452) <= b and not a;
    layer3_outputs(1453) <= not a or b;
    layer3_outputs(1454) <= b;
    layer3_outputs(1455) <= b;
    layer3_outputs(1456) <= not b or a;
    layer3_outputs(1457) <= a or b;
    layer3_outputs(1458) <= not (a xor b);
    layer3_outputs(1459) <= '1';
    layer3_outputs(1460) <= '0';
    layer3_outputs(1461) <= a or b;
    layer3_outputs(1462) <= not (a and b);
    layer3_outputs(1463) <= not b or a;
    layer3_outputs(1464) <= b;
    layer3_outputs(1465) <= a xor b;
    layer3_outputs(1466) <= not b;
    layer3_outputs(1467) <= not (a or b);
    layer3_outputs(1468) <= not (a or b);
    layer3_outputs(1469) <= b;
    layer3_outputs(1470) <= not b;
    layer3_outputs(1471) <= a and b;
    layer3_outputs(1472) <= a and not b;
    layer3_outputs(1473) <= not (a or b);
    layer3_outputs(1474) <= b and not a;
    layer3_outputs(1475) <= not b;
    layer3_outputs(1476) <= not a;
    layer3_outputs(1477) <= a and not b;
    layer3_outputs(1478) <= not a;
    layer3_outputs(1479) <= a;
    layer3_outputs(1480) <= a and b;
    layer3_outputs(1481) <= not b;
    layer3_outputs(1482) <= not b;
    layer3_outputs(1483) <= not (a and b);
    layer3_outputs(1484) <= not b;
    layer3_outputs(1485) <= not (a and b);
    layer3_outputs(1486) <= '1';
    layer3_outputs(1487) <= not b or a;
    layer3_outputs(1488) <= a or b;
    layer3_outputs(1489) <= b;
    layer3_outputs(1490) <= a and b;
    layer3_outputs(1491) <= not b;
    layer3_outputs(1492) <= not a;
    layer3_outputs(1493) <= not (a and b);
    layer3_outputs(1494) <= '1';
    layer3_outputs(1495) <= a or b;
    layer3_outputs(1496) <= a;
    layer3_outputs(1497) <= not b;
    layer3_outputs(1498) <= a xor b;
    layer3_outputs(1499) <= a xor b;
    layer3_outputs(1500) <= not (a or b);
    layer3_outputs(1501) <= b;
    layer3_outputs(1502) <= not b or a;
    layer3_outputs(1503) <= b and not a;
    layer3_outputs(1504) <= not (a or b);
    layer3_outputs(1505) <= not b;
    layer3_outputs(1506) <= a or b;
    layer3_outputs(1507) <= b;
    layer3_outputs(1508) <= a and not b;
    layer3_outputs(1509) <= not b;
    layer3_outputs(1510) <= not b or a;
    layer3_outputs(1511) <= not b;
    layer3_outputs(1512) <= a xor b;
    layer3_outputs(1513) <= a xor b;
    layer3_outputs(1514) <= not a;
    layer3_outputs(1515) <= not a or b;
    layer3_outputs(1516) <= not b or a;
    layer3_outputs(1517) <= not b;
    layer3_outputs(1518) <= a;
    layer3_outputs(1519) <= not b;
    layer3_outputs(1520) <= a and b;
    layer3_outputs(1521) <= not (a xor b);
    layer3_outputs(1522) <= '0';
    layer3_outputs(1523) <= a and b;
    layer3_outputs(1524) <= not a;
    layer3_outputs(1525) <= b and not a;
    layer3_outputs(1526) <= a and b;
    layer3_outputs(1527) <= a and b;
    layer3_outputs(1528) <= a and not b;
    layer3_outputs(1529) <= a or b;
    layer3_outputs(1530) <= b;
    layer3_outputs(1531) <= a;
    layer3_outputs(1532) <= a or b;
    layer3_outputs(1533) <= b;
    layer3_outputs(1534) <= not (a and b);
    layer3_outputs(1535) <= '1';
    layer3_outputs(1536) <= b;
    layer3_outputs(1537) <= a;
    layer3_outputs(1538) <= a and not b;
    layer3_outputs(1539) <= not a;
    layer3_outputs(1540) <= not b or a;
    layer3_outputs(1541) <= b;
    layer3_outputs(1542) <= b and not a;
    layer3_outputs(1543) <= b;
    layer3_outputs(1544) <= a and not b;
    layer3_outputs(1545) <= not b;
    layer3_outputs(1546) <= not (a or b);
    layer3_outputs(1547) <= a;
    layer3_outputs(1548) <= not b or a;
    layer3_outputs(1549) <= not b or a;
    layer3_outputs(1550) <= not a;
    layer3_outputs(1551) <= not b;
    layer3_outputs(1552) <= '0';
    layer3_outputs(1553) <= not a;
    layer3_outputs(1554) <= not (a or b);
    layer3_outputs(1555) <= not (a or b);
    layer3_outputs(1556) <= not b or a;
    layer3_outputs(1557) <= a;
    layer3_outputs(1558) <= a and b;
    layer3_outputs(1559) <= b;
    layer3_outputs(1560) <= not b;
    layer3_outputs(1561) <= not a or b;
    layer3_outputs(1562) <= '1';
    layer3_outputs(1563) <= a or b;
    layer3_outputs(1564) <= not (a or b);
    layer3_outputs(1565) <= not a or b;
    layer3_outputs(1566) <= a or b;
    layer3_outputs(1567) <= '1';
    layer3_outputs(1568) <= not a;
    layer3_outputs(1569) <= not b or a;
    layer3_outputs(1570) <= not (a xor b);
    layer3_outputs(1571) <= not (a or b);
    layer3_outputs(1572) <= a and b;
    layer3_outputs(1573) <= b;
    layer3_outputs(1574) <= a xor b;
    layer3_outputs(1575) <= not (a or b);
    layer3_outputs(1576) <= a;
    layer3_outputs(1577) <= not (a or b);
    layer3_outputs(1578) <= b and not a;
    layer3_outputs(1579) <= a;
    layer3_outputs(1580) <= a;
    layer3_outputs(1581) <= not b;
    layer3_outputs(1582) <= not a or b;
    layer3_outputs(1583) <= '1';
    layer3_outputs(1584) <= a and b;
    layer3_outputs(1585) <= not b;
    layer3_outputs(1586) <= a;
    layer3_outputs(1587) <= not a or b;
    layer3_outputs(1588) <= not (a and b);
    layer3_outputs(1589) <= '1';
    layer3_outputs(1590) <= not (a and b);
    layer3_outputs(1591) <= not b;
    layer3_outputs(1592) <= a and not b;
    layer3_outputs(1593) <= not a;
    layer3_outputs(1594) <= not (a xor b);
    layer3_outputs(1595) <= a and b;
    layer3_outputs(1596) <= not (a xor b);
    layer3_outputs(1597) <= not a;
    layer3_outputs(1598) <= a or b;
    layer3_outputs(1599) <= a or b;
    layer3_outputs(1600) <= a;
    layer3_outputs(1601) <= a or b;
    layer3_outputs(1602) <= not a or b;
    layer3_outputs(1603) <= not (a and b);
    layer3_outputs(1604) <= not b or a;
    layer3_outputs(1605) <= a;
    layer3_outputs(1606) <= not (a and b);
    layer3_outputs(1607) <= not (a or b);
    layer3_outputs(1608) <= not (a or b);
    layer3_outputs(1609) <= not (a and b);
    layer3_outputs(1610) <= a;
    layer3_outputs(1611) <= a and not b;
    layer3_outputs(1612) <= not (a and b);
    layer3_outputs(1613) <= not (a and b);
    layer3_outputs(1614) <= '0';
    layer3_outputs(1615) <= a and b;
    layer3_outputs(1616) <= a and b;
    layer3_outputs(1617) <= a or b;
    layer3_outputs(1618) <= not a;
    layer3_outputs(1619) <= not a;
    layer3_outputs(1620) <= a and not b;
    layer3_outputs(1621) <= not (a or b);
    layer3_outputs(1622) <= b and not a;
    layer3_outputs(1623) <= not a;
    layer3_outputs(1624) <= not (a and b);
    layer3_outputs(1625) <= b;
    layer3_outputs(1626) <= not b;
    layer3_outputs(1627) <= not a or b;
    layer3_outputs(1628) <= b and not a;
    layer3_outputs(1629) <= b and not a;
    layer3_outputs(1630) <= a or b;
    layer3_outputs(1631) <= a and not b;
    layer3_outputs(1632) <= not a;
    layer3_outputs(1633) <= '1';
    layer3_outputs(1634) <= not (a xor b);
    layer3_outputs(1635) <= not a or b;
    layer3_outputs(1636) <= not (a xor b);
    layer3_outputs(1637) <= not a;
    layer3_outputs(1638) <= '1';
    layer3_outputs(1639) <= not (a xor b);
    layer3_outputs(1640) <= not (a xor b);
    layer3_outputs(1641) <= '1';
    layer3_outputs(1642) <= a;
    layer3_outputs(1643) <= a;
    layer3_outputs(1644) <= not a or b;
    layer3_outputs(1645) <= not b;
    layer3_outputs(1646) <= a and b;
    layer3_outputs(1647) <= '1';
    layer3_outputs(1648) <= not a;
    layer3_outputs(1649) <= not (a and b);
    layer3_outputs(1650) <= '1';
    layer3_outputs(1651) <= not b or a;
    layer3_outputs(1652) <= a and b;
    layer3_outputs(1653) <= '0';
    layer3_outputs(1654) <= not (a and b);
    layer3_outputs(1655) <= not (a or b);
    layer3_outputs(1656) <= b and not a;
    layer3_outputs(1657) <= a xor b;
    layer3_outputs(1658) <= not a;
    layer3_outputs(1659) <= a and not b;
    layer3_outputs(1660) <= not b;
    layer3_outputs(1661) <= b and not a;
    layer3_outputs(1662) <= '1';
    layer3_outputs(1663) <= a;
    layer3_outputs(1664) <= not a;
    layer3_outputs(1665) <= a;
    layer3_outputs(1666) <= '1';
    layer3_outputs(1667) <= not a;
    layer3_outputs(1668) <= a or b;
    layer3_outputs(1669) <= b and not a;
    layer3_outputs(1670) <= '1';
    layer3_outputs(1671) <= a xor b;
    layer3_outputs(1672) <= a and b;
    layer3_outputs(1673) <= not (a and b);
    layer3_outputs(1674) <= a;
    layer3_outputs(1675) <= a and b;
    layer3_outputs(1676) <= not b;
    layer3_outputs(1677) <= not b;
    layer3_outputs(1678) <= '0';
    layer3_outputs(1679) <= not (a and b);
    layer3_outputs(1680) <= not a;
    layer3_outputs(1681) <= not b;
    layer3_outputs(1682) <= not b;
    layer3_outputs(1683) <= a and not b;
    layer3_outputs(1684) <= a and b;
    layer3_outputs(1685) <= a or b;
    layer3_outputs(1686) <= a;
    layer3_outputs(1687) <= not b;
    layer3_outputs(1688) <= b;
    layer3_outputs(1689) <= not b;
    layer3_outputs(1690) <= b;
    layer3_outputs(1691) <= not (a or b);
    layer3_outputs(1692) <= a;
    layer3_outputs(1693) <= a or b;
    layer3_outputs(1694) <= a and not b;
    layer3_outputs(1695) <= not b or a;
    layer3_outputs(1696) <= a xor b;
    layer3_outputs(1697) <= not a or b;
    layer3_outputs(1698) <= not a;
    layer3_outputs(1699) <= not b;
    layer3_outputs(1700) <= a and b;
    layer3_outputs(1701) <= a;
    layer3_outputs(1702) <= '1';
    layer3_outputs(1703) <= not b;
    layer3_outputs(1704) <= not a;
    layer3_outputs(1705) <= not a;
    layer3_outputs(1706) <= not a;
    layer3_outputs(1707) <= not (a and b);
    layer3_outputs(1708) <= b and not a;
    layer3_outputs(1709) <= not a;
    layer3_outputs(1710) <= a xor b;
    layer3_outputs(1711) <= '1';
    layer3_outputs(1712) <= not b;
    layer3_outputs(1713) <= b;
    layer3_outputs(1714) <= a;
    layer3_outputs(1715) <= not (a and b);
    layer3_outputs(1716) <= not (a and b);
    layer3_outputs(1717) <= a and b;
    layer3_outputs(1718) <= a;
    layer3_outputs(1719) <= not (a and b);
    layer3_outputs(1720) <= a;
    layer3_outputs(1721) <= b;
    layer3_outputs(1722) <= a and b;
    layer3_outputs(1723) <= a xor b;
    layer3_outputs(1724) <= b and not a;
    layer3_outputs(1725) <= not b or a;
    layer3_outputs(1726) <= a and b;
    layer3_outputs(1727) <= a and b;
    layer3_outputs(1728) <= not (a or b);
    layer3_outputs(1729) <= '0';
    layer3_outputs(1730) <= not b;
    layer3_outputs(1731) <= a or b;
    layer3_outputs(1732) <= a;
    layer3_outputs(1733) <= not b;
    layer3_outputs(1734) <= not a or b;
    layer3_outputs(1735) <= b;
    layer3_outputs(1736) <= not (a and b);
    layer3_outputs(1737) <= a;
    layer3_outputs(1738) <= not a;
    layer3_outputs(1739) <= not a or b;
    layer3_outputs(1740) <= not (a or b);
    layer3_outputs(1741) <= not b;
    layer3_outputs(1742) <= a or b;
    layer3_outputs(1743) <= not (a and b);
    layer3_outputs(1744) <= '1';
    layer3_outputs(1745) <= '0';
    layer3_outputs(1746) <= b;
    layer3_outputs(1747) <= b;
    layer3_outputs(1748) <= not (a and b);
    layer3_outputs(1749) <= not b or a;
    layer3_outputs(1750) <= not b;
    layer3_outputs(1751) <= not (a or b);
    layer3_outputs(1752) <= a and b;
    layer3_outputs(1753) <= '1';
    layer3_outputs(1754) <= a;
    layer3_outputs(1755) <= not (a and b);
    layer3_outputs(1756) <= not (a or b);
    layer3_outputs(1757) <= not b;
    layer3_outputs(1758) <= not (a or b);
    layer3_outputs(1759) <= not b or a;
    layer3_outputs(1760) <= not (a and b);
    layer3_outputs(1761) <= a xor b;
    layer3_outputs(1762) <= not b;
    layer3_outputs(1763) <= b and not a;
    layer3_outputs(1764) <= b;
    layer3_outputs(1765) <= a and not b;
    layer3_outputs(1766) <= a;
    layer3_outputs(1767) <= not (a and b);
    layer3_outputs(1768) <= a and not b;
    layer3_outputs(1769) <= not a;
    layer3_outputs(1770) <= not b;
    layer3_outputs(1771) <= b and not a;
    layer3_outputs(1772) <= a;
    layer3_outputs(1773) <= a;
    layer3_outputs(1774) <= '1';
    layer3_outputs(1775) <= not b;
    layer3_outputs(1776) <= not a or b;
    layer3_outputs(1777) <= not (a and b);
    layer3_outputs(1778) <= a and b;
    layer3_outputs(1779) <= not a or b;
    layer3_outputs(1780) <= not b;
    layer3_outputs(1781) <= a;
    layer3_outputs(1782) <= a and b;
    layer3_outputs(1783) <= not b or a;
    layer3_outputs(1784) <= not a;
    layer3_outputs(1785) <= not a or b;
    layer3_outputs(1786) <= a and not b;
    layer3_outputs(1787) <= not a;
    layer3_outputs(1788) <= not a;
    layer3_outputs(1789) <= not (a xor b);
    layer3_outputs(1790) <= not a or b;
    layer3_outputs(1791) <= '1';
    layer3_outputs(1792) <= '0';
    layer3_outputs(1793) <= not a;
    layer3_outputs(1794) <= not a;
    layer3_outputs(1795) <= b and not a;
    layer3_outputs(1796) <= not a;
    layer3_outputs(1797) <= not (a and b);
    layer3_outputs(1798) <= b and not a;
    layer3_outputs(1799) <= not (a and b);
    layer3_outputs(1800) <= not b or a;
    layer3_outputs(1801) <= a;
    layer3_outputs(1802) <= not a;
    layer3_outputs(1803) <= not (a and b);
    layer3_outputs(1804) <= not (a or b);
    layer3_outputs(1805) <= not b or a;
    layer3_outputs(1806) <= not b or a;
    layer3_outputs(1807) <= not b;
    layer3_outputs(1808) <= a;
    layer3_outputs(1809) <= not (a or b);
    layer3_outputs(1810) <= not (a and b);
    layer3_outputs(1811) <= '0';
    layer3_outputs(1812) <= not (a and b);
    layer3_outputs(1813) <= a;
    layer3_outputs(1814) <= a and b;
    layer3_outputs(1815) <= a and not b;
    layer3_outputs(1816) <= a and b;
    layer3_outputs(1817) <= not a or b;
    layer3_outputs(1818) <= a;
    layer3_outputs(1819) <= not (a xor b);
    layer3_outputs(1820) <= not a or b;
    layer3_outputs(1821) <= not b;
    layer3_outputs(1822) <= a and b;
    layer3_outputs(1823) <= not a or b;
    layer3_outputs(1824) <= '1';
    layer3_outputs(1825) <= not b;
    layer3_outputs(1826) <= not b;
    layer3_outputs(1827) <= b;
    layer3_outputs(1828) <= b;
    layer3_outputs(1829) <= not (a or b);
    layer3_outputs(1830) <= not (a and b);
    layer3_outputs(1831) <= not a or b;
    layer3_outputs(1832) <= a xor b;
    layer3_outputs(1833) <= not (a xor b);
    layer3_outputs(1834) <= '0';
    layer3_outputs(1835) <= a and b;
    layer3_outputs(1836) <= a;
    layer3_outputs(1837) <= not b;
    layer3_outputs(1838) <= not a;
    layer3_outputs(1839) <= not b or a;
    layer3_outputs(1840) <= not a or b;
    layer3_outputs(1841) <= b;
    layer3_outputs(1842) <= a;
    layer3_outputs(1843) <= a;
    layer3_outputs(1844) <= a;
    layer3_outputs(1845) <= not a;
    layer3_outputs(1846) <= b and not a;
    layer3_outputs(1847) <= a or b;
    layer3_outputs(1848) <= b;
    layer3_outputs(1849) <= not (a xor b);
    layer3_outputs(1850) <= not (a or b);
    layer3_outputs(1851) <= b;
    layer3_outputs(1852) <= a;
    layer3_outputs(1853) <= not b;
    layer3_outputs(1854) <= b;
    layer3_outputs(1855) <= not b;
    layer3_outputs(1856) <= '0';
    layer3_outputs(1857) <= not (a and b);
    layer3_outputs(1858) <= not b or a;
    layer3_outputs(1859) <= b;
    layer3_outputs(1860) <= a or b;
    layer3_outputs(1861) <= not a;
    layer3_outputs(1862) <= a;
    layer3_outputs(1863) <= not a;
    layer3_outputs(1864) <= not b;
    layer3_outputs(1865) <= a or b;
    layer3_outputs(1866) <= a xor b;
    layer3_outputs(1867) <= b;
    layer3_outputs(1868) <= not (a xor b);
    layer3_outputs(1869) <= not (a xor b);
    layer3_outputs(1870) <= a and not b;
    layer3_outputs(1871) <= a;
    layer3_outputs(1872) <= not a or b;
    layer3_outputs(1873) <= a and b;
    layer3_outputs(1874) <= b;
    layer3_outputs(1875) <= not a;
    layer3_outputs(1876) <= b and not a;
    layer3_outputs(1877) <= a or b;
    layer3_outputs(1878) <= b;
    layer3_outputs(1879) <= not a;
    layer3_outputs(1880) <= not b;
    layer3_outputs(1881) <= not b;
    layer3_outputs(1882) <= b;
    layer3_outputs(1883) <= not b;
    layer3_outputs(1884) <= '1';
    layer3_outputs(1885) <= not (a and b);
    layer3_outputs(1886) <= a or b;
    layer3_outputs(1887) <= not (a xor b);
    layer3_outputs(1888) <= a or b;
    layer3_outputs(1889) <= b;
    layer3_outputs(1890) <= not a or b;
    layer3_outputs(1891) <= not (a xor b);
    layer3_outputs(1892) <= b;
    layer3_outputs(1893) <= not b or a;
    layer3_outputs(1894) <= not a;
    layer3_outputs(1895) <= b;
    layer3_outputs(1896) <= a and b;
    layer3_outputs(1897) <= not (a and b);
    layer3_outputs(1898) <= a xor b;
    layer3_outputs(1899) <= '0';
    layer3_outputs(1900) <= a;
    layer3_outputs(1901) <= a or b;
    layer3_outputs(1902) <= '1';
    layer3_outputs(1903) <= a;
    layer3_outputs(1904) <= not b or a;
    layer3_outputs(1905) <= b;
    layer3_outputs(1906) <= a;
    layer3_outputs(1907) <= a and not b;
    layer3_outputs(1908) <= not a or b;
    layer3_outputs(1909) <= not a or b;
    layer3_outputs(1910) <= '0';
    layer3_outputs(1911) <= '1';
    layer3_outputs(1912) <= not (a or b);
    layer3_outputs(1913) <= not b or a;
    layer3_outputs(1914) <= not (a or b);
    layer3_outputs(1915) <= a and not b;
    layer3_outputs(1916) <= not a or b;
    layer3_outputs(1917) <= '1';
    layer3_outputs(1918) <= not (a or b);
    layer3_outputs(1919) <= not a;
    layer3_outputs(1920) <= not (a or b);
    layer3_outputs(1921) <= not a or b;
    layer3_outputs(1922) <= a or b;
    layer3_outputs(1923) <= b and not a;
    layer3_outputs(1924) <= '1';
    layer3_outputs(1925) <= a or b;
    layer3_outputs(1926) <= not a or b;
    layer3_outputs(1927) <= a;
    layer3_outputs(1928) <= not a or b;
    layer3_outputs(1929) <= a;
    layer3_outputs(1930) <= a and not b;
    layer3_outputs(1931) <= not b;
    layer3_outputs(1932) <= not (a and b);
    layer3_outputs(1933) <= '1';
    layer3_outputs(1934) <= a xor b;
    layer3_outputs(1935) <= not b or a;
    layer3_outputs(1936) <= not (a or b);
    layer3_outputs(1937) <= a or b;
    layer3_outputs(1938) <= not a;
    layer3_outputs(1939) <= a;
    layer3_outputs(1940) <= a or b;
    layer3_outputs(1941) <= a;
    layer3_outputs(1942) <= a and not b;
    layer3_outputs(1943) <= b;
    layer3_outputs(1944) <= a xor b;
    layer3_outputs(1945) <= not (a or b);
    layer3_outputs(1946) <= not (a xor b);
    layer3_outputs(1947) <= b;
    layer3_outputs(1948) <= a and not b;
    layer3_outputs(1949) <= '0';
    layer3_outputs(1950) <= a;
    layer3_outputs(1951) <= a;
    layer3_outputs(1952) <= not (a and b);
    layer3_outputs(1953) <= not b;
    layer3_outputs(1954) <= b;
    layer3_outputs(1955) <= '1';
    layer3_outputs(1956) <= not a;
    layer3_outputs(1957) <= not (a and b);
    layer3_outputs(1958) <= not (a and b);
    layer3_outputs(1959) <= a xor b;
    layer3_outputs(1960) <= '1';
    layer3_outputs(1961) <= not a;
    layer3_outputs(1962) <= a or b;
    layer3_outputs(1963) <= b;
    layer3_outputs(1964) <= '0';
    layer3_outputs(1965) <= a;
    layer3_outputs(1966) <= not (a and b);
    layer3_outputs(1967) <= not (a and b);
    layer3_outputs(1968) <= a;
    layer3_outputs(1969) <= not a;
    layer3_outputs(1970) <= '0';
    layer3_outputs(1971) <= a and b;
    layer3_outputs(1972) <= b and not a;
    layer3_outputs(1973) <= '0';
    layer3_outputs(1974) <= not a or b;
    layer3_outputs(1975) <= b;
    layer3_outputs(1976) <= a or b;
    layer3_outputs(1977) <= b and not a;
    layer3_outputs(1978) <= a and b;
    layer3_outputs(1979) <= b;
    layer3_outputs(1980) <= '0';
    layer3_outputs(1981) <= not b;
    layer3_outputs(1982) <= not a;
    layer3_outputs(1983) <= b and not a;
    layer3_outputs(1984) <= not (a and b);
    layer3_outputs(1985) <= a or b;
    layer3_outputs(1986) <= not (a or b);
    layer3_outputs(1987) <= not a;
    layer3_outputs(1988) <= not b;
    layer3_outputs(1989) <= '1';
    layer3_outputs(1990) <= a and b;
    layer3_outputs(1991) <= not a or b;
    layer3_outputs(1992) <= a;
    layer3_outputs(1993) <= not b or a;
    layer3_outputs(1994) <= '1';
    layer3_outputs(1995) <= not (a xor b);
    layer3_outputs(1996) <= not b;
    layer3_outputs(1997) <= not a;
    layer3_outputs(1998) <= a or b;
    layer3_outputs(1999) <= not (a and b);
    layer3_outputs(2000) <= not a;
    layer3_outputs(2001) <= a;
    layer3_outputs(2002) <= a and not b;
    layer3_outputs(2003) <= not a or b;
    layer3_outputs(2004) <= not b;
    layer3_outputs(2005) <= a and b;
    layer3_outputs(2006) <= not (a and b);
    layer3_outputs(2007) <= a;
    layer3_outputs(2008) <= not a or b;
    layer3_outputs(2009) <= not a or b;
    layer3_outputs(2010) <= not (a xor b);
    layer3_outputs(2011) <= '0';
    layer3_outputs(2012) <= not (a and b);
    layer3_outputs(2013) <= '1';
    layer3_outputs(2014) <= not b;
    layer3_outputs(2015) <= b and not a;
    layer3_outputs(2016) <= a and b;
    layer3_outputs(2017) <= a;
    layer3_outputs(2018) <= a;
    layer3_outputs(2019) <= a and b;
    layer3_outputs(2020) <= a and not b;
    layer3_outputs(2021) <= a or b;
    layer3_outputs(2022) <= not a or b;
    layer3_outputs(2023) <= a xor b;
    layer3_outputs(2024) <= not b;
    layer3_outputs(2025) <= b;
    layer3_outputs(2026) <= a or b;
    layer3_outputs(2027) <= not (a or b);
    layer3_outputs(2028) <= not a or b;
    layer3_outputs(2029) <= not (a and b);
    layer3_outputs(2030) <= '1';
    layer3_outputs(2031) <= not a;
    layer3_outputs(2032) <= not a;
    layer3_outputs(2033) <= a and b;
    layer3_outputs(2034) <= not (a and b);
    layer3_outputs(2035) <= a or b;
    layer3_outputs(2036) <= b and not a;
    layer3_outputs(2037) <= not (a and b);
    layer3_outputs(2038) <= not b;
    layer3_outputs(2039) <= not b;
    layer3_outputs(2040) <= a and b;
    layer3_outputs(2041) <= not (a and b);
    layer3_outputs(2042) <= not (a and b);
    layer3_outputs(2043) <= a or b;
    layer3_outputs(2044) <= not a;
    layer3_outputs(2045) <= a;
    layer3_outputs(2046) <= '1';
    layer3_outputs(2047) <= '0';
    layer3_outputs(2048) <= a and not b;
    layer3_outputs(2049) <= not b;
    layer3_outputs(2050) <= a and b;
    layer3_outputs(2051) <= not b;
    layer3_outputs(2052) <= not b;
    layer3_outputs(2053) <= not (a and b);
    layer3_outputs(2054) <= b;
    layer3_outputs(2055) <= a xor b;
    layer3_outputs(2056) <= a or b;
    layer3_outputs(2057) <= a and not b;
    layer3_outputs(2058) <= not (a and b);
    layer3_outputs(2059) <= not a or b;
    layer3_outputs(2060) <= not a;
    layer3_outputs(2061) <= not a or b;
    layer3_outputs(2062) <= a xor b;
    layer3_outputs(2063) <= '1';
    layer3_outputs(2064) <= b;
    layer3_outputs(2065) <= b;
    layer3_outputs(2066) <= not b;
    layer3_outputs(2067) <= a and not b;
    layer3_outputs(2068) <= a;
    layer3_outputs(2069) <= a;
    layer3_outputs(2070) <= b and not a;
    layer3_outputs(2071) <= b;
    layer3_outputs(2072) <= not a;
    layer3_outputs(2073) <= not (a and b);
    layer3_outputs(2074) <= a xor b;
    layer3_outputs(2075) <= not b or a;
    layer3_outputs(2076) <= '1';
    layer3_outputs(2077) <= not a or b;
    layer3_outputs(2078) <= a or b;
    layer3_outputs(2079) <= not b;
    layer3_outputs(2080) <= b and not a;
    layer3_outputs(2081) <= a xor b;
    layer3_outputs(2082) <= '0';
    layer3_outputs(2083) <= a and not b;
    layer3_outputs(2084) <= not (a or b);
    layer3_outputs(2085) <= not (a and b);
    layer3_outputs(2086) <= b and not a;
    layer3_outputs(2087) <= a or b;
    layer3_outputs(2088) <= b;
    layer3_outputs(2089) <= not b;
    layer3_outputs(2090) <= '0';
    layer3_outputs(2091) <= b and not a;
    layer3_outputs(2092) <= a or b;
    layer3_outputs(2093) <= '0';
    layer3_outputs(2094) <= not b;
    layer3_outputs(2095) <= a;
    layer3_outputs(2096) <= not b or a;
    layer3_outputs(2097) <= '0';
    layer3_outputs(2098) <= not (a xor b);
    layer3_outputs(2099) <= not a or b;
    layer3_outputs(2100) <= not b;
    layer3_outputs(2101) <= a and not b;
    layer3_outputs(2102) <= not a or b;
    layer3_outputs(2103) <= not (a or b);
    layer3_outputs(2104) <= not b;
    layer3_outputs(2105) <= b and not a;
    layer3_outputs(2106) <= not (a or b);
    layer3_outputs(2107) <= a;
    layer3_outputs(2108) <= not (a or b);
    layer3_outputs(2109) <= a and not b;
    layer3_outputs(2110) <= a and b;
    layer3_outputs(2111) <= not (a and b);
    layer3_outputs(2112) <= not (a or b);
    layer3_outputs(2113) <= b;
    layer3_outputs(2114) <= not a;
    layer3_outputs(2115) <= not b or a;
    layer3_outputs(2116) <= not a;
    layer3_outputs(2117) <= b and not a;
    layer3_outputs(2118) <= not a;
    layer3_outputs(2119) <= not a;
    layer3_outputs(2120) <= not a or b;
    layer3_outputs(2121) <= a and not b;
    layer3_outputs(2122) <= '1';
    layer3_outputs(2123) <= b;
    layer3_outputs(2124) <= b;
    layer3_outputs(2125) <= not b;
    layer3_outputs(2126) <= not b;
    layer3_outputs(2127) <= not a or b;
    layer3_outputs(2128) <= not (a and b);
    layer3_outputs(2129) <= a;
    layer3_outputs(2130) <= a or b;
    layer3_outputs(2131) <= not b or a;
    layer3_outputs(2132) <= not b;
    layer3_outputs(2133) <= not a or b;
    layer3_outputs(2134) <= '1';
    layer3_outputs(2135) <= not (a or b);
    layer3_outputs(2136) <= b;
    layer3_outputs(2137) <= b and not a;
    layer3_outputs(2138) <= a xor b;
    layer3_outputs(2139) <= a and b;
    layer3_outputs(2140) <= b;
    layer3_outputs(2141) <= not (a and b);
    layer3_outputs(2142) <= not (a or b);
    layer3_outputs(2143) <= a;
    layer3_outputs(2144) <= '0';
    layer3_outputs(2145) <= not a;
    layer3_outputs(2146) <= b;
    layer3_outputs(2147) <= not a;
    layer3_outputs(2148) <= b;
    layer3_outputs(2149) <= not b;
    layer3_outputs(2150) <= not (a or b);
    layer3_outputs(2151) <= a;
    layer3_outputs(2152) <= not (a or b);
    layer3_outputs(2153) <= not (a or b);
    layer3_outputs(2154) <= not a;
    layer3_outputs(2155) <= '1';
    layer3_outputs(2156) <= not b or a;
    layer3_outputs(2157) <= not (a and b);
    layer3_outputs(2158) <= not (a and b);
    layer3_outputs(2159) <= b;
    layer3_outputs(2160) <= a;
    layer3_outputs(2161) <= not b or a;
    layer3_outputs(2162) <= a and not b;
    layer3_outputs(2163) <= not (a or b);
    layer3_outputs(2164) <= a or b;
    layer3_outputs(2165) <= not (a or b);
    layer3_outputs(2166) <= not a;
    layer3_outputs(2167) <= a and b;
    layer3_outputs(2168) <= not b or a;
    layer3_outputs(2169) <= not a or b;
    layer3_outputs(2170) <= b;
    layer3_outputs(2171) <= not b;
    layer3_outputs(2172) <= a xor b;
    layer3_outputs(2173) <= not b or a;
    layer3_outputs(2174) <= a or b;
    layer3_outputs(2175) <= not b;
    layer3_outputs(2176) <= not (a and b);
    layer3_outputs(2177) <= b;
    layer3_outputs(2178) <= a and not b;
    layer3_outputs(2179) <= a and b;
    layer3_outputs(2180) <= b;
    layer3_outputs(2181) <= a and not b;
    layer3_outputs(2182) <= not (a and b);
    layer3_outputs(2183) <= not a;
    layer3_outputs(2184) <= not (a xor b);
    layer3_outputs(2185) <= '0';
    layer3_outputs(2186) <= a and not b;
    layer3_outputs(2187) <= a and not b;
    layer3_outputs(2188) <= not a or b;
    layer3_outputs(2189) <= b and not a;
    layer3_outputs(2190) <= not (a and b);
    layer3_outputs(2191) <= a and b;
    layer3_outputs(2192) <= not b or a;
    layer3_outputs(2193) <= b;
    layer3_outputs(2194) <= a and not b;
    layer3_outputs(2195) <= not b or a;
    layer3_outputs(2196) <= '1';
    layer3_outputs(2197) <= a xor b;
    layer3_outputs(2198) <= a or b;
    layer3_outputs(2199) <= a;
    layer3_outputs(2200) <= not a;
    layer3_outputs(2201) <= not a;
    layer3_outputs(2202) <= not (a or b);
    layer3_outputs(2203) <= a;
    layer3_outputs(2204) <= not (a and b);
    layer3_outputs(2205) <= a and b;
    layer3_outputs(2206) <= not b or a;
    layer3_outputs(2207) <= '0';
    layer3_outputs(2208) <= not a or b;
    layer3_outputs(2209) <= '1';
    layer3_outputs(2210) <= not (a and b);
    layer3_outputs(2211) <= '1';
    layer3_outputs(2212) <= a or b;
    layer3_outputs(2213) <= not a;
    layer3_outputs(2214) <= not a or b;
    layer3_outputs(2215) <= a;
    layer3_outputs(2216) <= not a or b;
    layer3_outputs(2217) <= a xor b;
    layer3_outputs(2218) <= a and b;
    layer3_outputs(2219) <= not (a xor b);
    layer3_outputs(2220) <= '0';
    layer3_outputs(2221) <= a;
    layer3_outputs(2222) <= not a;
    layer3_outputs(2223) <= b;
    layer3_outputs(2224) <= not a;
    layer3_outputs(2225) <= b;
    layer3_outputs(2226) <= a;
    layer3_outputs(2227) <= not b;
    layer3_outputs(2228) <= '1';
    layer3_outputs(2229) <= not (a or b);
    layer3_outputs(2230) <= not (a or b);
    layer3_outputs(2231) <= not b;
    layer3_outputs(2232) <= b;
    layer3_outputs(2233) <= a;
    layer3_outputs(2234) <= a xor b;
    layer3_outputs(2235) <= a or b;
    layer3_outputs(2236) <= not a;
    layer3_outputs(2237) <= a;
    layer3_outputs(2238) <= not a;
    layer3_outputs(2239) <= b;
    layer3_outputs(2240) <= not a;
    layer3_outputs(2241) <= b;
    layer3_outputs(2242) <= a;
    layer3_outputs(2243) <= a;
    layer3_outputs(2244) <= a;
    layer3_outputs(2245) <= b;
    layer3_outputs(2246) <= not b or a;
    layer3_outputs(2247) <= not b;
    layer3_outputs(2248) <= not b;
    layer3_outputs(2249) <= not (a xor b);
    layer3_outputs(2250) <= not (a and b);
    layer3_outputs(2251) <= not (a or b);
    layer3_outputs(2252) <= not a;
    layer3_outputs(2253) <= a;
    layer3_outputs(2254) <= not a or b;
    layer3_outputs(2255) <= a and not b;
    layer3_outputs(2256) <= not a;
    layer3_outputs(2257) <= not (a xor b);
    layer3_outputs(2258) <= not a or b;
    layer3_outputs(2259) <= not a or b;
    layer3_outputs(2260) <= not b or a;
    layer3_outputs(2261) <= '1';
    layer3_outputs(2262) <= not a or b;
    layer3_outputs(2263) <= b and not a;
    layer3_outputs(2264) <= not b;
    layer3_outputs(2265) <= b;
    layer3_outputs(2266) <= not a;
    layer3_outputs(2267) <= not a;
    layer3_outputs(2268) <= not (a and b);
    layer3_outputs(2269) <= not (a or b);
    layer3_outputs(2270) <= not b or a;
    layer3_outputs(2271) <= a and not b;
    layer3_outputs(2272) <= a xor b;
    layer3_outputs(2273) <= not b or a;
    layer3_outputs(2274) <= not a or b;
    layer3_outputs(2275) <= not (a or b);
    layer3_outputs(2276) <= not b;
    layer3_outputs(2277) <= not b;
    layer3_outputs(2278) <= not b;
    layer3_outputs(2279) <= '1';
    layer3_outputs(2280) <= not (a or b);
    layer3_outputs(2281) <= b and not a;
    layer3_outputs(2282) <= not (a xor b);
    layer3_outputs(2283) <= not (a and b);
    layer3_outputs(2284) <= a;
    layer3_outputs(2285) <= b;
    layer3_outputs(2286) <= not a;
    layer3_outputs(2287) <= '0';
    layer3_outputs(2288) <= '1';
    layer3_outputs(2289) <= not (a and b);
    layer3_outputs(2290) <= '1';
    layer3_outputs(2291) <= '1';
    layer3_outputs(2292) <= not b;
    layer3_outputs(2293) <= a or b;
    layer3_outputs(2294) <= a or b;
    layer3_outputs(2295) <= b and not a;
    layer3_outputs(2296) <= not b;
    layer3_outputs(2297) <= b and not a;
    layer3_outputs(2298) <= a and b;
    layer3_outputs(2299) <= not (a xor b);
    layer3_outputs(2300) <= b;
    layer3_outputs(2301) <= not (a or b);
    layer3_outputs(2302) <= not b or a;
    layer3_outputs(2303) <= not (a and b);
    layer3_outputs(2304) <= a and not b;
    layer3_outputs(2305) <= b;
    layer3_outputs(2306) <= a or b;
    layer3_outputs(2307) <= b;
    layer3_outputs(2308) <= not a or b;
    layer3_outputs(2309) <= not (a or b);
    layer3_outputs(2310) <= a;
    layer3_outputs(2311) <= not b;
    layer3_outputs(2312) <= not a;
    layer3_outputs(2313) <= a and b;
    layer3_outputs(2314) <= not b;
    layer3_outputs(2315) <= a xor b;
    layer3_outputs(2316) <= a and b;
    layer3_outputs(2317) <= '0';
    layer3_outputs(2318) <= not b;
    layer3_outputs(2319) <= not a;
    layer3_outputs(2320) <= not a or b;
    layer3_outputs(2321) <= b;
    layer3_outputs(2322) <= a;
    layer3_outputs(2323) <= not a;
    layer3_outputs(2324) <= a;
    layer3_outputs(2325) <= not a;
    layer3_outputs(2326) <= b and not a;
    layer3_outputs(2327) <= a xor b;
    layer3_outputs(2328) <= not (a xor b);
    layer3_outputs(2329) <= a xor b;
    layer3_outputs(2330) <= a;
    layer3_outputs(2331) <= a;
    layer3_outputs(2332) <= '0';
    layer3_outputs(2333) <= not b;
    layer3_outputs(2334) <= not (a or b);
    layer3_outputs(2335) <= not b or a;
    layer3_outputs(2336) <= not a or b;
    layer3_outputs(2337) <= not a or b;
    layer3_outputs(2338) <= a;
    layer3_outputs(2339) <= not (a and b);
    layer3_outputs(2340) <= not b;
    layer3_outputs(2341) <= not b or a;
    layer3_outputs(2342) <= not a or b;
    layer3_outputs(2343) <= a and b;
    layer3_outputs(2344) <= a and not b;
    layer3_outputs(2345) <= not (a xor b);
    layer3_outputs(2346) <= a and b;
    layer3_outputs(2347) <= not a;
    layer3_outputs(2348) <= not a;
    layer3_outputs(2349) <= not (a and b);
    layer3_outputs(2350) <= a and not b;
    layer3_outputs(2351) <= b and not a;
    layer3_outputs(2352) <= not (a xor b);
    layer3_outputs(2353) <= not a;
    layer3_outputs(2354) <= not a;
    layer3_outputs(2355) <= a or b;
    layer3_outputs(2356) <= not b or a;
    layer3_outputs(2357) <= not (a xor b);
    layer3_outputs(2358) <= not (a and b);
    layer3_outputs(2359) <= '0';
    layer3_outputs(2360) <= not b;
    layer3_outputs(2361) <= a;
    layer3_outputs(2362) <= not (a xor b);
    layer3_outputs(2363) <= not a or b;
    layer3_outputs(2364) <= not a;
    layer3_outputs(2365) <= not (a and b);
    layer3_outputs(2366) <= b and not a;
    layer3_outputs(2367) <= not (a and b);
    layer3_outputs(2368) <= a and not b;
    layer3_outputs(2369) <= not b;
    layer3_outputs(2370) <= not b;
    layer3_outputs(2371) <= not a;
    layer3_outputs(2372) <= a or b;
    layer3_outputs(2373) <= b;
    layer3_outputs(2374) <= a and b;
    layer3_outputs(2375) <= not a or b;
    layer3_outputs(2376) <= not b or a;
    layer3_outputs(2377) <= a;
    layer3_outputs(2378) <= a;
    layer3_outputs(2379) <= a and not b;
    layer3_outputs(2380) <= '0';
    layer3_outputs(2381) <= a;
    layer3_outputs(2382) <= not b or a;
    layer3_outputs(2383) <= a and not b;
    layer3_outputs(2384) <= b and not a;
    layer3_outputs(2385) <= a and b;
    layer3_outputs(2386) <= not a;
    layer3_outputs(2387) <= '0';
    layer3_outputs(2388) <= a;
    layer3_outputs(2389) <= not b;
    layer3_outputs(2390) <= not b;
    layer3_outputs(2391) <= b and not a;
    layer3_outputs(2392) <= a and b;
    layer3_outputs(2393) <= not a;
    layer3_outputs(2394) <= a and b;
    layer3_outputs(2395) <= not (a xor b);
    layer3_outputs(2396) <= not (a or b);
    layer3_outputs(2397) <= not b or a;
    layer3_outputs(2398) <= a xor b;
    layer3_outputs(2399) <= a or b;
    layer3_outputs(2400) <= not b;
    layer3_outputs(2401) <= a and b;
    layer3_outputs(2402) <= a;
    layer3_outputs(2403) <= b;
    layer3_outputs(2404) <= not b;
    layer3_outputs(2405) <= not b;
    layer3_outputs(2406) <= a and b;
    layer3_outputs(2407) <= b and not a;
    layer3_outputs(2408) <= b and not a;
    layer3_outputs(2409) <= '1';
    layer3_outputs(2410) <= not (a and b);
    layer3_outputs(2411) <= '0';
    layer3_outputs(2412) <= a and not b;
    layer3_outputs(2413) <= not b or a;
    layer3_outputs(2414) <= not (a and b);
    layer3_outputs(2415) <= a or b;
    layer3_outputs(2416) <= a or b;
    layer3_outputs(2417) <= not a or b;
    layer3_outputs(2418) <= b;
    layer3_outputs(2419) <= not a;
    layer3_outputs(2420) <= not a or b;
    layer3_outputs(2421) <= not (a or b);
    layer3_outputs(2422) <= a or b;
    layer3_outputs(2423) <= not a;
    layer3_outputs(2424) <= not a or b;
    layer3_outputs(2425) <= b;
    layer3_outputs(2426) <= b;
    layer3_outputs(2427) <= not (a or b);
    layer3_outputs(2428) <= a and b;
    layer3_outputs(2429) <= not a;
    layer3_outputs(2430) <= not a;
    layer3_outputs(2431) <= not a;
    layer3_outputs(2432) <= a and not b;
    layer3_outputs(2433) <= not (a or b);
    layer3_outputs(2434) <= a;
    layer3_outputs(2435) <= a and b;
    layer3_outputs(2436) <= a and not b;
    layer3_outputs(2437) <= a or b;
    layer3_outputs(2438) <= a and b;
    layer3_outputs(2439) <= a and b;
    layer3_outputs(2440) <= a or b;
    layer3_outputs(2441) <= b;
    layer3_outputs(2442) <= a;
    layer3_outputs(2443) <= not b;
    layer3_outputs(2444) <= a;
    layer3_outputs(2445) <= a and not b;
    layer3_outputs(2446) <= a and b;
    layer3_outputs(2447) <= b;
    layer3_outputs(2448) <= b;
    layer3_outputs(2449) <= not a or b;
    layer3_outputs(2450) <= a and b;
    layer3_outputs(2451) <= b;
    layer3_outputs(2452) <= '0';
    layer3_outputs(2453) <= not (a xor b);
    layer3_outputs(2454) <= not (a or b);
    layer3_outputs(2455) <= a;
    layer3_outputs(2456) <= not a;
    layer3_outputs(2457) <= a;
    layer3_outputs(2458) <= not (a or b);
    layer3_outputs(2459) <= not (a and b);
    layer3_outputs(2460) <= a xor b;
    layer3_outputs(2461) <= a or b;
    layer3_outputs(2462) <= not b;
    layer3_outputs(2463) <= '0';
    layer3_outputs(2464) <= b;
    layer3_outputs(2465) <= a xor b;
    layer3_outputs(2466) <= not (a and b);
    layer3_outputs(2467) <= not b or a;
    layer3_outputs(2468) <= not (a and b);
    layer3_outputs(2469) <= b and not a;
    layer3_outputs(2470) <= a and b;
    layer3_outputs(2471) <= a;
    layer3_outputs(2472) <= not a or b;
    layer3_outputs(2473) <= b;
    layer3_outputs(2474) <= not (a xor b);
    layer3_outputs(2475) <= not (a and b);
    layer3_outputs(2476) <= not a or b;
    layer3_outputs(2477) <= a and b;
    layer3_outputs(2478) <= a or b;
    layer3_outputs(2479) <= a or b;
    layer3_outputs(2480) <= not a or b;
    layer3_outputs(2481) <= b;
    layer3_outputs(2482) <= '0';
    layer3_outputs(2483) <= b;
    layer3_outputs(2484) <= a and not b;
    layer3_outputs(2485) <= b;
    layer3_outputs(2486) <= b;
    layer3_outputs(2487) <= not (a or b);
    layer3_outputs(2488) <= not b;
    layer3_outputs(2489) <= a xor b;
    layer3_outputs(2490) <= not (a and b);
    layer3_outputs(2491) <= a or b;
    layer3_outputs(2492) <= not a or b;
    layer3_outputs(2493) <= not a or b;
    layer3_outputs(2494) <= not (a xor b);
    layer3_outputs(2495) <= not b or a;
    layer3_outputs(2496) <= '0';
    layer3_outputs(2497) <= a or b;
    layer3_outputs(2498) <= b;
    layer3_outputs(2499) <= b and not a;
    layer3_outputs(2500) <= b;
    layer3_outputs(2501) <= not b or a;
    layer3_outputs(2502) <= a and b;
    layer3_outputs(2503) <= a;
    layer3_outputs(2504) <= not b;
    layer3_outputs(2505) <= a;
    layer3_outputs(2506) <= not b;
    layer3_outputs(2507) <= not b;
    layer3_outputs(2508) <= not a;
    layer3_outputs(2509) <= b;
    layer3_outputs(2510) <= a and b;
    layer3_outputs(2511) <= not b or a;
    layer3_outputs(2512) <= not a;
    layer3_outputs(2513) <= b;
    layer3_outputs(2514) <= not b;
    layer3_outputs(2515) <= b;
    layer3_outputs(2516) <= a;
    layer3_outputs(2517) <= b;
    layer3_outputs(2518) <= not b or a;
    layer3_outputs(2519) <= not (a or b);
    layer3_outputs(2520) <= b;
    layer3_outputs(2521) <= a and not b;
    layer3_outputs(2522) <= not a;
    layer3_outputs(2523) <= not (a or b);
    layer3_outputs(2524) <= b and not a;
    layer3_outputs(2525) <= not (a or b);
    layer3_outputs(2526) <= not b or a;
    layer3_outputs(2527) <= a xor b;
    layer3_outputs(2528) <= not a;
    layer3_outputs(2529) <= a and not b;
    layer3_outputs(2530) <= b;
    layer3_outputs(2531) <= not a;
    layer3_outputs(2532) <= not (a and b);
    layer3_outputs(2533) <= a or b;
    layer3_outputs(2534) <= not a or b;
    layer3_outputs(2535) <= b and not a;
    layer3_outputs(2536) <= '0';
    layer3_outputs(2537) <= not a or b;
    layer3_outputs(2538) <= a;
    layer3_outputs(2539) <= not b;
    layer3_outputs(2540) <= not b;
    layer3_outputs(2541) <= b;
    layer3_outputs(2542) <= not a or b;
    layer3_outputs(2543) <= not (a and b);
    layer3_outputs(2544) <= a or b;
    layer3_outputs(2545) <= a and b;
    layer3_outputs(2546) <= a or b;
    layer3_outputs(2547) <= b;
    layer3_outputs(2548) <= b;
    layer3_outputs(2549) <= '0';
    layer3_outputs(2550) <= a;
    layer3_outputs(2551) <= not a or b;
    layer3_outputs(2552) <= a and b;
    layer3_outputs(2553) <= '0';
    layer3_outputs(2554) <= not (a and b);
    layer3_outputs(2555) <= not (a xor b);
    layer3_outputs(2556) <= b and not a;
    layer3_outputs(2557) <= not (a and b);
    layer3_outputs(2558) <= not b;
    layer3_outputs(2559) <= not b;
    layer3_outputs(2560) <= '0';
    layer3_outputs(2561) <= a or b;
    layer3_outputs(2562) <= a or b;
    layer3_outputs(2563) <= not a;
    layer3_outputs(2564) <= not (a xor b);
    layer3_outputs(2565) <= not a;
    layer3_outputs(2566) <= b;
    layer3_outputs(2567) <= '0';
    layer3_outputs(2568) <= a;
    layer3_outputs(2569) <= a and b;
    layer3_outputs(2570) <= b;
    layer3_outputs(2571) <= a and not b;
    layer3_outputs(2572) <= a and b;
    layer3_outputs(2573) <= b and not a;
    layer3_outputs(2574) <= a or b;
    layer3_outputs(2575) <= a;
    layer3_outputs(2576) <= a;
    layer3_outputs(2577) <= a and not b;
    layer3_outputs(2578) <= a or b;
    layer3_outputs(2579) <= b;
    layer3_outputs(2580) <= b;
    layer3_outputs(2581) <= a or b;
    layer3_outputs(2582) <= not b or a;
    layer3_outputs(2583) <= not (a or b);
    layer3_outputs(2584) <= not (a and b);
    layer3_outputs(2585) <= b;
    layer3_outputs(2586) <= not a;
    layer3_outputs(2587) <= not a;
    layer3_outputs(2588) <= not b;
    layer3_outputs(2589) <= not (a xor b);
    layer3_outputs(2590) <= a and b;
    layer3_outputs(2591) <= not b;
    layer3_outputs(2592) <= not (a and b);
    layer3_outputs(2593) <= '1';
    layer3_outputs(2594) <= not a;
    layer3_outputs(2595) <= not a;
    layer3_outputs(2596) <= not b;
    layer3_outputs(2597) <= b;
    layer3_outputs(2598) <= not b or a;
    layer3_outputs(2599) <= a and not b;
    layer3_outputs(2600) <= not (a or b);
    layer3_outputs(2601) <= not a;
    layer3_outputs(2602) <= not a;
    layer3_outputs(2603) <= a or b;
    layer3_outputs(2604) <= not (a or b);
    layer3_outputs(2605) <= a or b;
    layer3_outputs(2606) <= not b or a;
    layer3_outputs(2607) <= a or b;
    layer3_outputs(2608) <= not (a or b);
    layer3_outputs(2609) <= not (a and b);
    layer3_outputs(2610) <= not (a or b);
    layer3_outputs(2611) <= '1';
    layer3_outputs(2612) <= '0';
    layer3_outputs(2613) <= a xor b;
    layer3_outputs(2614) <= not (a and b);
    layer3_outputs(2615) <= not (a and b);
    layer3_outputs(2616) <= not a;
    layer3_outputs(2617) <= a and not b;
    layer3_outputs(2618) <= not a;
    layer3_outputs(2619) <= b;
    layer3_outputs(2620) <= b;
    layer3_outputs(2621) <= a and b;
    layer3_outputs(2622) <= not (a or b);
    layer3_outputs(2623) <= a;
    layer3_outputs(2624) <= a and b;
    layer3_outputs(2625) <= a or b;
    layer3_outputs(2626) <= not (a or b);
    layer3_outputs(2627) <= not (a or b);
    layer3_outputs(2628) <= not b or a;
    layer3_outputs(2629) <= a;
    layer3_outputs(2630) <= not a or b;
    layer3_outputs(2631) <= not (a or b);
    layer3_outputs(2632) <= not b or a;
    layer3_outputs(2633) <= not b or a;
    layer3_outputs(2634) <= not (a xor b);
    layer3_outputs(2635) <= not a or b;
    layer3_outputs(2636) <= not b;
    layer3_outputs(2637) <= a and b;
    layer3_outputs(2638) <= not b or a;
    layer3_outputs(2639) <= not a;
    layer3_outputs(2640) <= not (a or b);
    layer3_outputs(2641) <= b;
    layer3_outputs(2642) <= not (a or b);
    layer3_outputs(2643) <= a and b;
    layer3_outputs(2644) <= a and b;
    layer3_outputs(2645) <= a and b;
    layer3_outputs(2646) <= '0';
    layer3_outputs(2647) <= a and b;
    layer3_outputs(2648) <= a;
    layer3_outputs(2649) <= '0';
    layer3_outputs(2650) <= b and not a;
    layer3_outputs(2651) <= not a;
    layer3_outputs(2652) <= not b or a;
    layer3_outputs(2653) <= '0';
    layer3_outputs(2654) <= not b or a;
    layer3_outputs(2655) <= a;
    layer3_outputs(2656) <= not b;
    layer3_outputs(2657) <= not a;
    layer3_outputs(2658) <= a or b;
    layer3_outputs(2659) <= not b;
    layer3_outputs(2660) <= not b or a;
    layer3_outputs(2661) <= a xor b;
    layer3_outputs(2662) <= '0';
    layer3_outputs(2663) <= not (a and b);
    layer3_outputs(2664) <= not a;
    layer3_outputs(2665) <= a xor b;
    layer3_outputs(2666) <= a or b;
    layer3_outputs(2667) <= not b;
    layer3_outputs(2668) <= not b or a;
    layer3_outputs(2669) <= a or b;
    layer3_outputs(2670) <= a and not b;
    layer3_outputs(2671) <= not (a or b);
    layer3_outputs(2672) <= not (a or b);
    layer3_outputs(2673) <= a and not b;
    layer3_outputs(2674) <= not b or a;
    layer3_outputs(2675) <= not (a xor b);
    layer3_outputs(2676) <= a or b;
    layer3_outputs(2677) <= a and b;
    layer3_outputs(2678) <= b;
    layer3_outputs(2679) <= a or b;
    layer3_outputs(2680) <= a;
    layer3_outputs(2681) <= a or b;
    layer3_outputs(2682) <= not (a and b);
    layer3_outputs(2683) <= not b;
    layer3_outputs(2684) <= a;
    layer3_outputs(2685) <= b;
    layer3_outputs(2686) <= not (a or b);
    layer3_outputs(2687) <= a;
    layer3_outputs(2688) <= not (a or b);
    layer3_outputs(2689) <= not b or a;
    layer3_outputs(2690) <= not a or b;
    layer3_outputs(2691) <= not b or a;
    layer3_outputs(2692) <= b and not a;
    layer3_outputs(2693) <= not (a or b);
    layer3_outputs(2694) <= a xor b;
    layer3_outputs(2695) <= not b;
    layer3_outputs(2696) <= b and not a;
    layer3_outputs(2697) <= not b;
    layer3_outputs(2698) <= a and not b;
    layer3_outputs(2699) <= not (a and b);
    layer3_outputs(2700) <= not a;
    layer3_outputs(2701) <= not b or a;
    layer3_outputs(2702) <= a and b;
    layer3_outputs(2703) <= a and b;
    layer3_outputs(2704) <= not b or a;
    layer3_outputs(2705) <= not (a or b);
    layer3_outputs(2706) <= not b;
    layer3_outputs(2707) <= not b;
    layer3_outputs(2708) <= a and b;
    layer3_outputs(2709) <= not (a and b);
    layer3_outputs(2710) <= not b or a;
    layer3_outputs(2711) <= not (a and b);
    layer3_outputs(2712) <= a or b;
    layer3_outputs(2713) <= a;
    layer3_outputs(2714) <= not a;
    layer3_outputs(2715) <= not a or b;
    layer3_outputs(2716) <= not (a and b);
    layer3_outputs(2717) <= a xor b;
    layer3_outputs(2718) <= not a;
    layer3_outputs(2719) <= not (a xor b);
    layer3_outputs(2720) <= a or b;
    layer3_outputs(2721) <= a and not b;
    layer3_outputs(2722) <= a;
    layer3_outputs(2723) <= a and b;
    layer3_outputs(2724) <= not b;
    layer3_outputs(2725) <= a or b;
    layer3_outputs(2726) <= not a;
    layer3_outputs(2727) <= not a or b;
    layer3_outputs(2728) <= b and not a;
    layer3_outputs(2729) <= not a or b;
    layer3_outputs(2730) <= not a or b;
    layer3_outputs(2731) <= a;
    layer3_outputs(2732) <= a and not b;
    layer3_outputs(2733) <= a and b;
    layer3_outputs(2734) <= a xor b;
    layer3_outputs(2735) <= '0';
    layer3_outputs(2736) <= not (a xor b);
    layer3_outputs(2737) <= b;
    layer3_outputs(2738) <= not b;
    layer3_outputs(2739) <= not b;
    layer3_outputs(2740) <= not a or b;
    layer3_outputs(2741) <= not a or b;
    layer3_outputs(2742) <= not a;
    layer3_outputs(2743) <= b;
    layer3_outputs(2744) <= b;
    layer3_outputs(2745) <= a or b;
    layer3_outputs(2746) <= a and not b;
    layer3_outputs(2747) <= a or b;
    layer3_outputs(2748) <= '1';
    layer3_outputs(2749) <= not b;
    layer3_outputs(2750) <= not b or a;
    layer3_outputs(2751) <= not (a xor b);
    layer3_outputs(2752) <= a xor b;
    layer3_outputs(2753) <= a;
    layer3_outputs(2754) <= b and not a;
    layer3_outputs(2755) <= not (a and b);
    layer3_outputs(2756) <= '0';
    layer3_outputs(2757) <= not b or a;
    layer3_outputs(2758) <= not (a and b);
    layer3_outputs(2759) <= a and b;
    layer3_outputs(2760) <= b and not a;
    layer3_outputs(2761) <= not b or a;
    layer3_outputs(2762) <= b;
    layer3_outputs(2763) <= a and not b;
    layer3_outputs(2764) <= a xor b;
    layer3_outputs(2765) <= not a;
    layer3_outputs(2766) <= a or b;
    layer3_outputs(2767) <= not b;
    layer3_outputs(2768) <= b;
    layer3_outputs(2769) <= '0';
    layer3_outputs(2770) <= '0';
    layer3_outputs(2771) <= not (a and b);
    layer3_outputs(2772) <= a and b;
    layer3_outputs(2773) <= not b;
    layer3_outputs(2774) <= a;
    layer3_outputs(2775) <= not (a and b);
    layer3_outputs(2776) <= a;
    layer3_outputs(2777) <= b and not a;
    layer3_outputs(2778) <= '0';
    layer3_outputs(2779) <= not b;
    layer3_outputs(2780) <= not b;
    layer3_outputs(2781) <= b;
    layer3_outputs(2782) <= '0';
    layer3_outputs(2783) <= a and b;
    layer3_outputs(2784) <= not b;
    layer3_outputs(2785) <= a or b;
    layer3_outputs(2786) <= not a or b;
    layer3_outputs(2787) <= a;
    layer3_outputs(2788) <= b and not a;
    layer3_outputs(2789) <= b and not a;
    layer3_outputs(2790) <= a or b;
    layer3_outputs(2791) <= a or b;
    layer3_outputs(2792) <= not b;
    layer3_outputs(2793) <= b;
    layer3_outputs(2794) <= not (a or b);
    layer3_outputs(2795) <= not b;
    layer3_outputs(2796) <= not (a and b);
    layer3_outputs(2797) <= not a or b;
    layer3_outputs(2798) <= not b;
    layer3_outputs(2799) <= a and not b;
    layer3_outputs(2800) <= a or b;
    layer3_outputs(2801) <= b;
    layer3_outputs(2802) <= a and not b;
    layer3_outputs(2803) <= not (a xor b);
    layer3_outputs(2804) <= not a;
    layer3_outputs(2805) <= not a;
    layer3_outputs(2806) <= a and not b;
    layer3_outputs(2807) <= a or b;
    layer3_outputs(2808) <= not b;
    layer3_outputs(2809) <= not (a or b);
    layer3_outputs(2810) <= b;
    layer3_outputs(2811) <= b;
    layer3_outputs(2812) <= '0';
    layer3_outputs(2813) <= a xor b;
    layer3_outputs(2814) <= not a;
    layer3_outputs(2815) <= a;
    layer3_outputs(2816) <= a xor b;
    layer3_outputs(2817) <= '1';
    layer3_outputs(2818) <= '0';
    layer3_outputs(2819) <= not (a and b);
    layer3_outputs(2820) <= a;
    layer3_outputs(2821) <= not a;
    layer3_outputs(2822) <= not (a or b);
    layer3_outputs(2823) <= not b or a;
    layer3_outputs(2824) <= not a or b;
    layer3_outputs(2825) <= '1';
    layer3_outputs(2826) <= not a;
    layer3_outputs(2827) <= not a;
    layer3_outputs(2828) <= '0';
    layer3_outputs(2829) <= not a;
    layer3_outputs(2830) <= not (a and b);
    layer3_outputs(2831) <= not (a and b);
    layer3_outputs(2832) <= not a;
    layer3_outputs(2833) <= not a;
    layer3_outputs(2834) <= b and not a;
    layer3_outputs(2835) <= a;
    layer3_outputs(2836) <= a;
    layer3_outputs(2837) <= not b;
    layer3_outputs(2838) <= not a or b;
    layer3_outputs(2839) <= a;
    layer3_outputs(2840) <= not a;
    layer3_outputs(2841) <= a and b;
    layer3_outputs(2842) <= b;
    layer3_outputs(2843) <= a or b;
    layer3_outputs(2844) <= not (a or b);
    layer3_outputs(2845) <= a and b;
    layer3_outputs(2846) <= not a;
    layer3_outputs(2847) <= b;
    layer3_outputs(2848) <= not a;
    layer3_outputs(2849) <= a;
    layer3_outputs(2850) <= not a;
    layer3_outputs(2851) <= b;
    layer3_outputs(2852) <= a or b;
    layer3_outputs(2853) <= not b or a;
    layer3_outputs(2854) <= a and b;
    layer3_outputs(2855) <= b and not a;
    layer3_outputs(2856) <= not (a or b);
    layer3_outputs(2857) <= a xor b;
    layer3_outputs(2858) <= not (a or b);
    layer3_outputs(2859) <= b;
    layer3_outputs(2860) <= not (a and b);
    layer3_outputs(2861) <= not (a or b);
    layer3_outputs(2862) <= '1';
    layer3_outputs(2863) <= not (a or b);
    layer3_outputs(2864) <= not a or b;
    layer3_outputs(2865) <= not b or a;
    layer3_outputs(2866) <= a and not b;
    layer3_outputs(2867) <= not b or a;
    layer3_outputs(2868) <= not (a and b);
    layer3_outputs(2869) <= '0';
    layer3_outputs(2870) <= a or b;
    layer3_outputs(2871) <= b;
    layer3_outputs(2872) <= not b;
    layer3_outputs(2873) <= b;
    layer3_outputs(2874) <= a and not b;
    layer3_outputs(2875) <= not a;
    layer3_outputs(2876) <= b;
    layer3_outputs(2877) <= b;
    layer3_outputs(2878) <= not (a and b);
    layer3_outputs(2879) <= a;
    layer3_outputs(2880) <= not b or a;
    layer3_outputs(2881) <= a and b;
    layer3_outputs(2882) <= a or b;
    layer3_outputs(2883) <= b and not a;
    layer3_outputs(2884) <= not b;
    layer3_outputs(2885) <= a;
    layer3_outputs(2886) <= b;
    layer3_outputs(2887) <= a xor b;
    layer3_outputs(2888) <= not a;
    layer3_outputs(2889) <= not (a xor b);
    layer3_outputs(2890) <= not a;
    layer3_outputs(2891) <= a and b;
    layer3_outputs(2892) <= a or b;
    layer3_outputs(2893) <= not b;
    layer3_outputs(2894) <= a or b;
    layer3_outputs(2895) <= not (a or b);
    layer3_outputs(2896) <= '0';
    layer3_outputs(2897) <= not (a or b);
    layer3_outputs(2898) <= not (a or b);
    layer3_outputs(2899) <= not a;
    layer3_outputs(2900) <= not a;
    layer3_outputs(2901) <= '1';
    layer3_outputs(2902) <= not (a xor b);
    layer3_outputs(2903) <= '1';
    layer3_outputs(2904) <= a;
    layer3_outputs(2905) <= a;
    layer3_outputs(2906) <= a and not b;
    layer3_outputs(2907) <= a and not b;
    layer3_outputs(2908) <= b;
    layer3_outputs(2909) <= not (a or b);
    layer3_outputs(2910) <= a;
    layer3_outputs(2911) <= a xor b;
    layer3_outputs(2912) <= a and not b;
    layer3_outputs(2913) <= not b or a;
    layer3_outputs(2914) <= b and not a;
    layer3_outputs(2915) <= a and b;
    layer3_outputs(2916) <= not a;
    layer3_outputs(2917) <= not (a xor b);
    layer3_outputs(2918) <= a and b;
    layer3_outputs(2919) <= not (a or b);
    layer3_outputs(2920) <= a and b;
    layer3_outputs(2921) <= not a or b;
    layer3_outputs(2922) <= b;
    layer3_outputs(2923) <= b and not a;
    layer3_outputs(2924) <= not (a and b);
    layer3_outputs(2925) <= not b or a;
    layer3_outputs(2926) <= not b;
    layer3_outputs(2927) <= a and not b;
    layer3_outputs(2928) <= not a;
    layer3_outputs(2929) <= a and b;
    layer3_outputs(2930) <= not b;
    layer3_outputs(2931) <= a and b;
    layer3_outputs(2932) <= '0';
    layer3_outputs(2933) <= b;
    layer3_outputs(2934) <= a and not b;
    layer3_outputs(2935) <= a and b;
    layer3_outputs(2936) <= '1';
    layer3_outputs(2937) <= not a;
    layer3_outputs(2938) <= not b or a;
    layer3_outputs(2939) <= '1';
    layer3_outputs(2940) <= a or b;
    layer3_outputs(2941) <= a or b;
    layer3_outputs(2942) <= a and b;
    layer3_outputs(2943) <= a and b;
    layer3_outputs(2944) <= b;
    layer3_outputs(2945) <= b and not a;
    layer3_outputs(2946) <= not b or a;
    layer3_outputs(2947) <= a and b;
    layer3_outputs(2948) <= not a;
    layer3_outputs(2949) <= '0';
    layer3_outputs(2950) <= a;
    layer3_outputs(2951) <= not b;
    layer3_outputs(2952) <= b;
    layer3_outputs(2953) <= a and b;
    layer3_outputs(2954) <= b and not a;
    layer3_outputs(2955) <= not a or b;
    layer3_outputs(2956) <= '1';
    layer3_outputs(2957) <= a;
    layer3_outputs(2958) <= not (a or b);
    layer3_outputs(2959) <= not (a or b);
    layer3_outputs(2960) <= a or b;
    layer3_outputs(2961) <= a and not b;
    layer3_outputs(2962) <= not b;
    layer3_outputs(2963) <= not b;
    layer3_outputs(2964) <= '0';
    layer3_outputs(2965) <= not b;
    layer3_outputs(2966) <= a;
    layer3_outputs(2967) <= b;
    layer3_outputs(2968) <= not (a and b);
    layer3_outputs(2969) <= not (a or b);
    layer3_outputs(2970) <= a or b;
    layer3_outputs(2971) <= not (a or b);
    layer3_outputs(2972) <= a or b;
    layer3_outputs(2973) <= not a;
    layer3_outputs(2974) <= not a or b;
    layer3_outputs(2975) <= not b;
    layer3_outputs(2976) <= not b;
    layer3_outputs(2977) <= not (a and b);
    layer3_outputs(2978) <= a;
    layer3_outputs(2979) <= not (a and b);
    layer3_outputs(2980) <= a and not b;
    layer3_outputs(2981) <= not a;
    layer3_outputs(2982) <= a or b;
    layer3_outputs(2983) <= not b;
    layer3_outputs(2984) <= not (a and b);
    layer3_outputs(2985) <= a and not b;
    layer3_outputs(2986) <= a;
    layer3_outputs(2987) <= not b;
    layer3_outputs(2988) <= a xor b;
    layer3_outputs(2989) <= not (a or b);
    layer3_outputs(2990) <= b;
    layer3_outputs(2991) <= b;
    layer3_outputs(2992) <= not a or b;
    layer3_outputs(2993) <= not a;
    layer3_outputs(2994) <= not b or a;
    layer3_outputs(2995) <= not (a or b);
    layer3_outputs(2996) <= not b;
    layer3_outputs(2997) <= '0';
    layer3_outputs(2998) <= not a;
    layer3_outputs(2999) <= b and not a;
    layer3_outputs(3000) <= not a;
    layer3_outputs(3001) <= not a or b;
    layer3_outputs(3002) <= a and not b;
    layer3_outputs(3003) <= not (a or b);
    layer3_outputs(3004) <= not (a or b);
    layer3_outputs(3005) <= a and not b;
    layer3_outputs(3006) <= a and not b;
    layer3_outputs(3007) <= b and not a;
    layer3_outputs(3008) <= not a or b;
    layer3_outputs(3009) <= not (a xor b);
    layer3_outputs(3010) <= not b;
    layer3_outputs(3011) <= not a;
    layer3_outputs(3012) <= not b or a;
    layer3_outputs(3013) <= b and not a;
    layer3_outputs(3014) <= b and not a;
    layer3_outputs(3015) <= not (a xor b);
    layer3_outputs(3016) <= a or b;
    layer3_outputs(3017) <= b;
    layer3_outputs(3018) <= a xor b;
    layer3_outputs(3019) <= b and not a;
    layer3_outputs(3020) <= '0';
    layer3_outputs(3021) <= b;
    layer3_outputs(3022) <= not (a or b);
    layer3_outputs(3023) <= b and not a;
    layer3_outputs(3024) <= a or b;
    layer3_outputs(3025) <= a and b;
    layer3_outputs(3026) <= a or b;
    layer3_outputs(3027) <= not a;
    layer3_outputs(3028) <= not (a or b);
    layer3_outputs(3029) <= a or b;
    layer3_outputs(3030) <= not a;
    layer3_outputs(3031) <= not (a or b);
    layer3_outputs(3032) <= a and b;
    layer3_outputs(3033) <= a xor b;
    layer3_outputs(3034) <= '0';
    layer3_outputs(3035) <= not (a and b);
    layer3_outputs(3036) <= a xor b;
    layer3_outputs(3037) <= a;
    layer3_outputs(3038) <= not b or a;
    layer3_outputs(3039) <= b and not a;
    layer3_outputs(3040) <= not (a and b);
    layer3_outputs(3041) <= '0';
    layer3_outputs(3042) <= not (a and b);
    layer3_outputs(3043) <= not b;
    layer3_outputs(3044) <= a;
    layer3_outputs(3045) <= not a or b;
    layer3_outputs(3046) <= a xor b;
    layer3_outputs(3047) <= b;
    layer3_outputs(3048) <= not (a and b);
    layer3_outputs(3049) <= '0';
    layer3_outputs(3050) <= a and b;
    layer3_outputs(3051) <= not a;
    layer3_outputs(3052) <= b;
    layer3_outputs(3053) <= b;
    layer3_outputs(3054) <= b and not a;
    layer3_outputs(3055) <= not a or b;
    layer3_outputs(3056) <= not a or b;
    layer3_outputs(3057) <= a and not b;
    layer3_outputs(3058) <= not (a or b);
    layer3_outputs(3059) <= a;
    layer3_outputs(3060) <= not (a or b);
    layer3_outputs(3061) <= not b or a;
    layer3_outputs(3062) <= not (a or b);
    layer3_outputs(3063) <= a;
    layer3_outputs(3064) <= not b;
    layer3_outputs(3065) <= not a or b;
    layer3_outputs(3066) <= not (a or b);
    layer3_outputs(3067) <= a or b;
    layer3_outputs(3068) <= a and b;
    layer3_outputs(3069) <= '0';
    layer3_outputs(3070) <= a;
    layer3_outputs(3071) <= not (a and b);
    layer3_outputs(3072) <= b and not a;
    layer3_outputs(3073) <= not (a xor b);
    layer3_outputs(3074) <= '0';
    layer3_outputs(3075) <= not a;
    layer3_outputs(3076) <= a or b;
    layer3_outputs(3077) <= not b or a;
    layer3_outputs(3078) <= not a;
    layer3_outputs(3079) <= a;
    layer3_outputs(3080) <= b;
    layer3_outputs(3081) <= not b;
    layer3_outputs(3082) <= '1';
    layer3_outputs(3083) <= '1';
    layer3_outputs(3084) <= '1';
    layer3_outputs(3085) <= '1';
    layer3_outputs(3086) <= '1';
    layer3_outputs(3087) <= not (a and b);
    layer3_outputs(3088) <= '0';
    layer3_outputs(3089) <= b;
    layer3_outputs(3090) <= a or b;
    layer3_outputs(3091) <= not a;
    layer3_outputs(3092) <= not (a or b);
    layer3_outputs(3093) <= a;
    layer3_outputs(3094) <= a xor b;
    layer3_outputs(3095) <= a and b;
    layer3_outputs(3096) <= a and b;
    layer3_outputs(3097) <= a;
    layer3_outputs(3098) <= a and b;
    layer3_outputs(3099) <= '0';
    layer3_outputs(3100) <= a;
    layer3_outputs(3101) <= a or b;
    layer3_outputs(3102) <= not (a or b);
    layer3_outputs(3103) <= a and not b;
    layer3_outputs(3104) <= '0';
    layer3_outputs(3105) <= a or b;
    layer3_outputs(3106) <= a or b;
    layer3_outputs(3107) <= not b or a;
    layer3_outputs(3108) <= b;
    layer3_outputs(3109) <= b;
    layer3_outputs(3110) <= not a or b;
    layer3_outputs(3111) <= not b or a;
    layer3_outputs(3112) <= b;
    layer3_outputs(3113) <= a;
    layer3_outputs(3114) <= a xor b;
    layer3_outputs(3115) <= a;
    layer3_outputs(3116) <= not (a or b);
    layer3_outputs(3117) <= b and not a;
    layer3_outputs(3118) <= not b;
    layer3_outputs(3119) <= a and not b;
    layer3_outputs(3120) <= not b or a;
    layer3_outputs(3121) <= not b;
    layer3_outputs(3122) <= a and not b;
    layer3_outputs(3123) <= b and not a;
    layer3_outputs(3124) <= not b or a;
    layer3_outputs(3125) <= not (a or b);
    layer3_outputs(3126) <= b and not a;
    layer3_outputs(3127) <= not (a or b);
    layer3_outputs(3128) <= b;
    layer3_outputs(3129) <= not (a or b);
    layer3_outputs(3130) <= b and not a;
    layer3_outputs(3131) <= a xor b;
    layer3_outputs(3132) <= not (a and b);
    layer3_outputs(3133) <= not a or b;
    layer3_outputs(3134) <= not (a or b);
    layer3_outputs(3135) <= '0';
    layer3_outputs(3136) <= not b;
    layer3_outputs(3137) <= '0';
    layer3_outputs(3138) <= b;
    layer3_outputs(3139) <= a;
    layer3_outputs(3140) <= a and b;
    layer3_outputs(3141) <= '1';
    layer3_outputs(3142) <= not a;
    layer3_outputs(3143) <= not b;
    layer3_outputs(3144) <= '0';
    layer3_outputs(3145) <= not (a and b);
    layer3_outputs(3146) <= not (a or b);
    layer3_outputs(3147) <= b;
    layer3_outputs(3148) <= not a;
    layer3_outputs(3149) <= a and b;
    layer3_outputs(3150) <= not b;
    layer3_outputs(3151) <= a and b;
    layer3_outputs(3152) <= a;
    layer3_outputs(3153) <= a and b;
    layer3_outputs(3154) <= b and not a;
    layer3_outputs(3155) <= a and not b;
    layer3_outputs(3156) <= b;
    layer3_outputs(3157) <= not (a and b);
    layer3_outputs(3158) <= a;
    layer3_outputs(3159) <= not a;
    layer3_outputs(3160) <= '0';
    layer3_outputs(3161) <= not (a xor b);
    layer3_outputs(3162) <= not b or a;
    layer3_outputs(3163) <= b;
    layer3_outputs(3164) <= a or b;
    layer3_outputs(3165) <= not a or b;
    layer3_outputs(3166) <= not b;
    layer3_outputs(3167) <= a and not b;
    layer3_outputs(3168) <= b;
    layer3_outputs(3169) <= not (a or b);
    layer3_outputs(3170) <= a;
    layer3_outputs(3171) <= not b;
    layer3_outputs(3172) <= b and not a;
    layer3_outputs(3173) <= not (a and b);
    layer3_outputs(3174) <= not (a xor b);
    layer3_outputs(3175) <= '1';
    layer3_outputs(3176) <= a and b;
    layer3_outputs(3177) <= a and not b;
    layer3_outputs(3178) <= b;
    layer3_outputs(3179) <= a;
    layer3_outputs(3180) <= a;
    layer3_outputs(3181) <= b;
    layer3_outputs(3182) <= not b or a;
    layer3_outputs(3183) <= not a or b;
    layer3_outputs(3184) <= not (a xor b);
    layer3_outputs(3185) <= a and not b;
    layer3_outputs(3186) <= not b or a;
    layer3_outputs(3187) <= b and not a;
    layer3_outputs(3188) <= b;
    layer3_outputs(3189) <= not b or a;
    layer3_outputs(3190) <= not (a and b);
    layer3_outputs(3191) <= a;
    layer3_outputs(3192) <= '1';
    layer3_outputs(3193) <= not a or b;
    layer3_outputs(3194) <= b;
    layer3_outputs(3195) <= a;
    layer3_outputs(3196) <= not a;
    layer3_outputs(3197) <= not a;
    layer3_outputs(3198) <= '0';
    layer3_outputs(3199) <= a and not b;
    layer3_outputs(3200) <= not (a and b);
    layer3_outputs(3201) <= not b;
    layer3_outputs(3202) <= a or b;
    layer3_outputs(3203) <= b;
    layer3_outputs(3204) <= b;
    layer3_outputs(3205) <= not b or a;
    layer3_outputs(3206) <= a and b;
    layer3_outputs(3207) <= not b;
    layer3_outputs(3208) <= a and b;
    layer3_outputs(3209) <= a and not b;
    layer3_outputs(3210) <= a and not b;
    layer3_outputs(3211) <= not b;
    layer3_outputs(3212) <= not a;
    layer3_outputs(3213) <= not a or b;
    layer3_outputs(3214) <= not b or a;
    layer3_outputs(3215) <= not (a or b);
    layer3_outputs(3216) <= a;
    layer3_outputs(3217) <= a and not b;
    layer3_outputs(3218) <= not a;
    layer3_outputs(3219) <= b;
    layer3_outputs(3220) <= a xor b;
    layer3_outputs(3221) <= a or b;
    layer3_outputs(3222) <= not (a and b);
    layer3_outputs(3223) <= not b;
    layer3_outputs(3224) <= not b;
    layer3_outputs(3225) <= not a;
    layer3_outputs(3226) <= not b;
    layer3_outputs(3227) <= a;
    layer3_outputs(3228) <= not (a and b);
    layer3_outputs(3229) <= not b;
    layer3_outputs(3230) <= a;
    layer3_outputs(3231) <= '0';
    layer3_outputs(3232) <= not b or a;
    layer3_outputs(3233) <= a and b;
    layer3_outputs(3234) <= not (a xor b);
    layer3_outputs(3235) <= a and not b;
    layer3_outputs(3236) <= b and not a;
    layer3_outputs(3237) <= not b or a;
    layer3_outputs(3238) <= not a or b;
    layer3_outputs(3239) <= not a or b;
    layer3_outputs(3240) <= a and not b;
    layer3_outputs(3241) <= b and not a;
    layer3_outputs(3242) <= not a or b;
    layer3_outputs(3243) <= a;
    layer3_outputs(3244) <= b;
    layer3_outputs(3245) <= b and not a;
    layer3_outputs(3246) <= not a;
    layer3_outputs(3247) <= b;
    layer3_outputs(3248) <= '1';
    layer3_outputs(3249) <= not (a xor b);
    layer3_outputs(3250) <= not b;
    layer3_outputs(3251) <= a;
    layer3_outputs(3252) <= a;
    layer3_outputs(3253) <= a;
    layer3_outputs(3254) <= not b;
    layer3_outputs(3255) <= not (a and b);
    layer3_outputs(3256) <= '1';
    layer3_outputs(3257) <= not b or a;
    layer3_outputs(3258) <= b and not a;
    layer3_outputs(3259) <= a and not b;
    layer3_outputs(3260) <= '1';
    layer3_outputs(3261) <= not a or b;
    layer3_outputs(3262) <= a and not b;
    layer3_outputs(3263) <= not (a or b);
    layer3_outputs(3264) <= a xor b;
    layer3_outputs(3265) <= a and b;
    layer3_outputs(3266) <= not a;
    layer3_outputs(3267) <= not b;
    layer3_outputs(3268) <= not (a xor b);
    layer3_outputs(3269) <= not (a xor b);
    layer3_outputs(3270) <= not b;
    layer3_outputs(3271) <= '1';
    layer3_outputs(3272) <= not b or a;
    layer3_outputs(3273) <= not a;
    layer3_outputs(3274) <= '0';
    layer3_outputs(3275) <= a;
    layer3_outputs(3276) <= '0';
    layer3_outputs(3277) <= not (a and b);
    layer3_outputs(3278) <= not a or b;
    layer3_outputs(3279) <= not (a xor b);
    layer3_outputs(3280) <= a;
    layer3_outputs(3281) <= a;
    layer3_outputs(3282) <= not b or a;
    layer3_outputs(3283) <= a or b;
    layer3_outputs(3284) <= a and not b;
    layer3_outputs(3285) <= not b;
    layer3_outputs(3286) <= '1';
    layer3_outputs(3287) <= not a;
    layer3_outputs(3288) <= not (a or b);
    layer3_outputs(3289) <= not b or a;
    layer3_outputs(3290) <= a and b;
    layer3_outputs(3291) <= not a;
    layer3_outputs(3292) <= a or b;
    layer3_outputs(3293) <= a or b;
    layer3_outputs(3294) <= b;
    layer3_outputs(3295) <= a and not b;
    layer3_outputs(3296) <= a or b;
    layer3_outputs(3297) <= not b;
    layer3_outputs(3298) <= a or b;
    layer3_outputs(3299) <= not (a and b);
    layer3_outputs(3300) <= not (a xor b);
    layer3_outputs(3301) <= a;
    layer3_outputs(3302) <= b;
    layer3_outputs(3303) <= b and not a;
    layer3_outputs(3304) <= b and not a;
    layer3_outputs(3305) <= not b or a;
    layer3_outputs(3306) <= not b or a;
    layer3_outputs(3307) <= not a;
    layer3_outputs(3308) <= '0';
    layer3_outputs(3309) <= not (a xor b);
    layer3_outputs(3310) <= '1';
    layer3_outputs(3311) <= not a;
    layer3_outputs(3312) <= a and b;
    layer3_outputs(3313) <= not (a and b);
    layer3_outputs(3314) <= a and b;
    layer3_outputs(3315) <= not (a xor b);
    layer3_outputs(3316) <= not b or a;
    layer3_outputs(3317) <= not a or b;
    layer3_outputs(3318) <= b;
    layer3_outputs(3319) <= a;
    layer3_outputs(3320) <= a or b;
    layer3_outputs(3321) <= a and b;
    layer3_outputs(3322) <= not a or b;
    layer3_outputs(3323) <= not b;
    layer3_outputs(3324) <= a and b;
    layer3_outputs(3325) <= not b or a;
    layer3_outputs(3326) <= not b;
    layer3_outputs(3327) <= not b;
    layer3_outputs(3328) <= not (a xor b);
    layer3_outputs(3329) <= not (a or b);
    layer3_outputs(3330) <= '0';
    layer3_outputs(3331) <= b;
    layer3_outputs(3332) <= a and not b;
    layer3_outputs(3333) <= not (a and b);
    layer3_outputs(3334) <= '0';
    layer3_outputs(3335) <= not b;
    layer3_outputs(3336) <= b;
    layer3_outputs(3337) <= not a or b;
    layer3_outputs(3338) <= not a;
    layer3_outputs(3339) <= a xor b;
    layer3_outputs(3340) <= a and not b;
    layer3_outputs(3341) <= a or b;
    layer3_outputs(3342) <= '0';
    layer3_outputs(3343) <= not a or b;
    layer3_outputs(3344) <= not (a xor b);
    layer3_outputs(3345) <= a or b;
    layer3_outputs(3346) <= not (a xor b);
    layer3_outputs(3347) <= not a;
    layer3_outputs(3348) <= not (a or b);
    layer3_outputs(3349) <= not (a or b);
    layer3_outputs(3350) <= not b or a;
    layer3_outputs(3351) <= a;
    layer3_outputs(3352) <= b and not a;
    layer3_outputs(3353) <= a and not b;
    layer3_outputs(3354) <= not a or b;
    layer3_outputs(3355) <= not (a or b);
    layer3_outputs(3356) <= a or b;
    layer3_outputs(3357) <= not a or b;
    layer3_outputs(3358) <= a and b;
    layer3_outputs(3359) <= b;
    layer3_outputs(3360) <= not b or a;
    layer3_outputs(3361) <= not b or a;
    layer3_outputs(3362) <= a and not b;
    layer3_outputs(3363) <= a xor b;
    layer3_outputs(3364) <= not a;
    layer3_outputs(3365) <= b;
    layer3_outputs(3366) <= a and b;
    layer3_outputs(3367) <= not b;
    layer3_outputs(3368) <= not (a and b);
    layer3_outputs(3369) <= a;
    layer3_outputs(3370) <= a and b;
    layer3_outputs(3371) <= a and b;
    layer3_outputs(3372) <= b and not a;
    layer3_outputs(3373) <= a and b;
    layer3_outputs(3374) <= a or b;
    layer3_outputs(3375) <= not a;
    layer3_outputs(3376) <= not b;
    layer3_outputs(3377) <= b and not a;
    layer3_outputs(3378) <= a;
    layer3_outputs(3379) <= not b;
    layer3_outputs(3380) <= not (a or b);
    layer3_outputs(3381) <= a and b;
    layer3_outputs(3382) <= not (a and b);
    layer3_outputs(3383) <= b;
    layer3_outputs(3384) <= not a;
    layer3_outputs(3385) <= not (a and b);
    layer3_outputs(3386) <= a;
    layer3_outputs(3387) <= a;
    layer3_outputs(3388) <= not b;
    layer3_outputs(3389) <= b;
    layer3_outputs(3390) <= b and not a;
    layer3_outputs(3391) <= not a or b;
    layer3_outputs(3392) <= a or b;
    layer3_outputs(3393) <= a and not b;
    layer3_outputs(3394) <= '1';
    layer3_outputs(3395) <= not a;
    layer3_outputs(3396) <= not (a and b);
    layer3_outputs(3397) <= b;
    layer3_outputs(3398) <= not a;
    layer3_outputs(3399) <= b;
    layer3_outputs(3400) <= not (a and b);
    layer3_outputs(3401) <= a;
    layer3_outputs(3402) <= a;
    layer3_outputs(3403) <= not a;
    layer3_outputs(3404) <= a and not b;
    layer3_outputs(3405) <= not b;
    layer3_outputs(3406) <= b;
    layer3_outputs(3407) <= b;
    layer3_outputs(3408) <= '0';
    layer3_outputs(3409) <= not b;
    layer3_outputs(3410) <= not (a and b);
    layer3_outputs(3411) <= not (a and b);
    layer3_outputs(3412) <= not a;
    layer3_outputs(3413) <= not b or a;
    layer3_outputs(3414) <= a or b;
    layer3_outputs(3415) <= not (a and b);
    layer3_outputs(3416) <= a xor b;
    layer3_outputs(3417) <= b and not a;
    layer3_outputs(3418) <= not b or a;
    layer3_outputs(3419) <= '1';
    layer3_outputs(3420) <= not a;
    layer3_outputs(3421) <= not b or a;
    layer3_outputs(3422) <= a or b;
    layer3_outputs(3423) <= b;
    layer3_outputs(3424) <= not a or b;
    layer3_outputs(3425) <= a and b;
    layer3_outputs(3426) <= not a or b;
    layer3_outputs(3427) <= a;
    layer3_outputs(3428) <= not a or b;
    layer3_outputs(3429) <= a;
    layer3_outputs(3430) <= not b or a;
    layer3_outputs(3431) <= '0';
    layer3_outputs(3432) <= '0';
    layer3_outputs(3433) <= a or b;
    layer3_outputs(3434) <= not (a and b);
    layer3_outputs(3435) <= b and not a;
    layer3_outputs(3436) <= not a;
    layer3_outputs(3437) <= a and not b;
    layer3_outputs(3438) <= a and b;
    layer3_outputs(3439) <= a;
    layer3_outputs(3440) <= a;
    layer3_outputs(3441) <= not b;
    layer3_outputs(3442) <= b and not a;
    layer3_outputs(3443) <= not (a and b);
    layer3_outputs(3444) <= a and not b;
    layer3_outputs(3445) <= not (a or b);
    layer3_outputs(3446) <= not a;
    layer3_outputs(3447) <= not b or a;
    layer3_outputs(3448) <= a;
    layer3_outputs(3449) <= '1';
    layer3_outputs(3450) <= '0';
    layer3_outputs(3451) <= not (a xor b);
    layer3_outputs(3452) <= not b;
    layer3_outputs(3453) <= a;
    layer3_outputs(3454) <= not a or b;
    layer3_outputs(3455) <= a xor b;
    layer3_outputs(3456) <= not (a or b);
    layer3_outputs(3457) <= not a or b;
    layer3_outputs(3458) <= a;
    layer3_outputs(3459) <= b;
    layer3_outputs(3460) <= a and b;
    layer3_outputs(3461) <= a or b;
    layer3_outputs(3462) <= not b;
    layer3_outputs(3463) <= a;
    layer3_outputs(3464) <= a or b;
    layer3_outputs(3465) <= not b;
    layer3_outputs(3466) <= a;
    layer3_outputs(3467) <= b;
    layer3_outputs(3468) <= a;
    layer3_outputs(3469) <= not a or b;
    layer3_outputs(3470) <= a and not b;
    layer3_outputs(3471) <= not b or a;
    layer3_outputs(3472) <= b;
    layer3_outputs(3473) <= a and not b;
    layer3_outputs(3474) <= not b or a;
    layer3_outputs(3475) <= a;
    layer3_outputs(3476) <= a;
    layer3_outputs(3477) <= not (a and b);
    layer3_outputs(3478) <= not b or a;
    layer3_outputs(3479) <= b;
    layer3_outputs(3480) <= a xor b;
    layer3_outputs(3481) <= not b;
    layer3_outputs(3482) <= a and b;
    layer3_outputs(3483) <= a;
    layer3_outputs(3484) <= a and not b;
    layer3_outputs(3485) <= not a or b;
    layer3_outputs(3486) <= not (a or b);
    layer3_outputs(3487) <= not (a or b);
    layer3_outputs(3488) <= not a;
    layer3_outputs(3489) <= not (a or b);
    layer3_outputs(3490) <= a;
    layer3_outputs(3491) <= a;
    layer3_outputs(3492) <= not b;
    layer3_outputs(3493) <= not (a and b);
    layer3_outputs(3494) <= not a;
    layer3_outputs(3495) <= not (a xor b);
    layer3_outputs(3496) <= b and not a;
    layer3_outputs(3497) <= not b;
    layer3_outputs(3498) <= a;
    layer3_outputs(3499) <= not (a or b);
    layer3_outputs(3500) <= not b;
    layer3_outputs(3501) <= a and b;
    layer3_outputs(3502) <= not b;
    layer3_outputs(3503) <= not a;
    layer3_outputs(3504) <= not b or a;
    layer3_outputs(3505) <= not (a and b);
    layer3_outputs(3506) <= b;
    layer3_outputs(3507) <= a or b;
    layer3_outputs(3508) <= b and not a;
    layer3_outputs(3509) <= a;
    layer3_outputs(3510) <= not a;
    layer3_outputs(3511) <= b;
    layer3_outputs(3512) <= not a;
    layer3_outputs(3513) <= not a or b;
    layer3_outputs(3514) <= a and not b;
    layer3_outputs(3515) <= not (a and b);
    layer3_outputs(3516) <= a xor b;
    layer3_outputs(3517) <= not a;
    layer3_outputs(3518) <= a and not b;
    layer3_outputs(3519) <= a;
    layer3_outputs(3520) <= not (a and b);
    layer3_outputs(3521) <= b;
    layer3_outputs(3522) <= b and not a;
    layer3_outputs(3523) <= not (a and b);
    layer3_outputs(3524) <= not b or a;
    layer3_outputs(3525) <= not a;
    layer3_outputs(3526) <= not (a xor b);
    layer3_outputs(3527) <= a;
    layer3_outputs(3528) <= a;
    layer3_outputs(3529) <= a and b;
    layer3_outputs(3530) <= not a or b;
    layer3_outputs(3531) <= a and b;
    layer3_outputs(3532) <= not (a or b);
    layer3_outputs(3533) <= not (a or b);
    layer3_outputs(3534) <= b;
    layer3_outputs(3535) <= b;
    layer3_outputs(3536) <= '1';
    layer3_outputs(3537) <= '0';
    layer3_outputs(3538) <= b;
    layer3_outputs(3539) <= b;
    layer3_outputs(3540) <= b;
    layer3_outputs(3541) <= b and not a;
    layer3_outputs(3542) <= '1';
    layer3_outputs(3543) <= '1';
    layer3_outputs(3544) <= not b;
    layer3_outputs(3545) <= b;
    layer3_outputs(3546) <= b;
    layer3_outputs(3547) <= not (a and b);
    layer3_outputs(3548) <= not (a and b);
    layer3_outputs(3549) <= not a;
    layer3_outputs(3550) <= a and b;
    layer3_outputs(3551) <= not b;
    layer3_outputs(3552) <= b and not a;
    layer3_outputs(3553) <= a and b;
    layer3_outputs(3554) <= '0';
    layer3_outputs(3555) <= not (a or b);
    layer3_outputs(3556) <= not a or b;
    layer3_outputs(3557) <= not (a or b);
    layer3_outputs(3558) <= b and not a;
    layer3_outputs(3559) <= not a;
    layer3_outputs(3560) <= not a;
    layer3_outputs(3561) <= not a;
    layer3_outputs(3562) <= '0';
    layer3_outputs(3563) <= b;
    layer3_outputs(3564) <= a or b;
    layer3_outputs(3565) <= not a or b;
    layer3_outputs(3566) <= b and not a;
    layer3_outputs(3567) <= not (a and b);
    layer3_outputs(3568) <= a and not b;
    layer3_outputs(3569) <= not (a or b);
    layer3_outputs(3570) <= a and b;
    layer3_outputs(3571) <= b;
    layer3_outputs(3572) <= not a;
    layer3_outputs(3573) <= a or b;
    layer3_outputs(3574) <= not (a or b);
    layer3_outputs(3575) <= a or b;
    layer3_outputs(3576) <= a and not b;
    layer3_outputs(3577) <= a;
    layer3_outputs(3578) <= b and not a;
    layer3_outputs(3579) <= a;
    layer3_outputs(3580) <= not (a and b);
    layer3_outputs(3581) <= a;
    layer3_outputs(3582) <= a and b;
    layer3_outputs(3583) <= not a or b;
    layer3_outputs(3584) <= b and not a;
    layer3_outputs(3585) <= not b;
    layer3_outputs(3586) <= not a;
    layer3_outputs(3587) <= not (a and b);
    layer3_outputs(3588) <= not (a or b);
    layer3_outputs(3589) <= a;
    layer3_outputs(3590) <= not a;
    layer3_outputs(3591) <= not a or b;
    layer3_outputs(3592) <= not (a and b);
    layer3_outputs(3593) <= not a;
    layer3_outputs(3594) <= not (a or b);
    layer3_outputs(3595) <= b;
    layer3_outputs(3596) <= a or b;
    layer3_outputs(3597) <= b;
    layer3_outputs(3598) <= not b;
    layer3_outputs(3599) <= not b or a;
    layer3_outputs(3600) <= b and not a;
    layer3_outputs(3601) <= b;
    layer3_outputs(3602) <= b;
    layer3_outputs(3603) <= not b or a;
    layer3_outputs(3604) <= a and b;
    layer3_outputs(3605) <= not (a and b);
    layer3_outputs(3606) <= b;
    layer3_outputs(3607) <= a and b;
    layer3_outputs(3608) <= b;
    layer3_outputs(3609) <= not (a or b);
    layer3_outputs(3610) <= not (a or b);
    layer3_outputs(3611) <= a and not b;
    layer3_outputs(3612) <= a and not b;
    layer3_outputs(3613) <= not (a and b);
    layer3_outputs(3614) <= a and b;
    layer3_outputs(3615) <= not (a or b);
    layer3_outputs(3616) <= a and not b;
    layer3_outputs(3617) <= not b;
    layer3_outputs(3618) <= a and not b;
    layer3_outputs(3619) <= b and not a;
    layer3_outputs(3620) <= a xor b;
    layer3_outputs(3621) <= a xor b;
    layer3_outputs(3622) <= a and b;
    layer3_outputs(3623) <= not a;
    layer3_outputs(3624) <= not (a or b);
    layer3_outputs(3625) <= b and not a;
    layer3_outputs(3626) <= not b;
    layer3_outputs(3627) <= a or b;
    layer3_outputs(3628) <= a;
    layer3_outputs(3629) <= b;
    layer3_outputs(3630) <= a and b;
    layer3_outputs(3631) <= not a;
    layer3_outputs(3632) <= b;
    layer3_outputs(3633) <= b;
    layer3_outputs(3634) <= b;
    layer3_outputs(3635) <= not b;
    layer3_outputs(3636) <= b and not a;
    layer3_outputs(3637) <= a;
    layer3_outputs(3638) <= not a;
    layer3_outputs(3639) <= a;
    layer3_outputs(3640) <= not b;
    layer3_outputs(3641) <= b and not a;
    layer3_outputs(3642) <= not a;
    layer3_outputs(3643) <= b;
    layer3_outputs(3644) <= a or b;
    layer3_outputs(3645) <= not (a or b);
    layer3_outputs(3646) <= '0';
    layer3_outputs(3647) <= a xor b;
    layer3_outputs(3648) <= a and not b;
    layer3_outputs(3649) <= '0';
    layer3_outputs(3650) <= not b or a;
    layer3_outputs(3651) <= not b;
    layer3_outputs(3652) <= not b or a;
    layer3_outputs(3653) <= b;
    layer3_outputs(3654) <= not a;
    layer3_outputs(3655) <= not (a xor b);
    layer3_outputs(3656) <= not (a or b);
    layer3_outputs(3657) <= b;
    layer3_outputs(3658) <= not (a and b);
    layer3_outputs(3659) <= not b or a;
    layer3_outputs(3660) <= not (a or b);
    layer3_outputs(3661) <= not (a xor b);
    layer3_outputs(3662) <= not b;
    layer3_outputs(3663) <= not b;
    layer3_outputs(3664) <= not a;
    layer3_outputs(3665) <= not b;
    layer3_outputs(3666) <= not (a or b);
    layer3_outputs(3667) <= a xor b;
    layer3_outputs(3668) <= not a;
    layer3_outputs(3669) <= b;
    layer3_outputs(3670) <= not a;
    layer3_outputs(3671) <= b and not a;
    layer3_outputs(3672) <= not (a and b);
    layer3_outputs(3673) <= '0';
    layer3_outputs(3674) <= not (a xor b);
    layer3_outputs(3675) <= not b;
    layer3_outputs(3676) <= a and b;
    layer3_outputs(3677) <= not b;
    layer3_outputs(3678) <= not b or a;
    layer3_outputs(3679) <= '0';
    layer3_outputs(3680) <= '1';
    layer3_outputs(3681) <= not b;
    layer3_outputs(3682) <= a or b;
    layer3_outputs(3683) <= not b or a;
    layer3_outputs(3684) <= not b;
    layer3_outputs(3685) <= a;
    layer3_outputs(3686) <= a and not b;
    layer3_outputs(3687) <= a;
    layer3_outputs(3688) <= '0';
    layer3_outputs(3689) <= b;
    layer3_outputs(3690) <= not b or a;
    layer3_outputs(3691) <= not a;
    layer3_outputs(3692) <= not a or b;
    layer3_outputs(3693) <= not (a or b);
    layer3_outputs(3694) <= not b;
    layer3_outputs(3695) <= '1';
    layer3_outputs(3696) <= '0';
    layer3_outputs(3697) <= a;
    layer3_outputs(3698) <= a;
    layer3_outputs(3699) <= not (a or b);
    layer3_outputs(3700) <= a;
    layer3_outputs(3701) <= not a;
    layer3_outputs(3702) <= a or b;
    layer3_outputs(3703) <= not b;
    layer3_outputs(3704) <= a;
    layer3_outputs(3705) <= not b;
    layer3_outputs(3706) <= not a;
    layer3_outputs(3707) <= '1';
    layer3_outputs(3708) <= not b or a;
    layer3_outputs(3709) <= not (a and b);
    layer3_outputs(3710) <= a and b;
    layer3_outputs(3711) <= a;
    layer3_outputs(3712) <= not (a or b);
    layer3_outputs(3713) <= '1';
    layer3_outputs(3714) <= a or b;
    layer3_outputs(3715) <= '0';
    layer3_outputs(3716) <= not b;
    layer3_outputs(3717) <= a;
    layer3_outputs(3718) <= not a or b;
    layer3_outputs(3719) <= a xor b;
    layer3_outputs(3720) <= b;
    layer3_outputs(3721) <= a;
    layer3_outputs(3722) <= not (a and b);
    layer3_outputs(3723) <= not b;
    layer3_outputs(3724) <= a and b;
    layer3_outputs(3725) <= b and not a;
    layer3_outputs(3726) <= '0';
    layer3_outputs(3727) <= not a or b;
    layer3_outputs(3728) <= not b;
    layer3_outputs(3729) <= a;
    layer3_outputs(3730) <= b and not a;
    layer3_outputs(3731) <= b;
    layer3_outputs(3732) <= not a;
    layer3_outputs(3733) <= a;
    layer3_outputs(3734) <= a and not b;
    layer3_outputs(3735) <= a xor b;
    layer3_outputs(3736) <= '1';
    layer3_outputs(3737) <= not b;
    layer3_outputs(3738) <= not (a xor b);
    layer3_outputs(3739) <= '0';
    layer3_outputs(3740) <= not (a or b);
    layer3_outputs(3741) <= not a;
    layer3_outputs(3742) <= not a or b;
    layer3_outputs(3743) <= not b;
    layer3_outputs(3744) <= a xor b;
    layer3_outputs(3745) <= b;
    layer3_outputs(3746) <= not b or a;
    layer3_outputs(3747) <= not a;
    layer3_outputs(3748) <= not (a xor b);
    layer3_outputs(3749) <= a or b;
    layer3_outputs(3750) <= b;
    layer3_outputs(3751) <= a and b;
    layer3_outputs(3752) <= b and not a;
    layer3_outputs(3753) <= a and not b;
    layer3_outputs(3754) <= not a or b;
    layer3_outputs(3755) <= a xor b;
    layer3_outputs(3756) <= not b;
    layer3_outputs(3757) <= not a or b;
    layer3_outputs(3758) <= not (a and b);
    layer3_outputs(3759) <= not (a and b);
    layer3_outputs(3760) <= not a or b;
    layer3_outputs(3761) <= b;
    layer3_outputs(3762) <= not (a and b);
    layer3_outputs(3763) <= b and not a;
    layer3_outputs(3764) <= not b or a;
    layer3_outputs(3765) <= not a or b;
    layer3_outputs(3766) <= not b or a;
    layer3_outputs(3767) <= a and b;
    layer3_outputs(3768) <= a or b;
    layer3_outputs(3769) <= not a;
    layer3_outputs(3770) <= not (a or b);
    layer3_outputs(3771) <= not b;
    layer3_outputs(3772) <= not a or b;
    layer3_outputs(3773) <= not b;
    layer3_outputs(3774) <= b;
    layer3_outputs(3775) <= b and not a;
    layer3_outputs(3776) <= a xor b;
    layer3_outputs(3777) <= not b;
    layer3_outputs(3778) <= not b or a;
    layer3_outputs(3779) <= a or b;
    layer3_outputs(3780) <= not (a and b);
    layer3_outputs(3781) <= not a or b;
    layer3_outputs(3782) <= not a or b;
    layer3_outputs(3783) <= not a;
    layer3_outputs(3784) <= not a;
    layer3_outputs(3785) <= not (a xor b);
    layer3_outputs(3786) <= b and not a;
    layer3_outputs(3787) <= not b or a;
    layer3_outputs(3788) <= '1';
    layer3_outputs(3789) <= a;
    layer3_outputs(3790) <= b and not a;
    layer3_outputs(3791) <= not a;
    layer3_outputs(3792) <= b;
    layer3_outputs(3793) <= not a or b;
    layer3_outputs(3794) <= b;
    layer3_outputs(3795) <= b and not a;
    layer3_outputs(3796) <= b and not a;
    layer3_outputs(3797) <= a and b;
    layer3_outputs(3798) <= a;
    layer3_outputs(3799) <= a and not b;
    layer3_outputs(3800) <= not (a and b);
    layer3_outputs(3801) <= a and b;
    layer3_outputs(3802) <= not b;
    layer3_outputs(3803) <= not (a and b);
    layer3_outputs(3804) <= not b;
    layer3_outputs(3805) <= not (a xor b);
    layer3_outputs(3806) <= not (a or b);
    layer3_outputs(3807) <= a or b;
    layer3_outputs(3808) <= not a;
    layer3_outputs(3809) <= '0';
    layer3_outputs(3810) <= a and b;
    layer3_outputs(3811) <= not (a or b);
    layer3_outputs(3812) <= '1';
    layer3_outputs(3813) <= b and not a;
    layer3_outputs(3814) <= b and not a;
    layer3_outputs(3815) <= not (a or b);
    layer3_outputs(3816) <= a and b;
    layer3_outputs(3817) <= b and not a;
    layer3_outputs(3818) <= not (a and b);
    layer3_outputs(3819) <= not (a or b);
    layer3_outputs(3820) <= a or b;
    layer3_outputs(3821) <= b and not a;
    layer3_outputs(3822) <= a or b;
    layer3_outputs(3823) <= not a or b;
    layer3_outputs(3824) <= not (a or b);
    layer3_outputs(3825) <= not a;
    layer3_outputs(3826) <= not a;
    layer3_outputs(3827) <= not b or a;
    layer3_outputs(3828) <= not a;
    layer3_outputs(3829) <= not (a and b);
    layer3_outputs(3830) <= not b or a;
    layer3_outputs(3831) <= a;
    layer3_outputs(3832) <= '0';
    layer3_outputs(3833) <= a;
    layer3_outputs(3834) <= b;
    layer3_outputs(3835) <= not (a xor b);
    layer3_outputs(3836) <= a and not b;
    layer3_outputs(3837) <= a and not b;
    layer3_outputs(3838) <= not b;
    layer3_outputs(3839) <= a;
    layer3_outputs(3840) <= not (a and b);
    layer3_outputs(3841) <= not a or b;
    layer3_outputs(3842) <= not b;
    layer3_outputs(3843) <= not (a and b);
    layer3_outputs(3844) <= not b or a;
    layer3_outputs(3845) <= not a;
    layer3_outputs(3846) <= not (a and b);
    layer3_outputs(3847) <= a;
    layer3_outputs(3848) <= b;
    layer3_outputs(3849) <= a or b;
    layer3_outputs(3850) <= '1';
    layer3_outputs(3851) <= not (a or b);
    layer3_outputs(3852) <= a and not b;
    layer3_outputs(3853) <= a or b;
    layer3_outputs(3854) <= a xor b;
    layer3_outputs(3855) <= not a;
    layer3_outputs(3856) <= a;
    layer3_outputs(3857) <= not b or a;
    layer3_outputs(3858) <= not (a or b);
    layer3_outputs(3859) <= b and not a;
    layer3_outputs(3860) <= b;
    layer3_outputs(3861) <= not b;
    layer3_outputs(3862) <= b;
    layer3_outputs(3863) <= a and b;
    layer3_outputs(3864) <= not b;
    layer3_outputs(3865) <= a;
    layer3_outputs(3866) <= b and not a;
    layer3_outputs(3867) <= a or b;
    layer3_outputs(3868) <= a xor b;
    layer3_outputs(3869) <= '1';
    layer3_outputs(3870) <= not b;
    layer3_outputs(3871) <= not a;
    layer3_outputs(3872) <= a;
    layer3_outputs(3873) <= not (a and b);
    layer3_outputs(3874) <= b and not a;
    layer3_outputs(3875) <= a;
    layer3_outputs(3876) <= a;
    layer3_outputs(3877) <= not b or a;
    layer3_outputs(3878) <= a and b;
    layer3_outputs(3879) <= a or b;
    layer3_outputs(3880) <= '1';
    layer3_outputs(3881) <= a or b;
    layer3_outputs(3882) <= b;
    layer3_outputs(3883) <= a and not b;
    layer3_outputs(3884) <= not a;
    layer3_outputs(3885) <= not a or b;
    layer3_outputs(3886) <= b;
    layer3_outputs(3887) <= a or b;
    layer3_outputs(3888) <= a and b;
    layer3_outputs(3889) <= a or b;
    layer3_outputs(3890) <= a and b;
    layer3_outputs(3891) <= not a or b;
    layer3_outputs(3892) <= not b or a;
    layer3_outputs(3893) <= not b;
    layer3_outputs(3894) <= b and not a;
    layer3_outputs(3895) <= not (a xor b);
    layer3_outputs(3896) <= not b or a;
    layer3_outputs(3897) <= not a or b;
    layer3_outputs(3898) <= a and b;
    layer3_outputs(3899) <= not b;
    layer3_outputs(3900) <= a;
    layer3_outputs(3901) <= a and b;
    layer3_outputs(3902) <= b;
    layer3_outputs(3903) <= a xor b;
    layer3_outputs(3904) <= '0';
    layer3_outputs(3905) <= '1';
    layer3_outputs(3906) <= a and not b;
    layer3_outputs(3907) <= a or b;
    layer3_outputs(3908) <= not a or b;
    layer3_outputs(3909) <= not b or a;
    layer3_outputs(3910) <= a;
    layer3_outputs(3911) <= a and b;
    layer3_outputs(3912) <= a;
    layer3_outputs(3913) <= b;
    layer3_outputs(3914) <= not b;
    layer3_outputs(3915) <= not b or a;
    layer3_outputs(3916) <= not a or b;
    layer3_outputs(3917) <= not (a xor b);
    layer3_outputs(3918) <= not a;
    layer3_outputs(3919) <= not a or b;
    layer3_outputs(3920) <= a and not b;
    layer3_outputs(3921) <= not b;
    layer3_outputs(3922) <= b and not a;
    layer3_outputs(3923) <= a or b;
    layer3_outputs(3924) <= not a;
    layer3_outputs(3925) <= a and b;
    layer3_outputs(3926) <= not (a or b);
    layer3_outputs(3927) <= a;
    layer3_outputs(3928) <= a or b;
    layer3_outputs(3929) <= not (a and b);
    layer3_outputs(3930) <= a and b;
    layer3_outputs(3931) <= not b or a;
    layer3_outputs(3932) <= not b;
    layer3_outputs(3933) <= not b;
    layer3_outputs(3934) <= not b or a;
    layer3_outputs(3935) <= a xor b;
    layer3_outputs(3936) <= '1';
    layer3_outputs(3937) <= not (a and b);
    layer3_outputs(3938) <= '1';
    layer3_outputs(3939) <= not b;
    layer3_outputs(3940) <= a;
    layer3_outputs(3941) <= '0';
    layer3_outputs(3942) <= not (a or b);
    layer3_outputs(3943) <= not a or b;
    layer3_outputs(3944) <= a;
    layer3_outputs(3945) <= b and not a;
    layer3_outputs(3946) <= a;
    layer3_outputs(3947) <= a and b;
    layer3_outputs(3948) <= not (a and b);
    layer3_outputs(3949) <= a xor b;
    layer3_outputs(3950) <= not b;
    layer3_outputs(3951) <= b;
    layer3_outputs(3952) <= not a;
    layer3_outputs(3953) <= not b;
    layer3_outputs(3954) <= not a;
    layer3_outputs(3955) <= not b;
    layer3_outputs(3956) <= not (a or b);
    layer3_outputs(3957) <= not a or b;
    layer3_outputs(3958) <= a xor b;
    layer3_outputs(3959) <= not (a or b);
    layer3_outputs(3960) <= not a;
    layer3_outputs(3961) <= a;
    layer3_outputs(3962) <= not (a and b);
    layer3_outputs(3963) <= not (a and b);
    layer3_outputs(3964) <= '0';
    layer3_outputs(3965) <= b;
    layer3_outputs(3966) <= not b or a;
    layer3_outputs(3967) <= a xor b;
    layer3_outputs(3968) <= b;
    layer3_outputs(3969) <= not (a and b);
    layer3_outputs(3970) <= b;
    layer3_outputs(3971) <= a and not b;
    layer3_outputs(3972) <= not a;
    layer3_outputs(3973) <= not a;
    layer3_outputs(3974) <= a or b;
    layer3_outputs(3975) <= b;
    layer3_outputs(3976) <= '1';
    layer3_outputs(3977) <= a;
    layer3_outputs(3978) <= not b;
    layer3_outputs(3979) <= not b;
    layer3_outputs(3980) <= '1';
    layer3_outputs(3981) <= a;
    layer3_outputs(3982) <= a and b;
    layer3_outputs(3983) <= a or b;
    layer3_outputs(3984) <= b;
    layer3_outputs(3985) <= not b;
    layer3_outputs(3986) <= a or b;
    layer3_outputs(3987) <= a;
    layer3_outputs(3988) <= not b;
    layer3_outputs(3989) <= not b or a;
    layer3_outputs(3990) <= b and not a;
    layer3_outputs(3991) <= not (a or b);
    layer3_outputs(3992) <= a and not b;
    layer3_outputs(3993) <= not (a and b);
    layer3_outputs(3994) <= '1';
    layer3_outputs(3995) <= a and not b;
    layer3_outputs(3996) <= a or b;
    layer3_outputs(3997) <= b;
    layer3_outputs(3998) <= b;
    layer3_outputs(3999) <= a xor b;
    layer3_outputs(4000) <= a;
    layer3_outputs(4001) <= not (a and b);
    layer3_outputs(4002) <= not (a xor b);
    layer3_outputs(4003) <= b;
    layer3_outputs(4004) <= b;
    layer3_outputs(4005) <= '0';
    layer3_outputs(4006) <= not a or b;
    layer3_outputs(4007) <= not (a xor b);
    layer3_outputs(4008) <= b;
    layer3_outputs(4009) <= not (a xor b);
    layer3_outputs(4010) <= a and not b;
    layer3_outputs(4011) <= a;
    layer3_outputs(4012) <= not (a or b);
    layer3_outputs(4013) <= b;
    layer3_outputs(4014) <= not (a or b);
    layer3_outputs(4015) <= not b or a;
    layer3_outputs(4016) <= a;
    layer3_outputs(4017) <= not a;
    layer3_outputs(4018) <= '1';
    layer3_outputs(4019) <= '1';
    layer3_outputs(4020) <= a and b;
    layer3_outputs(4021) <= not (a and b);
    layer3_outputs(4022) <= a;
    layer3_outputs(4023) <= a or b;
    layer3_outputs(4024) <= b and not a;
    layer3_outputs(4025) <= not a;
    layer3_outputs(4026) <= a;
    layer3_outputs(4027) <= '0';
    layer3_outputs(4028) <= '0';
    layer3_outputs(4029) <= not a;
    layer3_outputs(4030) <= not (a and b);
    layer3_outputs(4031) <= b;
    layer3_outputs(4032) <= a;
    layer3_outputs(4033) <= a;
    layer3_outputs(4034) <= not b or a;
    layer3_outputs(4035) <= b and not a;
    layer3_outputs(4036) <= a;
    layer3_outputs(4037) <= not (a xor b);
    layer3_outputs(4038) <= a or b;
    layer3_outputs(4039) <= b;
    layer3_outputs(4040) <= b;
    layer3_outputs(4041) <= a and not b;
    layer3_outputs(4042) <= not b or a;
    layer3_outputs(4043) <= not a;
    layer3_outputs(4044) <= b and not a;
    layer3_outputs(4045) <= a xor b;
    layer3_outputs(4046) <= not b;
    layer3_outputs(4047) <= not (a or b);
    layer3_outputs(4048) <= '0';
    layer3_outputs(4049) <= not b or a;
    layer3_outputs(4050) <= b;
    layer3_outputs(4051) <= a and b;
    layer3_outputs(4052) <= not (a or b);
    layer3_outputs(4053) <= not (a xor b);
    layer3_outputs(4054) <= not a;
    layer3_outputs(4055) <= a;
    layer3_outputs(4056) <= not b;
    layer3_outputs(4057) <= not (a xor b);
    layer3_outputs(4058) <= not (a and b);
    layer3_outputs(4059) <= not (a and b);
    layer3_outputs(4060) <= '1';
    layer3_outputs(4061) <= a xor b;
    layer3_outputs(4062) <= not b;
    layer3_outputs(4063) <= not b;
    layer3_outputs(4064) <= b;
    layer3_outputs(4065) <= not b or a;
    layer3_outputs(4066) <= a;
    layer3_outputs(4067) <= not (a or b);
    layer3_outputs(4068) <= not b;
    layer3_outputs(4069) <= a;
    layer3_outputs(4070) <= '0';
    layer3_outputs(4071) <= a and b;
    layer3_outputs(4072) <= '0';
    layer3_outputs(4073) <= not (a and b);
    layer3_outputs(4074) <= a;
    layer3_outputs(4075) <= a;
    layer3_outputs(4076) <= not b or a;
    layer3_outputs(4077) <= a and b;
    layer3_outputs(4078) <= not (a and b);
    layer3_outputs(4079) <= b;
    layer3_outputs(4080) <= not a or b;
    layer3_outputs(4081) <= not b or a;
    layer3_outputs(4082) <= a and not b;
    layer3_outputs(4083) <= a or b;
    layer3_outputs(4084) <= not a;
    layer3_outputs(4085) <= not b or a;
    layer3_outputs(4086) <= a;
    layer3_outputs(4087) <= a and b;
    layer3_outputs(4088) <= not (a and b);
    layer3_outputs(4089) <= not b or a;
    layer3_outputs(4090) <= b and not a;
    layer3_outputs(4091) <= b;
    layer3_outputs(4092) <= b;
    layer3_outputs(4093) <= not b;
    layer3_outputs(4094) <= '0';
    layer3_outputs(4095) <= not (a and b);
    layer3_outputs(4096) <= '1';
    layer3_outputs(4097) <= not a or b;
    layer3_outputs(4098) <= not a or b;
    layer3_outputs(4099) <= not b;
    layer3_outputs(4100) <= not b;
    layer3_outputs(4101) <= not b;
    layer3_outputs(4102) <= not a;
    layer3_outputs(4103) <= a or b;
    layer3_outputs(4104) <= not a or b;
    layer3_outputs(4105) <= a xor b;
    layer3_outputs(4106) <= a;
    layer3_outputs(4107) <= not a;
    layer3_outputs(4108) <= not (a and b);
    layer3_outputs(4109) <= not a or b;
    layer3_outputs(4110) <= not b;
    layer3_outputs(4111) <= not (a or b);
    layer3_outputs(4112) <= a xor b;
    layer3_outputs(4113) <= a xor b;
    layer3_outputs(4114) <= a and b;
    layer3_outputs(4115) <= not (a xor b);
    layer3_outputs(4116) <= not b or a;
    layer3_outputs(4117) <= a and not b;
    layer3_outputs(4118) <= not b or a;
    layer3_outputs(4119) <= not b;
    layer3_outputs(4120) <= a and b;
    layer3_outputs(4121) <= not b or a;
    layer3_outputs(4122) <= not a;
    layer3_outputs(4123) <= b;
    layer3_outputs(4124) <= a and not b;
    layer3_outputs(4125) <= a xor b;
    layer3_outputs(4126) <= b and not a;
    layer3_outputs(4127) <= not a or b;
    layer3_outputs(4128) <= not a;
    layer3_outputs(4129) <= a and not b;
    layer3_outputs(4130) <= not a or b;
    layer3_outputs(4131) <= not b;
    layer3_outputs(4132) <= a;
    layer3_outputs(4133) <= b and not a;
    layer3_outputs(4134) <= not b;
    layer3_outputs(4135) <= '0';
    layer3_outputs(4136) <= b and not a;
    layer3_outputs(4137) <= not (a and b);
    layer3_outputs(4138) <= not a or b;
    layer3_outputs(4139) <= not b or a;
    layer3_outputs(4140) <= b and not a;
    layer3_outputs(4141) <= not a or b;
    layer3_outputs(4142) <= a xor b;
    layer3_outputs(4143) <= a;
    layer3_outputs(4144) <= not a or b;
    layer3_outputs(4145) <= not (a or b);
    layer3_outputs(4146) <= a and b;
    layer3_outputs(4147) <= not (a or b);
    layer3_outputs(4148) <= not a or b;
    layer3_outputs(4149) <= not b;
    layer3_outputs(4150) <= not a;
    layer3_outputs(4151) <= not a;
    layer3_outputs(4152) <= not b;
    layer3_outputs(4153) <= a;
    layer3_outputs(4154) <= a xor b;
    layer3_outputs(4155) <= not a or b;
    layer3_outputs(4156) <= not (a and b);
    layer3_outputs(4157) <= b and not a;
    layer3_outputs(4158) <= not (a xor b);
    layer3_outputs(4159) <= a and not b;
    layer3_outputs(4160) <= a or b;
    layer3_outputs(4161) <= not (a or b);
    layer3_outputs(4162) <= not (a and b);
    layer3_outputs(4163) <= b and not a;
    layer3_outputs(4164) <= not b or a;
    layer3_outputs(4165) <= a and b;
    layer3_outputs(4166) <= not a or b;
    layer3_outputs(4167) <= '0';
    layer3_outputs(4168) <= not (a or b);
    layer3_outputs(4169) <= not (a or b);
    layer3_outputs(4170) <= not (a xor b);
    layer3_outputs(4171) <= a and not b;
    layer3_outputs(4172) <= not (a and b);
    layer3_outputs(4173) <= not b;
    layer3_outputs(4174) <= b;
    layer3_outputs(4175) <= not b or a;
    layer3_outputs(4176) <= b and not a;
    layer3_outputs(4177) <= not a;
    layer3_outputs(4178) <= not a;
    layer3_outputs(4179) <= b;
    layer3_outputs(4180) <= not b or a;
    layer3_outputs(4181) <= not (a and b);
    layer3_outputs(4182) <= not b or a;
    layer3_outputs(4183) <= a and b;
    layer3_outputs(4184) <= '0';
    layer3_outputs(4185) <= b;
    layer3_outputs(4186) <= '0';
    layer3_outputs(4187) <= not b;
    layer3_outputs(4188) <= not a;
    layer3_outputs(4189) <= b;
    layer3_outputs(4190) <= not b;
    layer3_outputs(4191) <= not b;
    layer3_outputs(4192) <= not a or b;
    layer3_outputs(4193) <= a and not b;
    layer3_outputs(4194) <= not b;
    layer3_outputs(4195) <= b;
    layer3_outputs(4196) <= not (a or b);
    layer3_outputs(4197) <= not a;
    layer3_outputs(4198) <= not a;
    layer3_outputs(4199) <= a;
    layer3_outputs(4200) <= a;
    layer3_outputs(4201) <= not (a and b);
    layer3_outputs(4202) <= b;
    layer3_outputs(4203) <= not a;
    layer3_outputs(4204) <= not a;
    layer3_outputs(4205) <= not b;
    layer3_outputs(4206) <= a and not b;
    layer3_outputs(4207) <= not (a xor b);
    layer3_outputs(4208) <= b and not a;
    layer3_outputs(4209) <= not a;
    layer3_outputs(4210) <= a;
    layer3_outputs(4211) <= b;
    layer3_outputs(4212) <= a and not b;
    layer3_outputs(4213) <= b and not a;
    layer3_outputs(4214) <= '0';
    layer3_outputs(4215) <= a or b;
    layer3_outputs(4216) <= not b or a;
    layer3_outputs(4217) <= not b or a;
    layer3_outputs(4218) <= not a;
    layer3_outputs(4219) <= a and not b;
    layer3_outputs(4220) <= '1';
    layer3_outputs(4221) <= not a or b;
    layer3_outputs(4222) <= not a or b;
    layer3_outputs(4223) <= a;
    layer3_outputs(4224) <= not b or a;
    layer3_outputs(4225) <= not a;
    layer3_outputs(4226) <= not (a xor b);
    layer3_outputs(4227) <= b;
    layer3_outputs(4228) <= not b or a;
    layer3_outputs(4229) <= not a or b;
    layer3_outputs(4230) <= '1';
    layer3_outputs(4231) <= not a or b;
    layer3_outputs(4232) <= a and b;
    layer3_outputs(4233) <= a or b;
    layer3_outputs(4234) <= a;
    layer3_outputs(4235) <= not b;
    layer3_outputs(4236) <= not (a and b);
    layer3_outputs(4237) <= not b or a;
    layer3_outputs(4238) <= a or b;
    layer3_outputs(4239) <= '1';
    layer3_outputs(4240) <= not a;
    layer3_outputs(4241) <= a;
    layer3_outputs(4242) <= b and not a;
    layer3_outputs(4243) <= not b or a;
    layer3_outputs(4244) <= not (a xor b);
    layer3_outputs(4245) <= b and not a;
    layer3_outputs(4246) <= a and not b;
    layer3_outputs(4247) <= a and not b;
    layer3_outputs(4248) <= not (a xor b);
    layer3_outputs(4249) <= a and b;
    layer3_outputs(4250) <= a;
    layer3_outputs(4251) <= not b;
    layer3_outputs(4252) <= '1';
    layer3_outputs(4253) <= '0';
    layer3_outputs(4254) <= not a;
    layer3_outputs(4255) <= not (a xor b);
    layer3_outputs(4256) <= not a;
    layer3_outputs(4257) <= a and not b;
    layer3_outputs(4258) <= not (a or b);
    layer3_outputs(4259) <= not b or a;
    layer3_outputs(4260) <= a;
    layer3_outputs(4261) <= not (a xor b);
    layer3_outputs(4262) <= a and not b;
    layer3_outputs(4263) <= a xor b;
    layer3_outputs(4264) <= not b or a;
    layer3_outputs(4265) <= not (a and b);
    layer3_outputs(4266) <= not (a xor b);
    layer3_outputs(4267) <= '1';
    layer3_outputs(4268) <= not (a or b);
    layer3_outputs(4269) <= a xor b;
    layer3_outputs(4270) <= b;
    layer3_outputs(4271) <= a;
    layer3_outputs(4272) <= a xor b;
    layer3_outputs(4273) <= b;
    layer3_outputs(4274) <= a;
    layer3_outputs(4275) <= '0';
    layer3_outputs(4276) <= a xor b;
    layer3_outputs(4277) <= '1';
    layer3_outputs(4278) <= a;
    layer3_outputs(4279) <= a and b;
    layer3_outputs(4280) <= not a;
    layer3_outputs(4281) <= not a;
    layer3_outputs(4282) <= b;
    layer3_outputs(4283) <= a;
    layer3_outputs(4284) <= '0';
    layer3_outputs(4285) <= not a;
    layer3_outputs(4286) <= b and not a;
    layer3_outputs(4287) <= b and not a;
    layer3_outputs(4288) <= a;
    layer3_outputs(4289) <= not b;
    layer3_outputs(4290) <= not b;
    layer3_outputs(4291) <= not a;
    layer3_outputs(4292) <= not (a or b);
    layer3_outputs(4293) <= not a;
    layer3_outputs(4294) <= a or b;
    layer3_outputs(4295) <= a;
    layer3_outputs(4296) <= a and not b;
    layer3_outputs(4297) <= '0';
    layer3_outputs(4298) <= not a;
    layer3_outputs(4299) <= '1';
    layer3_outputs(4300) <= not b;
    layer3_outputs(4301) <= '0';
    layer3_outputs(4302) <= not (a and b);
    layer3_outputs(4303) <= a;
    layer3_outputs(4304) <= not b or a;
    layer3_outputs(4305) <= not (a or b);
    layer3_outputs(4306) <= not b or a;
    layer3_outputs(4307) <= not (a and b);
    layer3_outputs(4308) <= not a or b;
    layer3_outputs(4309) <= b;
    layer3_outputs(4310) <= '0';
    layer3_outputs(4311) <= a and not b;
    layer3_outputs(4312) <= a and not b;
    layer3_outputs(4313) <= '1';
    layer3_outputs(4314) <= a;
    layer3_outputs(4315) <= not b;
    layer3_outputs(4316) <= b and not a;
    layer3_outputs(4317) <= '1';
    layer3_outputs(4318) <= a and b;
    layer3_outputs(4319) <= a and not b;
    layer3_outputs(4320) <= a xor b;
    layer3_outputs(4321) <= not a;
    layer3_outputs(4322) <= not a or b;
    layer3_outputs(4323) <= a or b;
    layer3_outputs(4324) <= a and b;
    layer3_outputs(4325) <= a and not b;
    layer3_outputs(4326) <= not b;
    layer3_outputs(4327) <= a;
    layer3_outputs(4328) <= a and not b;
    layer3_outputs(4329) <= '1';
    layer3_outputs(4330) <= not b;
    layer3_outputs(4331) <= not b or a;
    layer3_outputs(4332) <= b;
    layer3_outputs(4333) <= not b or a;
    layer3_outputs(4334) <= not b or a;
    layer3_outputs(4335) <= a xor b;
    layer3_outputs(4336) <= '1';
    layer3_outputs(4337) <= not (a or b);
    layer3_outputs(4338) <= not (a or b);
    layer3_outputs(4339) <= b;
    layer3_outputs(4340) <= not (a and b);
    layer3_outputs(4341) <= a;
    layer3_outputs(4342) <= not (a and b);
    layer3_outputs(4343) <= a;
    layer3_outputs(4344) <= not a;
    layer3_outputs(4345) <= not a or b;
    layer3_outputs(4346) <= a and not b;
    layer3_outputs(4347) <= not b;
    layer3_outputs(4348) <= a;
    layer3_outputs(4349) <= not a;
    layer3_outputs(4350) <= not b;
    layer3_outputs(4351) <= not b or a;
    layer3_outputs(4352) <= a;
    layer3_outputs(4353) <= not (a and b);
    layer3_outputs(4354) <= a xor b;
    layer3_outputs(4355) <= not (a or b);
    layer3_outputs(4356) <= not a or b;
    layer3_outputs(4357) <= b and not a;
    layer3_outputs(4358) <= not a or b;
    layer3_outputs(4359) <= not a or b;
    layer3_outputs(4360) <= not b or a;
    layer3_outputs(4361) <= not b;
    layer3_outputs(4362) <= b and not a;
    layer3_outputs(4363) <= not (a or b);
    layer3_outputs(4364) <= a and b;
    layer3_outputs(4365) <= not b;
    layer3_outputs(4366) <= not (a and b);
    layer3_outputs(4367) <= not (a or b);
    layer3_outputs(4368) <= not a;
    layer3_outputs(4369) <= not b;
    layer3_outputs(4370) <= '0';
    layer3_outputs(4371) <= '1';
    layer3_outputs(4372) <= b and not a;
    layer3_outputs(4373) <= a;
    layer3_outputs(4374) <= not (a xor b);
    layer3_outputs(4375) <= a or b;
    layer3_outputs(4376) <= a or b;
    layer3_outputs(4377) <= a and b;
    layer3_outputs(4378) <= not a;
    layer3_outputs(4379) <= not (a xor b);
    layer3_outputs(4380) <= a and not b;
    layer3_outputs(4381) <= a;
    layer3_outputs(4382) <= a;
    layer3_outputs(4383) <= a or b;
    layer3_outputs(4384) <= a or b;
    layer3_outputs(4385) <= not (a or b);
    layer3_outputs(4386) <= a;
    layer3_outputs(4387) <= not a or b;
    layer3_outputs(4388) <= not (a and b);
    layer3_outputs(4389) <= '0';
    layer3_outputs(4390) <= not a;
    layer3_outputs(4391) <= a and b;
    layer3_outputs(4392) <= a;
    layer3_outputs(4393) <= '0';
    layer3_outputs(4394) <= a and b;
    layer3_outputs(4395) <= not b;
    layer3_outputs(4396) <= a;
    layer3_outputs(4397) <= not b;
    layer3_outputs(4398) <= a;
    layer3_outputs(4399) <= '0';
    layer3_outputs(4400) <= not a or b;
    layer3_outputs(4401) <= a;
    layer3_outputs(4402) <= b;
    layer3_outputs(4403) <= not (a and b);
    layer3_outputs(4404) <= b and not a;
    layer3_outputs(4405) <= not (a and b);
    layer3_outputs(4406) <= not a or b;
    layer3_outputs(4407) <= a and not b;
    layer3_outputs(4408) <= a or b;
    layer3_outputs(4409) <= b and not a;
    layer3_outputs(4410) <= a and not b;
    layer3_outputs(4411) <= a;
    layer3_outputs(4412) <= not a;
    layer3_outputs(4413) <= b and not a;
    layer3_outputs(4414) <= a or b;
    layer3_outputs(4415) <= not (a or b);
    layer3_outputs(4416) <= not b;
    layer3_outputs(4417) <= b;
    layer3_outputs(4418) <= not a;
    layer3_outputs(4419) <= b;
    layer3_outputs(4420) <= a;
    layer3_outputs(4421) <= b;
    layer3_outputs(4422) <= b;
    layer3_outputs(4423) <= '0';
    layer3_outputs(4424) <= b;
    layer3_outputs(4425) <= not (a or b);
    layer3_outputs(4426) <= a;
    layer3_outputs(4427) <= not b;
    layer3_outputs(4428) <= not b or a;
    layer3_outputs(4429) <= a or b;
    layer3_outputs(4430) <= not b or a;
    layer3_outputs(4431) <= not a;
    layer3_outputs(4432) <= not a;
    layer3_outputs(4433) <= a xor b;
    layer3_outputs(4434) <= not b;
    layer3_outputs(4435) <= b;
    layer3_outputs(4436) <= a and b;
    layer3_outputs(4437) <= not b;
    layer3_outputs(4438) <= not (a or b);
    layer3_outputs(4439) <= not a;
    layer3_outputs(4440) <= not (a or b);
    layer3_outputs(4441) <= b;
    layer3_outputs(4442) <= b and not a;
    layer3_outputs(4443) <= a and b;
    layer3_outputs(4444) <= not (a xor b);
    layer3_outputs(4445) <= not (a and b);
    layer3_outputs(4446) <= b;
    layer3_outputs(4447) <= b and not a;
    layer3_outputs(4448) <= a xor b;
    layer3_outputs(4449) <= not a;
    layer3_outputs(4450) <= not a or b;
    layer3_outputs(4451) <= a;
    layer3_outputs(4452) <= not a;
    layer3_outputs(4453) <= not a;
    layer3_outputs(4454) <= a or b;
    layer3_outputs(4455) <= b;
    layer3_outputs(4456) <= not b;
    layer3_outputs(4457) <= a;
    layer3_outputs(4458) <= b;
    layer3_outputs(4459) <= b and not a;
    layer3_outputs(4460) <= a and b;
    layer3_outputs(4461) <= a and b;
    layer3_outputs(4462) <= b;
    layer3_outputs(4463) <= b;
    layer3_outputs(4464) <= not (a and b);
    layer3_outputs(4465) <= a and b;
    layer3_outputs(4466) <= a xor b;
    layer3_outputs(4467) <= a;
    layer3_outputs(4468) <= '1';
    layer3_outputs(4469) <= not a or b;
    layer3_outputs(4470) <= b and not a;
    layer3_outputs(4471) <= not b;
    layer3_outputs(4472) <= not (a or b);
    layer3_outputs(4473) <= not b or a;
    layer3_outputs(4474) <= a;
    layer3_outputs(4475) <= a xor b;
    layer3_outputs(4476) <= a;
    layer3_outputs(4477) <= not (a and b);
    layer3_outputs(4478) <= a and b;
    layer3_outputs(4479) <= b;
    layer3_outputs(4480) <= a;
    layer3_outputs(4481) <= not a;
    layer3_outputs(4482) <= a;
    layer3_outputs(4483) <= b;
    layer3_outputs(4484) <= not (a or b);
    layer3_outputs(4485) <= b;
    layer3_outputs(4486) <= b;
    layer3_outputs(4487) <= b and not a;
    layer3_outputs(4488) <= a;
    layer3_outputs(4489) <= not b;
    layer3_outputs(4490) <= not a;
    layer3_outputs(4491) <= a and b;
    layer3_outputs(4492) <= b;
    layer3_outputs(4493) <= not b or a;
    layer3_outputs(4494) <= not a or b;
    layer3_outputs(4495) <= not b;
    layer3_outputs(4496) <= not (a and b);
    layer3_outputs(4497) <= not (a xor b);
    layer3_outputs(4498) <= a;
    layer3_outputs(4499) <= a or b;
    layer3_outputs(4500) <= not a;
    layer3_outputs(4501) <= b;
    layer3_outputs(4502) <= not b or a;
    layer3_outputs(4503) <= not (a or b);
    layer3_outputs(4504) <= a;
    layer3_outputs(4505) <= not a;
    layer3_outputs(4506) <= not (a and b);
    layer3_outputs(4507) <= a or b;
    layer3_outputs(4508) <= b and not a;
    layer3_outputs(4509) <= not b or a;
    layer3_outputs(4510) <= a and b;
    layer3_outputs(4511) <= '1';
    layer3_outputs(4512) <= not b;
    layer3_outputs(4513) <= '0';
    layer3_outputs(4514) <= a and not b;
    layer3_outputs(4515) <= not (a and b);
    layer3_outputs(4516) <= a and b;
    layer3_outputs(4517) <= not (a and b);
    layer3_outputs(4518) <= not (a and b);
    layer3_outputs(4519) <= a;
    layer3_outputs(4520) <= '1';
    layer3_outputs(4521) <= a and not b;
    layer3_outputs(4522) <= a xor b;
    layer3_outputs(4523) <= not (a or b);
    layer3_outputs(4524) <= not b or a;
    layer3_outputs(4525) <= a xor b;
    layer3_outputs(4526) <= a and b;
    layer3_outputs(4527) <= not (a or b);
    layer3_outputs(4528) <= a or b;
    layer3_outputs(4529) <= '1';
    layer3_outputs(4530) <= '1';
    layer3_outputs(4531) <= '1';
    layer3_outputs(4532) <= a and b;
    layer3_outputs(4533) <= a and b;
    layer3_outputs(4534) <= b;
    layer3_outputs(4535) <= '1';
    layer3_outputs(4536) <= b and not a;
    layer3_outputs(4537) <= b and not a;
    layer3_outputs(4538) <= not b;
    layer3_outputs(4539) <= not (a or b);
    layer3_outputs(4540) <= a xor b;
    layer3_outputs(4541) <= not b;
    layer3_outputs(4542) <= a or b;
    layer3_outputs(4543) <= not (a or b);
    layer3_outputs(4544) <= not b or a;
    layer3_outputs(4545) <= a and not b;
    layer3_outputs(4546) <= not a;
    layer3_outputs(4547) <= not b;
    layer3_outputs(4548) <= b and not a;
    layer3_outputs(4549) <= a or b;
    layer3_outputs(4550) <= not b;
    layer3_outputs(4551) <= b;
    layer3_outputs(4552) <= not a;
    layer3_outputs(4553) <= a and b;
    layer3_outputs(4554) <= not (a or b);
    layer3_outputs(4555) <= a or b;
    layer3_outputs(4556) <= a;
    layer3_outputs(4557) <= a;
    layer3_outputs(4558) <= b and not a;
    layer3_outputs(4559) <= '0';
    layer3_outputs(4560) <= not a;
    layer3_outputs(4561) <= not b or a;
    layer3_outputs(4562) <= not (a or b);
    layer3_outputs(4563) <= b and not a;
    layer3_outputs(4564) <= not a or b;
    layer3_outputs(4565) <= '0';
    layer3_outputs(4566) <= not a or b;
    layer3_outputs(4567) <= a and not b;
    layer3_outputs(4568) <= a;
    layer3_outputs(4569) <= b and not a;
    layer3_outputs(4570) <= b and not a;
    layer3_outputs(4571) <= a and b;
    layer3_outputs(4572) <= a;
    layer3_outputs(4573) <= not (a and b);
    layer3_outputs(4574) <= not (a or b);
    layer3_outputs(4575) <= not a or b;
    layer3_outputs(4576) <= not a or b;
    layer3_outputs(4577) <= not (a or b);
    layer3_outputs(4578) <= a and not b;
    layer3_outputs(4579) <= not b or a;
    layer3_outputs(4580) <= b and not a;
    layer3_outputs(4581) <= b and not a;
    layer3_outputs(4582) <= a and not b;
    layer3_outputs(4583) <= b;
    layer3_outputs(4584) <= a;
    layer3_outputs(4585) <= a;
    layer3_outputs(4586) <= not b or a;
    layer3_outputs(4587) <= not b;
    layer3_outputs(4588) <= not a;
    layer3_outputs(4589) <= not a;
    layer3_outputs(4590) <= not (a and b);
    layer3_outputs(4591) <= a;
    layer3_outputs(4592) <= not (a or b);
    layer3_outputs(4593) <= a;
    layer3_outputs(4594) <= a and not b;
    layer3_outputs(4595) <= b;
    layer3_outputs(4596) <= a;
    layer3_outputs(4597) <= not (a and b);
    layer3_outputs(4598) <= '1';
    layer3_outputs(4599) <= b and not a;
    layer3_outputs(4600) <= '0';
    layer3_outputs(4601) <= not (a and b);
    layer3_outputs(4602) <= not a or b;
    layer3_outputs(4603) <= b;
    layer3_outputs(4604) <= b;
    layer3_outputs(4605) <= not b;
    layer3_outputs(4606) <= not (a xor b);
    layer3_outputs(4607) <= b;
    layer3_outputs(4608) <= a;
    layer3_outputs(4609) <= not (a xor b);
    layer3_outputs(4610) <= a and b;
    layer3_outputs(4611) <= a and b;
    layer3_outputs(4612) <= a or b;
    layer3_outputs(4613) <= a and b;
    layer3_outputs(4614) <= a and not b;
    layer3_outputs(4615) <= a;
    layer3_outputs(4616) <= '0';
    layer3_outputs(4617) <= a and not b;
    layer3_outputs(4618) <= '1';
    layer3_outputs(4619) <= a and b;
    layer3_outputs(4620) <= not (a or b);
    layer3_outputs(4621) <= a and b;
    layer3_outputs(4622) <= not a;
    layer3_outputs(4623) <= not (a and b);
    layer3_outputs(4624) <= not a or b;
    layer3_outputs(4625) <= not (a xor b);
    layer3_outputs(4626) <= a or b;
    layer3_outputs(4627) <= not b or a;
    layer3_outputs(4628) <= a and b;
    layer3_outputs(4629) <= not (a and b);
    layer3_outputs(4630) <= b and not a;
    layer3_outputs(4631) <= b and not a;
    layer3_outputs(4632) <= not (a or b);
    layer3_outputs(4633) <= not a;
    layer3_outputs(4634) <= not b;
    layer3_outputs(4635) <= b;
    layer3_outputs(4636) <= not (a or b);
    layer3_outputs(4637) <= b and not a;
    layer3_outputs(4638) <= not (a or b);
    layer3_outputs(4639) <= not (a or b);
    layer3_outputs(4640) <= not b;
    layer3_outputs(4641) <= not (a xor b);
    layer3_outputs(4642) <= b and not a;
    layer3_outputs(4643) <= a xor b;
    layer3_outputs(4644) <= b;
    layer3_outputs(4645) <= not (a or b);
    layer3_outputs(4646) <= a;
    layer3_outputs(4647) <= not a or b;
    layer3_outputs(4648) <= b;
    layer3_outputs(4649) <= a and b;
    layer3_outputs(4650) <= b;
    layer3_outputs(4651) <= '1';
    layer3_outputs(4652) <= a or b;
    layer3_outputs(4653) <= a xor b;
    layer3_outputs(4654) <= not a;
    layer3_outputs(4655) <= a and b;
    layer3_outputs(4656) <= a xor b;
    layer3_outputs(4657) <= a or b;
    layer3_outputs(4658) <= not b or a;
    layer3_outputs(4659) <= a;
    layer3_outputs(4660) <= not (a xor b);
    layer3_outputs(4661) <= a;
    layer3_outputs(4662) <= not (a or b);
    layer3_outputs(4663) <= not b;
    layer3_outputs(4664) <= not a or b;
    layer3_outputs(4665) <= b and not a;
    layer3_outputs(4666) <= not b;
    layer3_outputs(4667) <= not b or a;
    layer3_outputs(4668) <= not a;
    layer3_outputs(4669) <= not a or b;
    layer3_outputs(4670) <= a and b;
    layer3_outputs(4671) <= not b or a;
    layer3_outputs(4672) <= b;
    layer3_outputs(4673) <= not (a and b);
    layer3_outputs(4674) <= not b or a;
    layer3_outputs(4675) <= not a or b;
    layer3_outputs(4676) <= not a or b;
    layer3_outputs(4677) <= a or b;
    layer3_outputs(4678) <= '1';
    layer3_outputs(4679) <= not a;
    layer3_outputs(4680) <= a xor b;
    layer3_outputs(4681) <= not (a xor b);
    layer3_outputs(4682) <= not (a or b);
    layer3_outputs(4683) <= not a or b;
    layer3_outputs(4684) <= not a;
    layer3_outputs(4685) <= a;
    layer3_outputs(4686) <= not b;
    layer3_outputs(4687) <= a or b;
    layer3_outputs(4688) <= not a or b;
    layer3_outputs(4689) <= b and not a;
    layer3_outputs(4690) <= b and not a;
    layer3_outputs(4691) <= b;
    layer3_outputs(4692) <= not b or a;
    layer3_outputs(4693) <= a xor b;
    layer3_outputs(4694) <= not (a xor b);
    layer3_outputs(4695) <= a or b;
    layer3_outputs(4696) <= not a;
    layer3_outputs(4697) <= '0';
    layer3_outputs(4698) <= a;
    layer3_outputs(4699) <= '1';
    layer3_outputs(4700) <= b;
    layer3_outputs(4701) <= not b or a;
    layer3_outputs(4702) <= not b;
    layer3_outputs(4703) <= a;
    layer3_outputs(4704) <= a and not b;
    layer3_outputs(4705) <= not (a or b);
    layer3_outputs(4706) <= a and b;
    layer3_outputs(4707) <= a and not b;
    layer3_outputs(4708) <= a xor b;
    layer3_outputs(4709) <= '0';
    layer3_outputs(4710) <= a and not b;
    layer3_outputs(4711) <= a;
    layer3_outputs(4712) <= not a or b;
    layer3_outputs(4713) <= not b;
    layer3_outputs(4714) <= not a;
    layer3_outputs(4715) <= a or b;
    layer3_outputs(4716) <= not (a and b);
    layer3_outputs(4717) <= a;
    layer3_outputs(4718) <= a xor b;
    layer3_outputs(4719) <= a and b;
    layer3_outputs(4720) <= not b or a;
    layer3_outputs(4721) <= '1';
    layer3_outputs(4722) <= '0';
    layer3_outputs(4723) <= '1';
    layer3_outputs(4724) <= not a;
    layer3_outputs(4725) <= a;
    layer3_outputs(4726) <= not (a or b);
    layer3_outputs(4727) <= not b;
    layer3_outputs(4728) <= a and b;
    layer3_outputs(4729) <= a and b;
    layer3_outputs(4730) <= a xor b;
    layer3_outputs(4731) <= a and not b;
    layer3_outputs(4732) <= a;
    layer3_outputs(4733) <= not a or b;
    layer3_outputs(4734) <= not (a or b);
    layer3_outputs(4735) <= not b;
    layer3_outputs(4736) <= b and not a;
    layer3_outputs(4737) <= not b;
    layer3_outputs(4738) <= b and not a;
    layer3_outputs(4739) <= a;
    layer3_outputs(4740) <= not a or b;
    layer3_outputs(4741) <= not a;
    layer3_outputs(4742) <= a and b;
    layer3_outputs(4743) <= not b;
    layer3_outputs(4744) <= a or b;
    layer3_outputs(4745) <= b and not a;
    layer3_outputs(4746) <= not (a and b);
    layer3_outputs(4747) <= not b;
    layer3_outputs(4748) <= not (a and b);
    layer3_outputs(4749) <= not a;
    layer3_outputs(4750) <= b;
    layer3_outputs(4751) <= a and not b;
    layer3_outputs(4752) <= not a or b;
    layer3_outputs(4753) <= not (a xor b);
    layer3_outputs(4754) <= a and b;
    layer3_outputs(4755) <= not b;
    layer3_outputs(4756) <= '0';
    layer3_outputs(4757) <= not a;
    layer3_outputs(4758) <= '0';
    layer3_outputs(4759) <= a;
    layer3_outputs(4760) <= not b or a;
    layer3_outputs(4761) <= a;
    layer3_outputs(4762) <= not a or b;
    layer3_outputs(4763) <= a and b;
    layer3_outputs(4764) <= not a;
    layer3_outputs(4765) <= not (a and b);
    layer3_outputs(4766) <= '1';
    layer3_outputs(4767) <= not b;
    layer3_outputs(4768) <= b and not a;
    layer3_outputs(4769) <= not (a and b);
    layer3_outputs(4770) <= a xor b;
    layer3_outputs(4771) <= a xor b;
    layer3_outputs(4772) <= a or b;
    layer3_outputs(4773) <= '0';
    layer3_outputs(4774) <= b and not a;
    layer3_outputs(4775) <= not a or b;
    layer3_outputs(4776) <= not b or a;
    layer3_outputs(4777) <= a and b;
    layer3_outputs(4778) <= not (a xor b);
    layer3_outputs(4779) <= not (a or b);
    layer3_outputs(4780) <= b;
    layer3_outputs(4781) <= not a;
    layer3_outputs(4782) <= '0';
    layer3_outputs(4783) <= not b;
    layer3_outputs(4784) <= not b or a;
    layer3_outputs(4785) <= a xor b;
    layer3_outputs(4786) <= a;
    layer3_outputs(4787) <= a xor b;
    layer3_outputs(4788) <= not a or b;
    layer3_outputs(4789) <= not (a and b);
    layer3_outputs(4790) <= not (a or b);
    layer3_outputs(4791) <= not (a or b);
    layer3_outputs(4792) <= a and not b;
    layer3_outputs(4793) <= a and b;
    layer3_outputs(4794) <= not b;
    layer3_outputs(4795) <= a and b;
    layer3_outputs(4796) <= a or b;
    layer3_outputs(4797) <= a;
    layer3_outputs(4798) <= not a;
    layer3_outputs(4799) <= not a;
    layer3_outputs(4800) <= not a or b;
    layer3_outputs(4801) <= a and not b;
    layer3_outputs(4802) <= b;
    layer3_outputs(4803) <= not (a and b);
    layer3_outputs(4804) <= '1';
    layer3_outputs(4805) <= '1';
    layer3_outputs(4806) <= b;
    layer3_outputs(4807) <= a and not b;
    layer3_outputs(4808) <= a;
    layer3_outputs(4809) <= not b or a;
    layer3_outputs(4810) <= not (a xor b);
    layer3_outputs(4811) <= a xor b;
    layer3_outputs(4812) <= b and not a;
    layer3_outputs(4813) <= a;
    layer3_outputs(4814) <= a;
    layer3_outputs(4815) <= b;
    layer3_outputs(4816) <= not a;
    layer3_outputs(4817) <= a and not b;
    layer3_outputs(4818) <= a;
    layer3_outputs(4819) <= a and b;
    layer3_outputs(4820) <= not (a or b);
    layer3_outputs(4821) <= not b or a;
    layer3_outputs(4822) <= a;
    layer3_outputs(4823) <= b;
    layer3_outputs(4824) <= a;
    layer3_outputs(4825) <= a and b;
    layer3_outputs(4826) <= b;
    layer3_outputs(4827) <= a or b;
    layer3_outputs(4828) <= '0';
    layer3_outputs(4829) <= a;
    layer3_outputs(4830) <= a and b;
    layer3_outputs(4831) <= '0';
    layer3_outputs(4832) <= '0';
    layer3_outputs(4833) <= not a;
    layer3_outputs(4834) <= a or b;
    layer3_outputs(4835) <= '0';
    layer3_outputs(4836) <= b;
    layer3_outputs(4837) <= not (a xor b);
    layer3_outputs(4838) <= b;
    layer3_outputs(4839) <= b and not a;
    layer3_outputs(4840) <= not b;
    layer3_outputs(4841) <= not a;
    layer3_outputs(4842) <= a and not b;
    layer3_outputs(4843) <= a;
    layer3_outputs(4844) <= b and not a;
    layer3_outputs(4845) <= a xor b;
    layer3_outputs(4846) <= not (a or b);
    layer3_outputs(4847) <= not (a xor b);
    layer3_outputs(4848) <= not (a and b);
    layer3_outputs(4849) <= a or b;
    layer3_outputs(4850) <= a xor b;
    layer3_outputs(4851) <= not b or a;
    layer3_outputs(4852) <= b;
    layer3_outputs(4853) <= not a;
    layer3_outputs(4854) <= a and not b;
    layer3_outputs(4855) <= '1';
    layer3_outputs(4856) <= a;
    layer3_outputs(4857) <= a and b;
    layer3_outputs(4858) <= not (a or b);
    layer3_outputs(4859) <= not b;
    layer3_outputs(4860) <= b;
    layer3_outputs(4861) <= a;
    layer3_outputs(4862) <= not (a or b);
    layer3_outputs(4863) <= a and b;
    layer3_outputs(4864) <= not a;
    layer3_outputs(4865) <= not (a and b);
    layer3_outputs(4866) <= '0';
    layer3_outputs(4867) <= '1';
    layer3_outputs(4868) <= not (a or b);
    layer3_outputs(4869) <= not a;
    layer3_outputs(4870) <= '0';
    layer3_outputs(4871) <= a and not b;
    layer3_outputs(4872) <= not a;
    layer3_outputs(4873) <= a;
    layer3_outputs(4874) <= not b;
    layer3_outputs(4875) <= '1';
    layer3_outputs(4876) <= a or b;
    layer3_outputs(4877) <= not (a and b);
    layer3_outputs(4878) <= b;
    layer3_outputs(4879) <= not (a and b);
    layer3_outputs(4880) <= a;
    layer3_outputs(4881) <= '0';
    layer3_outputs(4882) <= '1';
    layer3_outputs(4883) <= a and b;
    layer3_outputs(4884) <= not b;
    layer3_outputs(4885) <= not a;
    layer3_outputs(4886) <= a xor b;
    layer3_outputs(4887) <= b and not a;
    layer3_outputs(4888) <= a xor b;
    layer3_outputs(4889) <= not b or a;
    layer3_outputs(4890) <= a;
    layer3_outputs(4891) <= b and not a;
    layer3_outputs(4892) <= not b;
    layer3_outputs(4893) <= not b;
    layer3_outputs(4894) <= not (a xor b);
    layer3_outputs(4895) <= a and b;
    layer3_outputs(4896) <= not a;
    layer3_outputs(4897) <= not (a xor b);
    layer3_outputs(4898) <= b and not a;
    layer3_outputs(4899) <= b;
    layer3_outputs(4900) <= a;
    layer3_outputs(4901) <= a and not b;
    layer3_outputs(4902) <= not a;
    layer3_outputs(4903) <= b;
    layer3_outputs(4904) <= a xor b;
    layer3_outputs(4905) <= not (a and b);
    layer3_outputs(4906) <= b;
    layer3_outputs(4907) <= a xor b;
    layer3_outputs(4908) <= not (a xor b);
    layer3_outputs(4909) <= a;
    layer3_outputs(4910) <= '1';
    layer3_outputs(4911) <= b and not a;
    layer3_outputs(4912) <= a or b;
    layer3_outputs(4913) <= a xor b;
    layer3_outputs(4914) <= b;
    layer3_outputs(4915) <= a;
    layer3_outputs(4916) <= not b;
    layer3_outputs(4917) <= b;
    layer3_outputs(4918) <= a or b;
    layer3_outputs(4919) <= b;
    layer3_outputs(4920) <= a;
    layer3_outputs(4921) <= b and not a;
    layer3_outputs(4922) <= not b;
    layer3_outputs(4923) <= b and not a;
    layer3_outputs(4924) <= not a;
    layer3_outputs(4925) <= not a or b;
    layer3_outputs(4926) <= not (a or b);
    layer3_outputs(4927) <= not b;
    layer3_outputs(4928) <= not b;
    layer3_outputs(4929) <= a;
    layer3_outputs(4930) <= not b or a;
    layer3_outputs(4931) <= not a;
    layer3_outputs(4932) <= not a;
    layer3_outputs(4933) <= a;
    layer3_outputs(4934) <= b and not a;
    layer3_outputs(4935) <= not (a or b);
    layer3_outputs(4936) <= '0';
    layer3_outputs(4937) <= not (a or b);
    layer3_outputs(4938) <= a xor b;
    layer3_outputs(4939) <= not (a or b);
    layer3_outputs(4940) <= not a;
    layer3_outputs(4941) <= not a;
    layer3_outputs(4942) <= not (a and b);
    layer3_outputs(4943) <= a and not b;
    layer3_outputs(4944) <= not (a and b);
    layer3_outputs(4945) <= not b or a;
    layer3_outputs(4946) <= not a;
    layer3_outputs(4947) <= not b or a;
    layer3_outputs(4948) <= b and not a;
    layer3_outputs(4949) <= a;
    layer3_outputs(4950) <= not b;
    layer3_outputs(4951) <= b;
    layer3_outputs(4952) <= a and not b;
    layer3_outputs(4953) <= not a;
    layer3_outputs(4954) <= not a or b;
    layer3_outputs(4955) <= a and b;
    layer3_outputs(4956) <= a and b;
    layer3_outputs(4957) <= not b or a;
    layer3_outputs(4958) <= b;
    layer3_outputs(4959) <= a xor b;
    layer3_outputs(4960) <= a;
    layer3_outputs(4961) <= a;
    layer3_outputs(4962) <= '0';
    layer3_outputs(4963) <= not b or a;
    layer3_outputs(4964) <= not a or b;
    layer3_outputs(4965) <= b and not a;
    layer3_outputs(4966) <= b and not a;
    layer3_outputs(4967) <= not b or a;
    layer3_outputs(4968) <= b;
    layer3_outputs(4969) <= b and not a;
    layer3_outputs(4970) <= a xor b;
    layer3_outputs(4971) <= a or b;
    layer3_outputs(4972) <= b;
    layer3_outputs(4973) <= a;
    layer3_outputs(4974) <= a xor b;
    layer3_outputs(4975) <= b;
    layer3_outputs(4976) <= not b;
    layer3_outputs(4977) <= not b;
    layer3_outputs(4978) <= b;
    layer3_outputs(4979) <= a;
    layer3_outputs(4980) <= b and not a;
    layer3_outputs(4981) <= a and b;
    layer3_outputs(4982) <= not a;
    layer3_outputs(4983) <= b;
    layer3_outputs(4984) <= '1';
    layer3_outputs(4985) <= a;
    layer3_outputs(4986) <= not a;
    layer3_outputs(4987) <= not b or a;
    layer3_outputs(4988) <= '1';
    layer3_outputs(4989) <= b;
    layer3_outputs(4990) <= not a;
    layer3_outputs(4991) <= '0';
    layer3_outputs(4992) <= not a;
    layer3_outputs(4993) <= b;
    layer3_outputs(4994) <= a;
    layer3_outputs(4995) <= not b;
    layer3_outputs(4996) <= '0';
    layer3_outputs(4997) <= not a;
    layer3_outputs(4998) <= '0';
    layer3_outputs(4999) <= not a;
    layer3_outputs(5000) <= not b or a;
    layer3_outputs(5001) <= not (a or b);
    layer3_outputs(5002) <= '1';
    layer3_outputs(5003) <= not (a or b);
    layer3_outputs(5004) <= '0';
    layer3_outputs(5005) <= not (a or b);
    layer3_outputs(5006) <= a;
    layer3_outputs(5007) <= a xor b;
    layer3_outputs(5008) <= '1';
    layer3_outputs(5009) <= a and b;
    layer3_outputs(5010) <= a and not b;
    layer3_outputs(5011) <= a xor b;
    layer3_outputs(5012) <= not (a or b);
    layer3_outputs(5013) <= not a;
    layer3_outputs(5014) <= b and not a;
    layer3_outputs(5015) <= a;
    layer3_outputs(5016) <= a or b;
    layer3_outputs(5017) <= '1';
    layer3_outputs(5018) <= not a or b;
    layer3_outputs(5019) <= not a or b;
    layer3_outputs(5020) <= b;
    layer3_outputs(5021) <= b and not a;
    layer3_outputs(5022) <= not b;
    layer3_outputs(5023) <= not (a or b);
    layer3_outputs(5024) <= not a;
    layer3_outputs(5025) <= '0';
    layer3_outputs(5026) <= b;
    layer3_outputs(5027) <= not b or a;
    layer3_outputs(5028) <= not b;
    layer3_outputs(5029) <= '1';
    layer3_outputs(5030) <= a;
    layer3_outputs(5031) <= '0';
    layer3_outputs(5032) <= not a;
    layer3_outputs(5033) <= a and b;
    layer3_outputs(5034) <= a;
    layer3_outputs(5035) <= '0';
    layer3_outputs(5036) <= a and b;
    layer3_outputs(5037) <= not (a xor b);
    layer3_outputs(5038) <= not (a xor b);
    layer3_outputs(5039) <= b;
    layer3_outputs(5040) <= not (a or b);
    layer3_outputs(5041) <= a;
    layer3_outputs(5042) <= a or b;
    layer3_outputs(5043) <= '0';
    layer3_outputs(5044) <= '1';
    layer3_outputs(5045) <= not (a or b);
    layer3_outputs(5046) <= not (a or b);
    layer3_outputs(5047) <= not (a xor b);
    layer3_outputs(5048) <= b;
    layer3_outputs(5049) <= a or b;
    layer3_outputs(5050) <= b;
    layer3_outputs(5051) <= not b;
    layer3_outputs(5052) <= not a;
    layer3_outputs(5053) <= not a;
    layer3_outputs(5054) <= not a or b;
    layer3_outputs(5055) <= a;
    layer3_outputs(5056) <= b;
    layer3_outputs(5057) <= not (a xor b);
    layer3_outputs(5058) <= not a;
    layer3_outputs(5059) <= a and b;
    layer3_outputs(5060) <= a and b;
    layer3_outputs(5061) <= a or b;
    layer3_outputs(5062) <= not b;
    layer3_outputs(5063) <= a or b;
    layer3_outputs(5064) <= not a;
    layer3_outputs(5065) <= a and b;
    layer3_outputs(5066) <= a;
    layer3_outputs(5067) <= a or b;
    layer3_outputs(5068) <= not a or b;
    layer3_outputs(5069) <= not a;
    layer3_outputs(5070) <= b and not a;
    layer3_outputs(5071) <= b and not a;
    layer3_outputs(5072) <= b;
    layer3_outputs(5073) <= a;
    layer3_outputs(5074) <= a;
    layer3_outputs(5075) <= a;
    layer3_outputs(5076) <= not a or b;
    layer3_outputs(5077) <= a or b;
    layer3_outputs(5078) <= b;
    layer3_outputs(5079) <= a and not b;
    layer3_outputs(5080) <= not a or b;
    layer3_outputs(5081) <= b;
    layer3_outputs(5082) <= not a or b;
    layer3_outputs(5083) <= a;
    layer3_outputs(5084) <= a and not b;
    layer3_outputs(5085) <= not b or a;
    layer3_outputs(5086) <= not a;
    layer3_outputs(5087) <= not (a and b);
    layer3_outputs(5088) <= not (a and b);
    layer3_outputs(5089) <= not a;
    layer3_outputs(5090) <= not b;
    layer3_outputs(5091) <= a;
    layer3_outputs(5092) <= '0';
    layer3_outputs(5093) <= a or b;
    layer3_outputs(5094) <= b and not a;
    layer3_outputs(5095) <= not b;
    layer3_outputs(5096) <= not b;
    layer3_outputs(5097) <= a or b;
    layer3_outputs(5098) <= not b or a;
    layer3_outputs(5099) <= not a or b;
    layer3_outputs(5100) <= a or b;
    layer3_outputs(5101) <= not b;
    layer3_outputs(5102) <= not b or a;
    layer3_outputs(5103) <= not (a or b);
    layer3_outputs(5104) <= b;
    layer3_outputs(5105) <= '1';
    layer3_outputs(5106) <= b;
    layer3_outputs(5107) <= a or b;
    layer3_outputs(5108) <= b;
    layer3_outputs(5109) <= not (a or b);
    layer3_outputs(5110) <= b and not a;
    layer3_outputs(5111) <= a and not b;
    layer3_outputs(5112) <= b;
    layer3_outputs(5113) <= a and not b;
    layer3_outputs(5114) <= '0';
    layer3_outputs(5115) <= not a or b;
    layer3_outputs(5116) <= b and not a;
    layer3_outputs(5117) <= a;
    layer3_outputs(5118) <= a;
    layer3_outputs(5119) <= not a or b;
    layer3_outputs(5120) <= not b;
    layer3_outputs(5121) <= not a or b;
    layer3_outputs(5122) <= not b or a;
    layer3_outputs(5123) <= not a;
    layer3_outputs(5124) <= a;
    layer3_outputs(5125) <= a;
    layer3_outputs(5126) <= not b or a;
    layer3_outputs(5127) <= b;
    layer3_outputs(5128) <= b;
    layer3_outputs(5129) <= not b or a;
    layer3_outputs(5130) <= a xor b;
    layer3_outputs(5131) <= not b;
    layer3_outputs(5132) <= not a or b;
    layer3_outputs(5133) <= a;
    layer3_outputs(5134) <= a and b;
    layer3_outputs(5135) <= not b;
    layer3_outputs(5136) <= a or b;
    layer3_outputs(5137) <= not a or b;
    layer3_outputs(5138) <= not (a or b);
    layer3_outputs(5139) <= not b;
    layer3_outputs(5140) <= a;
    layer3_outputs(5141) <= '0';
    layer3_outputs(5142) <= not (a and b);
    layer3_outputs(5143) <= b;
    layer3_outputs(5144) <= a and b;
    layer3_outputs(5145) <= a;
    layer3_outputs(5146) <= a and not b;
    layer3_outputs(5147) <= b;
    layer3_outputs(5148) <= b;
    layer3_outputs(5149) <= not a;
    layer3_outputs(5150) <= b and not a;
    layer3_outputs(5151) <= a;
    layer3_outputs(5152) <= a or b;
    layer3_outputs(5153) <= not (a or b);
    layer3_outputs(5154) <= not (a and b);
    layer3_outputs(5155) <= a or b;
    layer3_outputs(5156) <= '0';
    layer3_outputs(5157) <= '0';
    layer3_outputs(5158) <= a;
    layer3_outputs(5159) <= a;
    layer3_outputs(5160) <= not b or a;
    layer3_outputs(5161) <= '1';
    layer3_outputs(5162) <= not b or a;
    layer3_outputs(5163) <= a;
    layer3_outputs(5164) <= not a;
    layer3_outputs(5165) <= not (a or b);
    layer3_outputs(5166) <= a and not b;
    layer3_outputs(5167) <= b and not a;
    layer3_outputs(5168) <= a and not b;
    layer3_outputs(5169) <= not (a or b);
    layer3_outputs(5170) <= not a;
    layer3_outputs(5171) <= not a or b;
    layer3_outputs(5172) <= not (a and b);
    layer3_outputs(5173) <= not (a and b);
    layer3_outputs(5174) <= a;
    layer3_outputs(5175) <= not a;
    layer3_outputs(5176) <= not (a or b);
    layer3_outputs(5177) <= not b;
    layer3_outputs(5178) <= not (a or b);
    layer3_outputs(5179) <= not (a or b);
    layer3_outputs(5180) <= not (a xor b);
    layer3_outputs(5181) <= not a or b;
    layer3_outputs(5182) <= not b;
    layer3_outputs(5183) <= not b;
    layer3_outputs(5184) <= not a or b;
    layer3_outputs(5185) <= a;
    layer3_outputs(5186) <= a;
    layer3_outputs(5187) <= not a or b;
    layer3_outputs(5188) <= not a or b;
    layer3_outputs(5189) <= b and not a;
    layer3_outputs(5190) <= a and not b;
    layer3_outputs(5191) <= not (a and b);
    layer3_outputs(5192) <= not a or b;
    layer3_outputs(5193) <= a;
    layer3_outputs(5194) <= not b;
    layer3_outputs(5195) <= b and not a;
    layer3_outputs(5196) <= '1';
    layer3_outputs(5197) <= a;
    layer3_outputs(5198) <= '0';
    layer3_outputs(5199) <= not a;
    layer3_outputs(5200) <= b;
    layer3_outputs(5201) <= b and not a;
    layer3_outputs(5202) <= not a;
    layer3_outputs(5203) <= a and not b;
    layer3_outputs(5204) <= a;
    layer3_outputs(5205) <= not a;
    layer3_outputs(5206) <= not b or a;
    layer3_outputs(5207) <= a or b;
    layer3_outputs(5208) <= a xor b;
    layer3_outputs(5209) <= a;
    layer3_outputs(5210) <= not (a and b);
    layer3_outputs(5211) <= a and b;
    layer3_outputs(5212) <= '1';
    layer3_outputs(5213) <= a and not b;
    layer3_outputs(5214) <= b;
    layer3_outputs(5215) <= not b;
    layer3_outputs(5216) <= a xor b;
    layer3_outputs(5217) <= a xor b;
    layer3_outputs(5218) <= a;
    layer3_outputs(5219) <= not (a xor b);
    layer3_outputs(5220) <= not a or b;
    layer3_outputs(5221) <= b;
    layer3_outputs(5222) <= a and not b;
    layer3_outputs(5223) <= not a or b;
    layer3_outputs(5224) <= a and b;
    layer3_outputs(5225) <= a or b;
    layer3_outputs(5226) <= b;
    layer3_outputs(5227) <= a and not b;
    layer3_outputs(5228) <= a and not b;
    layer3_outputs(5229) <= b and not a;
    layer3_outputs(5230) <= not a;
    layer3_outputs(5231) <= b;
    layer3_outputs(5232) <= b;
    layer3_outputs(5233) <= a and b;
    layer3_outputs(5234) <= '1';
    layer3_outputs(5235) <= not b or a;
    layer3_outputs(5236) <= not (a and b);
    layer3_outputs(5237) <= a xor b;
    layer3_outputs(5238) <= not b;
    layer3_outputs(5239) <= not b or a;
    layer3_outputs(5240) <= a and not b;
    layer3_outputs(5241) <= not a;
    layer3_outputs(5242) <= a and not b;
    layer3_outputs(5243) <= b;
    layer3_outputs(5244) <= b;
    layer3_outputs(5245) <= not (a xor b);
    layer3_outputs(5246) <= not (a or b);
    layer3_outputs(5247) <= b and not a;
    layer3_outputs(5248) <= a;
    layer3_outputs(5249) <= b and not a;
    layer3_outputs(5250) <= b;
    layer3_outputs(5251) <= not a or b;
    layer3_outputs(5252) <= not (a and b);
    layer3_outputs(5253) <= b;
    layer3_outputs(5254) <= not b;
    layer3_outputs(5255) <= not a or b;
    layer3_outputs(5256) <= not a;
    layer3_outputs(5257) <= not b;
    layer3_outputs(5258) <= not b;
    layer3_outputs(5259) <= b;
    layer3_outputs(5260) <= '1';
    layer3_outputs(5261) <= b;
    layer3_outputs(5262) <= b;
    layer3_outputs(5263) <= not b or a;
    layer3_outputs(5264) <= not a;
    layer3_outputs(5265) <= a and not b;
    layer3_outputs(5266) <= not b;
    layer3_outputs(5267) <= b;
    layer3_outputs(5268) <= a;
    layer3_outputs(5269) <= a and not b;
    layer3_outputs(5270) <= not b or a;
    layer3_outputs(5271) <= not b;
    layer3_outputs(5272) <= not a;
    layer3_outputs(5273) <= not (a xor b);
    layer3_outputs(5274) <= not b;
    layer3_outputs(5275) <= not (a and b);
    layer3_outputs(5276) <= a xor b;
    layer3_outputs(5277) <= a or b;
    layer3_outputs(5278) <= '1';
    layer3_outputs(5279) <= a or b;
    layer3_outputs(5280) <= not (a xor b);
    layer3_outputs(5281) <= a;
    layer3_outputs(5282) <= not a;
    layer3_outputs(5283) <= not b or a;
    layer3_outputs(5284) <= not b;
    layer3_outputs(5285) <= not b or a;
    layer3_outputs(5286) <= not a;
    layer3_outputs(5287) <= b;
    layer3_outputs(5288) <= not b;
    layer3_outputs(5289) <= a or b;
    layer3_outputs(5290) <= not a;
    layer3_outputs(5291) <= '0';
    layer3_outputs(5292) <= b;
    layer3_outputs(5293) <= not a or b;
    layer3_outputs(5294) <= not a;
    layer3_outputs(5295) <= a;
    layer3_outputs(5296) <= not b or a;
    layer3_outputs(5297) <= not b;
    layer3_outputs(5298) <= a or b;
    layer3_outputs(5299) <= not a;
    layer3_outputs(5300) <= a;
    layer3_outputs(5301) <= not a or b;
    layer3_outputs(5302) <= not (a xor b);
    layer3_outputs(5303) <= a xor b;
    layer3_outputs(5304) <= not b;
    layer3_outputs(5305) <= not (a or b);
    layer3_outputs(5306) <= b;
    layer3_outputs(5307) <= not b;
    layer3_outputs(5308) <= not (a and b);
    layer3_outputs(5309) <= a or b;
    layer3_outputs(5310) <= not (a and b);
    layer3_outputs(5311) <= a and not b;
    layer3_outputs(5312) <= a;
    layer3_outputs(5313) <= not (a and b);
    layer3_outputs(5314) <= a xor b;
    layer3_outputs(5315) <= '0';
    layer3_outputs(5316) <= b;
    layer3_outputs(5317) <= not b;
    layer3_outputs(5318) <= a xor b;
    layer3_outputs(5319) <= not b;
    layer3_outputs(5320) <= a and not b;
    layer3_outputs(5321) <= b;
    layer3_outputs(5322) <= not (a or b);
    layer3_outputs(5323) <= not b;
    layer3_outputs(5324) <= a and not b;
    layer3_outputs(5325) <= not (a or b);
    layer3_outputs(5326) <= not a or b;
    layer3_outputs(5327) <= b;
    layer3_outputs(5328) <= b and not a;
    layer3_outputs(5329) <= a and not b;
    layer3_outputs(5330) <= a or b;
    layer3_outputs(5331) <= not a or b;
    layer3_outputs(5332) <= a xor b;
    layer3_outputs(5333) <= not (a or b);
    layer3_outputs(5334) <= not b;
    layer3_outputs(5335) <= a and b;
    layer3_outputs(5336) <= b and not a;
    layer3_outputs(5337) <= b and not a;
    layer3_outputs(5338) <= b;
    layer3_outputs(5339) <= a or b;
    layer3_outputs(5340) <= a or b;
    layer3_outputs(5341) <= not (a and b);
    layer3_outputs(5342) <= b and not a;
    layer3_outputs(5343) <= a or b;
    layer3_outputs(5344) <= a;
    layer3_outputs(5345) <= b;
    layer3_outputs(5346) <= a and b;
    layer3_outputs(5347) <= not b;
    layer3_outputs(5348) <= a;
    layer3_outputs(5349) <= not a or b;
    layer3_outputs(5350) <= b and not a;
    layer3_outputs(5351) <= '1';
    layer3_outputs(5352) <= a;
    layer3_outputs(5353) <= a and not b;
    layer3_outputs(5354) <= not (a or b);
    layer3_outputs(5355) <= '0';
    layer3_outputs(5356) <= '0';
    layer3_outputs(5357) <= not b;
    layer3_outputs(5358) <= not (a and b);
    layer3_outputs(5359) <= a and b;
    layer3_outputs(5360) <= '0';
    layer3_outputs(5361) <= b and not a;
    layer3_outputs(5362) <= not (a or b);
    layer3_outputs(5363) <= a;
    layer3_outputs(5364) <= a and not b;
    layer3_outputs(5365) <= not b or a;
    layer3_outputs(5366) <= not a or b;
    layer3_outputs(5367) <= not (a or b);
    layer3_outputs(5368) <= a xor b;
    layer3_outputs(5369) <= '1';
    layer3_outputs(5370) <= '0';
    layer3_outputs(5371) <= not a or b;
    layer3_outputs(5372) <= a;
    layer3_outputs(5373) <= b;
    layer3_outputs(5374) <= not a or b;
    layer3_outputs(5375) <= not b or a;
    layer3_outputs(5376) <= a or b;
    layer3_outputs(5377) <= a;
    layer3_outputs(5378) <= a or b;
    layer3_outputs(5379) <= not b or a;
    layer3_outputs(5380) <= a xor b;
    layer3_outputs(5381) <= not b;
    layer3_outputs(5382) <= not (a and b);
    layer3_outputs(5383) <= not b;
    layer3_outputs(5384) <= b;
    layer3_outputs(5385) <= not (a xor b);
    layer3_outputs(5386) <= a;
    layer3_outputs(5387) <= '0';
    layer3_outputs(5388) <= b;
    layer3_outputs(5389) <= a and b;
    layer3_outputs(5390) <= a and b;
    layer3_outputs(5391) <= a;
    layer3_outputs(5392) <= not (a or b);
    layer3_outputs(5393) <= not (a or b);
    layer3_outputs(5394) <= '0';
    layer3_outputs(5395) <= not b;
    layer3_outputs(5396) <= a or b;
    layer3_outputs(5397) <= not a or b;
    layer3_outputs(5398) <= not b;
    layer3_outputs(5399) <= b;
    layer3_outputs(5400) <= not b;
    layer3_outputs(5401) <= not b or a;
    layer3_outputs(5402) <= not (a and b);
    layer3_outputs(5403) <= a;
    layer3_outputs(5404) <= a and b;
    layer3_outputs(5405) <= a xor b;
    layer3_outputs(5406) <= not (a and b);
    layer3_outputs(5407) <= not (a or b);
    layer3_outputs(5408) <= '1';
    layer3_outputs(5409) <= not a;
    layer3_outputs(5410) <= not a;
    layer3_outputs(5411) <= '1';
    layer3_outputs(5412) <= not a;
    layer3_outputs(5413) <= b;
    layer3_outputs(5414) <= a xor b;
    layer3_outputs(5415) <= a or b;
    layer3_outputs(5416) <= not a or b;
    layer3_outputs(5417) <= '1';
    layer3_outputs(5418) <= b;
    layer3_outputs(5419) <= not b;
    layer3_outputs(5420) <= b and not a;
    layer3_outputs(5421) <= not (a and b);
    layer3_outputs(5422) <= b and not a;
    layer3_outputs(5423) <= not a or b;
    layer3_outputs(5424) <= '1';
    layer3_outputs(5425) <= '0';
    layer3_outputs(5426) <= not b or a;
    layer3_outputs(5427) <= '1';
    layer3_outputs(5428) <= a;
    layer3_outputs(5429) <= not a or b;
    layer3_outputs(5430) <= a and not b;
    layer3_outputs(5431) <= not b;
    layer3_outputs(5432) <= not (a xor b);
    layer3_outputs(5433) <= a and b;
    layer3_outputs(5434) <= a and b;
    layer3_outputs(5435) <= not a;
    layer3_outputs(5436) <= a xor b;
    layer3_outputs(5437) <= a;
    layer3_outputs(5438) <= not a;
    layer3_outputs(5439) <= b;
    layer3_outputs(5440) <= not b or a;
    layer3_outputs(5441) <= not (a and b);
    layer3_outputs(5442) <= '1';
    layer3_outputs(5443) <= not (a or b);
    layer3_outputs(5444) <= not b;
    layer3_outputs(5445) <= not b;
    layer3_outputs(5446) <= '1';
    layer3_outputs(5447) <= a and b;
    layer3_outputs(5448) <= b;
    layer3_outputs(5449) <= b;
    layer3_outputs(5450) <= b;
    layer3_outputs(5451) <= b;
    layer3_outputs(5452) <= a;
    layer3_outputs(5453) <= not a or b;
    layer3_outputs(5454) <= b;
    layer3_outputs(5455) <= not (a and b);
    layer3_outputs(5456) <= not (a or b);
    layer3_outputs(5457) <= not b or a;
    layer3_outputs(5458) <= not (a or b);
    layer3_outputs(5459) <= not a;
    layer3_outputs(5460) <= b and not a;
    layer3_outputs(5461) <= '1';
    layer3_outputs(5462) <= not a;
    layer3_outputs(5463) <= '1';
    layer3_outputs(5464) <= not (a or b);
    layer3_outputs(5465) <= a and not b;
    layer3_outputs(5466) <= not (a or b);
    layer3_outputs(5467) <= not (a or b);
    layer3_outputs(5468) <= a;
    layer3_outputs(5469) <= not (a xor b);
    layer3_outputs(5470) <= not (a and b);
    layer3_outputs(5471) <= not a;
    layer3_outputs(5472) <= '1';
    layer3_outputs(5473) <= not b;
    layer3_outputs(5474) <= a xor b;
    layer3_outputs(5475) <= a and not b;
    layer3_outputs(5476) <= a;
    layer3_outputs(5477) <= '1';
    layer3_outputs(5478) <= not a or b;
    layer3_outputs(5479) <= a or b;
    layer3_outputs(5480) <= not b;
    layer3_outputs(5481) <= a;
    layer3_outputs(5482) <= a xor b;
    layer3_outputs(5483) <= a and b;
    layer3_outputs(5484) <= not (a xor b);
    layer3_outputs(5485) <= not a;
    layer3_outputs(5486) <= b;
    layer3_outputs(5487) <= not b;
    layer3_outputs(5488) <= b;
    layer3_outputs(5489) <= b;
    layer3_outputs(5490) <= b;
    layer3_outputs(5491) <= a and not b;
    layer3_outputs(5492) <= b and not a;
    layer3_outputs(5493) <= a and b;
    layer3_outputs(5494) <= not (a xor b);
    layer3_outputs(5495) <= not (a or b);
    layer3_outputs(5496) <= a or b;
    layer3_outputs(5497) <= not (a or b);
    layer3_outputs(5498) <= a;
    layer3_outputs(5499) <= a and not b;
    layer3_outputs(5500) <= not b;
    layer3_outputs(5501) <= not a;
    layer3_outputs(5502) <= a xor b;
    layer3_outputs(5503) <= a;
    layer3_outputs(5504) <= not (a or b);
    layer3_outputs(5505) <= not (a and b);
    layer3_outputs(5506) <= not a or b;
    layer3_outputs(5507) <= a and not b;
    layer3_outputs(5508) <= not b or a;
    layer3_outputs(5509) <= '0';
    layer3_outputs(5510) <= a and not b;
    layer3_outputs(5511) <= a or b;
    layer3_outputs(5512) <= not a;
    layer3_outputs(5513) <= not a;
    layer3_outputs(5514) <= not (a xor b);
    layer3_outputs(5515) <= '0';
    layer3_outputs(5516) <= not (a xor b);
    layer3_outputs(5517) <= not a or b;
    layer3_outputs(5518) <= not a;
    layer3_outputs(5519) <= a;
    layer3_outputs(5520) <= not a;
    layer3_outputs(5521) <= b;
    layer3_outputs(5522) <= a and b;
    layer3_outputs(5523) <= not a;
    layer3_outputs(5524) <= a and not b;
    layer3_outputs(5525) <= '1';
    layer3_outputs(5526) <= not b;
    layer3_outputs(5527) <= b and not a;
    layer3_outputs(5528) <= '0';
    layer3_outputs(5529) <= not a or b;
    layer3_outputs(5530) <= a or b;
    layer3_outputs(5531) <= b;
    layer3_outputs(5532) <= not (a and b);
    layer3_outputs(5533) <= b;
    layer3_outputs(5534) <= not b;
    layer3_outputs(5535) <= a xor b;
    layer3_outputs(5536) <= not (a or b);
    layer3_outputs(5537) <= b and not a;
    layer3_outputs(5538) <= not b;
    layer3_outputs(5539) <= not b or a;
    layer3_outputs(5540) <= not a;
    layer3_outputs(5541) <= not a;
    layer3_outputs(5542) <= a and b;
    layer3_outputs(5543) <= a and not b;
    layer3_outputs(5544) <= not b;
    layer3_outputs(5545) <= not (a xor b);
    layer3_outputs(5546) <= not b;
    layer3_outputs(5547) <= not a;
    layer3_outputs(5548) <= not a;
    layer3_outputs(5549) <= b and not a;
    layer3_outputs(5550) <= a or b;
    layer3_outputs(5551) <= not a;
    layer3_outputs(5552) <= '0';
    layer3_outputs(5553) <= not a or b;
    layer3_outputs(5554) <= not (a or b);
    layer3_outputs(5555) <= not a;
    layer3_outputs(5556) <= not b;
    layer3_outputs(5557) <= not b;
    layer3_outputs(5558) <= not (a xor b);
    layer3_outputs(5559) <= '0';
    layer3_outputs(5560) <= not a;
    layer3_outputs(5561) <= not a;
    layer3_outputs(5562) <= not (a or b);
    layer3_outputs(5563) <= not b;
    layer3_outputs(5564) <= a or b;
    layer3_outputs(5565) <= a and b;
    layer3_outputs(5566) <= a;
    layer3_outputs(5567) <= '1';
    layer3_outputs(5568) <= a and not b;
    layer3_outputs(5569) <= not a;
    layer3_outputs(5570) <= not a;
    layer3_outputs(5571) <= not (a or b);
    layer3_outputs(5572) <= not (a and b);
    layer3_outputs(5573) <= b;
    layer3_outputs(5574) <= a xor b;
    layer3_outputs(5575) <= a;
    layer3_outputs(5576) <= a;
    layer3_outputs(5577) <= a or b;
    layer3_outputs(5578) <= not (a xor b);
    layer3_outputs(5579) <= not b or a;
    layer3_outputs(5580) <= not b;
    layer3_outputs(5581) <= not (a xor b);
    layer3_outputs(5582) <= not a;
    layer3_outputs(5583) <= b;
    layer3_outputs(5584) <= a;
    layer3_outputs(5585) <= not a or b;
    layer3_outputs(5586) <= not b;
    layer3_outputs(5587) <= a and not b;
    layer3_outputs(5588) <= not b or a;
    layer3_outputs(5589) <= b;
    layer3_outputs(5590) <= not a;
    layer3_outputs(5591) <= a and not b;
    layer3_outputs(5592) <= not a;
    layer3_outputs(5593) <= not b;
    layer3_outputs(5594) <= '1';
    layer3_outputs(5595) <= not b;
    layer3_outputs(5596) <= b;
    layer3_outputs(5597) <= not (a and b);
    layer3_outputs(5598) <= b;
    layer3_outputs(5599) <= b;
    layer3_outputs(5600) <= a and b;
    layer3_outputs(5601) <= not a or b;
    layer3_outputs(5602) <= a;
    layer3_outputs(5603) <= a;
    layer3_outputs(5604) <= not (a or b);
    layer3_outputs(5605) <= not (a or b);
    layer3_outputs(5606) <= not b;
    layer3_outputs(5607) <= not a;
    layer3_outputs(5608) <= b;
    layer3_outputs(5609) <= a;
    layer3_outputs(5610) <= b;
    layer3_outputs(5611) <= a and b;
    layer3_outputs(5612) <= b;
    layer3_outputs(5613) <= a or b;
    layer3_outputs(5614) <= '1';
    layer3_outputs(5615) <= a;
    layer3_outputs(5616) <= not a;
    layer3_outputs(5617) <= not (a xor b);
    layer3_outputs(5618) <= a xor b;
    layer3_outputs(5619) <= not (a xor b);
    layer3_outputs(5620) <= a xor b;
    layer3_outputs(5621) <= not a or b;
    layer3_outputs(5622) <= a and not b;
    layer3_outputs(5623) <= not b or a;
    layer3_outputs(5624) <= a;
    layer3_outputs(5625) <= '0';
    layer3_outputs(5626) <= not (a xor b);
    layer3_outputs(5627) <= not (a xor b);
    layer3_outputs(5628) <= not a;
    layer3_outputs(5629) <= b;
    layer3_outputs(5630) <= a xor b;
    layer3_outputs(5631) <= not b;
    layer3_outputs(5632) <= a or b;
    layer3_outputs(5633) <= a;
    layer3_outputs(5634) <= not b;
    layer3_outputs(5635) <= not a;
    layer3_outputs(5636) <= not a;
    layer3_outputs(5637) <= b;
    layer3_outputs(5638) <= not b;
    layer3_outputs(5639) <= a and not b;
    layer3_outputs(5640) <= '1';
    layer3_outputs(5641) <= not (a or b);
    layer3_outputs(5642) <= a and b;
    layer3_outputs(5643) <= not a or b;
    layer3_outputs(5644) <= b and not a;
    layer3_outputs(5645) <= b;
    layer3_outputs(5646) <= not b or a;
    layer3_outputs(5647) <= b and not a;
    layer3_outputs(5648) <= not a;
    layer3_outputs(5649) <= not (a xor b);
    layer3_outputs(5650) <= not b or a;
    layer3_outputs(5651) <= not a;
    layer3_outputs(5652) <= a xor b;
    layer3_outputs(5653) <= not a;
    layer3_outputs(5654) <= not a;
    layer3_outputs(5655) <= a and not b;
    layer3_outputs(5656) <= a xor b;
    layer3_outputs(5657) <= a and b;
    layer3_outputs(5658) <= a;
    layer3_outputs(5659) <= not b;
    layer3_outputs(5660) <= not a;
    layer3_outputs(5661) <= a and b;
    layer3_outputs(5662) <= not (a xor b);
    layer3_outputs(5663) <= a and not b;
    layer3_outputs(5664) <= not a;
    layer3_outputs(5665) <= '0';
    layer3_outputs(5666) <= not b or a;
    layer3_outputs(5667) <= not a;
    layer3_outputs(5668) <= not a;
    layer3_outputs(5669) <= not a or b;
    layer3_outputs(5670) <= b and not a;
    layer3_outputs(5671) <= a;
    layer3_outputs(5672) <= a or b;
    layer3_outputs(5673) <= a and b;
    layer3_outputs(5674) <= b;
    layer3_outputs(5675) <= a;
    layer3_outputs(5676) <= not (a and b);
    layer3_outputs(5677) <= a;
    layer3_outputs(5678) <= a;
    layer3_outputs(5679) <= b;
    layer3_outputs(5680) <= b;
    layer3_outputs(5681) <= a and not b;
    layer3_outputs(5682) <= b and not a;
    layer3_outputs(5683) <= a xor b;
    layer3_outputs(5684) <= not (a or b);
    layer3_outputs(5685) <= not (a xor b);
    layer3_outputs(5686) <= b;
    layer3_outputs(5687) <= '0';
    layer3_outputs(5688) <= '1';
    layer3_outputs(5689) <= '1';
    layer3_outputs(5690) <= '0';
    layer3_outputs(5691) <= '0';
    layer3_outputs(5692) <= b and not a;
    layer3_outputs(5693) <= a xor b;
    layer3_outputs(5694) <= b;
    layer3_outputs(5695) <= b;
    layer3_outputs(5696) <= not (a and b);
    layer3_outputs(5697) <= '1';
    layer3_outputs(5698) <= not (a and b);
    layer3_outputs(5699) <= a;
    layer3_outputs(5700) <= a and not b;
    layer3_outputs(5701) <= not a or b;
    layer3_outputs(5702) <= b and not a;
    layer3_outputs(5703) <= not (a and b);
    layer3_outputs(5704) <= not a or b;
    layer3_outputs(5705) <= b;
    layer3_outputs(5706) <= a and b;
    layer3_outputs(5707) <= not b or a;
    layer3_outputs(5708) <= a and b;
    layer3_outputs(5709) <= b and not a;
    layer3_outputs(5710) <= not b;
    layer3_outputs(5711) <= not b or a;
    layer3_outputs(5712) <= not b;
    layer3_outputs(5713) <= not a;
    layer3_outputs(5714) <= b and not a;
    layer3_outputs(5715) <= not (a and b);
    layer3_outputs(5716) <= a and not b;
    layer3_outputs(5717) <= b;
    layer3_outputs(5718) <= not a;
    layer3_outputs(5719) <= b and not a;
    layer3_outputs(5720) <= not b;
    layer3_outputs(5721) <= a;
    layer3_outputs(5722) <= a;
    layer3_outputs(5723) <= not b;
    layer3_outputs(5724) <= a xor b;
    layer3_outputs(5725) <= b and not a;
    layer3_outputs(5726) <= '1';
    layer3_outputs(5727) <= a and b;
    layer3_outputs(5728) <= a or b;
    layer3_outputs(5729) <= '1';
    layer3_outputs(5730) <= not b or a;
    layer3_outputs(5731) <= not (a or b);
    layer3_outputs(5732) <= a or b;
    layer3_outputs(5733) <= not (a xor b);
    layer3_outputs(5734) <= not (a xor b);
    layer3_outputs(5735) <= b and not a;
    layer3_outputs(5736) <= not a or b;
    layer3_outputs(5737) <= b;
    layer3_outputs(5738) <= b;
    layer3_outputs(5739) <= a;
    layer3_outputs(5740) <= a and b;
    layer3_outputs(5741) <= b and not a;
    layer3_outputs(5742) <= not (a and b);
    layer3_outputs(5743) <= not b or a;
    layer3_outputs(5744) <= not (a and b);
    layer3_outputs(5745) <= not b;
    layer3_outputs(5746) <= b;
    layer3_outputs(5747) <= not a;
    layer3_outputs(5748) <= a;
    layer3_outputs(5749) <= a and not b;
    layer3_outputs(5750) <= not (a and b);
    layer3_outputs(5751) <= a;
    layer3_outputs(5752) <= a;
    layer3_outputs(5753) <= a or b;
    layer3_outputs(5754) <= b;
    layer3_outputs(5755) <= not (a xor b);
    layer3_outputs(5756) <= not b or a;
    layer3_outputs(5757) <= b and not a;
    layer3_outputs(5758) <= not (a and b);
    layer3_outputs(5759) <= b;
    layer3_outputs(5760) <= not b;
    layer3_outputs(5761) <= not (a xor b);
    layer3_outputs(5762) <= b;
    layer3_outputs(5763) <= a;
    layer3_outputs(5764) <= '1';
    layer3_outputs(5765) <= '1';
    layer3_outputs(5766) <= not a or b;
    layer3_outputs(5767) <= b and not a;
    layer3_outputs(5768) <= not b or a;
    layer3_outputs(5769) <= a or b;
    layer3_outputs(5770) <= a and not b;
    layer3_outputs(5771) <= a;
    layer3_outputs(5772) <= a and b;
    layer3_outputs(5773) <= not (a xor b);
    layer3_outputs(5774) <= a and b;
    layer3_outputs(5775) <= a xor b;
    layer3_outputs(5776) <= '0';
    layer3_outputs(5777) <= not a;
    layer3_outputs(5778) <= b;
    layer3_outputs(5779) <= '1';
    layer3_outputs(5780) <= not (a or b);
    layer3_outputs(5781) <= not a;
    layer3_outputs(5782) <= a xor b;
    layer3_outputs(5783) <= a;
    layer3_outputs(5784) <= not b;
    layer3_outputs(5785) <= a or b;
    layer3_outputs(5786) <= not (a xor b);
    layer3_outputs(5787) <= a xor b;
    layer3_outputs(5788) <= a or b;
    layer3_outputs(5789) <= b;
    layer3_outputs(5790) <= b;
    layer3_outputs(5791) <= a and b;
    layer3_outputs(5792) <= not a;
    layer3_outputs(5793) <= a or b;
    layer3_outputs(5794) <= not b or a;
    layer3_outputs(5795) <= '1';
    layer3_outputs(5796) <= not b;
    layer3_outputs(5797) <= not b;
    layer3_outputs(5798) <= not a or b;
    layer3_outputs(5799) <= a and b;
    layer3_outputs(5800) <= a and b;
    layer3_outputs(5801) <= '0';
    layer3_outputs(5802) <= not (a and b);
    layer3_outputs(5803) <= a xor b;
    layer3_outputs(5804) <= not b;
    layer3_outputs(5805) <= '0';
    layer3_outputs(5806) <= a and b;
    layer3_outputs(5807) <= a;
    layer3_outputs(5808) <= not (a or b);
    layer3_outputs(5809) <= not a;
    layer3_outputs(5810) <= a;
    layer3_outputs(5811) <= not a;
    layer3_outputs(5812) <= not a or b;
    layer3_outputs(5813) <= not a;
    layer3_outputs(5814) <= a;
    layer3_outputs(5815) <= b;
    layer3_outputs(5816) <= a and b;
    layer3_outputs(5817) <= b and not a;
    layer3_outputs(5818) <= not a;
    layer3_outputs(5819) <= not (a or b);
    layer3_outputs(5820) <= b and not a;
    layer3_outputs(5821) <= b;
    layer3_outputs(5822) <= b and not a;
    layer3_outputs(5823) <= not (a or b);
    layer3_outputs(5824) <= a xor b;
    layer3_outputs(5825) <= not a;
    layer3_outputs(5826) <= a and not b;
    layer3_outputs(5827) <= not a;
    layer3_outputs(5828) <= not b or a;
    layer3_outputs(5829) <= a and not b;
    layer3_outputs(5830) <= not a;
    layer3_outputs(5831) <= not b or a;
    layer3_outputs(5832) <= not a or b;
    layer3_outputs(5833) <= not b;
    layer3_outputs(5834) <= a or b;
    layer3_outputs(5835) <= not b;
    layer3_outputs(5836) <= a and b;
    layer3_outputs(5837) <= not a or b;
    layer3_outputs(5838) <= a and not b;
    layer3_outputs(5839) <= b and not a;
    layer3_outputs(5840) <= not a;
    layer3_outputs(5841) <= a and not b;
    layer3_outputs(5842) <= a;
    layer3_outputs(5843) <= '1';
    layer3_outputs(5844) <= a or b;
    layer3_outputs(5845) <= not (a and b);
    layer3_outputs(5846) <= '0';
    layer3_outputs(5847) <= b and not a;
    layer3_outputs(5848) <= not b or a;
    layer3_outputs(5849) <= a or b;
    layer3_outputs(5850) <= not a;
    layer3_outputs(5851) <= b;
    layer3_outputs(5852) <= '0';
    layer3_outputs(5853) <= not (a or b);
    layer3_outputs(5854) <= not a;
    layer3_outputs(5855) <= not (a or b);
    layer3_outputs(5856) <= a xor b;
    layer3_outputs(5857) <= a and not b;
    layer3_outputs(5858) <= b;
    layer3_outputs(5859) <= '1';
    layer3_outputs(5860) <= not a or b;
    layer3_outputs(5861) <= not b;
    layer3_outputs(5862) <= a xor b;
    layer3_outputs(5863) <= a or b;
    layer3_outputs(5864) <= not (a and b);
    layer3_outputs(5865) <= not (a or b);
    layer3_outputs(5866) <= not (a xor b);
    layer3_outputs(5867) <= not b or a;
    layer3_outputs(5868) <= b and not a;
    layer3_outputs(5869) <= '0';
    layer3_outputs(5870) <= not (a or b);
    layer3_outputs(5871) <= not b;
    layer3_outputs(5872) <= '0';
    layer3_outputs(5873) <= a;
    layer3_outputs(5874) <= not (a or b);
    layer3_outputs(5875) <= b;
    layer3_outputs(5876) <= b and not a;
    layer3_outputs(5877) <= a or b;
    layer3_outputs(5878) <= not a;
    layer3_outputs(5879) <= not (a or b);
    layer3_outputs(5880) <= a or b;
    layer3_outputs(5881) <= not b;
    layer3_outputs(5882) <= '1';
    layer3_outputs(5883) <= b and not a;
    layer3_outputs(5884) <= b;
    layer3_outputs(5885) <= b;
    layer3_outputs(5886) <= not a;
    layer3_outputs(5887) <= b;
    layer3_outputs(5888) <= a;
    layer3_outputs(5889) <= not a;
    layer3_outputs(5890) <= not a or b;
    layer3_outputs(5891) <= b;
    layer3_outputs(5892) <= b;
    layer3_outputs(5893) <= a;
    layer3_outputs(5894) <= a;
    layer3_outputs(5895) <= not (a and b);
    layer3_outputs(5896) <= b;
    layer3_outputs(5897) <= not (a xor b);
    layer3_outputs(5898) <= '0';
    layer3_outputs(5899) <= a and b;
    layer3_outputs(5900) <= b and not a;
    layer3_outputs(5901) <= a;
    layer3_outputs(5902) <= a and b;
    layer3_outputs(5903) <= not (a xor b);
    layer3_outputs(5904) <= a xor b;
    layer3_outputs(5905) <= b;
    layer3_outputs(5906) <= a;
    layer3_outputs(5907) <= not b or a;
    layer3_outputs(5908) <= not b;
    layer3_outputs(5909) <= a;
    layer3_outputs(5910) <= b;
    layer3_outputs(5911) <= not (a xor b);
    layer3_outputs(5912) <= a and not b;
    layer3_outputs(5913) <= a and b;
    layer3_outputs(5914) <= '1';
    layer3_outputs(5915) <= a;
    layer3_outputs(5916) <= not b;
    layer3_outputs(5917) <= a or b;
    layer3_outputs(5918) <= a or b;
    layer3_outputs(5919) <= a and b;
    layer3_outputs(5920) <= b and not a;
    layer3_outputs(5921) <= not b;
    layer3_outputs(5922) <= not a or b;
    layer3_outputs(5923) <= a and not b;
    layer3_outputs(5924) <= '1';
    layer3_outputs(5925) <= not (a or b);
    layer3_outputs(5926) <= '0';
    layer3_outputs(5927) <= a xor b;
    layer3_outputs(5928) <= '0';
    layer3_outputs(5929) <= b and not a;
    layer3_outputs(5930) <= '1';
    layer3_outputs(5931) <= not a or b;
    layer3_outputs(5932) <= a or b;
    layer3_outputs(5933) <= b and not a;
    layer3_outputs(5934) <= not (a and b);
    layer3_outputs(5935) <= not b or a;
    layer3_outputs(5936) <= not (a and b);
    layer3_outputs(5937) <= not b or a;
    layer3_outputs(5938) <= a xor b;
    layer3_outputs(5939) <= not a or b;
    layer3_outputs(5940) <= not b;
    layer3_outputs(5941) <= '1';
    layer3_outputs(5942) <= a and not b;
    layer3_outputs(5943) <= a and b;
    layer3_outputs(5944) <= not a;
    layer3_outputs(5945) <= b and not a;
    layer3_outputs(5946) <= a and b;
    layer3_outputs(5947) <= not b or a;
    layer3_outputs(5948) <= a;
    layer3_outputs(5949) <= not b or a;
    layer3_outputs(5950) <= '1';
    layer3_outputs(5951) <= not a;
    layer3_outputs(5952) <= not (a or b);
    layer3_outputs(5953) <= not (a xor b);
    layer3_outputs(5954) <= a xor b;
    layer3_outputs(5955) <= not b;
    layer3_outputs(5956) <= not (a or b);
    layer3_outputs(5957) <= not a;
    layer3_outputs(5958) <= a;
    layer3_outputs(5959) <= a xor b;
    layer3_outputs(5960) <= b and not a;
    layer3_outputs(5961) <= a;
    layer3_outputs(5962) <= b and not a;
    layer3_outputs(5963) <= a and not b;
    layer3_outputs(5964) <= a;
    layer3_outputs(5965) <= b;
    layer3_outputs(5966) <= not (a xor b);
    layer3_outputs(5967) <= a xor b;
    layer3_outputs(5968) <= not a or b;
    layer3_outputs(5969) <= b;
    layer3_outputs(5970) <= not a;
    layer3_outputs(5971) <= not b;
    layer3_outputs(5972) <= not (a xor b);
    layer3_outputs(5973) <= not (a or b);
    layer3_outputs(5974) <= a and not b;
    layer3_outputs(5975) <= not (a and b);
    layer3_outputs(5976) <= b;
    layer3_outputs(5977) <= b;
    layer3_outputs(5978) <= a or b;
    layer3_outputs(5979) <= b;
    layer3_outputs(5980) <= b and not a;
    layer3_outputs(5981) <= a;
    layer3_outputs(5982) <= b;
    layer3_outputs(5983) <= a and not b;
    layer3_outputs(5984) <= not (a and b);
    layer3_outputs(5985) <= not (a or b);
    layer3_outputs(5986) <= not a;
    layer3_outputs(5987) <= b and not a;
    layer3_outputs(5988) <= '1';
    layer3_outputs(5989) <= a and not b;
    layer3_outputs(5990) <= not a or b;
    layer3_outputs(5991) <= a;
    layer3_outputs(5992) <= b;
    layer3_outputs(5993) <= '1';
    layer3_outputs(5994) <= a;
    layer3_outputs(5995) <= a;
    layer3_outputs(5996) <= a and b;
    layer3_outputs(5997) <= not a;
    layer3_outputs(5998) <= not a or b;
    layer3_outputs(5999) <= not (a or b);
    layer3_outputs(6000) <= a and not b;
    layer3_outputs(6001) <= not b or a;
    layer3_outputs(6002) <= not a;
    layer3_outputs(6003) <= b and not a;
    layer3_outputs(6004) <= not b or a;
    layer3_outputs(6005) <= '0';
    layer3_outputs(6006) <= a and b;
    layer3_outputs(6007) <= not b;
    layer3_outputs(6008) <= '1';
    layer3_outputs(6009) <= a and b;
    layer3_outputs(6010) <= b and not a;
    layer3_outputs(6011) <= not b;
    layer3_outputs(6012) <= '0';
    layer3_outputs(6013) <= not b;
    layer3_outputs(6014) <= not b;
    layer3_outputs(6015) <= not a;
    layer3_outputs(6016) <= b;
    layer3_outputs(6017) <= a;
    layer3_outputs(6018) <= not b;
    layer3_outputs(6019) <= not b;
    layer3_outputs(6020) <= not (a and b);
    layer3_outputs(6021) <= a;
    layer3_outputs(6022) <= not (a and b);
    layer3_outputs(6023) <= not a;
    layer3_outputs(6024) <= not b;
    layer3_outputs(6025) <= not (a and b);
    layer3_outputs(6026) <= not a;
    layer3_outputs(6027) <= '1';
    layer3_outputs(6028) <= a or b;
    layer3_outputs(6029) <= a;
    layer3_outputs(6030) <= not a or b;
    layer3_outputs(6031) <= b and not a;
    layer3_outputs(6032) <= a and b;
    layer3_outputs(6033) <= not (a and b);
    layer3_outputs(6034) <= '0';
    layer3_outputs(6035) <= b;
    layer3_outputs(6036) <= a or b;
    layer3_outputs(6037) <= b;
    layer3_outputs(6038) <= not (a and b);
    layer3_outputs(6039) <= '0';
    layer3_outputs(6040) <= not a;
    layer3_outputs(6041) <= a;
    layer3_outputs(6042) <= not a;
    layer3_outputs(6043) <= not b;
    layer3_outputs(6044) <= a and not b;
    layer3_outputs(6045) <= not a;
    layer3_outputs(6046) <= not a;
    layer3_outputs(6047) <= not b;
    layer3_outputs(6048) <= not (a xor b);
    layer3_outputs(6049) <= a xor b;
    layer3_outputs(6050) <= not (a and b);
    layer3_outputs(6051) <= not a;
    layer3_outputs(6052) <= b and not a;
    layer3_outputs(6053) <= not (a xor b);
    layer3_outputs(6054) <= a and not b;
    layer3_outputs(6055) <= not b;
    layer3_outputs(6056) <= a;
    layer3_outputs(6057) <= a and b;
    layer3_outputs(6058) <= a;
    layer3_outputs(6059) <= '0';
    layer3_outputs(6060) <= a or b;
    layer3_outputs(6061) <= not b;
    layer3_outputs(6062) <= b and not a;
    layer3_outputs(6063) <= not a or b;
    layer3_outputs(6064) <= not (a xor b);
    layer3_outputs(6065) <= not b;
    layer3_outputs(6066) <= '1';
    layer3_outputs(6067) <= a xor b;
    layer3_outputs(6068) <= not b or a;
    layer3_outputs(6069) <= b;
    layer3_outputs(6070) <= not (a and b);
    layer3_outputs(6071) <= b;
    layer3_outputs(6072) <= not (a xor b);
    layer3_outputs(6073) <= b;
    layer3_outputs(6074) <= not b;
    layer3_outputs(6075) <= a;
    layer3_outputs(6076) <= not (a or b);
    layer3_outputs(6077) <= a and b;
    layer3_outputs(6078) <= a or b;
    layer3_outputs(6079) <= a;
    layer3_outputs(6080) <= not a;
    layer3_outputs(6081) <= not (a and b);
    layer3_outputs(6082) <= not (a xor b);
    layer3_outputs(6083) <= not (a and b);
    layer3_outputs(6084) <= a;
    layer3_outputs(6085) <= not (a xor b);
    layer3_outputs(6086) <= '0';
    layer3_outputs(6087) <= a xor b;
    layer3_outputs(6088) <= a or b;
    layer3_outputs(6089) <= not a;
    layer3_outputs(6090) <= not b or a;
    layer3_outputs(6091) <= a xor b;
    layer3_outputs(6092) <= a and b;
    layer3_outputs(6093) <= not b or a;
    layer3_outputs(6094) <= b;
    layer3_outputs(6095) <= b and not a;
    layer3_outputs(6096) <= b and not a;
    layer3_outputs(6097) <= a or b;
    layer3_outputs(6098) <= not (a xor b);
    layer3_outputs(6099) <= not b or a;
    layer3_outputs(6100) <= not (a and b);
    layer3_outputs(6101) <= a or b;
    layer3_outputs(6102) <= b and not a;
    layer3_outputs(6103) <= a and b;
    layer3_outputs(6104) <= not b;
    layer3_outputs(6105) <= a;
    layer3_outputs(6106) <= not a or b;
    layer3_outputs(6107) <= not (a xor b);
    layer3_outputs(6108) <= a and not b;
    layer3_outputs(6109) <= not a;
    layer3_outputs(6110) <= a;
    layer3_outputs(6111) <= a or b;
    layer3_outputs(6112) <= b;
    layer3_outputs(6113) <= a xor b;
    layer3_outputs(6114) <= not a;
    layer3_outputs(6115) <= a xor b;
    layer3_outputs(6116) <= not a;
    layer3_outputs(6117) <= not (a xor b);
    layer3_outputs(6118) <= a xor b;
    layer3_outputs(6119) <= a;
    layer3_outputs(6120) <= not a or b;
    layer3_outputs(6121) <= a and b;
    layer3_outputs(6122) <= a and not b;
    layer3_outputs(6123) <= not (a and b);
    layer3_outputs(6124) <= not a;
    layer3_outputs(6125) <= not b;
    layer3_outputs(6126) <= b;
    layer3_outputs(6127) <= '1';
    layer3_outputs(6128) <= not b or a;
    layer3_outputs(6129) <= not (a or b);
    layer3_outputs(6130) <= not a;
    layer3_outputs(6131) <= not (a or b);
    layer3_outputs(6132) <= not (a or b);
    layer3_outputs(6133) <= b and not a;
    layer3_outputs(6134) <= not (a and b);
    layer3_outputs(6135) <= '1';
    layer3_outputs(6136) <= a and b;
    layer3_outputs(6137) <= '0';
    layer3_outputs(6138) <= not b;
    layer3_outputs(6139) <= not b;
    layer3_outputs(6140) <= not (a and b);
    layer3_outputs(6141) <= not b;
    layer3_outputs(6142) <= not b;
    layer3_outputs(6143) <= a and b;
    layer3_outputs(6144) <= not a or b;
    layer3_outputs(6145) <= a and not b;
    layer3_outputs(6146) <= not a;
    layer3_outputs(6147) <= not (a or b);
    layer3_outputs(6148) <= b and not a;
    layer3_outputs(6149) <= a or b;
    layer3_outputs(6150) <= not b or a;
    layer3_outputs(6151) <= not (a and b);
    layer3_outputs(6152) <= not b;
    layer3_outputs(6153) <= not a;
    layer3_outputs(6154) <= b and not a;
    layer3_outputs(6155) <= not a;
    layer3_outputs(6156) <= not (a and b);
    layer3_outputs(6157) <= b;
    layer3_outputs(6158) <= b;
    layer3_outputs(6159) <= not a;
    layer3_outputs(6160) <= a and not b;
    layer3_outputs(6161) <= not b or a;
    layer3_outputs(6162) <= not b;
    layer3_outputs(6163) <= a;
    layer3_outputs(6164) <= a;
    layer3_outputs(6165) <= not (a or b);
    layer3_outputs(6166) <= b and not a;
    layer3_outputs(6167) <= '1';
    layer3_outputs(6168) <= not b or a;
    layer3_outputs(6169) <= a;
    layer3_outputs(6170) <= not b or a;
    layer3_outputs(6171) <= b and not a;
    layer3_outputs(6172) <= not a;
    layer3_outputs(6173) <= not (a or b);
    layer3_outputs(6174) <= not a;
    layer3_outputs(6175) <= a;
    layer3_outputs(6176) <= b and not a;
    layer3_outputs(6177) <= a xor b;
    layer3_outputs(6178) <= not a;
    layer3_outputs(6179) <= b;
    layer3_outputs(6180) <= '0';
    layer3_outputs(6181) <= not b;
    layer3_outputs(6182) <= a and not b;
    layer3_outputs(6183) <= a;
    layer3_outputs(6184) <= not b or a;
    layer3_outputs(6185) <= a or b;
    layer3_outputs(6186) <= not (a and b);
    layer3_outputs(6187) <= a and b;
    layer3_outputs(6188) <= not b;
    layer3_outputs(6189) <= not a or b;
    layer3_outputs(6190) <= not (a or b);
    layer3_outputs(6191) <= not a or b;
    layer3_outputs(6192) <= not a or b;
    layer3_outputs(6193) <= a and b;
    layer3_outputs(6194) <= not (a and b);
    layer3_outputs(6195) <= a and b;
    layer3_outputs(6196) <= a and b;
    layer3_outputs(6197) <= '1';
    layer3_outputs(6198) <= a or b;
    layer3_outputs(6199) <= not a;
    layer3_outputs(6200) <= not b;
    layer3_outputs(6201) <= not b or a;
    layer3_outputs(6202) <= not a;
    layer3_outputs(6203) <= b;
    layer3_outputs(6204) <= '0';
    layer3_outputs(6205) <= not a;
    layer3_outputs(6206) <= b;
    layer3_outputs(6207) <= '1';
    layer3_outputs(6208) <= a or b;
    layer3_outputs(6209) <= not (a and b);
    layer3_outputs(6210) <= b;
    layer3_outputs(6211) <= a and b;
    layer3_outputs(6212) <= a;
    layer3_outputs(6213) <= b and not a;
    layer3_outputs(6214) <= a and b;
    layer3_outputs(6215) <= not (a and b);
    layer3_outputs(6216) <= not (a or b);
    layer3_outputs(6217) <= not b;
    layer3_outputs(6218) <= not (a and b);
    layer3_outputs(6219) <= not b;
    layer3_outputs(6220) <= b and not a;
    layer3_outputs(6221) <= a and not b;
    layer3_outputs(6222) <= b and not a;
    layer3_outputs(6223) <= not a;
    layer3_outputs(6224) <= a;
    layer3_outputs(6225) <= not b;
    layer3_outputs(6226) <= a or b;
    layer3_outputs(6227) <= not a;
    layer3_outputs(6228) <= a and not b;
    layer3_outputs(6229) <= a and not b;
    layer3_outputs(6230) <= not (a xor b);
    layer3_outputs(6231) <= not (a and b);
    layer3_outputs(6232) <= a;
    layer3_outputs(6233) <= b and not a;
    layer3_outputs(6234) <= a;
    layer3_outputs(6235) <= b;
    layer3_outputs(6236) <= a and not b;
    layer3_outputs(6237) <= not b;
    layer3_outputs(6238) <= not (a xor b);
    layer3_outputs(6239) <= not b or a;
    layer3_outputs(6240) <= b;
    layer3_outputs(6241) <= not (a or b);
    layer3_outputs(6242) <= a and b;
    layer3_outputs(6243) <= not b or a;
    layer3_outputs(6244) <= not b;
    layer3_outputs(6245) <= b and not a;
    layer3_outputs(6246) <= a;
    layer3_outputs(6247) <= not a or b;
    layer3_outputs(6248) <= b and not a;
    layer3_outputs(6249) <= a;
    layer3_outputs(6250) <= not (a or b);
    layer3_outputs(6251) <= a xor b;
    layer3_outputs(6252) <= not b;
    layer3_outputs(6253) <= not b;
    layer3_outputs(6254) <= b;
    layer3_outputs(6255) <= b and not a;
    layer3_outputs(6256) <= a or b;
    layer3_outputs(6257) <= not b or a;
    layer3_outputs(6258) <= '1';
    layer3_outputs(6259) <= not (a and b);
    layer3_outputs(6260) <= b and not a;
    layer3_outputs(6261) <= not b;
    layer3_outputs(6262) <= not b or a;
    layer3_outputs(6263) <= not a or b;
    layer3_outputs(6264) <= a and not b;
    layer3_outputs(6265) <= b;
    layer3_outputs(6266) <= b;
    layer3_outputs(6267) <= a;
    layer3_outputs(6268) <= a or b;
    layer3_outputs(6269) <= b;
    layer3_outputs(6270) <= not a;
    layer3_outputs(6271) <= not (a or b);
    layer3_outputs(6272) <= a;
    layer3_outputs(6273) <= a;
    layer3_outputs(6274) <= '1';
    layer3_outputs(6275) <= not b or a;
    layer3_outputs(6276) <= a xor b;
    layer3_outputs(6277) <= a and not b;
    layer3_outputs(6278) <= b;
    layer3_outputs(6279) <= not a;
    layer3_outputs(6280) <= a and b;
    layer3_outputs(6281) <= a and b;
    layer3_outputs(6282) <= b and not a;
    layer3_outputs(6283) <= not b or a;
    layer3_outputs(6284) <= b;
    layer3_outputs(6285) <= not (a or b);
    layer3_outputs(6286) <= not a or b;
    layer3_outputs(6287) <= b;
    layer3_outputs(6288) <= not (a or b);
    layer3_outputs(6289) <= a and b;
    layer3_outputs(6290) <= '1';
    layer3_outputs(6291) <= b and not a;
    layer3_outputs(6292) <= a or b;
    layer3_outputs(6293) <= not b;
    layer3_outputs(6294) <= not a or b;
    layer3_outputs(6295) <= not (a and b);
    layer3_outputs(6296) <= not b;
    layer3_outputs(6297) <= b and not a;
    layer3_outputs(6298) <= b and not a;
    layer3_outputs(6299) <= a and not b;
    layer3_outputs(6300) <= b;
    layer3_outputs(6301) <= '1';
    layer3_outputs(6302) <= b;
    layer3_outputs(6303) <= not (a and b);
    layer3_outputs(6304) <= '0';
    layer3_outputs(6305) <= not b;
    layer3_outputs(6306) <= b;
    layer3_outputs(6307) <= b and not a;
    layer3_outputs(6308) <= a or b;
    layer3_outputs(6309) <= not a or b;
    layer3_outputs(6310) <= not b;
    layer3_outputs(6311) <= a xor b;
    layer3_outputs(6312) <= a xor b;
    layer3_outputs(6313) <= a xor b;
    layer3_outputs(6314) <= a or b;
    layer3_outputs(6315) <= not b or a;
    layer3_outputs(6316) <= a and b;
    layer3_outputs(6317) <= not a or b;
    layer3_outputs(6318) <= not (a or b);
    layer3_outputs(6319) <= not (a and b);
    layer3_outputs(6320) <= b;
    layer3_outputs(6321) <= not a;
    layer3_outputs(6322) <= not b;
    layer3_outputs(6323) <= a and b;
    layer3_outputs(6324) <= not (a xor b);
    layer3_outputs(6325) <= a and not b;
    layer3_outputs(6326) <= not (a or b);
    layer3_outputs(6327) <= a;
    layer3_outputs(6328) <= a or b;
    layer3_outputs(6329) <= '0';
    layer3_outputs(6330) <= a or b;
    layer3_outputs(6331) <= a;
    layer3_outputs(6332) <= a or b;
    layer3_outputs(6333) <= not a;
    layer3_outputs(6334) <= not a;
    layer3_outputs(6335) <= not b or a;
    layer3_outputs(6336) <= a;
    layer3_outputs(6337) <= a;
    layer3_outputs(6338) <= not (a and b);
    layer3_outputs(6339) <= a and not b;
    layer3_outputs(6340) <= '0';
    layer3_outputs(6341) <= '0';
    layer3_outputs(6342) <= a or b;
    layer3_outputs(6343) <= not b;
    layer3_outputs(6344) <= not a or b;
    layer3_outputs(6345) <= not (a or b);
    layer3_outputs(6346) <= a xor b;
    layer3_outputs(6347) <= a and b;
    layer3_outputs(6348) <= b;
    layer3_outputs(6349) <= b;
    layer3_outputs(6350) <= not (a or b);
    layer3_outputs(6351) <= a and not b;
    layer3_outputs(6352) <= a and not b;
    layer3_outputs(6353) <= not (a and b);
    layer3_outputs(6354) <= not b;
    layer3_outputs(6355) <= b;
    layer3_outputs(6356) <= a and not b;
    layer3_outputs(6357) <= b;
    layer3_outputs(6358) <= a and b;
    layer3_outputs(6359) <= a and not b;
    layer3_outputs(6360) <= b and not a;
    layer3_outputs(6361) <= not b;
    layer3_outputs(6362) <= not (a and b);
    layer3_outputs(6363) <= not b or a;
    layer3_outputs(6364) <= not b or a;
    layer3_outputs(6365) <= not a;
    layer3_outputs(6366) <= '0';
    layer3_outputs(6367) <= not a;
    layer3_outputs(6368) <= a or b;
    layer3_outputs(6369) <= a;
    layer3_outputs(6370) <= '1';
    layer3_outputs(6371) <= a and b;
    layer3_outputs(6372) <= '1';
    layer3_outputs(6373) <= '0';
    layer3_outputs(6374) <= not b;
    layer3_outputs(6375) <= not b or a;
    layer3_outputs(6376) <= not b;
    layer3_outputs(6377) <= a;
    layer3_outputs(6378) <= not (a and b);
    layer3_outputs(6379) <= not a;
    layer3_outputs(6380) <= not b;
    layer3_outputs(6381) <= not b;
    layer3_outputs(6382) <= not (a or b);
    layer3_outputs(6383) <= not a;
    layer3_outputs(6384) <= a and b;
    layer3_outputs(6385) <= not a;
    layer3_outputs(6386) <= not a;
    layer3_outputs(6387) <= b and not a;
    layer3_outputs(6388) <= not (a and b);
    layer3_outputs(6389) <= a;
    layer3_outputs(6390) <= not b;
    layer3_outputs(6391) <= b;
    layer3_outputs(6392) <= not a;
    layer3_outputs(6393) <= not (a and b);
    layer3_outputs(6394) <= '1';
    layer3_outputs(6395) <= a or b;
    layer3_outputs(6396) <= not (a or b);
    layer3_outputs(6397) <= not b;
    layer3_outputs(6398) <= not a;
    layer3_outputs(6399) <= not b;
    layer3_outputs(6400) <= not a or b;
    layer3_outputs(6401) <= '1';
    layer3_outputs(6402) <= not b or a;
    layer3_outputs(6403) <= '1';
    layer3_outputs(6404) <= a or b;
    layer3_outputs(6405) <= not a;
    layer3_outputs(6406) <= not a or b;
    layer3_outputs(6407) <= not a;
    layer3_outputs(6408) <= not b;
    layer3_outputs(6409) <= not b;
    layer3_outputs(6410) <= '0';
    layer3_outputs(6411) <= b and not a;
    layer3_outputs(6412) <= not a or b;
    layer3_outputs(6413) <= a and not b;
    layer3_outputs(6414) <= not (a and b);
    layer3_outputs(6415) <= not (a xor b);
    layer3_outputs(6416) <= not b or a;
    layer3_outputs(6417) <= b and not a;
    layer3_outputs(6418) <= not a;
    layer3_outputs(6419) <= not b or a;
    layer3_outputs(6420) <= a xor b;
    layer3_outputs(6421) <= not b or a;
    layer3_outputs(6422) <= not b;
    layer3_outputs(6423) <= not b;
    layer3_outputs(6424) <= '1';
    layer3_outputs(6425) <= b and not a;
    layer3_outputs(6426) <= not b or a;
    layer3_outputs(6427) <= b;
    layer3_outputs(6428) <= not (a or b);
    layer3_outputs(6429) <= a xor b;
    layer3_outputs(6430) <= not a;
    layer3_outputs(6431) <= a and b;
    layer3_outputs(6432) <= a or b;
    layer3_outputs(6433) <= b;
    layer3_outputs(6434) <= not (a and b);
    layer3_outputs(6435) <= a xor b;
    layer3_outputs(6436) <= b;
    layer3_outputs(6437) <= not (a or b);
    layer3_outputs(6438) <= not (a or b);
    layer3_outputs(6439) <= b;
    layer3_outputs(6440) <= not a or b;
    layer3_outputs(6441) <= a;
    layer3_outputs(6442) <= not b or a;
    layer3_outputs(6443) <= not a;
    layer3_outputs(6444) <= not b or a;
    layer3_outputs(6445) <= a and b;
    layer3_outputs(6446) <= b and not a;
    layer3_outputs(6447) <= not (a or b);
    layer3_outputs(6448) <= not b;
    layer3_outputs(6449) <= b;
    layer3_outputs(6450) <= '1';
    layer3_outputs(6451) <= b;
    layer3_outputs(6452) <= a;
    layer3_outputs(6453) <= a and b;
    layer3_outputs(6454) <= '1';
    layer3_outputs(6455) <= not b or a;
    layer3_outputs(6456) <= a;
    layer3_outputs(6457) <= a and b;
    layer3_outputs(6458) <= not (a or b);
    layer3_outputs(6459) <= not a or b;
    layer3_outputs(6460) <= '1';
    layer3_outputs(6461) <= not (a xor b);
    layer3_outputs(6462) <= not a;
    layer3_outputs(6463) <= not (a xor b);
    layer3_outputs(6464) <= not b or a;
    layer3_outputs(6465) <= not (a and b);
    layer3_outputs(6466) <= not b or a;
    layer3_outputs(6467) <= a;
    layer3_outputs(6468) <= not (a or b);
    layer3_outputs(6469) <= not (a and b);
    layer3_outputs(6470) <= not (a and b);
    layer3_outputs(6471) <= a;
    layer3_outputs(6472) <= not b or a;
    layer3_outputs(6473) <= a xor b;
    layer3_outputs(6474) <= a;
    layer3_outputs(6475) <= '1';
    layer3_outputs(6476) <= a xor b;
    layer3_outputs(6477) <= not (a and b);
    layer3_outputs(6478) <= not b or a;
    layer3_outputs(6479) <= a and b;
    layer3_outputs(6480) <= not (a and b);
    layer3_outputs(6481) <= not a;
    layer3_outputs(6482) <= '0';
    layer3_outputs(6483) <= b and not a;
    layer3_outputs(6484) <= not a;
    layer3_outputs(6485) <= not (a xor b);
    layer3_outputs(6486) <= b and not a;
    layer3_outputs(6487) <= not b;
    layer3_outputs(6488) <= a and not b;
    layer3_outputs(6489) <= not b;
    layer3_outputs(6490) <= not (a or b);
    layer3_outputs(6491) <= not (a and b);
    layer3_outputs(6492) <= a and b;
    layer3_outputs(6493) <= a xor b;
    layer3_outputs(6494) <= b;
    layer3_outputs(6495) <= not (a and b);
    layer3_outputs(6496) <= not b;
    layer3_outputs(6497) <= '1';
    layer3_outputs(6498) <= not (a and b);
    layer3_outputs(6499) <= a xor b;
    layer3_outputs(6500) <= '0';
    layer3_outputs(6501) <= a;
    layer3_outputs(6502) <= not a or b;
    layer3_outputs(6503) <= a xor b;
    layer3_outputs(6504) <= not b;
    layer3_outputs(6505) <= a;
    layer3_outputs(6506) <= not (a or b);
    layer3_outputs(6507) <= a xor b;
    layer3_outputs(6508) <= a and not b;
    layer3_outputs(6509) <= not b;
    layer3_outputs(6510) <= a and not b;
    layer3_outputs(6511) <= not (a and b);
    layer3_outputs(6512) <= not a;
    layer3_outputs(6513) <= b;
    layer3_outputs(6514) <= b;
    layer3_outputs(6515) <= not a;
    layer3_outputs(6516) <= not (a or b);
    layer3_outputs(6517) <= not b or a;
    layer3_outputs(6518) <= not b;
    layer3_outputs(6519) <= not b;
    layer3_outputs(6520) <= not (a or b);
    layer3_outputs(6521) <= not (a or b);
    layer3_outputs(6522) <= a and b;
    layer3_outputs(6523) <= b and not a;
    layer3_outputs(6524) <= a or b;
    layer3_outputs(6525) <= b and not a;
    layer3_outputs(6526) <= a;
    layer3_outputs(6527) <= not a;
    layer3_outputs(6528) <= a and b;
    layer3_outputs(6529) <= b;
    layer3_outputs(6530) <= a and b;
    layer3_outputs(6531) <= not (a and b);
    layer3_outputs(6532) <= not (a and b);
    layer3_outputs(6533) <= not a or b;
    layer3_outputs(6534) <= a or b;
    layer3_outputs(6535) <= a and b;
    layer3_outputs(6536) <= not (a or b);
    layer3_outputs(6537) <= a;
    layer3_outputs(6538) <= not b or a;
    layer3_outputs(6539) <= not b;
    layer3_outputs(6540) <= not (a or b);
    layer3_outputs(6541) <= a;
    layer3_outputs(6542) <= b;
    layer3_outputs(6543) <= a or b;
    layer3_outputs(6544) <= a or b;
    layer3_outputs(6545) <= not (a xor b);
    layer3_outputs(6546) <= not (a xor b);
    layer3_outputs(6547) <= a;
    layer3_outputs(6548) <= b;
    layer3_outputs(6549) <= not a or b;
    layer3_outputs(6550) <= '1';
    layer3_outputs(6551) <= a;
    layer3_outputs(6552) <= b;
    layer3_outputs(6553) <= a or b;
    layer3_outputs(6554) <= not a;
    layer3_outputs(6555) <= not a;
    layer3_outputs(6556) <= not a;
    layer3_outputs(6557) <= not a or b;
    layer3_outputs(6558) <= not a;
    layer3_outputs(6559) <= a xor b;
    layer3_outputs(6560) <= not a or b;
    layer3_outputs(6561) <= a and not b;
    layer3_outputs(6562) <= '0';
    layer3_outputs(6563) <= a or b;
    layer3_outputs(6564) <= b and not a;
    layer3_outputs(6565) <= not a or b;
    layer3_outputs(6566) <= not (a or b);
    layer3_outputs(6567) <= not (a and b);
    layer3_outputs(6568) <= not (a xor b);
    layer3_outputs(6569) <= a and b;
    layer3_outputs(6570) <= not b;
    layer3_outputs(6571) <= a and not b;
    layer3_outputs(6572) <= not (a or b);
    layer3_outputs(6573) <= not (a and b);
    layer3_outputs(6574) <= a and b;
    layer3_outputs(6575) <= '1';
    layer3_outputs(6576) <= a xor b;
    layer3_outputs(6577) <= not a or b;
    layer3_outputs(6578) <= '0';
    layer3_outputs(6579) <= not (a and b);
    layer3_outputs(6580) <= a and not b;
    layer3_outputs(6581) <= not a or b;
    layer3_outputs(6582) <= not (a xor b);
    layer3_outputs(6583) <= a and b;
    layer3_outputs(6584) <= not b;
    layer3_outputs(6585) <= not (a or b);
    layer3_outputs(6586) <= b;
    layer3_outputs(6587) <= not b;
    layer3_outputs(6588) <= a and b;
    layer3_outputs(6589) <= b and not a;
    layer3_outputs(6590) <= a and not b;
    layer3_outputs(6591) <= not a;
    layer3_outputs(6592) <= a and not b;
    layer3_outputs(6593) <= a;
    layer3_outputs(6594) <= not b;
    layer3_outputs(6595) <= a and not b;
    layer3_outputs(6596) <= not (a or b);
    layer3_outputs(6597) <= a or b;
    layer3_outputs(6598) <= a or b;
    layer3_outputs(6599) <= a or b;
    layer3_outputs(6600) <= not b or a;
    layer3_outputs(6601) <= a xor b;
    layer3_outputs(6602) <= a or b;
    layer3_outputs(6603) <= not b;
    layer3_outputs(6604) <= not b;
    layer3_outputs(6605) <= not (a xor b);
    layer3_outputs(6606) <= not a;
    layer3_outputs(6607) <= not b or a;
    layer3_outputs(6608) <= a and b;
    layer3_outputs(6609) <= a and not b;
    layer3_outputs(6610) <= not b or a;
    layer3_outputs(6611) <= b and not a;
    layer3_outputs(6612) <= not a;
    layer3_outputs(6613) <= not b or a;
    layer3_outputs(6614) <= not b;
    layer3_outputs(6615) <= a;
    layer3_outputs(6616) <= b and not a;
    layer3_outputs(6617) <= b;
    layer3_outputs(6618) <= not a;
    layer3_outputs(6619) <= b;
    layer3_outputs(6620) <= not b;
    layer3_outputs(6621) <= not a or b;
    layer3_outputs(6622) <= a xor b;
    layer3_outputs(6623) <= '1';
    layer3_outputs(6624) <= not (a xor b);
    layer3_outputs(6625) <= b;
    layer3_outputs(6626) <= not (a and b);
    layer3_outputs(6627) <= not b or a;
    layer3_outputs(6628) <= b;
    layer3_outputs(6629) <= a xor b;
    layer3_outputs(6630) <= b;
    layer3_outputs(6631) <= not a;
    layer3_outputs(6632) <= not a;
    layer3_outputs(6633) <= not a;
    layer3_outputs(6634) <= not a or b;
    layer3_outputs(6635) <= not a;
    layer3_outputs(6636) <= a xor b;
    layer3_outputs(6637) <= a;
    layer3_outputs(6638) <= b;
    layer3_outputs(6639) <= '1';
    layer3_outputs(6640) <= not b;
    layer3_outputs(6641) <= not a;
    layer3_outputs(6642) <= not (a xor b);
    layer3_outputs(6643) <= not b or a;
    layer3_outputs(6644) <= not a or b;
    layer3_outputs(6645) <= b;
    layer3_outputs(6646) <= a;
    layer3_outputs(6647) <= not a;
    layer3_outputs(6648) <= not b;
    layer3_outputs(6649) <= not b or a;
    layer3_outputs(6650) <= not a;
    layer3_outputs(6651) <= a and b;
    layer3_outputs(6652) <= not b or a;
    layer3_outputs(6653) <= a and not b;
    layer3_outputs(6654) <= not (a or b);
    layer3_outputs(6655) <= a;
    layer3_outputs(6656) <= not (a or b);
    layer3_outputs(6657) <= a;
    layer3_outputs(6658) <= not (a and b);
    layer3_outputs(6659) <= not b or a;
    layer3_outputs(6660) <= not (a and b);
    layer3_outputs(6661) <= a or b;
    layer3_outputs(6662) <= b;
    layer3_outputs(6663) <= a and not b;
    layer3_outputs(6664) <= not b;
    layer3_outputs(6665) <= a;
    layer3_outputs(6666) <= a and not b;
    layer3_outputs(6667) <= not a;
    layer3_outputs(6668) <= '1';
    layer3_outputs(6669) <= b;
    layer3_outputs(6670) <= not a or b;
    layer3_outputs(6671) <= not (a and b);
    layer3_outputs(6672) <= a or b;
    layer3_outputs(6673) <= not (a xor b);
    layer3_outputs(6674) <= a and b;
    layer3_outputs(6675) <= b;
    layer3_outputs(6676) <= not (a or b);
    layer3_outputs(6677) <= b and not a;
    layer3_outputs(6678) <= a or b;
    layer3_outputs(6679) <= not b or a;
    layer3_outputs(6680) <= a or b;
    layer3_outputs(6681) <= a or b;
    layer3_outputs(6682) <= not a;
    layer3_outputs(6683) <= a;
    layer3_outputs(6684) <= not b;
    layer3_outputs(6685) <= a or b;
    layer3_outputs(6686) <= b;
    layer3_outputs(6687) <= not b or a;
    layer3_outputs(6688) <= not a or b;
    layer3_outputs(6689) <= not b or a;
    layer3_outputs(6690) <= a xor b;
    layer3_outputs(6691) <= not a;
    layer3_outputs(6692) <= a and not b;
    layer3_outputs(6693) <= not b;
    layer3_outputs(6694) <= not b;
    layer3_outputs(6695) <= b and not a;
    layer3_outputs(6696) <= not b;
    layer3_outputs(6697) <= b and not a;
    layer3_outputs(6698) <= a and b;
    layer3_outputs(6699) <= not a;
    layer3_outputs(6700) <= not a;
    layer3_outputs(6701) <= a and not b;
    layer3_outputs(6702) <= a xor b;
    layer3_outputs(6703) <= not b or a;
    layer3_outputs(6704) <= not b;
    layer3_outputs(6705) <= not a;
    layer3_outputs(6706) <= not a or b;
    layer3_outputs(6707) <= '0';
    layer3_outputs(6708) <= not a;
    layer3_outputs(6709) <= not a or b;
    layer3_outputs(6710) <= b;
    layer3_outputs(6711) <= '0';
    layer3_outputs(6712) <= not b or a;
    layer3_outputs(6713) <= not (a or b);
    layer3_outputs(6714) <= a and b;
    layer3_outputs(6715) <= a and not b;
    layer3_outputs(6716) <= a;
    layer3_outputs(6717) <= not b or a;
    layer3_outputs(6718) <= not b;
    layer3_outputs(6719) <= not (a or b);
    layer3_outputs(6720) <= not a;
    layer3_outputs(6721) <= a;
    layer3_outputs(6722) <= not b;
    layer3_outputs(6723) <= '1';
    layer3_outputs(6724) <= b;
    layer3_outputs(6725) <= a or b;
    layer3_outputs(6726) <= a and b;
    layer3_outputs(6727) <= b and not a;
    layer3_outputs(6728) <= not (a and b);
    layer3_outputs(6729) <= a and b;
    layer3_outputs(6730) <= not (a and b);
    layer3_outputs(6731) <= not a or b;
    layer3_outputs(6732) <= not a;
    layer3_outputs(6733) <= a;
    layer3_outputs(6734) <= b and not a;
    layer3_outputs(6735) <= a and b;
    layer3_outputs(6736) <= not b;
    layer3_outputs(6737) <= a and not b;
    layer3_outputs(6738) <= a and b;
    layer3_outputs(6739) <= '1';
    layer3_outputs(6740) <= b and not a;
    layer3_outputs(6741) <= not a or b;
    layer3_outputs(6742) <= not b or a;
    layer3_outputs(6743) <= a and not b;
    layer3_outputs(6744) <= not a or b;
    layer3_outputs(6745) <= b;
    layer3_outputs(6746) <= not (a or b);
    layer3_outputs(6747) <= not (a and b);
    layer3_outputs(6748) <= a xor b;
    layer3_outputs(6749) <= not (a and b);
    layer3_outputs(6750) <= not (a or b);
    layer3_outputs(6751) <= not (a and b);
    layer3_outputs(6752) <= not (a xor b);
    layer3_outputs(6753) <= not (a or b);
    layer3_outputs(6754) <= not a;
    layer3_outputs(6755) <= a xor b;
    layer3_outputs(6756) <= a and b;
    layer3_outputs(6757) <= not b;
    layer3_outputs(6758) <= not a;
    layer3_outputs(6759) <= a;
    layer3_outputs(6760) <= not (a xor b);
    layer3_outputs(6761) <= not b or a;
    layer3_outputs(6762) <= not (a or b);
    layer3_outputs(6763) <= not b;
    layer3_outputs(6764) <= not a;
    layer3_outputs(6765) <= b;
    layer3_outputs(6766) <= not b;
    layer3_outputs(6767) <= '0';
    layer3_outputs(6768) <= a and b;
    layer3_outputs(6769) <= a;
    layer3_outputs(6770) <= b and not a;
    layer3_outputs(6771) <= a;
    layer3_outputs(6772) <= a;
    layer3_outputs(6773) <= '1';
    layer3_outputs(6774) <= not a;
    layer3_outputs(6775) <= '0';
    layer3_outputs(6776) <= a and not b;
    layer3_outputs(6777) <= b;
    layer3_outputs(6778) <= a and not b;
    layer3_outputs(6779) <= a;
    layer3_outputs(6780) <= not a or b;
    layer3_outputs(6781) <= b;
    layer3_outputs(6782) <= a and b;
    layer3_outputs(6783) <= not b or a;
    layer3_outputs(6784) <= a and not b;
    layer3_outputs(6785) <= not a or b;
    layer3_outputs(6786) <= b;
    layer3_outputs(6787) <= not (a or b);
    layer3_outputs(6788) <= a or b;
    layer3_outputs(6789) <= not a;
    layer3_outputs(6790) <= not a;
    layer3_outputs(6791) <= b;
    layer3_outputs(6792) <= not a;
    layer3_outputs(6793) <= not b;
    layer3_outputs(6794) <= not (a xor b);
    layer3_outputs(6795) <= '0';
    layer3_outputs(6796) <= not a;
    layer3_outputs(6797) <= not b or a;
    layer3_outputs(6798) <= not a or b;
    layer3_outputs(6799) <= b;
    layer3_outputs(6800) <= a;
    layer3_outputs(6801) <= not (a or b);
    layer3_outputs(6802) <= b and not a;
    layer3_outputs(6803) <= b and not a;
    layer3_outputs(6804) <= '1';
    layer3_outputs(6805) <= not b;
    layer3_outputs(6806) <= not b or a;
    layer3_outputs(6807) <= not (a and b);
    layer3_outputs(6808) <= not b or a;
    layer3_outputs(6809) <= b;
    layer3_outputs(6810) <= not b or a;
    layer3_outputs(6811) <= not b;
    layer3_outputs(6812) <= a and not b;
    layer3_outputs(6813) <= b and not a;
    layer3_outputs(6814) <= not a;
    layer3_outputs(6815) <= b;
    layer3_outputs(6816) <= a and not b;
    layer3_outputs(6817) <= not (a and b);
    layer3_outputs(6818) <= not (a and b);
    layer3_outputs(6819) <= b and not a;
    layer3_outputs(6820) <= not b or a;
    layer3_outputs(6821) <= not (a and b);
    layer3_outputs(6822) <= b;
    layer3_outputs(6823) <= not b or a;
    layer3_outputs(6824) <= b;
    layer3_outputs(6825) <= a and b;
    layer3_outputs(6826) <= not a;
    layer3_outputs(6827) <= '1';
    layer3_outputs(6828) <= not (a and b);
    layer3_outputs(6829) <= not a;
    layer3_outputs(6830) <= b and not a;
    layer3_outputs(6831) <= not b or a;
    layer3_outputs(6832) <= '1';
    layer3_outputs(6833) <= b;
    layer3_outputs(6834) <= a and b;
    layer3_outputs(6835) <= a or b;
    layer3_outputs(6836) <= '1';
    layer3_outputs(6837) <= not b;
    layer3_outputs(6838) <= not b;
    layer3_outputs(6839) <= a and not b;
    layer3_outputs(6840) <= a xor b;
    layer3_outputs(6841) <= not a;
    layer3_outputs(6842) <= not a;
    layer3_outputs(6843) <= a and b;
    layer3_outputs(6844) <= not a or b;
    layer3_outputs(6845) <= a and b;
    layer3_outputs(6846) <= not (a or b);
    layer3_outputs(6847) <= b;
    layer3_outputs(6848) <= a;
    layer3_outputs(6849) <= b;
    layer3_outputs(6850) <= a or b;
    layer3_outputs(6851) <= not (a and b);
    layer3_outputs(6852) <= a and b;
    layer3_outputs(6853) <= not b;
    layer3_outputs(6854) <= '1';
    layer3_outputs(6855) <= a and not b;
    layer3_outputs(6856) <= not a;
    layer3_outputs(6857) <= a and b;
    layer3_outputs(6858) <= a;
    layer3_outputs(6859) <= b;
    layer3_outputs(6860) <= a;
    layer3_outputs(6861) <= '0';
    layer3_outputs(6862) <= not b;
    layer3_outputs(6863) <= a;
    layer3_outputs(6864) <= a;
    layer3_outputs(6865) <= '1';
    layer3_outputs(6866) <= not (a and b);
    layer3_outputs(6867) <= a;
    layer3_outputs(6868) <= not b;
    layer3_outputs(6869) <= not b;
    layer3_outputs(6870) <= not a or b;
    layer3_outputs(6871) <= a;
    layer3_outputs(6872) <= not b;
    layer3_outputs(6873) <= b and not a;
    layer3_outputs(6874) <= a;
    layer3_outputs(6875) <= not (a or b);
    layer3_outputs(6876) <= b;
    layer3_outputs(6877) <= b;
    layer3_outputs(6878) <= a;
    layer3_outputs(6879) <= not (a xor b);
    layer3_outputs(6880) <= not a or b;
    layer3_outputs(6881) <= not b;
    layer3_outputs(6882) <= not a;
    layer3_outputs(6883) <= a and b;
    layer3_outputs(6884) <= a and b;
    layer3_outputs(6885) <= b;
    layer3_outputs(6886) <= a;
    layer3_outputs(6887) <= not a or b;
    layer3_outputs(6888) <= not (a and b);
    layer3_outputs(6889) <= b;
    layer3_outputs(6890) <= not b or a;
    layer3_outputs(6891) <= not a or b;
    layer3_outputs(6892) <= a;
    layer3_outputs(6893) <= '0';
    layer3_outputs(6894) <= not a or b;
    layer3_outputs(6895) <= not (a and b);
    layer3_outputs(6896) <= not (a or b);
    layer3_outputs(6897) <= b;
    layer3_outputs(6898) <= not a or b;
    layer3_outputs(6899) <= not b;
    layer3_outputs(6900) <= not b;
    layer3_outputs(6901) <= a xor b;
    layer3_outputs(6902) <= not a;
    layer3_outputs(6903) <= a;
    layer3_outputs(6904) <= not a or b;
    layer3_outputs(6905) <= b;
    layer3_outputs(6906) <= not b or a;
    layer3_outputs(6907) <= a and not b;
    layer3_outputs(6908) <= not a;
    layer3_outputs(6909) <= b;
    layer3_outputs(6910) <= not a;
    layer3_outputs(6911) <= a and not b;
    layer3_outputs(6912) <= a;
    layer3_outputs(6913) <= not b;
    layer3_outputs(6914) <= a and b;
    layer3_outputs(6915) <= not (a xor b);
    layer3_outputs(6916) <= a and b;
    layer3_outputs(6917) <= not (a xor b);
    layer3_outputs(6918) <= not a;
    layer3_outputs(6919) <= a or b;
    layer3_outputs(6920) <= not b or a;
    layer3_outputs(6921) <= not b or a;
    layer3_outputs(6922) <= not b or a;
    layer3_outputs(6923) <= not b;
    layer3_outputs(6924) <= b and not a;
    layer3_outputs(6925) <= a or b;
    layer3_outputs(6926) <= not (a or b);
    layer3_outputs(6927) <= not a;
    layer3_outputs(6928) <= a;
    layer3_outputs(6929) <= not b;
    layer3_outputs(6930) <= not b;
    layer3_outputs(6931) <= not a;
    layer3_outputs(6932) <= b;
    layer3_outputs(6933) <= b;
    layer3_outputs(6934) <= b and not a;
    layer3_outputs(6935) <= '0';
    layer3_outputs(6936) <= not (a or b);
    layer3_outputs(6937) <= not b or a;
    layer3_outputs(6938) <= a;
    layer3_outputs(6939) <= not a or b;
    layer3_outputs(6940) <= a;
    layer3_outputs(6941) <= not b or a;
    layer3_outputs(6942) <= a and not b;
    layer3_outputs(6943) <= b;
    layer3_outputs(6944) <= a;
    layer3_outputs(6945) <= not (a xor b);
    layer3_outputs(6946) <= a;
    layer3_outputs(6947) <= a or b;
    layer3_outputs(6948) <= a xor b;
    layer3_outputs(6949) <= not a;
    layer3_outputs(6950) <= not (a and b);
    layer3_outputs(6951) <= not a or b;
    layer3_outputs(6952) <= a and not b;
    layer3_outputs(6953) <= not a or b;
    layer3_outputs(6954) <= not (a and b);
    layer3_outputs(6955) <= not (a or b);
    layer3_outputs(6956) <= not a;
    layer3_outputs(6957) <= a or b;
    layer3_outputs(6958) <= '1';
    layer3_outputs(6959) <= a and b;
    layer3_outputs(6960) <= a;
    layer3_outputs(6961) <= b;
    layer3_outputs(6962) <= b;
    layer3_outputs(6963) <= not (a or b);
    layer3_outputs(6964) <= not b;
    layer3_outputs(6965) <= b and not a;
    layer3_outputs(6966) <= not b or a;
    layer3_outputs(6967) <= not (a and b);
    layer3_outputs(6968) <= not (a xor b);
    layer3_outputs(6969) <= a and b;
    layer3_outputs(6970) <= not a or b;
    layer3_outputs(6971) <= a and b;
    layer3_outputs(6972) <= '0';
    layer3_outputs(6973) <= not a or b;
    layer3_outputs(6974) <= not b;
    layer3_outputs(6975) <= a and not b;
    layer3_outputs(6976) <= not b or a;
    layer3_outputs(6977) <= not (a or b);
    layer3_outputs(6978) <= a or b;
    layer3_outputs(6979) <= not a or b;
    layer3_outputs(6980) <= not a or b;
    layer3_outputs(6981) <= a or b;
    layer3_outputs(6982) <= not b;
    layer3_outputs(6983) <= a;
    layer3_outputs(6984) <= not b;
    layer3_outputs(6985) <= a and b;
    layer3_outputs(6986) <= not (a or b);
    layer3_outputs(6987) <= '1';
    layer3_outputs(6988) <= not (a and b);
    layer3_outputs(6989) <= not b;
    layer3_outputs(6990) <= not b;
    layer3_outputs(6991) <= '0';
    layer3_outputs(6992) <= not a or b;
    layer3_outputs(6993) <= a;
    layer3_outputs(6994) <= not (a and b);
    layer3_outputs(6995) <= '1';
    layer3_outputs(6996) <= not b or a;
    layer3_outputs(6997) <= not (a and b);
    layer3_outputs(6998) <= not b;
    layer3_outputs(6999) <= not a;
    layer3_outputs(7000) <= not (a and b);
    layer3_outputs(7001) <= a and not b;
    layer3_outputs(7002) <= a or b;
    layer3_outputs(7003) <= not a;
    layer3_outputs(7004) <= not (a or b);
    layer3_outputs(7005) <= a xor b;
    layer3_outputs(7006) <= a;
    layer3_outputs(7007) <= '1';
    layer3_outputs(7008) <= not a or b;
    layer3_outputs(7009) <= not (a and b);
    layer3_outputs(7010) <= not b;
    layer3_outputs(7011) <= a xor b;
    layer3_outputs(7012) <= b;
    layer3_outputs(7013) <= not (a or b);
    layer3_outputs(7014) <= not (a xor b);
    layer3_outputs(7015) <= not a or b;
    layer3_outputs(7016) <= not (a and b);
    layer3_outputs(7017) <= a and not b;
    layer3_outputs(7018) <= a;
    layer3_outputs(7019) <= not a;
    layer3_outputs(7020) <= not b;
    layer3_outputs(7021) <= not b;
    layer3_outputs(7022) <= not b;
    layer3_outputs(7023) <= not b;
    layer3_outputs(7024) <= a;
    layer3_outputs(7025) <= not (a and b);
    layer3_outputs(7026) <= '0';
    layer3_outputs(7027) <= '0';
    layer3_outputs(7028) <= a and b;
    layer3_outputs(7029) <= not a or b;
    layer3_outputs(7030) <= a;
    layer3_outputs(7031) <= b and not a;
    layer3_outputs(7032) <= not (a and b);
    layer3_outputs(7033) <= not (a or b);
    layer3_outputs(7034) <= a and not b;
    layer3_outputs(7035) <= not a or b;
    layer3_outputs(7036) <= not b or a;
    layer3_outputs(7037) <= not (a or b);
    layer3_outputs(7038) <= a and b;
    layer3_outputs(7039) <= not a;
    layer3_outputs(7040) <= a;
    layer3_outputs(7041) <= a xor b;
    layer3_outputs(7042) <= not a or b;
    layer3_outputs(7043) <= a;
    layer3_outputs(7044) <= not a;
    layer3_outputs(7045) <= not b;
    layer3_outputs(7046) <= b and not a;
    layer3_outputs(7047) <= not (a xor b);
    layer3_outputs(7048) <= b;
    layer3_outputs(7049) <= not (a and b);
    layer3_outputs(7050) <= not (a and b);
    layer3_outputs(7051) <= not (a xor b);
    layer3_outputs(7052) <= a and not b;
    layer3_outputs(7053) <= b;
    layer3_outputs(7054) <= a;
    layer3_outputs(7055) <= not b;
    layer3_outputs(7056) <= not (a and b);
    layer3_outputs(7057) <= a and b;
    layer3_outputs(7058) <= b and not a;
    layer3_outputs(7059) <= not b;
    layer3_outputs(7060) <= not (a and b);
    layer3_outputs(7061) <= a;
    layer3_outputs(7062) <= a or b;
    layer3_outputs(7063) <= a;
    layer3_outputs(7064) <= a and not b;
    layer3_outputs(7065) <= b;
    layer3_outputs(7066) <= a;
    layer3_outputs(7067) <= a and b;
    layer3_outputs(7068) <= '0';
    layer3_outputs(7069) <= a and not b;
    layer3_outputs(7070) <= not a;
    layer3_outputs(7071) <= not (a or b);
    layer3_outputs(7072) <= not a;
    layer3_outputs(7073) <= a xor b;
    layer3_outputs(7074) <= b and not a;
    layer3_outputs(7075) <= not b or a;
    layer3_outputs(7076) <= a or b;
    layer3_outputs(7077) <= a;
    layer3_outputs(7078) <= not a;
    layer3_outputs(7079) <= not (a or b);
    layer3_outputs(7080) <= '1';
    layer3_outputs(7081) <= a and b;
    layer3_outputs(7082) <= '0';
    layer3_outputs(7083) <= a and b;
    layer3_outputs(7084) <= not (a or b);
    layer3_outputs(7085) <= not a;
    layer3_outputs(7086) <= not a or b;
    layer3_outputs(7087) <= not b or a;
    layer3_outputs(7088) <= a;
    layer3_outputs(7089) <= not b;
    layer3_outputs(7090) <= not (a or b);
    layer3_outputs(7091) <= not a;
    layer3_outputs(7092) <= b and not a;
    layer3_outputs(7093) <= not b or a;
    layer3_outputs(7094) <= not (a and b);
    layer3_outputs(7095) <= not b or a;
    layer3_outputs(7096) <= a and not b;
    layer3_outputs(7097) <= b and not a;
    layer3_outputs(7098) <= '0';
    layer3_outputs(7099) <= not a;
    layer3_outputs(7100) <= b and not a;
    layer3_outputs(7101) <= '1';
    layer3_outputs(7102) <= not b;
    layer3_outputs(7103) <= a xor b;
    layer3_outputs(7104) <= not a or b;
    layer3_outputs(7105) <= not a or b;
    layer3_outputs(7106) <= not (a or b);
    layer3_outputs(7107) <= a and not b;
    layer3_outputs(7108) <= not a;
    layer3_outputs(7109) <= a;
    layer3_outputs(7110) <= not (a or b);
    layer3_outputs(7111) <= not (a or b);
    layer3_outputs(7112) <= a;
    layer3_outputs(7113) <= a;
    layer3_outputs(7114) <= not b;
    layer3_outputs(7115) <= not (a and b);
    layer3_outputs(7116) <= a or b;
    layer3_outputs(7117) <= a and not b;
    layer3_outputs(7118) <= a and not b;
    layer3_outputs(7119) <= b;
    layer3_outputs(7120) <= not a;
    layer3_outputs(7121) <= b;
    layer3_outputs(7122) <= b;
    layer3_outputs(7123) <= '1';
    layer3_outputs(7124) <= a and not b;
    layer3_outputs(7125) <= not b;
    layer3_outputs(7126) <= a and not b;
    layer3_outputs(7127) <= b;
    layer3_outputs(7128) <= b;
    layer3_outputs(7129) <= not b;
    layer3_outputs(7130) <= '0';
    layer3_outputs(7131) <= b;
    layer3_outputs(7132) <= not (a or b);
    layer3_outputs(7133) <= '1';
    layer3_outputs(7134) <= not b or a;
    layer3_outputs(7135) <= a and not b;
    layer3_outputs(7136) <= a or b;
    layer3_outputs(7137) <= a;
    layer3_outputs(7138) <= b;
    layer3_outputs(7139) <= a and not b;
    layer3_outputs(7140) <= not b;
    layer3_outputs(7141) <= not a or b;
    layer3_outputs(7142) <= not (a and b);
    layer3_outputs(7143) <= not a;
    layer3_outputs(7144) <= a xor b;
    layer3_outputs(7145) <= not b or a;
    layer3_outputs(7146) <= a and b;
    layer3_outputs(7147) <= a;
    layer3_outputs(7148) <= '0';
    layer3_outputs(7149) <= not (a and b);
    layer3_outputs(7150) <= '1';
    layer3_outputs(7151) <= a xor b;
    layer3_outputs(7152) <= b;
    layer3_outputs(7153) <= a;
    layer3_outputs(7154) <= a;
    layer3_outputs(7155) <= a or b;
    layer3_outputs(7156) <= not a or b;
    layer3_outputs(7157) <= b;
    layer3_outputs(7158) <= a or b;
    layer3_outputs(7159) <= b;
    layer3_outputs(7160) <= not a or b;
    layer3_outputs(7161) <= not b;
    layer3_outputs(7162) <= '0';
    layer3_outputs(7163) <= b;
    layer3_outputs(7164) <= not a;
    layer3_outputs(7165) <= not b or a;
    layer3_outputs(7166) <= a;
    layer3_outputs(7167) <= not a;
    layer3_outputs(7168) <= b and not a;
    layer3_outputs(7169) <= b and not a;
    layer3_outputs(7170) <= not (a and b);
    layer3_outputs(7171) <= not a or b;
    layer3_outputs(7172) <= b and not a;
    layer3_outputs(7173) <= not b;
    layer3_outputs(7174) <= a and b;
    layer3_outputs(7175) <= a or b;
    layer3_outputs(7176) <= a;
    layer3_outputs(7177) <= not b;
    layer3_outputs(7178) <= not a;
    layer3_outputs(7179) <= not a;
    layer3_outputs(7180) <= a and b;
    layer3_outputs(7181) <= b and not a;
    layer3_outputs(7182) <= a and b;
    layer3_outputs(7183) <= not b or a;
    layer3_outputs(7184) <= b;
    layer3_outputs(7185) <= not a;
    layer3_outputs(7186) <= not a;
    layer3_outputs(7187) <= not a;
    layer3_outputs(7188) <= b and not a;
    layer3_outputs(7189) <= a or b;
    layer3_outputs(7190) <= not b;
    layer3_outputs(7191) <= a and b;
    layer3_outputs(7192) <= not a;
    layer3_outputs(7193) <= not b;
    layer3_outputs(7194) <= b and not a;
    layer3_outputs(7195) <= a and b;
    layer3_outputs(7196) <= a xor b;
    layer3_outputs(7197) <= not (a or b);
    layer3_outputs(7198) <= a xor b;
    layer3_outputs(7199) <= a;
    layer3_outputs(7200) <= a;
    layer3_outputs(7201) <= not a or b;
    layer3_outputs(7202) <= a or b;
    layer3_outputs(7203) <= '1';
    layer3_outputs(7204) <= not a;
    layer3_outputs(7205) <= not b;
    layer3_outputs(7206) <= not a;
    layer3_outputs(7207) <= a xor b;
    layer3_outputs(7208) <= not (a or b);
    layer3_outputs(7209) <= b;
    layer3_outputs(7210) <= b and not a;
    layer3_outputs(7211) <= b and not a;
    layer3_outputs(7212) <= not a;
    layer3_outputs(7213) <= b;
    layer3_outputs(7214) <= a or b;
    layer3_outputs(7215) <= not a or b;
    layer3_outputs(7216) <= a;
    layer3_outputs(7217) <= not (a and b);
    layer3_outputs(7218) <= b;
    layer3_outputs(7219) <= a;
    layer3_outputs(7220) <= not b;
    layer3_outputs(7221) <= not (a xor b);
    layer3_outputs(7222) <= not b or a;
    layer3_outputs(7223) <= '0';
    layer3_outputs(7224) <= not a;
    layer3_outputs(7225) <= '1';
    layer3_outputs(7226) <= not (a or b);
    layer3_outputs(7227) <= b;
    layer3_outputs(7228) <= a or b;
    layer3_outputs(7229) <= a xor b;
    layer3_outputs(7230) <= a and not b;
    layer3_outputs(7231) <= not (a and b);
    layer3_outputs(7232) <= b;
    layer3_outputs(7233) <= a and b;
    layer3_outputs(7234) <= not (a and b);
    layer3_outputs(7235) <= not b or a;
    layer3_outputs(7236) <= not (a and b);
    layer3_outputs(7237) <= a and not b;
    layer3_outputs(7238) <= b;
    layer3_outputs(7239) <= not a or b;
    layer3_outputs(7240) <= '0';
    layer3_outputs(7241) <= not b;
    layer3_outputs(7242) <= a and b;
    layer3_outputs(7243) <= not b;
    layer3_outputs(7244) <= not a or b;
    layer3_outputs(7245) <= not a;
    layer3_outputs(7246) <= not b;
    layer3_outputs(7247) <= '0';
    layer3_outputs(7248) <= b;
    layer3_outputs(7249) <= b;
    layer3_outputs(7250) <= not b or a;
    layer3_outputs(7251) <= b;
    layer3_outputs(7252) <= b;
    layer3_outputs(7253) <= a or b;
    layer3_outputs(7254) <= a xor b;
    layer3_outputs(7255) <= not a;
    layer3_outputs(7256) <= b and not a;
    layer3_outputs(7257) <= b;
    layer3_outputs(7258) <= '1';
    layer3_outputs(7259) <= not b;
    layer3_outputs(7260) <= not (a xor b);
    layer3_outputs(7261) <= not (a and b);
    layer3_outputs(7262) <= not b;
    layer3_outputs(7263) <= not a or b;
    layer3_outputs(7264) <= not (a or b);
    layer3_outputs(7265) <= not a;
    layer3_outputs(7266) <= a and b;
    layer3_outputs(7267) <= b;
    layer3_outputs(7268) <= not b;
    layer3_outputs(7269) <= a and b;
    layer3_outputs(7270) <= not a;
    layer3_outputs(7271) <= a;
    layer3_outputs(7272) <= b;
    layer3_outputs(7273) <= a and not b;
    layer3_outputs(7274) <= not b;
    layer3_outputs(7275) <= a and not b;
    layer3_outputs(7276) <= b and not a;
    layer3_outputs(7277) <= not (a and b);
    layer3_outputs(7278) <= a and not b;
    layer3_outputs(7279) <= a;
    layer3_outputs(7280) <= '0';
    layer3_outputs(7281) <= not a;
    layer3_outputs(7282) <= a or b;
    layer3_outputs(7283) <= not (a and b);
    layer3_outputs(7284) <= not b or a;
    layer3_outputs(7285) <= not b or a;
    layer3_outputs(7286) <= a and not b;
    layer3_outputs(7287) <= b;
    layer3_outputs(7288) <= a xor b;
    layer3_outputs(7289) <= b and not a;
    layer3_outputs(7290) <= not b;
    layer3_outputs(7291) <= '1';
    layer3_outputs(7292) <= a or b;
    layer3_outputs(7293) <= '0';
    layer3_outputs(7294) <= not b;
    layer3_outputs(7295) <= not (a and b);
    layer3_outputs(7296) <= not a;
    layer3_outputs(7297) <= b and not a;
    layer3_outputs(7298) <= not (a and b);
    layer3_outputs(7299) <= not (a or b);
    layer3_outputs(7300) <= not b or a;
    layer3_outputs(7301) <= a and not b;
    layer3_outputs(7302) <= not a;
    layer3_outputs(7303) <= not b;
    layer3_outputs(7304) <= not a;
    layer3_outputs(7305) <= a and b;
    layer3_outputs(7306) <= a;
    layer3_outputs(7307) <= b;
    layer3_outputs(7308) <= not b or a;
    layer3_outputs(7309) <= a;
    layer3_outputs(7310) <= a xor b;
    layer3_outputs(7311) <= a or b;
    layer3_outputs(7312) <= b and not a;
    layer3_outputs(7313) <= not a or b;
    layer3_outputs(7314) <= not b;
    layer3_outputs(7315) <= not (a and b);
    layer3_outputs(7316) <= not a or b;
    layer3_outputs(7317) <= not b or a;
    layer3_outputs(7318) <= a xor b;
    layer3_outputs(7319) <= not a or b;
    layer3_outputs(7320) <= '1';
    layer3_outputs(7321) <= not b;
    layer3_outputs(7322) <= not (a or b);
    layer3_outputs(7323) <= not b;
    layer3_outputs(7324) <= b;
    layer3_outputs(7325) <= not b;
    layer3_outputs(7326) <= '0';
    layer3_outputs(7327) <= a and b;
    layer3_outputs(7328) <= not (a or b);
    layer3_outputs(7329) <= not b;
    layer3_outputs(7330) <= not b;
    layer3_outputs(7331) <= not b or a;
    layer3_outputs(7332) <= not a or b;
    layer3_outputs(7333) <= not b;
    layer3_outputs(7334) <= not a;
    layer3_outputs(7335) <= not b;
    layer3_outputs(7336) <= b;
    layer3_outputs(7337) <= not (a and b);
    layer3_outputs(7338) <= '0';
    layer3_outputs(7339) <= not b;
    layer3_outputs(7340) <= '0';
    layer3_outputs(7341) <= not a;
    layer3_outputs(7342) <= a;
    layer3_outputs(7343) <= '1';
    layer3_outputs(7344) <= not (a or b);
    layer3_outputs(7345) <= a and not b;
    layer3_outputs(7346) <= not (a xor b);
    layer3_outputs(7347) <= a;
    layer3_outputs(7348) <= '1';
    layer3_outputs(7349) <= a;
    layer3_outputs(7350) <= not a;
    layer3_outputs(7351) <= '0';
    layer3_outputs(7352) <= not b or a;
    layer3_outputs(7353) <= not (a and b);
    layer3_outputs(7354) <= a;
    layer3_outputs(7355) <= not (a xor b);
    layer3_outputs(7356) <= not a or b;
    layer3_outputs(7357) <= not b or a;
    layer3_outputs(7358) <= not b or a;
    layer3_outputs(7359) <= '1';
    layer3_outputs(7360) <= not (a or b);
    layer3_outputs(7361) <= a;
    layer3_outputs(7362) <= a or b;
    layer3_outputs(7363) <= not (a xor b);
    layer3_outputs(7364) <= a xor b;
    layer3_outputs(7365) <= not a;
    layer3_outputs(7366) <= b;
    layer3_outputs(7367) <= b;
    layer3_outputs(7368) <= a and b;
    layer3_outputs(7369) <= b;
    layer3_outputs(7370) <= not b;
    layer3_outputs(7371) <= b and not a;
    layer3_outputs(7372) <= not a;
    layer3_outputs(7373) <= not (a or b);
    layer3_outputs(7374) <= a or b;
    layer3_outputs(7375) <= a and b;
    layer3_outputs(7376) <= not (a or b);
    layer3_outputs(7377) <= b and not a;
    layer3_outputs(7378) <= a xor b;
    layer3_outputs(7379) <= '1';
    layer3_outputs(7380) <= a and not b;
    layer3_outputs(7381) <= b;
    layer3_outputs(7382) <= not (a and b);
    layer3_outputs(7383) <= not (a or b);
    layer3_outputs(7384) <= '0';
    layer3_outputs(7385) <= not b;
    layer3_outputs(7386) <= not b;
    layer3_outputs(7387) <= not (a and b);
    layer3_outputs(7388) <= not (a or b);
    layer3_outputs(7389) <= not (a xor b);
    layer3_outputs(7390) <= not a or b;
    layer3_outputs(7391) <= '1';
    layer3_outputs(7392) <= a xor b;
    layer3_outputs(7393) <= a and b;
    layer3_outputs(7394) <= not b or a;
    layer3_outputs(7395) <= '1';
    layer3_outputs(7396) <= not b;
    layer3_outputs(7397) <= a or b;
    layer3_outputs(7398) <= a and not b;
    layer3_outputs(7399) <= a and not b;
    layer3_outputs(7400) <= a or b;
    layer3_outputs(7401) <= '1';
    layer3_outputs(7402) <= not b or a;
    layer3_outputs(7403) <= not (a and b);
    layer3_outputs(7404) <= b and not a;
    layer3_outputs(7405) <= a and b;
    layer3_outputs(7406) <= '1';
    layer3_outputs(7407) <= b and not a;
    layer3_outputs(7408) <= not a;
    layer3_outputs(7409) <= a and not b;
    layer3_outputs(7410) <= '0';
    layer3_outputs(7411) <= a or b;
    layer3_outputs(7412) <= not a;
    layer3_outputs(7413) <= a and not b;
    layer3_outputs(7414) <= a;
    layer3_outputs(7415) <= a and b;
    layer3_outputs(7416) <= a and not b;
    layer3_outputs(7417) <= not a;
    layer3_outputs(7418) <= a or b;
    layer3_outputs(7419) <= a xor b;
    layer3_outputs(7420) <= not (a or b);
    layer3_outputs(7421) <= a and not b;
    layer3_outputs(7422) <= a xor b;
    layer3_outputs(7423) <= b;
    layer3_outputs(7424) <= not a or b;
    layer3_outputs(7425) <= '0';
    layer3_outputs(7426) <= a;
    layer3_outputs(7427) <= not a or b;
    layer3_outputs(7428) <= a or b;
    layer3_outputs(7429) <= b and not a;
    layer3_outputs(7430) <= a or b;
    layer3_outputs(7431) <= not a;
    layer3_outputs(7432) <= '0';
    layer3_outputs(7433) <= not a or b;
    layer3_outputs(7434) <= not b;
    layer3_outputs(7435) <= not b or a;
    layer3_outputs(7436) <= a;
    layer3_outputs(7437) <= a xor b;
    layer3_outputs(7438) <= a and b;
    layer3_outputs(7439) <= '0';
    layer3_outputs(7440) <= '1';
    layer3_outputs(7441) <= not a;
    layer3_outputs(7442) <= not a;
    layer3_outputs(7443) <= '1';
    layer3_outputs(7444) <= not a or b;
    layer3_outputs(7445) <= not b or a;
    layer3_outputs(7446) <= b and not a;
    layer3_outputs(7447) <= a and b;
    layer3_outputs(7448) <= not a or b;
    layer3_outputs(7449) <= not (a or b);
    layer3_outputs(7450) <= a and b;
    layer3_outputs(7451) <= a or b;
    layer3_outputs(7452) <= not (a or b);
    layer3_outputs(7453) <= not (a and b);
    layer3_outputs(7454) <= not a or b;
    layer3_outputs(7455) <= not a;
    layer3_outputs(7456) <= a and not b;
    layer3_outputs(7457) <= not b;
    layer3_outputs(7458) <= not (a and b);
    layer3_outputs(7459) <= b and not a;
    layer3_outputs(7460) <= a xor b;
    layer3_outputs(7461) <= not a or b;
    layer3_outputs(7462) <= b and not a;
    layer3_outputs(7463) <= a;
    layer3_outputs(7464) <= '1';
    layer3_outputs(7465) <= a or b;
    layer3_outputs(7466) <= not a;
    layer3_outputs(7467) <= not b or a;
    layer3_outputs(7468) <= not a;
    layer3_outputs(7469) <= a and b;
    layer3_outputs(7470) <= not a or b;
    layer3_outputs(7471) <= a and b;
    layer3_outputs(7472) <= a or b;
    layer3_outputs(7473) <= not b;
    layer3_outputs(7474) <= not b;
    layer3_outputs(7475) <= not a;
    layer3_outputs(7476) <= b;
    layer3_outputs(7477) <= a;
    layer3_outputs(7478) <= not a or b;
    layer3_outputs(7479) <= a and not b;
    layer3_outputs(7480) <= '1';
    layer3_outputs(7481) <= b;
    layer3_outputs(7482) <= not a;
    layer3_outputs(7483) <= b and not a;
    layer3_outputs(7484) <= not a;
    layer3_outputs(7485) <= b and not a;
    layer3_outputs(7486) <= not b;
    layer3_outputs(7487) <= not a or b;
    layer3_outputs(7488) <= a xor b;
    layer3_outputs(7489) <= not (a or b);
    layer3_outputs(7490) <= not (a and b);
    layer3_outputs(7491) <= not (a and b);
    layer3_outputs(7492) <= not (a xor b);
    layer3_outputs(7493) <= b;
    layer3_outputs(7494) <= a;
    layer3_outputs(7495) <= not (a or b);
    layer3_outputs(7496) <= '0';
    layer3_outputs(7497) <= a and not b;
    layer3_outputs(7498) <= b and not a;
    layer3_outputs(7499) <= a or b;
    layer3_outputs(7500) <= a;
    layer3_outputs(7501) <= b;
    layer3_outputs(7502) <= a;
    layer3_outputs(7503) <= '1';
    layer3_outputs(7504) <= not b or a;
    layer3_outputs(7505) <= b;
    layer3_outputs(7506) <= b;
    layer3_outputs(7507) <= not (a xor b);
    layer3_outputs(7508) <= a xor b;
    layer3_outputs(7509) <= a and b;
    layer3_outputs(7510) <= b and not a;
    layer3_outputs(7511) <= not (a xor b);
    layer3_outputs(7512) <= not (a and b);
    layer3_outputs(7513) <= not b or a;
    layer3_outputs(7514) <= a;
    layer3_outputs(7515) <= not b or a;
    layer3_outputs(7516) <= not (a or b);
    layer3_outputs(7517) <= not a;
    layer3_outputs(7518) <= not (a and b);
    layer3_outputs(7519) <= not b or a;
    layer3_outputs(7520) <= a and b;
    layer3_outputs(7521) <= a;
    layer3_outputs(7522) <= a and b;
    layer3_outputs(7523) <= a xor b;
    layer3_outputs(7524) <= a;
    layer3_outputs(7525) <= a or b;
    layer3_outputs(7526) <= '1';
    layer3_outputs(7527) <= b;
    layer3_outputs(7528) <= not b or a;
    layer3_outputs(7529) <= not a;
    layer3_outputs(7530) <= not (a or b);
    layer3_outputs(7531) <= not a;
    layer3_outputs(7532) <= not b or a;
    layer3_outputs(7533) <= not (a or b);
    layer3_outputs(7534) <= not b or a;
    layer3_outputs(7535) <= not b or a;
    layer3_outputs(7536) <= a;
    layer3_outputs(7537) <= a;
    layer3_outputs(7538) <= not a or b;
    layer3_outputs(7539) <= a;
    layer3_outputs(7540) <= b;
    layer3_outputs(7541) <= '0';
    layer3_outputs(7542) <= a or b;
    layer3_outputs(7543) <= not a;
    layer3_outputs(7544) <= not (a or b);
    layer3_outputs(7545) <= not b;
    layer3_outputs(7546) <= '1';
    layer3_outputs(7547) <= not a;
    layer3_outputs(7548) <= not (a and b);
    layer3_outputs(7549) <= a and b;
    layer3_outputs(7550) <= '0';
    layer3_outputs(7551) <= a xor b;
    layer3_outputs(7552) <= a or b;
    layer3_outputs(7553) <= a;
    layer3_outputs(7554) <= not b;
    layer3_outputs(7555) <= not (a xor b);
    layer3_outputs(7556) <= a;
    layer3_outputs(7557) <= not (a and b);
    layer3_outputs(7558) <= not (a or b);
    layer3_outputs(7559) <= not (a or b);
    layer3_outputs(7560) <= not a;
    layer3_outputs(7561) <= b;
    layer3_outputs(7562) <= a and b;
    layer3_outputs(7563) <= '1';
    layer3_outputs(7564) <= not b;
    layer3_outputs(7565) <= b;
    layer3_outputs(7566) <= '1';
    layer3_outputs(7567) <= '1';
    layer3_outputs(7568) <= not (a or b);
    layer3_outputs(7569) <= b;
    layer3_outputs(7570) <= not a;
    layer3_outputs(7571) <= '0';
    layer3_outputs(7572) <= a;
    layer3_outputs(7573) <= a xor b;
    layer3_outputs(7574) <= not (a and b);
    layer3_outputs(7575) <= a;
    layer3_outputs(7576) <= a and not b;
    layer3_outputs(7577) <= not a or b;
    layer3_outputs(7578) <= b and not a;
    layer3_outputs(7579) <= a or b;
    layer3_outputs(7580) <= a and b;
    layer3_outputs(7581) <= b;
    layer3_outputs(7582) <= a;
    layer3_outputs(7583) <= b and not a;
    layer3_outputs(7584) <= a or b;
    layer3_outputs(7585) <= a and not b;
    layer3_outputs(7586) <= '1';
    layer3_outputs(7587) <= '1';
    layer3_outputs(7588) <= '1';
    layer3_outputs(7589) <= not (a or b);
    layer3_outputs(7590) <= a;
    layer3_outputs(7591) <= a;
    layer3_outputs(7592) <= b;
    layer3_outputs(7593) <= a and b;
    layer3_outputs(7594) <= not b;
    layer3_outputs(7595) <= a;
    layer3_outputs(7596) <= not b or a;
    layer3_outputs(7597) <= a and b;
    layer3_outputs(7598) <= not b;
    layer3_outputs(7599) <= '1';
    layer3_outputs(7600) <= not (a xor b);
    layer3_outputs(7601) <= b;
    layer3_outputs(7602) <= '0';
    layer3_outputs(7603) <= not a or b;
    layer3_outputs(7604) <= b and not a;
    layer3_outputs(7605) <= not b or a;
    layer3_outputs(7606) <= not b;
    layer3_outputs(7607) <= b;
    layer3_outputs(7608) <= b;
    layer3_outputs(7609) <= a or b;
    layer3_outputs(7610) <= not (a and b);
    layer3_outputs(7611) <= not (a and b);
    layer3_outputs(7612) <= not (a or b);
    layer3_outputs(7613) <= a and not b;
    layer3_outputs(7614) <= b;
    layer3_outputs(7615) <= a;
    layer3_outputs(7616) <= not b;
    layer3_outputs(7617) <= not a or b;
    layer3_outputs(7618) <= a and not b;
    layer3_outputs(7619) <= not a;
    layer3_outputs(7620) <= not b or a;
    layer3_outputs(7621) <= not a;
    layer3_outputs(7622) <= '0';
    layer3_outputs(7623) <= not a or b;
    layer3_outputs(7624) <= not a;
    layer3_outputs(7625) <= not b;
    layer3_outputs(7626) <= not (a or b);
    layer3_outputs(7627) <= not (a or b);
    layer3_outputs(7628) <= not a;
    layer3_outputs(7629) <= b and not a;
    layer3_outputs(7630) <= not (a or b);
    layer3_outputs(7631) <= '0';
    layer3_outputs(7632) <= not a or b;
    layer3_outputs(7633) <= a and not b;
    layer3_outputs(7634) <= b and not a;
    layer3_outputs(7635) <= not (a and b);
    layer3_outputs(7636) <= not a or b;
    layer3_outputs(7637) <= a;
    layer3_outputs(7638) <= a or b;
    layer3_outputs(7639) <= not b;
    layer3_outputs(7640) <= b;
    layer3_outputs(7641) <= b;
    layer3_outputs(7642) <= not b;
    layer3_outputs(7643) <= b;
    layer3_outputs(7644) <= not (a or b);
    layer3_outputs(7645) <= not (a xor b);
    layer3_outputs(7646) <= not (a and b);
    layer3_outputs(7647) <= a and not b;
    layer3_outputs(7648) <= not a;
    layer3_outputs(7649) <= b and not a;
    layer3_outputs(7650) <= a;
    layer3_outputs(7651) <= not a;
    layer3_outputs(7652) <= not a;
    layer3_outputs(7653) <= not (a xor b);
    layer3_outputs(7654) <= b;
    layer3_outputs(7655) <= b;
    layer3_outputs(7656) <= not (a or b);
    layer3_outputs(7657) <= b and not a;
    layer3_outputs(7658) <= not b;
    layer3_outputs(7659) <= not (a or b);
    layer3_outputs(7660) <= a;
    layer3_outputs(7661) <= b;
    layer3_outputs(7662) <= a and b;
    layer3_outputs(7663) <= not b;
    layer3_outputs(7664) <= not a;
    layer3_outputs(7665) <= not b;
    layer3_outputs(7666) <= not a or b;
    layer3_outputs(7667) <= b and not a;
    layer3_outputs(7668) <= not a;
    layer3_outputs(7669) <= a;
    layer3_outputs(7670) <= not a;
    layer3_outputs(7671) <= a or b;
    layer3_outputs(7672) <= a or b;
    layer3_outputs(7673) <= b;
    layer3_outputs(7674) <= not (a or b);
    layer3_outputs(7675) <= not b;
    layer3_outputs(7676) <= a and not b;
    layer3_outputs(7677) <= a and b;
    layer3_outputs(7678) <= not a;
    layer3_outputs(7679) <= not b;
    layer3_outputs(7680) <= a and b;
    layer3_outputs(7681) <= not (a and b);
    layer3_outputs(7682) <= not (a or b);
    layer3_outputs(7683) <= not (a or b);
    layer3_outputs(7684) <= '0';
    layer3_outputs(7685) <= '0';
    layer3_outputs(7686) <= not b;
    layer3_outputs(7687) <= not (a or b);
    layer3_outputs(7688) <= not a or b;
    layer3_outputs(7689) <= '1';
    layer3_outputs(7690) <= a and b;
    layer3_outputs(7691) <= not a;
    layer3_outputs(7692) <= b;
    layer3_outputs(7693) <= a and not b;
    layer3_outputs(7694) <= not a;
    layer3_outputs(7695) <= not b or a;
    layer3_outputs(7696) <= a and b;
    layer3_outputs(7697) <= b and not a;
    layer3_outputs(7698) <= b and not a;
    layer3_outputs(7699) <= not (a and b);
    layer3_outputs(7700) <= not (a xor b);
    layer3_outputs(7701) <= not (a or b);
    layer3_outputs(7702) <= not b or a;
    layer3_outputs(7703) <= '0';
    layer3_outputs(7704) <= a or b;
    layer3_outputs(7705) <= not (a xor b);
    layer3_outputs(7706) <= b;
    layer3_outputs(7707) <= not (a and b);
    layer3_outputs(7708) <= not b;
    layer3_outputs(7709) <= not b or a;
    layer3_outputs(7710) <= '0';
    layer3_outputs(7711) <= not a;
    layer3_outputs(7712) <= a;
    layer3_outputs(7713) <= not (a and b);
    layer3_outputs(7714) <= not a;
    layer3_outputs(7715) <= a;
    layer3_outputs(7716) <= b;
    layer3_outputs(7717) <= a or b;
    layer3_outputs(7718) <= b;
    layer3_outputs(7719) <= not b or a;
    layer3_outputs(7720) <= not a;
    layer3_outputs(7721) <= not b;
    layer3_outputs(7722) <= not a;
    layer3_outputs(7723) <= a and not b;
    layer3_outputs(7724) <= a xor b;
    layer3_outputs(7725) <= not a;
    layer3_outputs(7726) <= not (a or b);
    layer3_outputs(7727) <= a and not b;
    layer3_outputs(7728) <= not b or a;
    layer3_outputs(7729) <= b;
    layer3_outputs(7730) <= a;
    layer3_outputs(7731) <= '0';
    layer3_outputs(7732) <= '0';
    layer3_outputs(7733) <= a xor b;
    layer3_outputs(7734) <= not a;
    layer3_outputs(7735) <= not b;
    layer3_outputs(7736) <= b;
    layer3_outputs(7737) <= not a;
    layer3_outputs(7738) <= a xor b;
    layer3_outputs(7739) <= b and not a;
    layer3_outputs(7740) <= not (a or b);
    layer3_outputs(7741) <= a;
    layer3_outputs(7742) <= not b or a;
    layer3_outputs(7743) <= a and b;
    layer3_outputs(7744) <= not (a or b);
    layer3_outputs(7745) <= not b;
    layer3_outputs(7746) <= not a;
    layer3_outputs(7747) <= a or b;
    layer3_outputs(7748) <= '1';
    layer3_outputs(7749) <= a;
    layer3_outputs(7750) <= not b;
    layer3_outputs(7751) <= not b;
    layer3_outputs(7752) <= a xor b;
    layer3_outputs(7753) <= b and not a;
    layer3_outputs(7754) <= not (a and b);
    layer3_outputs(7755) <= not a;
    layer3_outputs(7756) <= not (a or b);
    layer3_outputs(7757) <= not b or a;
    layer3_outputs(7758) <= a;
    layer3_outputs(7759) <= b;
    layer3_outputs(7760) <= a and b;
    layer3_outputs(7761) <= not a;
    layer3_outputs(7762) <= not a or b;
    layer3_outputs(7763) <= a or b;
    layer3_outputs(7764) <= not (a and b);
    layer3_outputs(7765) <= a or b;
    layer3_outputs(7766) <= b and not a;
    layer3_outputs(7767) <= '0';
    layer3_outputs(7768) <= not b;
    layer3_outputs(7769) <= not a;
    layer3_outputs(7770) <= a and not b;
    layer3_outputs(7771) <= not a or b;
    layer3_outputs(7772) <= b;
    layer3_outputs(7773) <= a xor b;
    layer3_outputs(7774) <= not (a and b);
    layer3_outputs(7775) <= b and not a;
    layer3_outputs(7776) <= not (a or b);
    layer3_outputs(7777) <= not (a or b);
    layer3_outputs(7778) <= a and b;
    layer3_outputs(7779) <= b and not a;
    layer3_outputs(7780) <= '0';
    layer3_outputs(7781) <= not (a xor b);
    layer3_outputs(7782) <= not (a or b);
    layer3_outputs(7783) <= b and not a;
    layer3_outputs(7784) <= a or b;
    layer3_outputs(7785) <= not b or a;
    layer3_outputs(7786) <= b and not a;
    layer3_outputs(7787) <= not (a and b);
    layer3_outputs(7788) <= a or b;
    layer3_outputs(7789) <= not a;
    layer3_outputs(7790) <= a and not b;
    layer3_outputs(7791) <= '0';
    layer3_outputs(7792) <= a;
    layer3_outputs(7793) <= not a;
    layer3_outputs(7794) <= b and not a;
    layer3_outputs(7795) <= a or b;
    layer3_outputs(7796) <= b and not a;
    layer3_outputs(7797) <= b and not a;
    layer3_outputs(7798) <= not a;
    layer3_outputs(7799) <= not (a or b);
    layer3_outputs(7800) <= not b or a;
    layer3_outputs(7801) <= '0';
    layer3_outputs(7802) <= a and b;
    layer3_outputs(7803) <= a xor b;
    layer3_outputs(7804) <= not a or b;
    layer3_outputs(7805) <= not (a and b);
    layer3_outputs(7806) <= b and not a;
    layer3_outputs(7807) <= '0';
    layer3_outputs(7808) <= b;
    layer3_outputs(7809) <= a and not b;
    layer3_outputs(7810) <= not a;
    layer3_outputs(7811) <= not (a and b);
    layer3_outputs(7812) <= a;
    layer3_outputs(7813) <= a;
    layer3_outputs(7814) <= a xor b;
    layer3_outputs(7815) <= not a;
    layer3_outputs(7816) <= not a;
    layer3_outputs(7817) <= b and not a;
    layer3_outputs(7818) <= not a;
    layer3_outputs(7819) <= a and b;
    layer3_outputs(7820) <= not a or b;
    layer3_outputs(7821) <= b;
    layer3_outputs(7822) <= not b;
    layer3_outputs(7823) <= a and not b;
    layer3_outputs(7824) <= not a or b;
    layer3_outputs(7825) <= b;
    layer3_outputs(7826) <= a or b;
    layer3_outputs(7827) <= not a;
    layer3_outputs(7828) <= a;
    layer3_outputs(7829) <= not b or a;
    layer3_outputs(7830) <= not a;
    layer3_outputs(7831) <= b;
    layer3_outputs(7832) <= not b or a;
    layer3_outputs(7833) <= not b;
    layer3_outputs(7834) <= '1';
    layer3_outputs(7835) <= b;
    layer3_outputs(7836) <= a;
    layer3_outputs(7837) <= a;
    layer3_outputs(7838) <= a xor b;
    layer3_outputs(7839) <= b;
    layer3_outputs(7840) <= not b or a;
    layer3_outputs(7841) <= b and not a;
    layer3_outputs(7842) <= b;
    layer3_outputs(7843) <= b;
    layer3_outputs(7844) <= a and b;
    layer3_outputs(7845) <= a or b;
    layer3_outputs(7846) <= not b or a;
    layer3_outputs(7847) <= not b or a;
    layer3_outputs(7848) <= a or b;
    layer3_outputs(7849) <= a;
    layer3_outputs(7850) <= '0';
    layer3_outputs(7851) <= not (a and b);
    layer3_outputs(7852) <= not (a xor b);
    layer3_outputs(7853) <= not a or b;
    layer3_outputs(7854) <= not b;
    layer3_outputs(7855) <= not b;
    layer3_outputs(7856) <= a and not b;
    layer3_outputs(7857) <= a xor b;
    layer3_outputs(7858) <= not (a or b);
    layer3_outputs(7859) <= not b;
    layer3_outputs(7860) <= b;
    layer3_outputs(7861) <= a and b;
    layer3_outputs(7862) <= not b;
    layer3_outputs(7863) <= a;
    layer3_outputs(7864) <= a and not b;
    layer3_outputs(7865) <= a and not b;
    layer3_outputs(7866) <= not b;
    layer3_outputs(7867) <= not (a or b);
    layer3_outputs(7868) <= not (a and b);
    layer3_outputs(7869) <= a or b;
    layer3_outputs(7870) <= a or b;
    layer3_outputs(7871) <= a and not b;
    layer3_outputs(7872) <= '0';
    layer3_outputs(7873) <= not (a xor b);
    layer3_outputs(7874) <= a and b;
    layer3_outputs(7875) <= a and not b;
    layer3_outputs(7876) <= not b;
    layer3_outputs(7877) <= a and b;
    layer3_outputs(7878) <= a xor b;
    layer3_outputs(7879) <= b and not a;
    layer3_outputs(7880) <= '1';
    layer3_outputs(7881) <= not (a xor b);
    layer3_outputs(7882) <= b;
    layer3_outputs(7883) <= a or b;
    layer3_outputs(7884) <= not (a xor b);
    layer3_outputs(7885) <= not (a and b);
    layer3_outputs(7886) <= not b or a;
    layer3_outputs(7887) <= a and b;
    layer3_outputs(7888) <= a and not b;
    layer3_outputs(7889) <= not b;
    layer3_outputs(7890) <= not b;
    layer3_outputs(7891) <= b and not a;
    layer3_outputs(7892) <= a;
    layer3_outputs(7893) <= a or b;
    layer3_outputs(7894) <= not (a or b);
    layer3_outputs(7895) <= not (a xor b);
    layer3_outputs(7896) <= not (a and b);
    layer3_outputs(7897) <= not a;
    layer3_outputs(7898) <= a or b;
    layer3_outputs(7899) <= a and b;
    layer3_outputs(7900) <= a;
    layer3_outputs(7901) <= not (a or b);
    layer3_outputs(7902) <= a xor b;
    layer3_outputs(7903) <= not (a xor b);
    layer3_outputs(7904) <= a and not b;
    layer3_outputs(7905) <= a;
    layer3_outputs(7906) <= not b;
    layer3_outputs(7907) <= not b;
    layer3_outputs(7908) <= a;
    layer3_outputs(7909) <= b;
    layer3_outputs(7910) <= '1';
    layer3_outputs(7911) <= a;
    layer3_outputs(7912) <= not b or a;
    layer3_outputs(7913) <= a or b;
    layer3_outputs(7914) <= a or b;
    layer3_outputs(7915) <= not (a xor b);
    layer3_outputs(7916) <= not a or b;
    layer3_outputs(7917) <= not b or a;
    layer3_outputs(7918) <= a;
    layer3_outputs(7919) <= not a or b;
    layer3_outputs(7920) <= '0';
    layer3_outputs(7921) <= '1';
    layer3_outputs(7922) <= '0';
    layer3_outputs(7923) <= a and not b;
    layer3_outputs(7924) <= '1';
    layer3_outputs(7925) <= a or b;
    layer3_outputs(7926) <= not (a or b);
    layer3_outputs(7927) <= a or b;
    layer3_outputs(7928) <= not a;
    layer3_outputs(7929) <= not (a xor b);
    layer3_outputs(7930) <= not b;
    layer3_outputs(7931) <= b and not a;
    layer3_outputs(7932) <= not b;
    layer3_outputs(7933) <= b and not a;
    layer3_outputs(7934) <= a and b;
    layer3_outputs(7935) <= not (a and b);
    layer3_outputs(7936) <= b;
    layer3_outputs(7937) <= a and b;
    layer3_outputs(7938) <= b and not a;
    layer3_outputs(7939) <= a;
    layer3_outputs(7940) <= not (a and b);
    layer3_outputs(7941) <= b;
    layer3_outputs(7942) <= not (a and b);
    layer3_outputs(7943) <= b and not a;
    layer3_outputs(7944) <= not (a or b);
    layer3_outputs(7945) <= not (a and b);
    layer3_outputs(7946) <= a or b;
    layer3_outputs(7947) <= not (a or b);
    layer3_outputs(7948) <= not (a or b);
    layer3_outputs(7949) <= not (a and b);
    layer3_outputs(7950) <= a and b;
    layer3_outputs(7951) <= '0';
    layer3_outputs(7952) <= not b;
    layer3_outputs(7953) <= a or b;
    layer3_outputs(7954) <= not b;
    layer3_outputs(7955) <= not b;
    layer3_outputs(7956) <= not b;
    layer3_outputs(7957) <= not a or b;
    layer3_outputs(7958) <= '1';
    layer3_outputs(7959) <= a;
    layer3_outputs(7960) <= b;
    layer3_outputs(7961) <= '0';
    layer3_outputs(7962) <= not b or a;
    layer3_outputs(7963) <= not (a xor b);
    layer3_outputs(7964) <= a and b;
    layer3_outputs(7965) <= not (a and b);
    layer3_outputs(7966) <= not (a xor b);
    layer3_outputs(7967) <= not b;
    layer3_outputs(7968) <= b;
    layer3_outputs(7969) <= a and not b;
    layer3_outputs(7970) <= '1';
    layer3_outputs(7971) <= a and b;
    layer3_outputs(7972) <= b;
    layer3_outputs(7973) <= not a or b;
    layer3_outputs(7974) <= a or b;
    layer3_outputs(7975) <= a and not b;
    layer3_outputs(7976) <= not a or b;
    layer3_outputs(7977) <= b and not a;
    layer3_outputs(7978) <= a and b;
    layer3_outputs(7979) <= b and not a;
    layer3_outputs(7980) <= not (a and b);
    layer3_outputs(7981) <= a;
    layer3_outputs(7982) <= not a or b;
    layer3_outputs(7983) <= not b;
    layer3_outputs(7984) <= a xor b;
    layer3_outputs(7985) <= not b;
    layer3_outputs(7986) <= not a or b;
    layer3_outputs(7987) <= a xor b;
    layer3_outputs(7988) <= a;
    layer3_outputs(7989) <= not b or a;
    layer3_outputs(7990) <= not a;
    layer3_outputs(7991) <= b;
    layer3_outputs(7992) <= a;
    layer3_outputs(7993) <= not a;
    layer3_outputs(7994) <= '0';
    layer3_outputs(7995) <= not b or a;
    layer3_outputs(7996) <= not b or a;
    layer3_outputs(7997) <= not b;
    layer3_outputs(7998) <= not b or a;
    layer3_outputs(7999) <= not (a and b);
    layer3_outputs(8000) <= a xor b;
    layer3_outputs(8001) <= b;
    layer3_outputs(8002) <= a or b;
    layer3_outputs(8003) <= a or b;
    layer3_outputs(8004) <= not a;
    layer3_outputs(8005) <= a;
    layer3_outputs(8006) <= not b;
    layer3_outputs(8007) <= not b or a;
    layer3_outputs(8008) <= not b or a;
    layer3_outputs(8009) <= a and not b;
    layer3_outputs(8010) <= not (a xor b);
    layer3_outputs(8011) <= '0';
    layer3_outputs(8012) <= not b or a;
    layer3_outputs(8013) <= not (a xor b);
    layer3_outputs(8014) <= not a or b;
    layer3_outputs(8015) <= a;
    layer3_outputs(8016) <= not (a xor b);
    layer3_outputs(8017) <= not b;
    layer3_outputs(8018) <= not a;
    layer3_outputs(8019) <= not (a or b);
    layer3_outputs(8020) <= '1';
    layer3_outputs(8021) <= not (a and b);
    layer3_outputs(8022) <= '1';
    layer3_outputs(8023) <= not (a xor b);
    layer3_outputs(8024) <= a and not b;
    layer3_outputs(8025) <= b and not a;
    layer3_outputs(8026) <= not (a and b);
    layer3_outputs(8027) <= not (a and b);
    layer3_outputs(8028) <= not a;
    layer3_outputs(8029) <= a xor b;
    layer3_outputs(8030) <= '1';
    layer3_outputs(8031) <= a or b;
    layer3_outputs(8032) <= not (a xor b);
    layer3_outputs(8033) <= a;
    layer3_outputs(8034) <= a;
    layer3_outputs(8035) <= not (a or b);
    layer3_outputs(8036) <= b;
    layer3_outputs(8037) <= not (a or b);
    layer3_outputs(8038) <= b and not a;
    layer3_outputs(8039) <= a and not b;
    layer3_outputs(8040) <= b and not a;
    layer3_outputs(8041) <= b;
    layer3_outputs(8042) <= not b;
    layer3_outputs(8043) <= a;
    layer3_outputs(8044) <= b and not a;
    layer3_outputs(8045) <= a or b;
    layer3_outputs(8046) <= '1';
    layer3_outputs(8047) <= b and not a;
    layer3_outputs(8048) <= not b;
    layer3_outputs(8049) <= b;
    layer3_outputs(8050) <= not a;
    layer3_outputs(8051) <= not a;
    layer3_outputs(8052) <= not b;
    layer3_outputs(8053) <= a and b;
    layer3_outputs(8054) <= a and not b;
    layer3_outputs(8055) <= a and b;
    layer3_outputs(8056) <= not b;
    layer3_outputs(8057) <= b and not a;
    layer3_outputs(8058) <= a xor b;
    layer3_outputs(8059) <= b and not a;
    layer3_outputs(8060) <= a and not b;
    layer3_outputs(8061) <= '1';
    layer3_outputs(8062) <= a and b;
    layer3_outputs(8063) <= b and not a;
    layer3_outputs(8064) <= not a;
    layer3_outputs(8065) <= not b;
    layer3_outputs(8066) <= a;
    layer3_outputs(8067) <= not a or b;
    layer3_outputs(8068) <= not (a and b);
    layer3_outputs(8069) <= a;
    layer3_outputs(8070) <= a or b;
    layer3_outputs(8071) <= a or b;
    layer3_outputs(8072) <= a or b;
    layer3_outputs(8073) <= not a;
    layer3_outputs(8074) <= '1';
    layer3_outputs(8075) <= a and b;
    layer3_outputs(8076) <= not a;
    layer3_outputs(8077) <= not (a and b);
    layer3_outputs(8078) <= b and not a;
    layer3_outputs(8079) <= not a;
    layer3_outputs(8080) <= a and b;
    layer3_outputs(8081) <= not a;
    layer3_outputs(8082) <= '1';
    layer3_outputs(8083) <= a and not b;
    layer3_outputs(8084) <= not b or a;
    layer3_outputs(8085) <= '1';
    layer3_outputs(8086) <= '0';
    layer3_outputs(8087) <= b and not a;
    layer3_outputs(8088) <= a;
    layer3_outputs(8089) <= not a;
    layer3_outputs(8090) <= not b;
    layer3_outputs(8091) <= not b;
    layer3_outputs(8092) <= a or b;
    layer3_outputs(8093) <= a and b;
    layer3_outputs(8094) <= a;
    layer3_outputs(8095) <= b;
    layer3_outputs(8096) <= not b or a;
    layer3_outputs(8097) <= not b;
    layer3_outputs(8098) <= not a or b;
    layer3_outputs(8099) <= '0';
    layer3_outputs(8100) <= a xor b;
    layer3_outputs(8101) <= b and not a;
    layer3_outputs(8102) <= '1';
    layer3_outputs(8103) <= a;
    layer3_outputs(8104) <= not b;
    layer3_outputs(8105) <= a and b;
    layer3_outputs(8106) <= not (a and b);
    layer3_outputs(8107) <= b;
    layer3_outputs(8108) <= a;
    layer3_outputs(8109) <= not a or b;
    layer3_outputs(8110) <= a and not b;
    layer3_outputs(8111) <= b;
    layer3_outputs(8112) <= b;
    layer3_outputs(8113) <= a or b;
    layer3_outputs(8114) <= not b;
    layer3_outputs(8115) <= not b;
    layer3_outputs(8116) <= a xor b;
    layer3_outputs(8117) <= a and not b;
    layer3_outputs(8118) <= not a or b;
    layer3_outputs(8119) <= not b;
    layer3_outputs(8120) <= a;
    layer3_outputs(8121) <= a and b;
    layer3_outputs(8122) <= not (a or b);
    layer3_outputs(8123) <= b and not a;
    layer3_outputs(8124) <= not (a and b);
    layer3_outputs(8125) <= not a;
    layer3_outputs(8126) <= b;
    layer3_outputs(8127) <= b and not a;
    layer3_outputs(8128) <= not a;
    layer3_outputs(8129) <= not b;
    layer3_outputs(8130) <= '1';
    layer3_outputs(8131) <= b;
    layer3_outputs(8132) <= not a;
    layer3_outputs(8133) <= a or b;
    layer3_outputs(8134) <= not b;
    layer3_outputs(8135) <= not (a or b);
    layer3_outputs(8136) <= not b or a;
    layer3_outputs(8137) <= b;
    layer3_outputs(8138) <= not a or b;
    layer3_outputs(8139) <= not b;
    layer3_outputs(8140) <= a and b;
    layer3_outputs(8141) <= not (a or b);
    layer3_outputs(8142) <= not b;
    layer3_outputs(8143) <= not (a or b);
    layer3_outputs(8144) <= not a;
    layer3_outputs(8145) <= b;
    layer3_outputs(8146) <= not b;
    layer3_outputs(8147) <= not (a and b);
    layer3_outputs(8148) <= a or b;
    layer3_outputs(8149) <= a and not b;
    layer3_outputs(8150) <= a and b;
    layer3_outputs(8151) <= b and not a;
    layer3_outputs(8152) <= not b;
    layer3_outputs(8153) <= not (a or b);
    layer3_outputs(8154) <= b;
    layer3_outputs(8155) <= '0';
    layer3_outputs(8156) <= not b or a;
    layer3_outputs(8157) <= not b or a;
    layer3_outputs(8158) <= not b;
    layer3_outputs(8159) <= not (a or b);
    layer3_outputs(8160) <= not b;
    layer3_outputs(8161) <= '0';
    layer3_outputs(8162) <= not b;
    layer3_outputs(8163) <= '0';
    layer3_outputs(8164) <= b;
    layer3_outputs(8165) <= b;
    layer3_outputs(8166) <= not b;
    layer3_outputs(8167) <= not a or b;
    layer3_outputs(8168) <= not a;
    layer3_outputs(8169) <= not (a or b);
    layer3_outputs(8170) <= not b;
    layer3_outputs(8171) <= a and b;
    layer3_outputs(8172) <= a or b;
    layer3_outputs(8173) <= b;
    layer3_outputs(8174) <= '0';
    layer3_outputs(8175) <= not a;
    layer3_outputs(8176) <= not a;
    layer3_outputs(8177) <= not b;
    layer3_outputs(8178) <= a and b;
    layer3_outputs(8179) <= not a;
    layer3_outputs(8180) <= b and not a;
    layer3_outputs(8181) <= a xor b;
    layer3_outputs(8182) <= a xor b;
    layer3_outputs(8183) <= b and not a;
    layer3_outputs(8184) <= not b;
    layer3_outputs(8185) <= b;
    layer3_outputs(8186) <= not a;
    layer3_outputs(8187) <= not b;
    layer3_outputs(8188) <= a xor b;
    layer3_outputs(8189) <= a;
    layer3_outputs(8190) <= a xor b;
    layer3_outputs(8191) <= '0';
    layer3_outputs(8192) <= a;
    layer3_outputs(8193) <= '1';
    layer3_outputs(8194) <= a;
    layer3_outputs(8195) <= a and b;
    layer3_outputs(8196) <= not b;
    layer3_outputs(8197) <= a and b;
    layer3_outputs(8198) <= '1';
    layer3_outputs(8199) <= not a;
    layer3_outputs(8200) <= b;
    layer3_outputs(8201) <= a and not b;
    layer3_outputs(8202) <= not (a xor b);
    layer3_outputs(8203) <= not a or b;
    layer3_outputs(8204) <= not b;
    layer3_outputs(8205) <= b;
    layer3_outputs(8206) <= not b;
    layer3_outputs(8207) <= '1';
    layer3_outputs(8208) <= b and not a;
    layer3_outputs(8209) <= b and not a;
    layer3_outputs(8210) <= not a or b;
    layer3_outputs(8211) <= a xor b;
    layer3_outputs(8212) <= a and b;
    layer3_outputs(8213) <= a and b;
    layer3_outputs(8214) <= b;
    layer3_outputs(8215) <= not b or a;
    layer3_outputs(8216) <= b and not a;
    layer3_outputs(8217) <= not (a and b);
    layer3_outputs(8218) <= not (a or b);
    layer3_outputs(8219) <= not b;
    layer3_outputs(8220) <= b and not a;
    layer3_outputs(8221) <= a;
    layer3_outputs(8222) <= '1';
    layer3_outputs(8223) <= not a;
    layer3_outputs(8224) <= a;
    layer3_outputs(8225) <= a or b;
    layer3_outputs(8226) <= a or b;
    layer3_outputs(8227) <= not b;
    layer3_outputs(8228) <= not (a and b);
    layer3_outputs(8229) <= not a;
    layer3_outputs(8230) <= not (a or b);
    layer3_outputs(8231) <= '0';
    layer3_outputs(8232) <= a and b;
    layer3_outputs(8233) <= a and not b;
    layer3_outputs(8234) <= a or b;
    layer3_outputs(8235) <= a or b;
    layer3_outputs(8236) <= not (a or b);
    layer3_outputs(8237) <= a or b;
    layer3_outputs(8238) <= a or b;
    layer3_outputs(8239) <= b and not a;
    layer3_outputs(8240) <= not b or a;
    layer3_outputs(8241) <= a and not b;
    layer3_outputs(8242) <= a;
    layer3_outputs(8243) <= a;
    layer3_outputs(8244) <= not (a or b);
    layer3_outputs(8245) <= '1';
    layer3_outputs(8246) <= not a;
    layer3_outputs(8247) <= a or b;
    layer3_outputs(8248) <= a and b;
    layer3_outputs(8249) <= a;
    layer3_outputs(8250) <= b and not a;
    layer3_outputs(8251) <= a and not b;
    layer3_outputs(8252) <= not (a xor b);
    layer3_outputs(8253) <= a and b;
    layer3_outputs(8254) <= not (a and b);
    layer3_outputs(8255) <= not b or a;
    layer3_outputs(8256) <= not a;
    layer3_outputs(8257) <= a or b;
    layer3_outputs(8258) <= a xor b;
    layer3_outputs(8259) <= a and not b;
    layer3_outputs(8260) <= b and not a;
    layer3_outputs(8261) <= a;
    layer3_outputs(8262) <= a;
    layer3_outputs(8263) <= not a;
    layer3_outputs(8264) <= not (a and b);
    layer3_outputs(8265) <= a and b;
    layer3_outputs(8266) <= a or b;
    layer3_outputs(8267) <= a;
    layer3_outputs(8268) <= not (a or b);
    layer3_outputs(8269) <= not (a or b);
    layer3_outputs(8270) <= not b or a;
    layer3_outputs(8271) <= a and not b;
    layer3_outputs(8272) <= not b or a;
    layer3_outputs(8273) <= not b or a;
    layer3_outputs(8274) <= not (a and b);
    layer3_outputs(8275) <= not a;
    layer3_outputs(8276) <= not (a or b);
    layer3_outputs(8277) <= a and not b;
    layer3_outputs(8278) <= not b;
    layer3_outputs(8279) <= not (a and b);
    layer3_outputs(8280) <= a and not b;
    layer3_outputs(8281) <= b and not a;
    layer3_outputs(8282) <= not (a or b);
    layer3_outputs(8283) <= '1';
    layer3_outputs(8284) <= b and not a;
    layer3_outputs(8285) <= not b or a;
    layer3_outputs(8286) <= not a or b;
    layer3_outputs(8287) <= a or b;
    layer3_outputs(8288) <= b and not a;
    layer3_outputs(8289) <= a and not b;
    layer3_outputs(8290) <= b;
    layer3_outputs(8291) <= '1';
    layer3_outputs(8292) <= a or b;
    layer3_outputs(8293) <= not a;
    layer3_outputs(8294) <= b and not a;
    layer3_outputs(8295) <= a;
    layer3_outputs(8296) <= not (a xor b);
    layer3_outputs(8297) <= not a or b;
    layer3_outputs(8298) <= a;
    layer3_outputs(8299) <= not (a or b);
    layer3_outputs(8300) <= a or b;
    layer3_outputs(8301) <= not b or a;
    layer3_outputs(8302) <= not a;
    layer3_outputs(8303) <= a;
    layer3_outputs(8304) <= not a or b;
    layer3_outputs(8305) <= a xor b;
    layer3_outputs(8306) <= a;
    layer3_outputs(8307) <= '1';
    layer3_outputs(8308) <= a xor b;
    layer3_outputs(8309) <= not a;
    layer3_outputs(8310) <= b;
    layer3_outputs(8311) <= '1';
    layer3_outputs(8312) <= not (a xor b);
    layer3_outputs(8313) <= b and not a;
    layer3_outputs(8314) <= a and not b;
    layer3_outputs(8315) <= a;
    layer3_outputs(8316) <= '0';
    layer3_outputs(8317) <= not b or a;
    layer3_outputs(8318) <= not b or a;
    layer3_outputs(8319) <= b;
    layer3_outputs(8320) <= not (a and b);
    layer3_outputs(8321) <= not b;
    layer3_outputs(8322) <= a xor b;
    layer3_outputs(8323) <= a and b;
    layer3_outputs(8324) <= a and not b;
    layer3_outputs(8325) <= a or b;
    layer3_outputs(8326) <= not a;
    layer3_outputs(8327) <= a or b;
    layer3_outputs(8328) <= not a or b;
    layer3_outputs(8329) <= not b;
    layer3_outputs(8330) <= a;
    layer3_outputs(8331) <= a or b;
    layer3_outputs(8332) <= a xor b;
    layer3_outputs(8333) <= a and not b;
    layer3_outputs(8334) <= not (a and b);
    layer3_outputs(8335) <= not (a and b);
    layer3_outputs(8336) <= a or b;
    layer3_outputs(8337) <= a and not b;
    layer3_outputs(8338) <= b;
    layer3_outputs(8339) <= not (a and b);
    layer3_outputs(8340) <= '1';
    layer3_outputs(8341) <= a xor b;
    layer3_outputs(8342) <= not b or a;
    layer3_outputs(8343) <= not b;
    layer3_outputs(8344) <= a;
    layer3_outputs(8345) <= not b;
    layer3_outputs(8346) <= a and not b;
    layer3_outputs(8347) <= a xor b;
    layer3_outputs(8348) <= a or b;
    layer3_outputs(8349) <= a and b;
    layer3_outputs(8350) <= a and b;
    layer3_outputs(8351) <= a;
    layer3_outputs(8352) <= not a;
    layer3_outputs(8353) <= a xor b;
    layer3_outputs(8354) <= b and not a;
    layer3_outputs(8355) <= not b or a;
    layer3_outputs(8356) <= b;
    layer3_outputs(8357) <= not b;
    layer3_outputs(8358) <= b and not a;
    layer3_outputs(8359) <= not a;
    layer3_outputs(8360) <= not a;
    layer3_outputs(8361) <= not b;
    layer3_outputs(8362) <= not a or b;
    layer3_outputs(8363) <= not a;
    layer3_outputs(8364) <= '1';
    layer3_outputs(8365) <= not a or b;
    layer3_outputs(8366) <= not a or b;
    layer3_outputs(8367) <= a xor b;
    layer3_outputs(8368) <= b;
    layer3_outputs(8369) <= '0';
    layer3_outputs(8370) <= not a;
    layer3_outputs(8371) <= not a;
    layer3_outputs(8372) <= a or b;
    layer3_outputs(8373) <= a or b;
    layer3_outputs(8374) <= not (a and b);
    layer3_outputs(8375) <= b and not a;
    layer3_outputs(8376) <= b and not a;
    layer3_outputs(8377) <= b;
    layer3_outputs(8378) <= a;
    layer3_outputs(8379) <= a and not b;
    layer3_outputs(8380) <= b and not a;
    layer3_outputs(8381) <= b;
    layer3_outputs(8382) <= b;
    layer3_outputs(8383) <= a or b;
    layer3_outputs(8384) <= not (a or b);
    layer3_outputs(8385) <= not b;
    layer3_outputs(8386) <= '0';
    layer3_outputs(8387) <= a;
    layer3_outputs(8388) <= b;
    layer3_outputs(8389) <= '0';
    layer3_outputs(8390) <= not a;
    layer3_outputs(8391) <= b and not a;
    layer3_outputs(8392) <= not a or b;
    layer3_outputs(8393) <= not b or a;
    layer3_outputs(8394) <= not (a and b);
    layer3_outputs(8395) <= '1';
    layer3_outputs(8396) <= not a or b;
    layer3_outputs(8397) <= b;
    layer3_outputs(8398) <= a and not b;
    layer3_outputs(8399) <= a and not b;
    layer3_outputs(8400) <= a xor b;
    layer3_outputs(8401) <= b;
    layer3_outputs(8402) <= a and not b;
    layer3_outputs(8403) <= a;
    layer3_outputs(8404) <= a and b;
    layer3_outputs(8405) <= a;
    layer3_outputs(8406) <= a or b;
    layer3_outputs(8407) <= not a;
    layer3_outputs(8408) <= a and b;
    layer3_outputs(8409) <= not a or b;
    layer3_outputs(8410) <= not b or a;
    layer3_outputs(8411) <= not a or b;
    layer3_outputs(8412) <= a;
    layer3_outputs(8413) <= not a;
    layer3_outputs(8414) <= a xor b;
    layer3_outputs(8415) <= not b;
    layer3_outputs(8416) <= a or b;
    layer3_outputs(8417) <= '1';
    layer3_outputs(8418) <= not (a or b);
    layer3_outputs(8419) <= a or b;
    layer3_outputs(8420) <= a or b;
    layer3_outputs(8421) <= not (a and b);
    layer3_outputs(8422) <= b and not a;
    layer3_outputs(8423) <= not a or b;
    layer3_outputs(8424) <= '1';
    layer3_outputs(8425) <= not a;
    layer3_outputs(8426) <= not b or a;
    layer3_outputs(8427) <= not b or a;
    layer3_outputs(8428) <= not b or a;
    layer3_outputs(8429) <= not b;
    layer3_outputs(8430) <= not (a and b);
    layer3_outputs(8431) <= a and not b;
    layer3_outputs(8432) <= not (a and b);
    layer3_outputs(8433) <= not b;
    layer3_outputs(8434) <= b;
    layer3_outputs(8435) <= not (a and b);
    layer3_outputs(8436) <= not b;
    layer3_outputs(8437) <= a;
    layer3_outputs(8438) <= not b or a;
    layer3_outputs(8439) <= b;
    layer3_outputs(8440) <= a and b;
    layer3_outputs(8441) <= a;
    layer3_outputs(8442) <= a and b;
    layer3_outputs(8443) <= a and b;
    layer3_outputs(8444) <= a and b;
    layer3_outputs(8445) <= not a or b;
    layer3_outputs(8446) <= b;
    layer3_outputs(8447) <= '0';
    layer3_outputs(8448) <= not b or a;
    layer3_outputs(8449) <= b;
    layer3_outputs(8450) <= a;
    layer3_outputs(8451) <= b;
    layer3_outputs(8452) <= not (a and b);
    layer3_outputs(8453) <= not a or b;
    layer3_outputs(8454) <= a and not b;
    layer3_outputs(8455) <= b;
    layer3_outputs(8456) <= not b or a;
    layer3_outputs(8457) <= not a;
    layer3_outputs(8458) <= not b or a;
    layer3_outputs(8459) <= not a or b;
    layer3_outputs(8460) <= a and not b;
    layer3_outputs(8461) <= not a;
    layer3_outputs(8462) <= not (a and b);
    layer3_outputs(8463) <= b;
    layer3_outputs(8464) <= not a;
    layer3_outputs(8465) <= not b or a;
    layer3_outputs(8466) <= a;
    layer3_outputs(8467) <= '0';
    layer3_outputs(8468) <= b;
    layer3_outputs(8469) <= not (a or b);
    layer3_outputs(8470) <= a or b;
    layer3_outputs(8471) <= b;
    layer3_outputs(8472) <= a;
    layer3_outputs(8473) <= not a;
    layer3_outputs(8474) <= b and not a;
    layer3_outputs(8475) <= a or b;
    layer3_outputs(8476) <= '1';
    layer3_outputs(8477) <= a or b;
    layer3_outputs(8478) <= not a or b;
    layer3_outputs(8479) <= not b;
    layer3_outputs(8480) <= a;
    layer3_outputs(8481) <= '0';
    layer3_outputs(8482) <= a;
    layer3_outputs(8483) <= b and not a;
    layer3_outputs(8484) <= not b;
    layer3_outputs(8485) <= a;
    layer3_outputs(8486) <= a;
    layer3_outputs(8487) <= not (a and b);
    layer3_outputs(8488) <= not b or a;
    layer3_outputs(8489) <= b and not a;
    layer3_outputs(8490) <= '0';
    layer3_outputs(8491) <= a or b;
    layer3_outputs(8492) <= not (a and b);
    layer3_outputs(8493) <= a or b;
    layer3_outputs(8494) <= a;
    layer3_outputs(8495) <= not a or b;
    layer3_outputs(8496) <= a;
    layer3_outputs(8497) <= b;
    layer3_outputs(8498) <= a xor b;
    layer3_outputs(8499) <= b and not a;
    layer3_outputs(8500) <= not a or b;
    layer3_outputs(8501) <= b;
    layer3_outputs(8502) <= a;
    layer3_outputs(8503) <= not b;
    layer3_outputs(8504) <= '1';
    layer3_outputs(8505) <= a and not b;
    layer3_outputs(8506) <= '1';
    layer3_outputs(8507) <= a;
    layer3_outputs(8508) <= not a;
    layer3_outputs(8509) <= not a;
    layer3_outputs(8510) <= a;
    layer3_outputs(8511) <= not (a and b);
    layer3_outputs(8512) <= not (a xor b);
    layer3_outputs(8513) <= a and b;
    layer3_outputs(8514) <= not a or b;
    layer3_outputs(8515) <= '0';
    layer3_outputs(8516) <= a or b;
    layer3_outputs(8517) <= not a or b;
    layer3_outputs(8518) <= not b;
    layer3_outputs(8519) <= a or b;
    layer3_outputs(8520) <= not (a xor b);
    layer3_outputs(8521) <= not (a or b);
    layer3_outputs(8522) <= not b;
    layer3_outputs(8523) <= not a;
    layer3_outputs(8524) <= a and b;
    layer3_outputs(8525) <= not (a xor b);
    layer3_outputs(8526) <= not (a xor b);
    layer3_outputs(8527) <= not b or a;
    layer3_outputs(8528) <= not (a and b);
    layer3_outputs(8529) <= b and not a;
    layer3_outputs(8530) <= not a or b;
    layer3_outputs(8531) <= not b;
    layer3_outputs(8532) <= not a;
    layer3_outputs(8533) <= a and b;
    layer3_outputs(8534) <= not b or a;
    layer3_outputs(8535) <= '0';
    layer3_outputs(8536) <= not a;
    layer3_outputs(8537) <= b;
    layer3_outputs(8538) <= b;
    layer3_outputs(8539) <= not b;
    layer3_outputs(8540) <= a;
    layer3_outputs(8541) <= a;
    layer3_outputs(8542) <= not b;
    layer3_outputs(8543) <= a and not b;
    layer3_outputs(8544) <= not b;
    layer3_outputs(8545) <= not a or b;
    layer3_outputs(8546) <= a;
    layer3_outputs(8547) <= b and not a;
    layer3_outputs(8548) <= not a;
    layer3_outputs(8549) <= not b or a;
    layer3_outputs(8550) <= a and not b;
    layer3_outputs(8551) <= not b;
    layer3_outputs(8552) <= not b or a;
    layer3_outputs(8553) <= a and not b;
    layer3_outputs(8554) <= not b;
    layer3_outputs(8555) <= a;
    layer3_outputs(8556) <= not b;
    layer3_outputs(8557) <= a or b;
    layer3_outputs(8558) <= not b;
    layer3_outputs(8559) <= not (a xor b);
    layer3_outputs(8560) <= a or b;
    layer3_outputs(8561) <= not a;
    layer3_outputs(8562) <= not b or a;
    layer3_outputs(8563) <= not b or a;
    layer3_outputs(8564) <= b and not a;
    layer3_outputs(8565) <= a or b;
    layer3_outputs(8566) <= not a;
    layer3_outputs(8567) <= not b or a;
    layer3_outputs(8568) <= '0';
    layer3_outputs(8569) <= a;
    layer3_outputs(8570) <= '1';
    layer3_outputs(8571) <= not b;
    layer3_outputs(8572) <= '0';
    layer3_outputs(8573) <= not a or b;
    layer3_outputs(8574) <= '1';
    layer3_outputs(8575) <= a;
    layer3_outputs(8576) <= '0';
    layer3_outputs(8577) <= a and b;
    layer3_outputs(8578) <= b;
    layer3_outputs(8579) <= not (a or b);
    layer3_outputs(8580) <= not b;
    layer3_outputs(8581) <= not b;
    layer3_outputs(8582) <= not (a and b);
    layer3_outputs(8583) <= b and not a;
    layer3_outputs(8584) <= a and not b;
    layer3_outputs(8585) <= '0';
    layer3_outputs(8586) <= not b;
    layer3_outputs(8587) <= not b;
    layer3_outputs(8588) <= not (a and b);
    layer3_outputs(8589) <= '1';
    layer3_outputs(8590) <= b;
    layer3_outputs(8591) <= b;
    layer3_outputs(8592) <= a and b;
    layer3_outputs(8593) <= b;
    layer3_outputs(8594) <= not (a and b);
    layer3_outputs(8595) <= not b or a;
    layer3_outputs(8596) <= a xor b;
    layer3_outputs(8597) <= a and not b;
    layer3_outputs(8598) <= a;
    layer3_outputs(8599) <= not b;
    layer3_outputs(8600) <= not a;
    layer3_outputs(8601) <= b;
    layer3_outputs(8602) <= not a;
    layer3_outputs(8603) <= a;
    layer3_outputs(8604) <= not (a xor b);
    layer3_outputs(8605) <= not a;
    layer3_outputs(8606) <= not b;
    layer3_outputs(8607) <= a and not b;
    layer3_outputs(8608) <= not a;
    layer3_outputs(8609) <= b;
    layer3_outputs(8610) <= a and b;
    layer3_outputs(8611) <= a and not b;
    layer3_outputs(8612) <= not b;
    layer3_outputs(8613) <= not a;
    layer3_outputs(8614) <= not a;
    layer3_outputs(8615) <= a;
    layer3_outputs(8616) <= b;
    layer3_outputs(8617) <= a;
    layer3_outputs(8618) <= b;
    layer3_outputs(8619) <= not b;
    layer3_outputs(8620) <= not b or a;
    layer3_outputs(8621) <= a and b;
    layer3_outputs(8622) <= a and not b;
    layer3_outputs(8623) <= b;
    layer3_outputs(8624) <= not a or b;
    layer3_outputs(8625) <= not b;
    layer3_outputs(8626) <= a or b;
    layer3_outputs(8627) <= a xor b;
    layer3_outputs(8628) <= '0';
    layer3_outputs(8629) <= '1';
    layer3_outputs(8630) <= a;
    layer3_outputs(8631) <= '0';
    layer3_outputs(8632) <= not (a or b);
    layer3_outputs(8633) <= not b;
    layer3_outputs(8634) <= '0';
    layer3_outputs(8635) <= not a;
    layer3_outputs(8636) <= b;
    layer3_outputs(8637) <= a and not b;
    layer3_outputs(8638) <= a or b;
    layer3_outputs(8639) <= '0';
    layer3_outputs(8640) <= not a;
    layer3_outputs(8641) <= b and not a;
    layer3_outputs(8642) <= '0';
    layer3_outputs(8643) <= a and b;
    layer3_outputs(8644) <= not a;
    layer3_outputs(8645) <= '1';
    layer3_outputs(8646) <= not (a and b);
    layer3_outputs(8647) <= not (a and b);
    layer3_outputs(8648) <= a and not b;
    layer3_outputs(8649) <= not a;
    layer3_outputs(8650) <= '0';
    layer3_outputs(8651) <= '1';
    layer3_outputs(8652) <= a;
    layer3_outputs(8653) <= b;
    layer3_outputs(8654) <= not b or a;
    layer3_outputs(8655) <= not b or a;
    layer3_outputs(8656) <= a and not b;
    layer3_outputs(8657) <= b;
    layer3_outputs(8658) <= not a or b;
    layer3_outputs(8659) <= not (a or b);
    layer3_outputs(8660) <= not b or a;
    layer3_outputs(8661) <= not (a and b);
    layer3_outputs(8662) <= b;
    layer3_outputs(8663) <= b;
    layer3_outputs(8664) <= not a or b;
    layer3_outputs(8665) <= not b or a;
    layer3_outputs(8666) <= not a;
    layer3_outputs(8667) <= a;
    layer3_outputs(8668) <= not b;
    layer3_outputs(8669) <= b and not a;
    layer3_outputs(8670) <= b and not a;
    layer3_outputs(8671) <= a;
    layer3_outputs(8672) <= not b;
    layer3_outputs(8673) <= a and b;
    layer3_outputs(8674) <= not (a or b);
    layer3_outputs(8675) <= a and not b;
    layer3_outputs(8676) <= '0';
    layer3_outputs(8677) <= not b;
    layer3_outputs(8678) <= not a or b;
    layer3_outputs(8679) <= a and not b;
    layer3_outputs(8680) <= not (a or b);
    layer3_outputs(8681) <= '0';
    layer3_outputs(8682) <= not a;
    layer3_outputs(8683) <= '0';
    layer3_outputs(8684) <= not (a or b);
    layer3_outputs(8685) <= b;
    layer3_outputs(8686) <= '1';
    layer3_outputs(8687) <= not a or b;
    layer3_outputs(8688) <= '0';
    layer3_outputs(8689) <= not a or b;
    layer3_outputs(8690) <= not b or a;
    layer3_outputs(8691) <= a;
    layer3_outputs(8692) <= b;
    layer3_outputs(8693) <= not (a and b);
    layer3_outputs(8694) <= not (a and b);
    layer3_outputs(8695) <= b and not a;
    layer3_outputs(8696) <= '1';
    layer3_outputs(8697) <= not b;
    layer3_outputs(8698) <= not a or b;
    layer3_outputs(8699) <= b;
    layer3_outputs(8700) <= a or b;
    layer3_outputs(8701) <= b;
    layer3_outputs(8702) <= a or b;
    layer3_outputs(8703) <= not b;
    layer3_outputs(8704) <= not b;
    layer3_outputs(8705) <= a and not b;
    layer3_outputs(8706) <= not b;
    layer3_outputs(8707) <= a;
    layer3_outputs(8708) <= not (a or b);
    layer3_outputs(8709) <= not (a xor b);
    layer3_outputs(8710) <= a and b;
    layer3_outputs(8711) <= not (a xor b);
    layer3_outputs(8712) <= b;
    layer3_outputs(8713) <= b and not a;
    layer3_outputs(8714) <= not b or a;
    layer3_outputs(8715) <= b;
    layer3_outputs(8716) <= b;
    layer3_outputs(8717) <= '1';
    layer3_outputs(8718) <= b and not a;
    layer3_outputs(8719) <= not b or a;
    layer3_outputs(8720) <= a and not b;
    layer3_outputs(8721) <= b;
    layer3_outputs(8722) <= not b;
    layer3_outputs(8723) <= not a;
    layer3_outputs(8724) <= b;
    layer3_outputs(8725) <= a and b;
    layer3_outputs(8726) <= not (a and b);
    layer3_outputs(8727) <= a and b;
    layer3_outputs(8728) <= a and b;
    layer3_outputs(8729) <= a and b;
    layer3_outputs(8730) <= b and not a;
    layer3_outputs(8731) <= not (a or b);
    layer3_outputs(8732) <= not b;
    layer3_outputs(8733) <= a;
    layer3_outputs(8734) <= not a;
    layer3_outputs(8735) <= b;
    layer3_outputs(8736) <= b;
    layer3_outputs(8737) <= a or b;
    layer3_outputs(8738) <= b;
    layer3_outputs(8739) <= not a or b;
    layer3_outputs(8740) <= b and not a;
    layer3_outputs(8741) <= a;
    layer3_outputs(8742) <= a and b;
    layer3_outputs(8743) <= not b or a;
    layer3_outputs(8744) <= not (a xor b);
    layer3_outputs(8745) <= b and not a;
    layer3_outputs(8746) <= a;
    layer3_outputs(8747) <= a and not b;
    layer3_outputs(8748) <= not b or a;
    layer3_outputs(8749) <= not a;
    layer3_outputs(8750) <= not (a and b);
    layer3_outputs(8751) <= a or b;
    layer3_outputs(8752) <= a and not b;
    layer3_outputs(8753) <= not a;
    layer3_outputs(8754) <= a xor b;
    layer3_outputs(8755) <= not b;
    layer3_outputs(8756) <= a;
    layer3_outputs(8757) <= not a;
    layer3_outputs(8758) <= not a;
    layer3_outputs(8759) <= a;
    layer3_outputs(8760) <= '1';
    layer3_outputs(8761) <= not b;
    layer3_outputs(8762) <= a or b;
    layer3_outputs(8763) <= a and b;
    layer3_outputs(8764) <= a and b;
    layer3_outputs(8765) <= a;
    layer3_outputs(8766) <= '0';
    layer3_outputs(8767) <= a;
    layer3_outputs(8768) <= not (a and b);
    layer3_outputs(8769) <= not b;
    layer3_outputs(8770) <= not (a and b);
    layer3_outputs(8771) <= a;
    layer3_outputs(8772) <= '0';
    layer3_outputs(8773) <= '0';
    layer3_outputs(8774) <= not a;
    layer3_outputs(8775) <= not b;
    layer3_outputs(8776) <= not a;
    layer3_outputs(8777) <= b;
    layer3_outputs(8778) <= a and b;
    layer3_outputs(8779) <= not b or a;
    layer3_outputs(8780) <= not b or a;
    layer3_outputs(8781) <= not a;
    layer3_outputs(8782) <= a and not b;
    layer3_outputs(8783) <= a or b;
    layer3_outputs(8784) <= a and b;
    layer3_outputs(8785) <= a;
    layer3_outputs(8786) <= b and not a;
    layer3_outputs(8787) <= a or b;
    layer3_outputs(8788) <= a and b;
    layer3_outputs(8789) <= a;
    layer3_outputs(8790) <= a;
    layer3_outputs(8791) <= '0';
    layer3_outputs(8792) <= not b;
    layer3_outputs(8793) <= not b;
    layer3_outputs(8794) <= a or b;
    layer3_outputs(8795) <= not (a or b);
    layer3_outputs(8796) <= b;
    layer3_outputs(8797) <= a and not b;
    layer3_outputs(8798) <= b;
    layer3_outputs(8799) <= a or b;
    layer3_outputs(8800) <= a and not b;
    layer3_outputs(8801) <= b and not a;
    layer3_outputs(8802) <= not b or a;
    layer3_outputs(8803) <= b and not a;
    layer3_outputs(8804) <= not b;
    layer3_outputs(8805) <= not b;
    layer3_outputs(8806) <= a xor b;
    layer3_outputs(8807) <= not b;
    layer3_outputs(8808) <= a;
    layer3_outputs(8809) <= not b or a;
    layer3_outputs(8810) <= not a or b;
    layer3_outputs(8811) <= b;
    layer3_outputs(8812) <= b and not a;
    layer3_outputs(8813) <= not a;
    layer3_outputs(8814) <= not b;
    layer3_outputs(8815) <= a;
    layer3_outputs(8816) <= not (a and b);
    layer3_outputs(8817) <= not a;
    layer3_outputs(8818) <= a and not b;
    layer3_outputs(8819) <= '1';
    layer3_outputs(8820) <= not (a and b);
    layer3_outputs(8821) <= b;
    layer3_outputs(8822) <= b;
    layer3_outputs(8823) <= a;
    layer3_outputs(8824) <= not b;
    layer3_outputs(8825) <= b and not a;
    layer3_outputs(8826) <= not b or a;
    layer3_outputs(8827) <= b;
    layer3_outputs(8828) <= a;
    layer3_outputs(8829) <= not a;
    layer3_outputs(8830) <= not (a xor b);
    layer3_outputs(8831) <= a;
    layer3_outputs(8832) <= a xor b;
    layer3_outputs(8833) <= b;
    layer3_outputs(8834) <= not b or a;
    layer3_outputs(8835) <= a;
    layer3_outputs(8836) <= not b;
    layer3_outputs(8837) <= not (a or b);
    layer3_outputs(8838) <= a or b;
    layer3_outputs(8839) <= not (a and b);
    layer3_outputs(8840) <= a and not b;
    layer3_outputs(8841) <= a and b;
    layer3_outputs(8842) <= not (a and b);
    layer3_outputs(8843) <= not (a and b);
    layer3_outputs(8844) <= '0';
    layer3_outputs(8845) <= not b;
    layer3_outputs(8846) <= not (a or b);
    layer3_outputs(8847) <= not a;
    layer3_outputs(8848) <= not a;
    layer3_outputs(8849) <= not (a and b);
    layer3_outputs(8850) <= not a;
    layer3_outputs(8851) <= '1';
    layer3_outputs(8852) <= not b or a;
    layer3_outputs(8853) <= b and not a;
    layer3_outputs(8854) <= a and not b;
    layer3_outputs(8855) <= a;
    layer3_outputs(8856) <= a and not b;
    layer3_outputs(8857) <= not (a and b);
    layer3_outputs(8858) <= not (a and b);
    layer3_outputs(8859) <= a;
    layer3_outputs(8860) <= '0';
    layer3_outputs(8861) <= not a or b;
    layer3_outputs(8862) <= not a;
    layer3_outputs(8863) <= a;
    layer3_outputs(8864) <= a or b;
    layer3_outputs(8865) <= not (a and b);
    layer3_outputs(8866) <= b and not a;
    layer3_outputs(8867) <= a;
    layer3_outputs(8868) <= not b;
    layer3_outputs(8869) <= a or b;
    layer3_outputs(8870) <= not b;
    layer3_outputs(8871) <= not b;
    layer3_outputs(8872) <= a;
    layer3_outputs(8873) <= b;
    layer3_outputs(8874) <= not b;
    layer3_outputs(8875) <= not (a or b);
    layer3_outputs(8876) <= not b or a;
    layer3_outputs(8877) <= not (a xor b);
    layer3_outputs(8878) <= a or b;
    layer3_outputs(8879) <= not (a and b);
    layer3_outputs(8880) <= not (a or b);
    layer3_outputs(8881) <= a and b;
    layer3_outputs(8882) <= not a;
    layer3_outputs(8883) <= a;
    layer3_outputs(8884) <= not b;
    layer3_outputs(8885) <= b;
    layer3_outputs(8886) <= b and not a;
    layer3_outputs(8887) <= a and not b;
    layer3_outputs(8888) <= b;
    layer3_outputs(8889) <= a and b;
    layer3_outputs(8890) <= not b;
    layer3_outputs(8891) <= a and b;
    layer3_outputs(8892) <= a or b;
    layer3_outputs(8893) <= not b;
    layer3_outputs(8894) <= not b;
    layer3_outputs(8895) <= b and not a;
    layer3_outputs(8896) <= a;
    layer3_outputs(8897) <= a;
    layer3_outputs(8898) <= a;
    layer3_outputs(8899) <= not (a xor b);
    layer3_outputs(8900) <= a and not b;
    layer3_outputs(8901) <= a and not b;
    layer3_outputs(8902) <= a and b;
    layer3_outputs(8903) <= b;
    layer3_outputs(8904) <= not b or a;
    layer3_outputs(8905) <= not a or b;
    layer3_outputs(8906) <= not a or b;
    layer3_outputs(8907) <= a xor b;
    layer3_outputs(8908) <= '1';
    layer3_outputs(8909) <= not b or a;
    layer3_outputs(8910) <= not b;
    layer3_outputs(8911) <= not b or a;
    layer3_outputs(8912) <= not a or b;
    layer3_outputs(8913) <= not a;
    layer3_outputs(8914) <= a and b;
    layer3_outputs(8915) <= not b or a;
    layer3_outputs(8916) <= a and not b;
    layer3_outputs(8917) <= not a;
    layer3_outputs(8918) <= not (a xor b);
    layer3_outputs(8919) <= a and not b;
    layer3_outputs(8920) <= not b;
    layer3_outputs(8921) <= b and not a;
    layer3_outputs(8922) <= '0';
    layer3_outputs(8923) <= a and b;
    layer3_outputs(8924) <= b and not a;
    layer3_outputs(8925) <= a and not b;
    layer3_outputs(8926) <= b;
    layer3_outputs(8927) <= a and b;
    layer3_outputs(8928) <= a;
    layer3_outputs(8929) <= a or b;
    layer3_outputs(8930) <= not a or b;
    layer3_outputs(8931) <= not (a or b);
    layer3_outputs(8932) <= b;
    layer3_outputs(8933) <= a and b;
    layer3_outputs(8934) <= '1';
    layer3_outputs(8935) <= not (a or b);
    layer3_outputs(8936) <= not a or b;
    layer3_outputs(8937) <= a and not b;
    layer3_outputs(8938) <= not b or a;
    layer3_outputs(8939) <= b and not a;
    layer3_outputs(8940) <= a;
    layer3_outputs(8941) <= a and not b;
    layer3_outputs(8942) <= not a;
    layer3_outputs(8943) <= not (a or b);
    layer3_outputs(8944) <= not b or a;
    layer3_outputs(8945) <= not (a or b);
    layer3_outputs(8946) <= a or b;
    layer3_outputs(8947) <= '1';
    layer3_outputs(8948) <= b and not a;
    layer3_outputs(8949) <= a and not b;
    layer3_outputs(8950) <= not a or b;
    layer3_outputs(8951) <= not b;
    layer3_outputs(8952) <= '1';
    layer3_outputs(8953) <= not a or b;
    layer3_outputs(8954) <= not (a xor b);
    layer3_outputs(8955) <= not (a or b);
    layer3_outputs(8956) <= a and not b;
    layer3_outputs(8957) <= not a;
    layer3_outputs(8958) <= b;
    layer3_outputs(8959) <= not b or a;
    layer3_outputs(8960) <= not b;
    layer3_outputs(8961) <= b;
    layer3_outputs(8962) <= not (a xor b);
    layer3_outputs(8963) <= b and not a;
    layer3_outputs(8964) <= b and not a;
    layer3_outputs(8965) <= a;
    layer3_outputs(8966) <= not (a and b);
    layer3_outputs(8967) <= not b or a;
    layer3_outputs(8968) <= a and b;
    layer3_outputs(8969) <= not b or a;
    layer3_outputs(8970) <= not a;
    layer3_outputs(8971) <= b;
    layer3_outputs(8972) <= a;
    layer3_outputs(8973) <= a;
    layer3_outputs(8974) <= '0';
    layer3_outputs(8975) <= b and not a;
    layer3_outputs(8976) <= not b;
    layer3_outputs(8977) <= a or b;
    layer3_outputs(8978) <= not (a or b);
    layer3_outputs(8979) <= a;
    layer3_outputs(8980) <= not (a xor b);
    layer3_outputs(8981) <= a;
    layer3_outputs(8982) <= '0';
    layer3_outputs(8983) <= a or b;
    layer3_outputs(8984) <= a and b;
    layer3_outputs(8985) <= not b;
    layer3_outputs(8986) <= not (a or b);
    layer3_outputs(8987) <= '0';
    layer3_outputs(8988) <= not b;
    layer3_outputs(8989) <= a;
    layer3_outputs(8990) <= a xor b;
    layer3_outputs(8991) <= a or b;
    layer3_outputs(8992) <= a or b;
    layer3_outputs(8993) <= b;
    layer3_outputs(8994) <= a;
    layer3_outputs(8995) <= not a or b;
    layer3_outputs(8996) <= not a or b;
    layer3_outputs(8997) <= not (a or b);
    layer3_outputs(8998) <= a xor b;
    layer3_outputs(8999) <= not b;
    layer3_outputs(9000) <= a or b;
    layer3_outputs(9001) <= not b;
    layer3_outputs(9002) <= not a or b;
    layer3_outputs(9003) <= a and not b;
    layer3_outputs(9004) <= '1';
    layer3_outputs(9005) <= a;
    layer3_outputs(9006) <= '0';
    layer3_outputs(9007) <= '1';
    layer3_outputs(9008) <= a;
    layer3_outputs(9009) <= a;
    layer3_outputs(9010) <= b;
    layer3_outputs(9011) <= '0';
    layer3_outputs(9012) <= not b;
    layer3_outputs(9013) <= a and b;
    layer3_outputs(9014) <= a xor b;
    layer3_outputs(9015) <= not b;
    layer3_outputs(9016) <= a;
    layer3_outputs(9017) <= not b or a;
    layer3_outputs(9018) <= not (a xor b);
    layer3_outputs(9019) <= b and not a;
    layer3_outputs(9020) <= a;
    layer3_outputs(9021) <= not b or a;
    layer3_outputs(9022) <= a and not b;
    layer3_outputs(9023) <= not (a or b);
    layer3_outputs(9024) <= not (a or b);
    layer3_outputs(9025) <= b and not a;
    layer3_outputs(9026) <= not (a xor b);
    layer3_outputs(9027) <= not b;
    layer3_outputs(9028) <= not b or a;
    layer3_outputs(9029) <= not (a and b);
    layer3_outputs(9030) <= not a or b;
    layer3_outputs(9031) <= a;
    layer3_outputs(9032) <= b;
    layer3_outputs(9033) <= not (a and b);
    layer3_outputs(9034) <= b;
    layer3_outputs(9035) <= '1';
    layer3_outputs(9036) <= a and b;
    layer3_outputs(9037) <= a and b;
    layer3_outputs(9038) <= b and not a;
    layer3_outputs(9039) <= a and b;
    layer3_outputs(9040) <= b;
    layer3_outputs(9041) <= not a;
    layer3_outputs(9042) <= not a or b;
    layer3_outputs(9043) <= not (a or b);
    layer3_outputs(9044) <= a and b;
    layer3_outputs(9045) <= not b or a;
    layer3_outputs(9046) <= '1';
    layer3_outputs(9047) <= a and not b;
    layer3_outputs(9048) <= not (a and b);
    layer3_outputs(9049) <= a and b;
    layer3_outputs(9050) <= a;
    layer3_outputs(9051) <= not (a and b);
    layer3_outputs(9052) <= a or b;
    layer3_outputs(9053) <= a or b;
    layer3_outputs(9054) <= a;
    layer3_outputs(9055) <= not a;
    layer3_outputs(9056) <= not (a xor b);
    layer3_outputs(9057) <= b and not a;
    layer3_outputs(9058) <= not b;
    layer3_outputs(9059) <= b;
    layer3_outputs(9060) <= not a or b;
    layer3_outputs(9061) <= not (a or b);
    layer3_outputs(9062) <= not (a or b);
    layer3_outputs(9063) <= not (a xor b);
    layer3_outputs(9064) <= not b or a;
    layer3_outputs(9065) <= a;
    layer3_outputs(9066) <= not a or b;
    layer3_outputs(9067) <= not a;
    layer3_outputs(9068) <= not (a xor b);
    layer3_outputs(9069) <= a or b;
    layer3_outputs(9070) <= not b;
    layer3_outputs(9071) <= a and b;
    layer3_outputs(9072) <= not (a and b);
    layer3_outputs(9073) <= not b;
    layer3_outputs(9074) <= not a or b;
    layer3_outputs(9075) <= b;
    layer3_outputs(9076) <= a and not b;
    layer3_outputs(9077) <= not b or a;
    layer3_outputs(9078) <= a;
    layer3_outputs(9079) <= b and not a;
    layer3_outputs(9080) <= not a or b;
    layer3_outputs(9081) <= not (a xor b);
    layer3_outputs(9082) <= a;
    layer3_outputs(9083) <= not a;
    layer3_outputs(9084) <= not (a and b);
    layer3_outputs(9085) <= not b or a;
    layer3_outputs(9086) <= a or b;
    layer3_outputs(9087) <= not a or b;
    layer3_outputs(9088) <= not a;
    layer3_outputs(9089) <= b;
    layer3_outputs(9090) <= a;
    layer3_outputs(9091) <= not a;
    layer3_outputs(9092) <= b;
    layer3_outputs(9093) <= a and not b;
    layer3_outputs(9094) <= a;
    layer3_outputs(9095) <= a and not b;
    layer3_outputs(9096) <= '0';
    layer3_outputs(9097) <= '0';
    layer3_outputs(9098) <= not b;
    layer3_outputs(9099) <= b and not a;
    layer3_outputs(9100) <= not a;
    layer3_outputs(9101) <= '0';
    layer3_outputs(9102) <= not (a xor b);
    layer3_outputs(9103) <= not a;
    layer3_outputs(9104) <= b;
    layer3_outputs(9105) <= not b;
    layer3_outputs(9106) <= not b;
    layer3_outputs(9107) <= not b;
    layer3_outputs(9108) <= not b or a;
    layer3_outputs(9109) <= not a or b;
    layer3_outputs(9110) <= not a;
    layer3_outputs(9111) <= b;
    layer3_outputs(9112) <= '1';
    layer3_outputs(9113) <= not a;
    layer3_outputs(9114) <= a;
    layer3_outputs(9115) <= a or b;
    layer3_outputs(9116) <= a and not b;
    layer3_outputs(9117) <= '1';
    layer3_outputs(9118) <= not a;
    layer3_outputs(9119) <= a and b;
    layer3_outputs(9120) <= a and b;
    layer3_outputs(9121) <= a;
    layer3_outputs(9122) <= a;
    layer3_outputs(9123) <= not b;
    layer3_outputs(9124) <= not a or b;
    layer3_outputs(9125) <= b;
    layer3_outputs(9126) <= not b or a;
    layer3_outputs(9127) <= a;
    layer3_outputs(9128) <= a xor b;
    layer3_outputs(9129) <= a and b;
    layer3_outputs(9130) <= not a or b;
    layer3_outputs(9131) <= b;
    layer3_outputs(9132) <= a xor b;
    layer3_outputs(9133) <= not (a or b);
    layer3_outputs(9134) <= not (a xor b);
    layer3_outputs(9135) <= a and not b;
    layer3_outputs(9136) <= not a;
    layer3_outputs(9137) <= a and not b;
    layer3_outputs(9138) <= not b or a;
    layer3_outputs(9139) <= not b;
    layer3_outputs(9140) <= not (a or b);
    layer3_outputs(9141) <= a and b;
    layer3_outputs(9142) <= not (a and b);
    layer3_outputs(9143) <= b and not a;
    layer3_outputs(9144) <= a;
    layer3_outputs(9145) <= a or b;
    layer3_outputs(9146) <= a and not b;
    layer3_outputs(9147) <= not b;
    layer3_outputs(9148) <= a xor b;
    layer3_outputs(9149) <= not (a or b);
    layer3_outputs(9150) <= not (a and b);
    layer3_outputs(9151) <= not b;
    layer3_outputs(9152) <= a xor b;
    layer3_outputs(9153) <= a and not b;
    layer3_outputs(9154) <= not (a and b);
    layer3_outputs(9155) <= not b;
    layer3_outputs(9156) <= not (a and b);
    layer3_outputs(9157) <= a and not b;
    layer3_outputs(9158) <= a or b;
    layer3_outputs(9159) <= a and not b;
    layer3_outputs(9160) <= a or b;
    layer3_outputs(9161) <= a;
    layer3_outputs(9162) <= b and not a;
    layer3_outputs(9163) <= a and not b;
    layer3_outputs(9164) <= not a;
    layer3_outputs(9165) <= a;
    layer3_outputs(9166) <= not a or b;
    layer3_outputs(9167) <= a and not b;
    layer3_outputs(9168) <= a and not b;
    layer3_outputs(9169) <= not a or b;
    layer3_outputs(9170) <= not a;
    layer3_outputs(9171) <= a;
    layer3_outputs(9172) <= not a;
    layer3_outputs(9173) <= not (a xor b);
    layer3_outputs(9174) <= not a;
    layer3_outputs(9175) <= not (a or b);
    layer3_outputs(9176) <= not a or b;
    layer3_outputs(9177) <= a and b;
    layer3_outputs(9178) <= not a;
    layer3_outputs(9179) <= a and b;
    layer3_outputs(9180) <= b;
    layer3_outputs(9181) <= not a;
    layer3_outputs(9182) <= a and b;
    layer3_outputs(9183) <= b and not a;
    layer3_outputs(9184) <= b and not a;
    layer3_outputs(9185) <= not (a or b);
    layer3_outputs(9186) <= not b or a;
    layer3_outputs(9187) <= not b or a;
    layer3_outputs(9188) <= not (a and b);
    layer3_outputs(9189) <= a;
    layer3_outputs(9190) <= '0';
    layer3_outputs(9191) <= b;
    layer3_outputs(9192) <= not a or b;
    layer3_outputs(9193) <= not a;
    layer3_outputs(9194) <= not b or a;
    layer3_outputs(9195) <= not b;
    layer3_outputs(9196) <= not b or a;
    layer3_outputs(9197) <= b;
    layer3_outputs(9198) <= a;
    layer3_outputs(9199) <= b;
    layer3_outputs(9200) <= a xor b;
    layer3_outputs(9201) <= not b;
    layer3_outputs(9202) <= a and b;
    layer3_outputs(9203) <= not (a or b);
    layer3_outputs(9204) <= not a;
    layer3_outputs(9205) <= a and b;
    layer3_outputs(9206) <= not a;
    layer3_outputs(9207) <= b;
    layer3_outputs(9208) <= b;
    layer3_outputs(9209) <= not a;
    layer3_outputs(9210) <= not b or a;
    layer3_outputs(9211) <= not a;
    layer3_outputs(9212) <= '0';
    layer3_outputs(9213) <= not b or a;
    layer3_outputs(9214) <= b and not a;
    layer3_outputs(9215) <= not b;
    layer3_outputs(9216) <= a or b;
    layer3_outputs(9217) <= not a;
    layer3_outputs(9218) <= a and not b;
    layer3_outputs(9219) <= a and b;
    layer3_outputs(9220) <= not a or b;
    layer3_outputs(9221) <= '1';
    layer3_outputs(9222) <= '0';
    layer3_outputs(9223) <= not b;
    layer3_outputs(9224) <= '1';
    layer3_outputs(9225) <= '1';
    layer3_outputs(9226) <= not a;
    layer3_outputs(9227) <= not b or a;
    layer3_outputs(9228) <= a and b;
    layer3_outputs(9229) <= b;
    layer3_outputs(9230) <= a or b;
    layer3_outputs(9231) <= b;
    layer3_outputs(9232) <= a;
    layer3_outputs(9233) <= not b;
    layer3_outputs(9234) <= a or b;
    layer3_outputs(9235) <= not (a and b);
    layer3_outputs(9236) <= a;
    layer3_outputs(9237) <= not (a and b);
    layer3_outputs(9238) <= not (a and b);
    layer3_outputs(9239) <= a;
    layer3_outputs(9240) <= not (a and b);
    layer3_outputs(9241) <= b and not a;
    layer3_outputs(9242) <= b;
    layer3_outputs(9243) <= a;
    layer3_outputs(9244) <= a or b;
    layer3_outputs(9245) <= not b or a;
    layer3_outputs(9246) <= a;
    layer3_outputs(9247) <= not a;
    layer3_outputs(9248) <= not (a and b);
    layer3_outputs(9249) <= b and not a;
    layer3_outputs(9250) <= not b;
    layer3_outputs(9251) <= not a;
    layer3_outputs(9252) <= not a or b;
    layer3_outputs(9253) <= b;
    layer3_outputs(9254) <= a or b;
    layer3_outputs(9255) <= a or b;
    layer3_outputs(9256) <= b and not a;
    layer3_outputs(9257) <= a or b;
    layer3_outputs(9258) <= a and b;
    layer3_outputs(9259) <= a and b;
    layer3_outputs(9260) <= a and b;
    layer3_outputs(9261) <= b;
    layer3_outputs(9262) <= not b;
    layer3_outputs(9263) <= a;
    layer3_outputs(9264) <= not a or b;
    layer3_outputs(9265) <= a xor b;
    layer3_outputs(9266) <= b;
    layer3_outputs(9267) <= not b;
    layer3_outputs(9268) <= a or b;
    layer3_outputs(9269) <= a;
    layer3_outputs(9270) <= a and not b;
    layer3_outputs(9271) <= a;
    layer3_outputs(9272) <= a or b;
    layer3_outputs(9273) <= a;
    layer3_outputs(9274) <= b;
    layer3_outputs(9275) <= not b;
    layer3_outputs(9276) <= not b or a;
    layer3_outputs(9277) <= '0';
    layer3_outputs(9278) <= not (a xor b);
    layer3_outputs(9279) <= a xor b;
    layer3_outputs(9280) <= not (a xor b);
    layer3_outputs(9281) <= b;
    layer3_outputs(9282) <= a;
    layer3_outputs(9283) <= b and not a;
    layer3_outputs(9284) <= a;
    layer3_outputs(9285) <= a xor b;
    layer3_outputs(9286) <= a or b;
    layer3_outputs(9287) <= b;
    layer3_outputs(9288) <= not (a or b);
    layer3_outputs(9289) <= not a or b;
    layer3_outputs(9290) <= a;
    layer3_outputs(9291) <= not b or a;
    layer3_outputs(9292) <= a and b;
    layer3_outputs(9293) <= a xor b;
    layer3_outputs(9294) <= not a or b;
    layer3_outputs(9295) <= a or b;
    layer3_outputs(9296) <= b and not a;
    layer3_outputs(9297) <= '0';
    layer3_outputs(9298) <= not b or a;
    layer3_outputs(9299) <= not a or b;
    layer3_outputs(9300) <= not (a and b);
    layer3_outputs(9301) <= b and not a;
    layer3_outputs(9302) <= '0';
    layer3_outputs(9303) <= a;
    layer3_outputs(9304) <= '0';
    layer3_outputs(9305) <= a;
    layer3_outputs(9306) <= not (a or b);
    layer3_outputs(9307) <= a;
    layer3_outputs(9308) <= a;
    layer3_outputs(9309) <= not (a or b);
    layer3_outputs(9310) <= a;
    layer3_outputs(9311) <= not b or a;
    layer3_outputs(9312) <= not b;
    layer3_outputs(9313) <= not (a or b);
    layer3_outputs(9314) <= not a;
    layer3_outputs(9315) <= not (a xor b);
    layer3_outputs(9316) <= not (a or b);
    layer3_outputs(9317) <= b and not a;
    layer3_outputs(9318) <= not b or a;
    layer3_outputs(9319) <= a xor b;
    layer3_outputs(9320) <= a xor b;
    layer3_outputs(9321) <= not (a and b);
    layer3_outputs(9322) <= b and not a;
    layer3_outputs(9323) <= not (a xor b);
    layer3_outputs(9324) <= a and not b;
    layer3_outputs(9325) <= not (a or b);
    layer3_outputs(9326) <= not b or a;
    layer3_outputs(9327) <= not a or b;
    layer3_outputs(9328) <= '0';
    layer3_outputs(9329) <= not b or a;
    layer3_outputs(9330) <= not b or a;
    layer3_outputs(9331) <= a and b;
    layer3_outputs(9332) <= '0';
    layer3_outputs(9333) <= a;
    layer3_outputs(9334) <= not (a or b);
    layer3_outputs(9335) <= '0';
    layer3_outputs(9336) <= a and not b;
    layer3_outputs(9337) <= a xor b;
    layer3_outputs(9338) <= a xor b;
    layer3_outputs(9339) <= not b or a;
    layer3_outputs(9340) <= not b or a;
    layer3_outputs(9341) <= '1';
    layer3_outputs(9342) <= a xor b;
    layer3_outputs(9343) <= a xor b;
    layer3_outputs(9344) <= a and not b;
    layer3_outputs(9345) <= not (a or b);
    layer3_outputs(9346) <= not b;
    layer3_outputs(9347) <= not b;
    layer3_outputs(9348) <= a or b;
    layer3_outputs(9349) <= not b;
    layer3_outputs(9350) <= b;
    layer3_outputs(9351) <= a;
    layer3_outputs(9352) <= not a;
    layer3_outputs(9353) <= '0';
    layer3_outputs(9354) <= a xor b;
    layer3_outputs(9355) <= '0';
    layer3_outputs(9356) <= not (a xor b);
    layer3_outputs(9357) <= a or b;
    layer3_outputs(9358) <= a;
    layer3_outputs(9359) <= not b;
    layer3_outputs(9360) <= not a;
    layer3_outputs(9361) <= a;
    layer3_outputs(9362) <= '1';
    layer3_outputs(9363) <= not a;
    layer3_outputs(9364) <= a or b;
    layer3_outputs(9365) <= a and not b;
    layer3_outputs(9366) <= '0';
    layer3_outputs(9367) <= b;
    layer3_outputs(9368) <= b and not a;
    layer3_outputs(9369) <= a and not b;
    layer3_outputs(9370) <= not b or a;
    layer3_outputs(9371) <= a;
    layer3_outputs(9372) <= not (a and b);
    layer3_outputs(9373) <= a or b;
    layer3_outputs(9374) <= b and not a;
    layer3_outputs(9375) <= not b;
    layer3_outputs(9376) <= not (a and b);
    layer3_outputs(9377) <= not a or b;
    layer3_outputs(9378) <= '0';
    layer3_outputs(9379) <= b;
    layer3_outputs(9380) <= not a or b;
    layer3_outputs(9381) <= '0';
    layer3_outputs(9382) <= not (a and b);
    layer3_outputs(9383) <= not (a or b);
    layer3_outputs(9384) <= a xor b;
    layer3_outputs(9385) <= b;
    layer3_outputs(9386) <= not b or a;
    layer3_outputs(9387) <= not b or a;
    layer3_outputs(9388) <= a or b;
    layer3_outputs(9389) <= b and not a;
    layer3_outputs(9390) <= b and not a;
    layer3_outputs(9391) <= not b;
    layer3_outputs(9392) <= not b;
    layer3_outputs(9393) <= a and b;
    layer3_outputs(9394) <= b;
    layer3_outputs(9395) <= not a;
    layer3_outputs(9396) <= a;
    layer3_outputs(9397) <= a and not b;
    layer3_outputs(9398) <= not (a and b);
    layer3_outputs(9399) <= '1';
    layer3_outputs(9400) <= not a;
    layer3_outputs(9401) <= not (a or b);
    layer3_outputs(9402) <= not a or b;
    layer3_outputs(9403) <= a;
    layer3_outputs(9404) <= not a;
    layer3_outputs(9405) <= a;
    layer3_outputs(9406) <= not (a xor b);
    layer3_outputs(9407) <= not b;
    layer3_outputs(9408) <= not a;
    layer3_outputs(9409) <= '1';
    layer3_outputs(9410) <= b;
    layer3_outputs(9411) <= not (a or b);
    layer3_outputs(9412) <= '1';
    layer3_outputs(9413) <= not (a and b);
    layer3_outputs(9414) <= b;
    layer3_outputs(9415) <= '0';
    layer3_outputs(9416) <= not a;
    layer3_outputs(9417) <= a xor b;
    layer3_outputs(9418) <= not (a and b);
    layer3_outputs(9419) <= not a or b;
    layer3_outputs(9420) <= not a;
    layer3_outputs(9421) <= not (a and b);
    layer3_outputs(9422) <= b;
    layer3_outputs(9423) <= a or b;
    layer3_outputs(9424) <= not b or a;
    layer3_outputs(9425) <= not b or a;
    layer3_outputs(9426) <= not b or a;
    layer3_outputs(9427) <= b and not a;
    layer3_outputs(9428) <= not (a and b);
    layer3_outputs(9429) <= a and not b;
    layer3_outputs(9430) <= b and not a;
    layer3_outputs(9431) <= not (a or b);
    layer3_outputs(9432) <= '0';
    layer3_outputs(9433) <= not b;
    layer3_outputs(9434) <= a or b;
    layer3_outputs(9435) <= not a;
    layer3_outputs(9436) <= b and not a;
    layer3_outputs(9437) <= not (a or b);
    layer3_outputs(9438) <= a;
    layer3_outputs(9439) <= a and b;
    layer3_outputs(9440) <= not (a or b);
    layer3_outputs(9441) <= not b;
    layer3_outputs(9442) <= not (a or b);
    layer3_outputs(9443) <= not b;
    layer3_outputs(9444) <= not a;
    layer3_outputs(9445) <= not (a and b);
    layer3_outputs(9446) <= not a or b;
    layer3_outputs(9447) <= not (a and b);
    layer3_outputs(9448) <= b;
    layer3_outputs(9449) <= not b or a;
    layer3_outputs(9450) <= a and b;
    layer3_outputs(9451) <= a or b;
    layer3_outputs(9452) <= not a or b;
    layer3_outputs(9453) <= not b;
    layer3_outputs(9454) <= a xor b;
    layer3_outputs(9455) <= not a or b;
    layer3_outputs(9456) <= b;
    layer3_outputs(9457) <= not b or a;
    layer3_outputs(9458) <= not a or b;
    layer3_outputs(9459) <= not a;
    layer3_outputs(9460) <= not b;
    layer3_outputs(9461) <= a and b;
    layer3_outputs(9462) <= not (a xor b);
    layer3_outputs(9463) <= a or b;
    layer3_outputs(9464) <= not a;
    layer3_outputs(9465) <= b;
    layer3_outputs(9466) <= a and b;
    layer3_outputs(9467) <= not a or b;
    layer3_outputs(9468) <= a xor b;
    layer3_outputs(9469) <= not a or b;
    layer3_outputs(9470) <= not b;
    layer3_outputs(9471) <= not b;
    layer3_outputs(9472) <= a xor b;
    layer3_outputs(9473) <= not a or b;
    layer3_outputs(9474) <= a and not b;
    layer3_outputs(9475) <= '1';
    layer3_outputs(9476) <= b and not a;
    layer3_outputs(9477) <= not a;
    layer3_outputs(9478) <= a and b;
    layer3_outputs(9479) <= not b;
    layer3_outputs(9480) <= a and not b;
    layer3_outputs(9481) <= b;
    layer3_outputs(9482) <= b and not a;
    layer3_outputs(9483) <= '1';
    layer3_outputs(9484) <= a and b;
    layer3_outputs(9485) <= a and b;
    layer3_outputs(9486) <= a or b;
    layer3_outputs(9487) <= not a;
    layer3_outputs(9488) <= b;
    layer3_outputs(9489) <= a;
    layer3_outputs(9490) <= b;
    layer3_outputs(9491) <= b and not a;
    layer3_outputs(9492) <= b and not a;
    layer3_outputs(9493) <= not b;
    layer3_outputs(9494) <= b;
    layer3_outputs(9495) <= not b;
    layer3_outputs(9496) <= b;
    layer3_outputs(9497) <= not (a and b);
    layer3_outputs(9498) <= a and not b;
    layer3_outputs(9499) <= not b;
    layer3_outputs(9500) <= a;
    layer3_outputs(9501) <= not b;
    layer3_outputs(9502) <= not (a or b);
    layer3_outputs(9503) <= not (a or b);
    layer3_outputs(9504) <= not (a xor b);
    layer3_outputs(9505) <= a and b;
    layer3_outputs(9506) <= a;
    layer3_outputs(9507) <= a;
    layer3_outputs(9508) <= not (a and b);
    layer3_outputs(9509) <= not (a and b);
    layer3_outputs(9510) <= a;
    layer3_outputs(9511) <= a or b;
    layer3_outputs(9512) <= not b;
    layer3_outputs(9513) <= b and not a;
    layer3_outputs(9514) <= a and b;
    layer3_outputs(9515) <= b;
    layer3_outputs(9516) <= b and not a;
    layer3_outputs(9517) <= b;
    layer3_outputs(9518) <= b and not a;
    layer3_outputs(9519) <= not b or a;
    layer3_outputs(9520) <= not b;
    layer3_outputs(9521) <= a or b;
    layer3_outputs(9522) <= not (a xor b);
    layer3_outputs(9523) <= not a;
    layer3_outputs(9524) <= a xor b;
    layer3_outputs(9525) <= a;
    layer3_outputs(9526) <= not a;
    layer3_outputs(9527) <= a and b;
    layer3_outputs(9528) <= not b;
    layer3_outputs(9529) <= a and b;
    layer3_outputs(9530) <= not (a and b);
    layer3_outputs(9531) <= not b;
    layer3_outputs(9532) <= '0';
    layer3_outputs(9533) <= not b or a;
    layer3_outputs(9534) <= not a or b;
    layer3_outputs(9535) <= a and not b;
    layer3_outputs(9536) <= not (a and b);
    layer3_outputs(9537) <= not b;
    layer3_outputs(9538) <= '1';
    layer3_outputs(9539) <= not b;
    layer3_outputs(9540) <= b and not a;
    layer3_outputs(9541) <= '1';
    layer3_outputs(9542) <= b and not a;
    layer3_outputs(9543) <= not a or b;
    layer3_outputs(9544) <= not a or b;
    layer3_outputs(9545) <= not a;
    layer3_outputs(9546) <= not (a or b);
    layer3_outputs(9547) <= not a;
    layer3_outputs(9548) <= not (a or b);
    layer3_outputs(9549) <= not b;
    layer3_outputs(9550) <= not a or b;
    layer3_outputs(9551) <= a and not b;
    layer3_outputs(9552) <= a xor b;
    layer3_outputs(9553) <= a and b;
    layer3_outputs(9554) <= a and not b;
    layer3_outputs(9555) <= a xor b;
    layer3_outputs(9556) <= not (a and b);
    layer3_outputs(9557) <= not (a and b);
    layer3_outputs(9558) <= a and not b;
    layer3_outputs(9559) <= a;
    layer3_outputs(9560) <= not b;
    layer3_outputs(9561) <= not (a or b);
    layer3_outputs(9562) <= not b;
    layer3_outputs(9563) <= a or b;
    layer3_outputs(9564) <= not b;
    layer3_outputs(9565) <= a;
    layer3_outputs(9566) <= not a or b;
    layer3_outputs(9567) <= a;
    layer3_outputs(9568) <= b;
    layer3_outputs(9569) <= not (a and b);
    layer3_outputs(9570) <= not (a and b);
    layer3_outputs(9571) <= a xor b;
    layer3_outputs(9572) <= a or b;
    layer3_outputs(9573) <= b;
    layer3_outputs(9574) <= b and not a;
    layer3_outputs(9575) <= a;
    layer3_outputs(9576) <= not b or a;
    layer3_outputs(9577) <= a or b;
    layer3_outputs(9578) <= b;
    layer3_outputs(9579) <= b;
    layer3_outputs(9580) <= not a;
    layer3_outputs(9581) <= not (a and b);
    layer3_outputs(9582) <= not (a xor b);
    layer3_outputs(9583) <= a and not b;
    layer3_outputs(9584) <= not b;
    layer3_outputs(9585) <= '1';
    layer3_outputs(9586) <= a and b;
    layer3_outputs(9587) <= a xor b;
    layer3_outputs(9588) <= a and b;
    layer3_outputs(9589) <= not a;
    layer3_outputs(9590) <= not a;
    layer3_outputs(9591) <= a or b;
    layer3_outputs(9592) <= b;
    layer3_outputs(9593) <= not (a xor b);
    layer3_outputs(9594) <= not (a and b);
    layer3_outputs(9595) <= b;
    layer3_outputs(9596) <= not a;
    layer3_outputs(9597) <= b;
    layer3_outputs(9598) <= not b;
    layer3_outputs(9599) <= a and not b;
    layer3_outputs(9600) <= '0';
    layer3_outputs(9601) <= a;
    layer3_outputs(9602) <= not a or b;
    layer3_outputs(9603) <= a and not b;
    layer3_outputs(9604) <= b;
    layer3_outputs(9605) <= not b;
    layer3_outputs(9606) <= not a or b;
    layer3_outputs(9607) <= a;
    layer3_outputs(9608) <= not (a and b);
    layer3_outputs(9609) <= not b or a;
    layer3_outputs(9610) <= not b;
    layer3_outputs(9611) <= b;
    layer3_outputs(9612) <= not (a xor b);
    layer3_outputs(9613) <= not b or a;
    layer3_outputs(9614) <= b;
    layer3_outputs(9615) <= a xor b;
    layer3_outputs(9616) <= not a or b;
    layer3_outputs(9617) <= b;
    layer3_outputs(9618) <= b and not a;
    layer3_outputs(9619) <= not b;
    layer3_outputs(9620) <= not (a and b);
    layer3_outputs(9621) <= not b or a;
    layer3_outputs(9622) <= a and b;
    layer3_outputs(9623) <= '1';
    layer3_outputs(9624) <= b;
    layer3_outputs(9625) <= b and not a;
    layer3_outputs(9626) <= not a;
    layer3_outputs(9627) <= a;
    layer3_outputs(9628) <= a or b;
    layer3_outputs(9629) <= not b or a;
    layer3_outputs(9630) <= a and not b;
    layer3_outputs(9631) <= not (a or b);
    layer3_outputs(9632) <= not (a xor b);
    layer3_outputs(9633) <= a;
    layer3_outputs(9634) <= not (a xor b);
    layer3_outputs(9635) <= not b;
    layer3_outputs(9636) <= not b or a;
    layer3_outputs(9637) <= a;
    layer3_outputs(9638) <= not b;
    layer3_outputs(9639) <= b;
    layer3_outputs(9640) <= a;
    layer3_outputs(9641) <= not (a xor b);
    layer3_outputs(9642) <= a;
    layer3_outputs(9643) <= a;
    layer3_outputs(9644) <= not (a or b);
    layer3_outputs(9645) <= not a;
    layer3_outputs(9646) <= a;
    layer3_outputs(9647) <= not a or b;
    layer3_outputs(9648) <= a xor b;
    layer3_outputs(9649) <= a;
    layer3_outputs(9650) <= a and b;
    layer3_outputs(9651) <= a and b;
    layer3_outputs(9652) <= not a or b;
    layer3_outputs(9653) <= not b;
    layer3_outputs(9654) <= not a or b;
    layer3_outputs(9655) <= b and not a;
    layer3_outputs(9656) <= a and b;
    layer3_outputs(9657) <= not a or b;
    layer3_outputs(9658) <= not b or a;
    layer3_outputs(9659) <= not (a or b);
    layer3_outputs(9660) <= a and b;
    layer3_outputs(9661) <= not (a or b);
    layer3_outputs(9662) <= not b or a;
    layer3_outputs(9663) <= not a;
    layer3_outputs(9664) <= not b;
    layer3_outputs(9665) <= not b;
    layer3_outputs(9666) <= not b;
    layer3_outputs(9667) <= b and not a;
    layer3_outputs(9668) <= b and not a;
    layer3_outputs(9669) <= not b;
    layer3_outputs(9670) <= not b;
    layer3_outputs(9671) <= not (a or b);
    layer3_outputs(9672) <= not (a xor b);
    layer3_outputs(9673) <= not (a xor b);
    layer3_outputs(9674) <= a and b;
    layer3_outputs(9675) <= a or b;
    layer3_outputs(9676) <= a or b;
    layer3_outputs(9677) <= not (a or b);
    layer3_outputs(9678) <= not b or a;
    layer3_outputs(9679) <= not b or a;
    layer3_outputs(9680) <= not (a or b);
    layer3_outputs(9681) <= not a;
    layer3_outputs(9682) <= not (a and b);
    layer3_outputs(9683) <= not a;
    layer3_outputs(9684) <= b;
    layer3_outputs(9685) <= a;
    layer3_outputs(9686) <= not (a and b);
    layer3_outputs(9687) <= a or b;
    layer3_outputs(9688) <= not a or b;
    layer3_outputs(9689) <= not b or a;
    layer3_outputs(9690) <= '1';
    layer3_outputs(9691) <= '1';
    layer3_outputs(9692) <= not (a and b);
    layer3_outputs(9693) <= not (a and b);
    layer3_outputs(9694) <= a or b;
    layer3_outputs(9695) <= b;
    layer3_outputs(9696) <= b and not a;
    layer3_outputs(9697) <= b and not a;
    layer3_outputs(9698) <= not b;
    layer3_outputs(9699) <= not b;
    layer3_outputs(9700) <= b and not a;
    layer3_outputs(9701) <= a and b;
    layer3_outputs(9702) <= a or b;
    layer3_outputs(9703) <= not (a and b);
    layer3_outputs(9704) <= b;
    layer3_outputs(9705) <= b;
    layer3_outputs(9706) <= b;
    layer3_outputs(9707) <= a or b;
    layer3_outputs(9708) <= a or b;
    layer3_outputs(9709) <= a and not b;
    layer3_outputs(9710) <= a;
    layer3_outputs(9711) <= not (a and b);
    layer3_outputs(9712) <= a;
    layer3_outputs(9713) <= a or b;
    layer3_outputs(9714) <= not (a or b);
    layer3_outputs(9715) <= not b;
    layer3_outputs(9716) <= '1';
    layer3_outputs(9717) <= b;
    layer3_outputs(9718) <= not a or b;
    layer3_outputs(9719) <= a;
    layer3_outputs(9720) <= not b;
    layer3_outputs(9721) <= not (a or b);
    layer3_outputs(9722) <= not a or b;
    layer3_outputs(9723) <= a;
    layer3_outputs(9724) <= not (a or b);
    layer3_outputs(9725) <= b;
    layer3_outputs(9726) <= b;
    layer3_outputs(9727) <= b;
    layer3_outputs(9728) <= b and not a;
    layer3_outputs(9729) <= b and not a;
    layer3_outputs(9730) <= b;
    layer3_outputs(9731) <= not (a or b);
    layer3_outputs(9732) <= b;
    layer3_outputs(9733) <= not b;
    layer3_outputs(9734) <= not b or a;
    layer3_outputs(9735) <= '0';
    layer3_outputs(9736) <= '1';
    layer3_outputs(9737) <= a xor b;
    layer3_outputs(9738) <= not a or b;
    layer3_outputs(9739) <= a and not b;
    layer3_outputs(9740) <= a or b;
    layer3_outputs(9741) <= b;
    layer3_outputs(9742) <= not (a or b);
    layer3_outputs(9743) <= not (a and b);
    layer3_outputs(9744) <= not (a and b);
    layer3_outputs(9745) <= b;
    layer3_outputs(9746) <= not a;
    layer3_outputs(9747) <= '0';
    layer3_outputs(9748) <= not b;
    layer3_outputs(9749) <= a or b;
    layer3_outputs(9750) <= a xor b;
    layer3_outputs(9751) <= not (a or b);
    layer3_outputs(9752) <= b;
    layer3_outputs(9753) <= not (a or b);
    layer3_outputs(9754) <= a;
    layer3_outputs(9755) <= not b;
    layer3_outputs(9756) <= a;
    layer3_outputs(9757) <= not (a and b);
    layer3_outputs(9758) <= not a;
    layer3_outputs(9759) <= a and b;
    layer3_outputs(9760) <= a and not b;
    layer3_outputs(9761) <= not (a or b);
    layer3_outputs(9762) <= not a;
    layer3_outputs(9763) <= not (a and b);
    layer3_outputs(9764) <= b and not a;
    layer3_outputs(9765) <= a xor b;
    layer3_outputs(9766) <= a or b;
    layer3_outputs(9767) <= not (a and b);
    layer3_outputs(9768) <= a or b;
    layer3_outputs(9769) <= b and not a;
    layer3_outputs(9770) <= a xor b;
    layer3_outputs(9771) <= not (a or b);
    layer3_outputs(9772) <= a;
    layer3_outputs(9773) <= not a;
    layer3_outputs(9774) <= a;
    layer3_outputs(9775) <= b and not a;
    layer3_outputs(9776) <= not (a or b);
    layer3_outputs(9777) <= not a;
    layer3_outputs(9778) <= a;
    layer3_outputs(9779) <= not (a and b);
    layer3_outputs(9780) <= not a;
    layer3_outputs(9781) <= not b;
    layer3_outputs(9782) <= b and not a;
    layer3_outputs(9783) <= b;
    layer3_outputs(9784) <= not a;
    layer3_outputs(9785) <= a or b;
    layer3_outputs(9786) <= a;
    layer3_outputs(9787) <= b and not a;
    layer3_outputs(9788) <= a;
    layer3_outputs(9789) <= a and not b;
    layer3_outputs(9790) <= a and not b;
    layer3_outputs(9791) <= not (a or b);
    layer3_outputs(9792) <= not a;
    layer3_outputs(9793) <= a and not b;
    layer3_outputs(9794) <= a and not b;
    layer3_outputs(9795) <= b;
    layer3_outputs(9796) <= '1';
    layer3_outputs(9797) <= not (a and b);
    layer3_outputs(9798) <= not a;
    layer3_outputs(9799) <= '0';
    layer3_outputs(9800) <= not a;
    layer3_outputs(9801) <= not b or a;
    layer3_outputs(9802) <= a and b;
    layer3_outputs(9803) <= not (a xor b);
    layer3_outputs(9804) <= a;
    layer3_outputs(9805) <= not b or a;
    layer3_outputs(9806) <= not b;
    layer3_outputs(9807) <= not a;
    layer3_outputs(9808) <= not a;
    layer3_outputs(9809) <= b;
    layer3_outputs(9810) <= a or b;
    layer3_outputs(9811) <= a and b;
    layer3_outputs(9812) <= '1';
    layer3_outputs(9813) <= not (a and b);
    layer3_outputs(9814) <= not b or a;
    layer3_outputs(9815) <= not a;
    layer3_outputs(9816) <= not a;
    layer3_outputs(9817) <= not b or a;
    layer3_outputs(9818) <= a;
    layer3_outputs(9819) <= not b;
    layer3_outputs(9820) <= not b;
    layer3_outputs(9821) <= b;
    layer3_outputs(9822) <= b and not a;
    layer3_outputs(9823) <= not b or a;
    layer3_outputs(9824) <= not (a or b);
    layer3_outputs(9825) <= a;
    layer3_outputs(9826) <= b and not a;
    layer3_outputs(9827) <= not (a and b);
    layer3_outputs(9828) <= '0';
    layer3_outputs(9829) <= b;
    layer3_outputs(9830) <= not a or b;
    layer3_outputs(9831) <= a and b;
    layer3_outputs(9832) <= not (a xor b);
    layer3_outputs(9833) <= '1';
    layer3_outputs(9834) <= not a or b;
    layer3_outputs(9835) <= a and not b;
    layer3_outputs(9836) <= '1';
    layer3_outputs(9837) <= not a;
    layer3_outputs(9838) <= b;
    layer3_outputs(9839) <= b;
    layer3_outputs(9840) <= a and not b;
    layer3_outputs(9841) <= not b or a;
    layer3_outputs(9842) <= b;
    layer3_outputs(9843) <= b;
    layer3_outputs(9844) <= not b;
    layer3_outputs(9845) <= a and b;
    layer3_outputs(9846) <= b;
    layer3_outputs(9847) <= not b or a;
    layer3_outputs(9848) <= not b;
    layer3_outputs(9849) <= not (a or b);
    layer3_outputs(9850) <= a and b;
    layer3_outputs(9851) <= a;
    layer3_outputs(9852) <= a and not b;
    layer3_outputs(9853) <= not a;
    layer3_outputs(9854) <= a and not b;
    layer3_outputs(9855) <= '0';
    layer3_outputs(9856) <= not a or b;
    layer3_outputs(9857) <= b;
    layer3_outputs(9858) <= b;
    layer3_outputs(9859) <= not b;
    layer3_outputs(9860) <= a;
    layer3_outputs(9861) <= a;
    layer3_outputs(9862) <= not a or b;
    layer3_outputs(9863) <= a;
    layer3_outputs(9864) <= not b;
    layer3_outputs(9865) <= a and not b;
    layer3_outputs(9866) <= '0';
    layer3_outputs(9867) <= b;
    layer3_outputs(9868) <= b;
    layer3_outputs(9869) <= b and not a;
    layer3_outputs(9870) <= a;
    layer3_outputs(9871) <= not b or a;
    layer3_outputs(9872) <= a;
    layer3_outputs(9873) <= '1';
    layer3_outputs(9874) <= a and not b;
    layer3_outputs(9875) <= not b or a;
    layer3_outputs(9876) <= a and b;
    layer3_outputs(9877) <= not b;
    layer3_outputs(9878) <= a and b;
    layer3_outputs(9879) <= a and not b;
    layer3_outputs(9880) <= not b;
    layer3_outputs(9881) <= b and not a;
    layer3_outputs(9882) <= not b;
    layer3_outputs(9883) <= a and not b;
    layer3_outputs(9884) <= not b;
    layer3_outputs(9885) <= a;
    layer3_outputs(9886) <= not (a xor b);
    layer3_outputs(9887) <= b;
    layer3_outputs(9888) <= b and not a;
    layer3_outputs(9889) <= not (a and b);
    layer3_outputs(9890) <= a and not b;
    layer3_outputs(9891) <= '0';
    layer3_outputs(9892) <= '1';
    layer3_outputs(9893) <= not a or b;
    layer3_outputs(9894) <= a;
    layer3_outputs(9895) <= '0';
    layer3_outputs(9896) <= b;
    layer3_outputs(9897) <= a;
    layer3_outputs(9898) <= a and not b;
    layer3_outputs(9899) <= a xor b;
    layer3_outputs(9900) <= a or b;
    layer3_outputs(9901) <= not b or a;
    layer3_outputs(9902) <= a xor b;
    layer3_outputs(9903) <= not a;
    layer3_outputs(9904) <= b and not a;
    layer3_outputs(9905) <= b and not a;
    layer3_outputs(9906) <= not b;
    layer3_outputs(9907) <= not b;
    layer3_outputs(9908) <= not a or b;
    layer3_outputs(9909) <= not b;
    layer3_outputs(9910) <= not b;
    layer3_outputs(9911) <= a and b;
    layer3_outputs(9912) <= a;
    layer3_outputs(9913) <= not a or b;
    layer3_outputs(9914) <= not b;
    layer3_outputs(9915) <= not a;
    layer3_outputs(9916) <= not b or a;
    layer3_outputs(9917) <= a;
    layer3_outputs(9918) <= b;
    layer3_outputs(9919) <= '1';
    layer3_outputs(9920) <= not (a or b);
    layer3_outputs(9921) <= a xor b;
    layer3_outputs(9922) <= '1';
    layer3_outputs(9923) <= not a or b;
    layer3_outputs(9924) <= a and not b;
    layer3_outputs(9925) <= not (a and b);
    layer3_outputs(9926) <= b and not a;
    layer3_outputs(9927) <= a or b;
    layer3_outputs(9928) <= not a;
    layer3_outputs(9929) <= b;
    layer3_outputs(9930) <= '0';
    layer3_outputs(9931) <= a and not b;
    layer3_outputs(9932) <= not (a and b);
    layer3_outputs(9933) <= not a;
    layer3_outputs(9934) <= b;
    layer3_outputs(9935) <= b and not a;
    layer3_outputs(9936) <= a and b;
    layer3_outputs(9937) <= not (a or b);
    layer3_outputs(9938) <= a and b;
    layer3_outputs(9939) <= a or b;
    layer3_outputs(9940) <= a xor b;
    layer3_outputs(9941) <= not (a and b);
    layer3_outputs(9942) <= not a;
    layer3_outputs(9943) <= b;
    layer3_outputs(9944) <= a;
    layer3_outputs(9945) <= a and b;
    layer3_outputs(9946) <= not b;
    layer3_outputs(9947) <= b and not a;
    layer3_outputs(9948) <= a;
    layer3_outputs(9949) <= not b;
    layer3_outputs(9950) <= '0';
    layer3_outputs(9951) <= a and b;
    layer3_outputs(9952) <= a;
    layer3_outputs(9953) <= not a or b;
    layer3_outputs(9954) <= '0';
    layer3_outputs(9955) <= not (a and b);
    layer3_outputs(9956) <= a;
    layer3_outputs(9957) <= a and b;
    layer3_outputs(9958) <= a and b;
    layer3_outputs(9959) <= not (a xor b);
    layer3_outputs(9960) <= not b;
    layer3_outputs(9961) <= not b;
    layer3_outputs(9962) <= a or b;
    layer3_outputs(9963) <= a;
    layer3_outputs(9964) <= not a or b;
    layer3_outputs(9965) <= not b;
    layer3_outputs(9966) <= a;
    layer3_outputs(9967) <= not (a or b);
    layer3_outputs(9968) <= not b;
    layer3_outputs(9969) <= a;
    layer3_outputs(9970) <= not a;
    layer3_outputs(9971) <= a and b;
    layer3_outputs(9972) <= a and b;
    layer3_outputs(9973) <= not a;
    layer3_outputs(9974) <= '0';
    layer3_outputs(9975) <= b;
    layer3_outputs(9976) <= '0';
    layer3_outputs(9977) <= a and b;
    layer3_outputs(9978) <= b;
    layer3_outputs(9979) <= b and not a;
    layer3_outputs(9980) <= a or b;
    layer3_outputs(9981) <= not a;
    layer3_outputs(9982) <= b;
    layer3_outputs(9983) <= a and b;
    layer3_outputs(9984) <= a and b;
    layer3_outputs(9985) <= a and b;
    layer3_outputs(9986) <= a;
    layer3_outputs(9987) <= not b;
    layer3_outputs(9988) <= a and b;
    layer3_outputs(9989) <= a;
    layer3_outputs(9990) <= not (a xor b);
    layer3_outputs(9991) <= a;
    layer3_outputs(9992) <= not a;
    layer3_outputs(9993) <= not b or a;
    layer3_outputs(9994) <= '1';
    layer3_outputs(9995) <= b;
    layer3_outputs(9996) <= b;
    layer3_outputs(9997) <= a and b;
    layer3_outputs(9998) <= not b;
    layer3_outputs(9999) <= b;
    layer3_outputs(10000) <= not b;
    layer3_outputs(10001) <= not (a xor b);
    layer3_outputs(10002) <= '0';
    layer3_outputs(10003) <= b and not a;
    layer3_outputs(10004) <= not (a and b);
    layer3_outputs(10005) <= not (a or b);
    layer3_outputs(10006) <= a and not b;
    layer3_outputs(10007) <= b;
    layer3_outputs(10008) <= not b;
    layer3_outputs(10009) <= not a or b;
    layer3_outputs(10010) <= not (a or b);
    layer3_outputs(10011) <= a;
    layer3_outputs(10012) <= b and not a;
    layer3_outputs(10013) <= a or b;
    layer3_outputs(10014) <= not (a and b);
    layer3_outputs(10015) <= a xor b;
    layer3_outputs(10016) <= b and not a;
    layer3_outputs(10017) <= not b;
    layer3_outputs(10018) <= b and not a;
    layer3_outputs(10019) <= not (a and b);
    layer3_outputs(10020) <= not b or a;
    layer3_outputs(10021) <= b;
    layer3_outputs(10022) <= not b or a;
    layer3_outputs(10023) <= b and not a;
    layer3_outputs(10024) <= b;
    layer3_outputs(10025) <= not a;
    layer3_outputs(10026) <= b and not a;
    layer3_outputs(10027) <= a;
    layer3_outputs(10028) <= a or b;
    layer3_outputs(10029) <= a and not b;
    layer3_outputs(10030) <= not a or b;
    layer3_outputs(10031) <= a xor b;
    layer3_outputs(10032) <= not a;
    layer3_outputs(10033) <= a and not b;
    layer3_outputs(10034) <= b;
    layer3_outputs(10035) <= a and not b;
    layer3_outputs(10036) <= a;
    layer3_outputs(10037) <= not (a and b);
    layer3_outputs(10038) <= a and not b;
    layer3_outputs(10039) <= b and not a;
    layer3_outputs(10040) <= not (a or b);
    layer3_outputs(10041) <= a;
    layer3_outputs(10042) <= a or b;
    layer3_outputs(10043) <= b;
    layer3_outputs(10044) <= a or b;
    layer3_outputs(10045) <= not a or b;
    layer3_outputs(10046) <= not b or a;
    layer3_outputs(10047) <= not (a or b);
    layer3_outputs(10048) <= a xor b;
    layer3_outputs(10049) <= not b;
    layer3_outputs(10050) <= not b or a;
    layer3_outputs(10051) <= not b;
    layer3_outputs(10052) <= not a;
    layer3_outputs(10053) <= not a or b;
    layer3_outputs(10054) <= a;
    layer3_outputs(10055) <= a or b;
    layer3_outputs(10056) <= not (a xor b);
    layer3_outputs(10057) <= a;
    layer3_outputs(10058) <= b;
    layer3_outputs(10059) <= a;
    layer3_outputs(10060) <= not (a xor b);
    layer3_outputs(10061) <= b;
    layer3_outputs(10062) <= not a or b;
    layer3_outputs(10063) <= '1';
    layer3_outputs(10064) <= a;
    layer3_outputs(10065) <= not b;
    layer3_outputs(10066) <= a and not b;
    layer3_outputs(10067) <= not (a or b);
    layer3_outputs(10068) <= a and b;
    layer3_outputs(10069) <= a;
    layer3_outputs(10070) <= not (a and b);
    layer3_outputs(10071) <= not b;
    layer3_outputs(10072) <= not b;
    layer3_outputs(10073) <= not (a xor b);
    layer3_outputs(10074) <= not (a and b);
    layer3_outputs(10075) <= b and not a;
    layer3_outputs(10076) <= not b;
    layer3_outputs(10077) <= a or b;
    layer3_outputs(10078) <= not b;
    layer3_outputs(10079) <= b and not a;
    layer3_outputs(10080) <= not a;
    layer3_outputs(10081) <= not b;
    layer3_outputs(10082) <= not a;
    layer3_outputs(10083) <= not (a and b);
    layer3_outputs(10084) <= not a;
    layer3_outputs(10085) <= not (a and b);
    layer3_outputs(10086) <= b and not a;
    layer3_outputs(10087) <= not a;
    layer3_outputs(10088) <= b;
    layer3_outputs(10089) <= a xor b;
    layer3_outputs(10090) <= not a or b;
    layer3_outputs(10091) <= a;
    layer3_outputs(10092) <= '0';
    layer3_outputs(10093) <= a and not b;
    layer3_outputs(10094) <= a or b;
    layer3_outputs(10095) <= b and not a;
    layer3_outputs(10096) <= '0';
    layer3_outputs(10097) <= '0';
    layer3_outputs(10098) <= not (a and b);
    layer3_outputs(10099) <= not b or a;
    layer3_outputs(10100) <= a and b;
    layer3_outputs(10101) <= not b;
    layer3_outputs(10102) <= not a;
    layer3_outputs(10103) <= not (a or b);
    layer3_outputs(10104) <= not a or b;
    layer3_outputs(10105) <= '1';
    layer3_outputs(10106) <= not (a and b);
    layer3_outputs(10107) <= not (a or b);
    layer3_outputs(10108) <= not b or a;
    layer3_outputs(10109) <= not (a or b);
    layer3_outputs(10110) <= not (a xor b);
    layer3_outputs(10111) <= not a;
    layer3_outputs(10112) <= a and not b;
    layer3_outputs(10113) <= not a or b;
    layer3_outputs(10114) <= a and not b;
    layer3_outputs(10115) <= a;
    layer3_outputs(10116) <= not (a and b);
    layer3_outputs(10117) <= a and not b;
    layer3_outputs(10118) <= not a or b;
    layer3_outputs(10119) <= not b;
    layer3_outputs(10120) <= a or b;
    layer3_outputs(10121) <= not a or b;
    layer3_outputs(10122) <= b and not a;
    layer3_outputs(10123) <= '1';
    layer3_outputs(10124) <= not b or a;
    layer3_outputs(10125) <= a and not b;
    layer3_outputs(10126) <= a and b;
    layer3_outputs(10127) <= not b or a;
    layer3_outputs(10128) <= b;
    layer3_outputs(10129) <= not a;
    layer3_outputs(10130) <= not (a or b);
    layer3_outputs(10131) <= not a;
    layer3_outputs(10132) <= b and not a;
    layer3_outputs(10133) <= not b;
    layer3_outputs(10134) <= not a;
    layer3_outputs(10135) <= not b;
    layer3_outputs(10136) <= a and b;
    layer3_outputs(10137) <= a or b;
    layer3_outputs(10138) <= not b;
    layer3_outputs(10139) <= not b;
    layer3_outputs(10140) <= a;
    layer3_outputs(10141) <= a;
    layer3_outputs(10142) <= not a or b;
    layer3_outputs(10143) <= not (a and b);
    layer3_outputs(10144) <= not a;
    layer3_outputs(10145) <= b and not a;
    layer3_outputs(10146) <= b;
    layer3_outputs(10147) <= b;
    layer3_outputs(10148) <= not a or b;
    layer3_outputs(10149) <= a and b;
    layer3_outputs(10150) <= a or b;
    layer3_outputs(10151) <= '0';
    layer3_outputs(10152) <= not (a and b);
    layer3_outputs(10153) <= not (a or b);
    layer3_outputs(10154) <= '1';
    layer3_outputs(10155) <= a or b;
    layer3_outputs(10156) <= not (a and b);
    layer3_outputs(10157) <= not (a or b);
    layer3_outputs(10158) <= not (a xor b);
    layer3_outputs(10159) <= a and not b;
    layer3_outputs(10160) <= a and b;
    layer3_outputs(10161) <= a;
    layer3_outputs(10162) <= a and not b;
    layer3_outputs(10163) <= not a;
    layer3_outputs(10164) <= not (a or b);
    layer3_outputs(10165) <= not a;
    layer3_outputs(10166) <= a or b;
    layer3_outputs(10167) <= not a;
    layer3_outputs(10168) <= a;
    layer3_outputs(10169) <= not b;
    layer3_outputs(10170) <= a;
    layer3_outputs(10171) <= not a or b;
    layer3_outputs(10172) <= b and not a;
    layer3_outputs(10173) <= a;
    layer3_outputs(10174) <= b;
    layer3_outputs(10175) <= not a or b;
    layer3_outputs(10176) <= a;
    layer3_outputs(10177) <= a or b;
    layer3_outputs(10178) <= a and not b;
    layer3_outputs(10179) <= a;
    layer3_outputs(10180) <= not b;
    layer3_outputs(10181) <= not a;
    layer3_outputs(10182) <= not b;
    layer3_outputs(10183) <= not (a and b);
    layer3_outputs(10184) <= a;
    layer3_outputs(10185) <= not b;
    layer3_outputs(10186) <= b and not a;
    layer3_outputs(10187) <= not (a and b);
    layer3_outputs(10188) <= b and not a;
    layer3_outputs(10189) <= not b or a;
    layer3_outputs(10190) <= not b;
    layer3_outputs(10191) <= '0';
    layer3_outputs(10192) <= not (a xor b);
    layer3_outputs(10193) <= not b or a;
    layer3_outputs(10194) <= not (a and b);
    layer3_outputs(10195) <= not a or b;
    layer3_outputs(10196) <= not b;
    layer3_outputs(10197) <= not (a and b);
    layer3_outputs(10198) <= b;
    layer3_outputs(10199) <= '1';
    layer3_outputs(10200) <= b and not a;
    layer3_outputs(10201) <= not b or a;
    layer3_outputs(10202) <= not (a or b);
    layer3_outputs(10203) <= b and not a;
    layer3_outputs(10204) <= not b;
    layer3_outputs(10205) <= not b;
    layer3_outputs(10206) <= a and not b;
    layer3_outputs(10207) <= a or b;
    layer3_outputs(10208) <= a;
    layer3_outputs(10209) <= not (a and b);
    layer3_outputs(10210) <= a;
    layer3_outputs(10211) <= b;
    layer3_outputs(10212) <= b;
    layer3_outputs(10213) <= a or b;
    layer3_outputs(10214) <= not a or b;
    layer3_outputs(10215) <= not (a xor b);
    layer3_outputs(10216) <= b and not a;
    layer3_outputs(10217) <= not b or a;
    layer3_outputs(10218) <= b and not a;
    layer3_outputs(10219) <= '0';
    layer3_outputs(10220) <= not (a or b);
    layer3_outputs(10221) <= not a;
    layer3_outputs(10222) <= a;
    layer3_outputs(10223) <= not (a or b);
    layer3_outputs(10224) <= '1';
    layer3_outputs(10225) <= not (a or b);
    layer3_outputs(10226) <= a or b;
    layer3_outputs(10227) <= '1';
    layer3_outputs(10228) <= a xor b;
    layer3_outputs(10229) <= not b;
    layer3_outputs(10230) <= b and not a;
    layer3_outputs(10231) <= not a;
    layer3_outputs(10232) <= not b or a;
    layer3_outputs(10233) <= '1';
    layer3_outputs(10234) <= b;
    layer3_outputs(10235) <= not b;
    layer3_outputs(10236) <= not a;
    layer3_outputs(10237) <= a;
    layer3_outputs(10238) <= not b;
    layer3_outputs(10239) <= '1';
    layer4_outputs(0) <= a or b;
    layer4_outputs(1) <= not a;
    layer4_outputs(2) <= not a or b;
    layer4_outputs(3) <= a;
    layer4_outputs(4) <= a;
    layer4_outputs(5) <= b and not a;
    layer4_outputs(6) <= not a;
    layer4_outputs(7) <= a or b;
    layer4_outputs(8) <= a or b;
    layer4_outputs(9) <= b;
    layer4_outputs(10) <= a;
    layer4_outputs(11) <= b and not a;
    layer4_outputs(12) <= not b;
    layer4_outputs(13) <= a and b;
    layer4_outputs(14) <= a or b;
    layer4_outputs(15) <= not b or a;
    layer4_outputs(16) <= not b;
    layer4_outputs(17) <= a;
    layer4_outputs(18) <= a and not b;
    layer4_outputs(19) <= a;
    layer4_outputs(20) <= not b;
    layer4_outputs(21) <= a;
    layer4_outputs(22) <= a;
    layer4_outputs(23) <= not (a or b);
    layer4_outputs(24) <= a;
    layer4_outputs(25) <= not b;
    layer4_outputs(26) <= a;
    layer4_outputs(27) <= b;
    layer4_outputs(28) <= '1';
    layer4_outputs(29) <= not a or b;
    layer4_outputs(30) <= a and b;
    layer4_outputs(31) <= a or b;
    layer4_outputs(32) <= not a;
    layer4_outputs(33) <= a xor b;
    layer4_outputs(34) <= not a;
    layer4_outputs(35) <= b and not a;
    layer4_outputs(36) <= a and not b;
    layer4_outputs(37) <= b;
    layer4_outputs(38) <= not a;
    layer4_outputs(39) <= a and not b;
    layer4_outputs(40) <= not b or a;
    layer4_outputs(41) <= not a;
    layer4_outputs(42) <= a;
    layer4_outputs(43) <= a and b;
    layer4_outputs(44) <= not a or b;
    layer4_outputs(45) <= a or b;
    layer4_outputs(46) <= b;
    layer4_outputs(47) <= not (a or b);
    layer4_outputs(48) <= not (a and b);
    layer4_outputs(49) <= b;
    layer4_outputs(50) <= not (a and b);
    layer4_outputs(51) <= '0';
    layer4_outputs(52) <= not (a and b);
    layer4_outputs(53) <= b;
    layer4_outputs(54) <= a and not b;
    layer4_outputs(55) <= a and b;
    layer4_outputs(56) <= b and not a;
    layer4_outputs(57) <= not a;
    layer4_outputs(58) <= b;
    layer4_outputs(59) <= a and b;
    layer4_outputs(60) <= a and not b;
    layer4_outputs(61) <= '1';
    layer4_outputs(62) <= not b;
    layer4_outputs(63) <= not b;
    layer4_outputs(64) <= not (a xor b);
    layer4_outputs(65) <= not b or a;
    layer4_outputs(66) <= not (a or b);
    layer4_outputs(67) <= a and b;
    layer4_outputs(68) <= b and not a;
    layer4_outputs(69) <= not b;
    layer4_outputs(70) <= not a;
    layer4_outputs(71) <= not (a xor b);
    layer4_outputs(72) <= not b;
    layer4_outputs(73) <= not a or b;
    layer4_outputs(74) <= not (a or b);
    layer4_outputs(75) <= a xor b;
    layer4_outputs(76) <= not (a xor b);
    layer4_outputs(77) <= not (a xor b);
    layer4_outputs(78) <= not a;
    layer4_outputs(79) <= a xor b;
    layer4_outputs(80) <= not (a xor b);
    layer4_outputs(81) <= not (a and b);
    layer4_outputs(82) <= not a;
    layer4_outputs(83) <= b;
    layer4_outputs(84) <= not b;
    layer4_outputs(85) <= not b;
    layer4_outputs(86) <= a;
    layer4_outputs(87) <= a;
    layer4_outputs(88) <= a and not b;
    layer4_outputs(89) <= a xor b;
    layer4_outputs(90) <= not (a or b);
    layer4_outputs(91) <= a and not b;
    layer4_outputs(92) <= a and b;
    layer4_outputs(93) <= a and not b;
    layer4_outputs(94) <= not (a or b);
    layer4_outputs(95) <= a or b;
    layer4_outputs(96) <= not b or a;
    layer4_outputs(97) <= a;
    layer4_outputs(98) <= not b;
    layer4_outputs(99) <= b;
    layer4_outputs(100) <= not b or a;
    layer4_outputs(101) <= not b;
    layer4_outputs(102) <= not a;
    layer4_outputs(103) <= a or b;
    layer4_outputs(104) <= b and not a;
    layer4_outputs(105) <= a and not b;
    layer4_outputs(106) <= not b;
    layer4_outputs(107) <= not (a xor b);
    layer4_outputs(108) <= not b or a;
    layer4_outputs(109) <= not b or a;
    layer4_outputs(110) <= a;
    layer4_outputs(111) <= not a or b;
    layer4_outputs(112) <= not (a or b);
    layer4_outputs(113) <= not (a and b);
    layer4_outputs(114) <= a;
    layer4_outputs(115) <= not a;
    layer4_outputs(116) <= a xor b;
    layer4_outputs(117) <= a and not b;
    layer4_outputs(118) <= not b;
    layer4_outputs(119) <= not (a or b);
    layer4_outputs(120) <= not b;
    layer4_outputs(121) <= not b or a;
    layer4_outputs(122) <= a;
    layer4_outputs(123) <= a and b;
    layer4_outputs(124) <= a and b;
    layer4_outputs(125) <= not (a xor b);
    layer4_outputs(126) <= not a or b;
    layer4_outputs(127) <= '0';
    layer4_outputs(128) <= not b or a;
    layer4_outputs(129) <= not (a and b);
    layer4_outputs(130) <= not a;
    layer4_outputs(131) <= not a;
    layer4_outputs(132) <= not (a or b);
    layer4_outputs(133) <= b;
    layer4_outputs(134) <= a or b;
    layer4_outputs(135) <= not (a or b);
    layer4_outputs(136) <= not a;
    layer4_outputs(137) <= not b;
    layer4_outputs(138) <= not b;
    layer4_outputs(139) <= a;
    layer4_outputs(140) <= not (a or b);
    layer4_outputs(141) <= not a;
    layer4_outputs(142) <= a;
    layer4_outputs(143) <= '0';
    layer4_outputs(144) <= a;
    layer4_outputs(145) <= b;
    layer4_outputs(146) <= a xor b;
    layer4_outputs(147) <= a;
    layer4_outputs(148) <= not (a or b);
    layer4_outputs(149) <= not (a or b);
    layer4_outputs(150) <= not b;
    layer4_outputs(151) <= a and b;
    layer4_outputs(152) <= not (a or b);
    layer4_outputs(153) <= a;
    layer4_outputs(154) <= a and not b;
    layer4_outputs(155) <= b and not a;
    layer4_outputs(156) <= b;
    layer4_outputs(157) <= not b;
    layer4_outputs(158) <= not (a or b);
    layer4_outputs(159) <= not (a or b);
    layer4_outputs(160) <= a or b;
    layer4_outputs(161) <= not a;
    layer4_outputs(162) <= not b or a;
    layer4_outputs(163) <= not (a or b);
    layer4_outputs(164) <= not b;
    layer4_outputs(165) <= a and not b;
    layer4_outputs(166) <= not (a or b);
    layer4_outputs(167) <= b and not a;
    layer4_outputs(168) <= not b or a;
    layer4_outputs(169) <= b and not a;
    layer4_outputs(170) <= b and not a;
    layer4_outputs(171) <= b and not a;
    layer4_outputs(172) <= a;
    layer4_outputs(173) <= not (a and b);
    layer4_outputs(174) <= a;
    layer4_outputs(175) <= b and not a;
    layer4_outputs(176) <= a and not b;
    layer4_outputs(177) <= a xor b;
    layer4_outputs(178) <= a and not b;
    layer4_outputs(179) <= a or b;
    layer4_outputs(180) <= a;
    layer4_outputs(181) <= not b or a;
    layer4_outputs(182) <= a xor b;
    layer4_outputs(183) <= a;
    layer4_outputs(184) <= not (a xor b);
    layer4_outputs(185) <= a or b;
    layer4_outputs(186) <= not a or b;
    layer4_outputs(187) <= not b;
    layer4_outputs(188) <= not b;
    layer4_outputs(189) <= not b;
    layer4_outputs(190) <= a xor b;
    layer4_outputs(191) <= a and b;
    layer4_outputs(192) <= not a;
    layer4_outputs(193) <= a;
    layer4_outputs(194) <= a xor b;
    layer4_outputs(195) <= b;
    layer4_outputs(196) <= b;
    layer4_outputs(197) <= b;
    layer4_outputs(198) <= a;
    layer4_outputs(199) <= not a or b;
    layer4_outputs(200) <= a or b;
    layer4_outputs(201) <= not a;
    layer4_outputs(202) <= not (a xor b);
    layer4_outputs(203) <= not b or a;
    layer4_outputs(204) <= b;
    layer4_outputs(205) <= not b;
    layer4_outputs(206) <= not (a and b);
    layer4_outputs(207) <= not (a xor b);
    layer4_outputs(208) <= not (a or b);
    layer4_outputs(209) <= not a or b;
    layer4_outputs(210) <= not (a or b);
    layer4_outputs(211) <= a;
    layer4_outputs(212) <= a;
    layer4_outputs(213) <= b;
    layer4_outputs(214) <= a and b;
    layer4_outputs(215) <= not b or a;
    layer4_outputs(216) <= not (a and b);
    layer4_outputs(217) <= '0';
    layer4_outputs(218) <= not a or b;
    layer4_outputs(219) <= b and not a;
    layer4_outputs(220) <= b;
    layer4_outputs(221) <= not (a or b);
    layer4_outputs(222) <= b and not a;
    layer4_outputs(223) <= a;
    layer4_outputs(224) <= a and not b;
    layer4_outputs(225) <= not (a and b);
    layer4_outputs(226) <= not (a or b);
    layer4_outputs(227) <= not (a or b);
    layer4_outputs(228) <= a;
    layer4_outputs(229) <= not b;
    layer4_outputs(230) <= a and b;
    layer4_outputs(231) <= not b;
    layer4_outputs(232) <= not (a and b);
    layer4_outputs(233) <= not a;
    layer4_outputs(234) <= '0';
    layer4_outputs(235) <= '0';
    layer4_outputs(236) <= a or b;
    layer4_outputs(237) <= a or b;
    layer4_outputs(238) <= a and not b;
    layer4_outputs(239) <= a;
    layer4_outputs(240) <= a xor b;
    layer4_outputs(241) <= '1';
    layer4_outputs(242) <= not (a xor b);
    layer4_outputs(243) <= '1';
    layer4_outputs(244) <= b and not a;
    layer4_outputs(245) <= a and not b;
    layer4_outputs(246) <= not b;
    layer4_outputs(247) <= a or b;
    layer4_outputs(248) <= a and b;
    layer4_outputs(249) <= b and not a;
    layer4_outputs(250) <= a and b;
    layer4_outputs(251) <= a and b;
    layer4_outputs(252) <= not a or b;
    layer4_outputs(253) <= not a or b;
    layer4_outputs(254) <= a or b;
    layer4_outputs(255) <= not (a and b);
    layer4_outputs(256) <= a;
    layer4_outputs(257) <= not (a and b);
    layer4_outputs(258) <= '1';
    layer4_outputs(259) <= b and not a;
    layer4_outputs(260) <= not (a xor b);
    layer4_outputs(261) <= not (a xor b);
    layer4_outputs(262) <= b and not a;
    layer4_outputs(263) <= b and not a;
    layer4_outputs(264) <= not b or a;
    layer4_outputs(265) <= not (a xor b);
    layer4_outputs(266) <= a;
    layer4_outputs(267) <= a and b;
    layer4_outputs(268) <= a or b;
    layer4_outputs(269) <= b and not a;
    layer4_outputs(270) <= a xor b;
    layer4_outputs(271) <= not b;
    layer4_outputs(272) <= not (a xor b);
    layer4_outputs(273) <= not a;
    layer4_outputs(274) <= a or b;
    layer4_outputs(275) <= '0';
    layer4_outputs(276) <= a or b;
    layer4_outputs(277) <= not b or a;
    layer4_outputs(278) <= a;
    layer4_outputs(279) <= not a;
    layer4_outputs(280) <= a;
    layer4_outputs(281) <= a or b;
    layer4_outputs(282) <= not a;
    layer4_outputs(283) <= a or b;
    layer4_outputs(284) <= b and not a;
    layer4_outputs(285) <= not a or b;
    layer4_outputs(286) <= not b;
    layer4_outputs(287) <= not a;
    layer4_outputs(288) <= not (a xor b);
    layer4_outputs(289) <= not a;
    layer4_outputs(290) <= a and b;
    layer4_outputs(291) <= not a or b;
    layer4_outputs(292) <= '0';
    layer4_outputs(293) <= a and b;
    layer4_outputs(294) <= not a or b;
    layer4_outputs(295) <= b;
    layer4_outputs(296) <= not b or a;
    layer4_outputs(297) <= b and not a;
    layer4_outputs(298) <= not a or b;
    layer4_outputs(299) <= not b or a;
    layer4_outputs(300) <= not (a and b);
    layer4_outputs(301) <= '1';
    layer4_outputs(302) <= not a;
    layer4_outputs(303) <= '0';
    layer4_outputs(304) <= not a;
    layer4_outputs(305) <= b;
    layer4_outputs(306) <= b;
    layer4_outputs(307) <= not b;
    layer4_outputs(308) <= not b;
    layer4_outputs(309) <= a;
    layer4_outputs(310) <= not (a and b);
    layer4_outputs(311) <= not b;
    layer4_outputs(312) <= not b;
    layer4_outputs(313) <= a xor b;
    layer4_outputs(314) <= '0';
    layer4_outputs(315) <= a;
    layer4_outputs(316) <= not a;
    layer4_outputs(317) <= a xor b;
    layer4_outputs(318) <= a and b;
    layer4_outputs(319) <= a and not b;
    layer4_outputs(320) <= not b;
    layer4_outputs(321) <= a xor b;
    layer4_outputs(322) <= b;
    layer4_outputs(323) <= a and not b;
    layer4_outputs(324) <= not (a and b);
    layer4_outputs(325) <= not a;
    layer4_outputs(326) <= not a or b;
    layer4_outputs(327) <= not (a and b);
    layer4_outputs(328) <= not (a xor b);
    layer4_outputs(329) <= not a;
    layer4_outputs(330) <= a and b;
    layer4_outputs(331) <= a or b;
    layer4_outputs(332) <= not b;
    layer4_outputs(333) <= not b;
    layer4_outputs(334) <= a;
    layer4_outputs(335) <= a and not b;
    layer4_outputs(336) <= not b or a;
    layer4_outputs(337) <= a or b;
    layer4_outputs(338) <= b and not a;
    layer4_outputs(339) <= not b;
    layer4_outputs(340) <= b;
    layer4_outputs(341) <= a;
    layer4_outputs(342) <= a;
    layer4_outputs(343) <= not a;
    layer4_outputs(344) <= not (a xor b);
    layer4_outputs(345) <= not a;
    layer4_outputs(346) <= not (a and b);
    layer4_outputs(347) <= a and not b;
    layer4_outputs(348) <= a xor b;
    layer4_outputs(349) <= not b;
    layer4_outputs(350) <= a xor b;
    layer4_outputs(351) <= a and not b;
    layer4_outputs(352) <= not a;
    layer4_outputs(353) <= not b;
    layer4_outputs(354) <= not (a or b);
    layer4_outputs(355) <= not a;
    layer4_outputs(356) <= b;
    layer4_outputs(357) <= a;
    layer4_outputs(358) <= b;
    layer4_outputs(359) <= b and not a;
    layer4_outputs(360) <= a and not b;
    layer4_outputs(361) <= '0';
    layer4_outputs(362) <= a and b;
    layer4_outputs(363) <= a and b;
    layer4_outputs(364) <= not b or a;
    layer4_outputs(365) <= not (a and b);
    layer4_outputs(366) <= not (a and b);
    layer4_outputs(367) <= not b or a;
    layer4_outputs(368) <= not a;
    layer4_outputs(369) <= a and b;
    layer4_outputs(370) <= a;
    layer4_outputs(371) <= b and not a;
    layer4_outputs(372) <= b and not a;
    layer4_outputs(373) <= a or b;
    layer4_outputs(374) <= b;
    layer4_outputs(375) <= b;
    layer4_outputs(376) <= b;
    layer4_outputs(377) <= a and not b;
    layer4_outputs(378) <= b;
    layer4_outputs(379) <= not b;
    layer4_outputs(380) <= not a or b;
    layer4_outputs(381) <= a and b;
    layer4_outputs(382) <= not (a or b);
    layer4_outputs(383) <= not (a or b);
    layer4_outputs(384) <= not b;
    layer4_outputs(385) <= not b;
    layer4_outputs(386) <= b;
    layer4_outputs(387) <= a xor b;
    layer4_outputs(388) <= b;
    layer4_outputs(389) <= not (a or b);
    layer4_outputs(390) <= b and not a;
    layer4_outputs(391) <= b;
    layer4_outputs(392) <= not a;
    layer4_outputs(393) <= not a;
    layer4_outputs(394) <= not a;
    layer4_outputs(395) <= a;
    layer4_outputs(396) <= a and b;
    layer4_outputs(397) <= not a;
    layer4_outputs(398) <= not a;
    layer4_outputs(399) <= a;
    layer4_outputs(400) <= not a or b;
    layer4_outputs(401) <= not (a xor b);
    layer4_outputs(402) <= '1';
    layer4_outputs(403) <= b;
    layer4_outputs(404) <= not (a or b);
    layer4_outputs(405) <= a and b;
    layer4_outputs(406) <= not b or a;
    layer4_outputs(407) <= a;
    layer4_outputs(408) <= a xor b;
    layer4_outputs(409) <= not a or b;
    layer4_outputs(410) <= '1';
    layer4_outputs(411) <= not a;
    layer4_outputs(412) <= a and b;
    layer4_outputs(413) <= a;
    layer4_outputs(414) <= b;
    layer4_outputs(415) <= a xor b;
    layer4_outputs(416) <= a and b;
    layer4_outputs(417) <= not b or a;
    layer4_outputs(418) <= not b;
    layer4_outputs(419) <= not (a or b);
    layer4_outputs(420) <= a and b;
    layer4_outputs(421) <= '1';
    layer4_outputs(422) <= '0';
    layer4_outputs(423) <= not (a xor b);
    layer4_outputs(424) <= b;
    layer4_outputs(425) <= not a;
    layer4_outputs(426) <= not (a or b);
    layer4_outputs(427) <= b;
    layer4_outputs(428) <= a;
    layer4_outputs(429) <= b and not a;
    layer4_outputs(430) <= not a or b;
    layer4_outputs(431) <= a;
    layer4_outputs(432) <= not a;
    layer4_outputs(433) <= not (a xor b);
    layer4_outputs(434) <= not (a xor b);
    layer4_outputs(435) <= a xor b;
    layer4_outputs(436) <= a and not b;
    layer4_outputs(437) <= not (a and b);
    layer4_outputs(438) <= not a or b;
    layer4_outputs(439) <= b and not a;
    layer4_outputs(440) <= a and not b;
    layer4_outputs(441) <= a xor b;
    layer4_outputs(442) <= not b;
    layer4_outputs(443) <= b;
    layer4_outputs(444) <= not (a and b);
    layer4_outputs(445) <= b;
    layer4_outputs(446) <= not b or a;
    layer4_outputs(447) <= not b;
    layer4_outputs(448) <= a xor b;
    layer4_outputs(449) <= a and b;
    layer4_outputs(450) <= not b;
    layer4_outputs(451) <= a;
    layer4_outputs(452) <= not b;
    layer4_outputs(453) <= b;
    layer4_outputs(454) <= b;
    layer4_outputs(455) <= not a;
    layer4_outputs(456) <= '1';
    layer4_outputs(457) <= a;
    layer4_outputs(458) <= '0';
    layer4_outputs(459) <= not (a and b);
    layer4_outputs(460) <= b;
    layer4_outputs(461) <= a and b;
    layer4_outputs(462) <= '0';
    layer4_outputs(463) <= a and b;
    layer4_outputs(464) <= not a;
    layer4_outputs(465) <= a;
    layer4_outputs(466) <= not (a or b);
    layer4_outputs(467) <= not a or b;
    layer4_outputs(468) <= b;
    layer4_outputs(469) <= not b;
    layer4_outputs(470) <= '0';
    layer4_outputs(471) <= not (a and b);
    layer4_outputs(472) <= not a or b;
    layer4_outputs(473) <= not a or b;
    layer4_outputs(474) <= a;
    layer4_outputs(475) <= not a;
    layer4_outputs(476) <= not (a xor b);
    layer4_outputs(477) <= not b or a;
    layer4_outputs(478) <= not a;
    layer4_outputs(479) <= a or b;
    layer4_outputs(480) <= a and not b;
    layer4_outputs(481) <= not (a and b);
    layer4_outputs(482) <= b;
    layer4_outputs(483) <= not b;
    layer4_outputs(484) <= a and b;
    layer4_outputs(485) <= not b;
    layer4_outputs(486) <= a and not b;
    layer4_outputs(487) <= not (a and b);
    layer4_outputs(488) <= not b;
    layer4_outputs(489) <= not (a and b);
    layer4_outputs(490) <= not b or a;
    layer4_outputs(491) <= a xor b;
    layer4_outputs(492) <= not b;
    layer4_outputs(493) <= b;
    layer4_outputs(494) <= a or b;
    layer4_outputs(495) <= a or b;
    layer4_outputs(496) <= a and b;
    layer4_outputs(497) <= not (a and b);
    layer4_outputs(498) <= not b;
    layer4_outputs(499) <= not a;
    layer4_outputs(500) <= not (a and b);
    layer4_outputs(501) <= not a or b;
    layer4_outputs(502) <= a;
    layer4_outputs(503) <= not a;
    layer4_outputs(504) <= a xor b;
    layer4_outputs(505) <= a and not b;
    layer4_outputs(506) <= not b;
    layer4_outputs(507) <= a;
    layer4_outputs(508) <= b and not a;
    layer4_outputs(509) <= not a;
    layer4_outputs(510) <= b and not a;
    layer4_outputs(511) <= a xor b;
    layer4_outputs(512) <= not a;
    layer4_outputs(513) <= not (a and b);
    layer4_outputs(514) <= a;
    layer4_outputs(515) <= a;
    layer4_outputs(516) <= a or b;
    layer4_outputs(517) <= not b;
    layer4_outputs(518) <= not b;
    layer4_outputs(519) <= a and b;
    layer4_outputs(520) <= not a;
    layer4_outputs(521) <= '1';
    layer4_outputs(522) <= not (a and b);
    layer4_outputs(523) <= a and not b;
    layer4_outputs(524) <= a xor b;
    layer4_outputs(525) <= not b or a;
    layer4_outputs(526) <= '0';
    layer4_outputs(527) <= a;
    layer4_outputs(528) <= not a or b;
    layer4_outputs(529) <= b;
    layer4_outputs(530) <= a and not b;
    layer4_outputs(531) <= not a;
    layer4_outputs(532) <= a;
    layer4_outputs(533) <= b;
    layer4_outputs(534) <= a and not b;
    layer4_outputs(535) <= b and not a;
    layer4_outputs(536) <= not (a and b);
    layer4_outputs(537) <= not a;
    layer4_outputs(538) <= not a;
    layer4_outputs(539) <= a xor b;
    layer4_outputs(540) <= '0';
    layer4_outputs(541) <= not (a and b);
    layer4_outputs(542) <= b and not a;
    layer4_outputs(543) <= a xor b;
    layer4_outputs(544) <= not a;
    layer4_outputs(545) <= not (a xor b);
    layer4_outputs(546) <= not b;
    layer4_outputs(547) <= not a;
    layer4_outputs(548) <= not a or b;
    layer4_outputs(549) <= not (a or b);
    layer4_outputs(550) <= a;
    layer4_outputs(551) <= not b;
    layer4_outputs(552) <= not a or b;
    layer4_outputs(553) <= b and not a;
    layer4_outputs(554) <= not (a or b);
    layer4_outputs(555) <= a;
    layer4_outputs(556) <= not (a and b);
    layer4_outputs(557) <= not (a or b);
    layer4_outputs(558) <= b and not a;
    layer4_outputs(559) <= a xor b;
    layer4_outputs(560) <= not a or b;
    layer4_outputs(561) <= a xor b;
    layer4_outputs(562) <= not (a xor b);
    layer4_outputs(563) <= not a;
    layer4_outputs(564) <= b;
    layer4_outputs(565) <= '0';
    layer4_outputs(566) <= not b or a;
    layer4_outputs(567) <= a and not b;
    layer4_outputs(568) <= not a or b;
    layer4_outputs(569) <= b;
    layer4_outputs(570) <= not b or a;
    layer4_outputs(571) <= a xor b;
    layer4_outputs(572) <= a xor b;
    layer4_outputs(573) <= b;
    layer4_outputs(574) <= a;
    layer4_outputs(575) <= not (a xor b);
    layer4_outputs(576) <= b;
    layer4_outputs(577) <= a and b;
    layer4_outputs(578) <= a;
    layer4_outputs(579) <= not a or b;
    layer4_outputs(580) <= b;
    layer4_outputs(581) <= a and not b;
    layer4_outputs(582) <= not a;
    layer4_outputs(583) <= a xor b;
    layer4_outputs(584) <= not b or a;
    layer4_outputs(585) <= not a;
    layer4_outputs(586) <= not a;
    layer4_outputs(587) <= a and b;
    layer4_outputs(588) <= not a;
    layer4_outputs(589) <= not a or b;
    layer4_outputs(590) <= not b;
    layer4_outputs(591) <= not b or a;
    layer4_outputs(592) <= b and not a;
    layer4_outputs(593) <= not b;
    layer4_outputs(594) <= not b;
    layer4_outputs(595) <= not b;
    layer4_outputs(596) <= not b;
    layer4_outputs(597) <= not a;
    layer4_outputs(598) <= b and not a;
    layer4_outputs(599) <= a;
    layer4_outputs(600) <= a xor b;
    layer4_outputs(601) <= not (a xor b);
    layer4_outputs(602) <= not (a and b);
    layer4_outputs(603) <= not a;
    layer4_outputs(604) <= not b;
    layer4_outputs(605) <= a or b;
    layer4_outputs(606) <= a or b;
    layer4_outputs(607) <= not a;
    layer4_outputs(608) <= b and not a;
    layer4_outputs(609) <= a and not b;
    layer4_outputs(610) <= not a;
    layer4_outputs(611) <= b;
    layer4_outputs(612) <= not (a xor b);
    layer4_outputs(613) <= '1';
    layer4_outputs(614) <= '0';
    layer4_outputs(615) <= '1';
    layer4_outputs(616) <= not b or a;
    layer4_outputs(617) <= a or b;
    layer4_outputs(618) <= not (a or b);
    layer4_outputs(619) <= not (a xor b);
    layer4_outputs(620) <= '1';
    layer4_outputs(621) <= b;
    layer4_outputs(622) <= a or b;
    layer4_outputs(623) <= a;
    layer4_outputs(624) <= not b;
    layer4_outputs(625) <= a;
    layer4_outputs(626) <= not (a and b);
    layer4_outputs(627) <= not b;
    layer4_outputs(628) <= not a or b;
    layer4_outputs(629) <= a;
    layer4_outputs(630) <= a;
    layer4_outputs(631) <= not (a and b);
    layer4_outputs(632) <= not (a and b);
    layer4_outputs(633) <= '0';
    layer4_outputs(634) <= a;
    layer4_outputs(635) <= b and not a;
    layer4_outputs(636) <= not a;
    layer4_outputs(637) <= not (a or b);
    layer4_outputs(638) <= a xor b;
    layer4_outputs(639) <= not (a and b);
    layer4_outputs(640) <= a or b;
    layer4_outputs(641) <= a xor b;
    layer4_outputs(642) <= not a;
    layer4_outputs(643) <= b and not a;
    layer4_outputs(644) <= not b;
    layer4_outputs(645) <= a and not b;
    layer4_outputs(646) <= not (a or b);
    layer4_outputs(647) <= not a or b;
    layer4_outputs(648) <= not b;
    layer4_outputs(649) <= not a or b;
    layer4_outputs(650) <= '0';
    layer4_outputs(651) <= not (a and b);
    layer4_outputs(652) <= b;
    layer4_outputs(653) <= a xor b;
    layer4_outputs(654) <= '1';
    layer4_outputs(655) <= a;
    layer4_outputs(656) <= a;
    layer4_outputs(657) <= b and not a;
    layer4_outputs(658) <= not (a or b);
    layer4_outputs(659) <= a xor b;
    layer4_outputs(660) <= not a;
    layer4_outputs(661) <= not b;
    layer4_outputs(662) <= not (a or b);
    layer4_outputs(663) <= a;
    layer4_outputs(664) <= a or b;
    layer4_outputs(665) <= a;
    layer4_outputs(666) <= a;
    layer4_outputs(667) <= not b or a;
    layer4_outputs(668) <= not a;
    layer4_outputs(669) <= b;
    layer4_outputs(670) <= b;
    layer4_outputs(671) <= a and b;
    layer4_outputs(672) <= not a or b;
    layer4_outputs(673) <= '0';
    layer4_outputs(674) <= b;
    layer4_outputs(675) <= not a;
    layer4_outputs(676) <= not (a or b);
    layer4_outputs(677) <= a or b;
    layer4_outputs(678) <= '1';
    layer4_outputs(679) <= not a;
    layer4_outputs(680) <= a and not b;
    layer4_outputs(681) <= a xor b;
    layer4_outputs(682) <= not b or a;
    layer4_outputs(683) <= not b;
    layer4_outputs(684) <= not b;
    layer4_outputs(685) <= '0';
    layer4_outputs(686) <= not a or b;
    layer4_outputs(687) <= not (a xor b);
    layer4_outputs(688) <= b;
    layer4_outputs(689) <= '0';
    layer4_outputs(690) <= not (a or b);
    layer4_outputs(691) <= a;
    layer4_outputs(692) <= a and b;
    layer4_outputs(693) <= b;
    layer4_outputs(694) <= a or b;
    layer4_outputs(695) <= not (a or b);
    layer4_outputs(696) <= not (a xor b);
    layer4_outputs(697) <= b;
    layer4_outputs(698) <= not (a and b);
    layer4_outputs(699) <= not a;
    layer4_outputs(700) <= not (a or b);
    layer4_outputs(701) <= a;
    layer4_outputs(702) <= b and not a;
    layer4_outputs(703) <= not (a and b);
    layer4_outputs(704) <= not b;
    layer4_outputs(705) <= not b or a;
    layer4_outputs(706) <= b;
    layer4_outputs(707) <= not (a or b);
    layer4_outputs(708) <= a and b;
    layer4_outputs(709) <= a;
    layer4_outputs(710) <= a and not b;
    layer4_outputs(711) <= a;
    layer4_outputs(712) <= not b;
    layer4_outputs(713) <= not b;
    layer4_outputs(714) <= a or b;
    layer4_outputs(715) <= not a;
    layer4_outputs(716) <= a and b;
    layer4_outputs(717) <= a and b;
    layer4_outputs(718) <= not a;
    layer4_outputs(719) <= a and b;
    layer4_outputs(720) <= a and b;
    layer4_outputs(721) <= not (a and b);
    layer4_outputs(722) <= a;
    layer4_outputs(723) <= a;
    layer4_outputs(724) <= a xor b;
    layer4_outputs(725) <= not a or b;
    layer4_outputs(726) <= b and not a;
    layer4_outputs(727) <= b;
    layer4_outputs(728) <= not b;
    layer4_outputs(729) <= not b;
    layer4_outputs(730) <= not (a and b);
    layer4_outputs(731) <= a;
    layer4_outputs(732) <= not a;
    layer4_outputs(733) <= b and not a;
    layer4_outputs(734) <= a;
    layer4_outputs(735) <= '1';
    layer4_outputs(736) <= not (a or b);
    layer4_outputs(737) <= not (a xor b);
    layer4_outputs(738) <= not (a xor b);
    layer4_outputs(739) <= a and b;
    layer4_outputs(740) <= not b;
    layer4_outputs(741) <= not a;
    layer4_outputs(742) <= not b;
    layer4_outputs(743) <= a;
    layer4_outputs(744) <= not (a xor b);
    layer4_outputs(745) <= not (a or b);
    layer4_outputs(746) <= '1';
    layer4_outputs(747) <= a xor b;
    layer4_outputs(748) <= a;
    layer4_outputs(749) <= a and b;
    layer4_outputs(750) <= a;
    layer4_outputs(751) <= not (a and b);
    layer4_outputs(752) <= not a;
    layer4_outputs(753) <= a;
    layer4_outputs(754) <= not b;
    layer4_outputs(755) <= not a or b;
    layer4_outputs(756) <= not b;
    layer4_outputs(757) <= a and b;
    layer4_outputs(758) <= a;
    layer4_outputs(759) <= b and not a;
    layer4_outputs(760) <= not (a xor b);
    layer4_outputs(761) <= not b;
    layer4_outputs(762) <= b;
    layer4_outputs(763) <= a;
    layer4_outputs(764) <= not (a or b);
    layer4_outputs(765) <= not (a and b);
    layer4_outputs(766) <= not (a or b);
    layer4_outputs(767) <= not (a or b);
    layer4_outputs(768) <= a;
    layer4_outputs(769) <= b and not a;
    layer4_outputs(770) <= b;
    layer4_outputs(771) <= not b;
    layer4_outputs(772) <= b;
    layer4_outputs(773) <= a xor b;
    layer4_outputs(774) <= not a or b;
    layer4_outputs(775) <= b;
    layer4_outputs(776) <= b;
    layer4_outputs(777) <= not b;
    layer4_outputs(778) <= '1';
    layer4_outputs(779) <= a;
    layer4_outputs(780) <= not a or b;
    layer4_outputs(781) <= a and not b;
    layer4_outputs(782) <= not (a and b);
    layer4_outputs(783) <= a;
    layer4_outputs(784) <= a;
    layer4_outputs(785) <= not a;
    layer4_outputs(786) <= not (a and b);
    layer4_outputs(787) <= not a;
    layer4_outputs(788) <= not b;
    layer4_outputs(789) <= a and b;
    layer4_outputs(790) <= a or b;
    layer4_outputs(791) <= not b or a;
    layer4_outputs(792) <= b;
    layer4_outputs(793) <= not b;
    layer4_outputs(794) <= not (a xor b);
    layer4_outputs(795) <= not (a xor b);
    layer4_outputs(796) <= a xor b;
    layer4_outputs(797) <= b and not a;
    layer4_outputs(798) <= b;
    layer4_outputs(799) <= not a;
    layer4_outputs(800) <= not b;
    layer4_outputs(801) <= a;
    layer4_outputs(802) <= a xor b;
    layer4_outputs(803) <= a;
    layer4_outputs(804) <= b;
    layer4_outputs(805) <= a xor b;
    layer4_outputs(806) <= b;
    layer4_outputs(807) <= a;
    layer4_outputs(808) <= not b;
    layer4_outputs(809) <= not a;
    layer4_outputs(810) <= not a or b;
    layer4_outputs(811) <= not a or b;
    layer4_outputs(812) <= b and not a;
    layer4_outputs(813) <= b and not a;
    layer4_outputs(814) <= not a or b;
    layer4_outputs(815) <= b;
    layer4_outputs(816) <= not b;
    layer4_outputs(817) <= not b;
    layer4_outputs(818) <= not a;
    layer4_outputs(819) <= not (a and b);
    layer4_outputs(820) <= not (a xor b);
    layer4_outputs(821) <= a or b;
    layer4_outputs(822) <= b;
    layer4_outputs(823) <= a;
    layer4_outputs(824) <= a xor b;
    layer4_outputs(825) <= not a or b;
    layer4_outputs(826) <= not a;
    layer4_outputs(827) <= not b or a;
    layer4_outputs(828) <= a or b;
    layer4_outputs(829) <= not b or a;
    layer4_outputs(830) <= a;
    layer4_outputs(831) <= b and not a;
    layer4_outputs(832) <= not b;
    layer4_outputs(833) <= not b or a;
    layer4_outputs(834) <= b;
    layer4_outputs(835) <= not (a xor b);
    layer4_outputs(836) <= not (a and b);
    layer4_outputs(837) <= not (a or b);
    layer4_outputs(838) <= a;
    layer4_outputs(839) <= not (a or b);
    layer4_outputs(840) <= a;
    layer4_outputs(841) <= b;
    layer4_outputs(842) <= not a;
    layer4_outputs(843) <= a;
    layer4_outputs(844) <= a;
    layer4_outputs(845) <= not (a or b);
    layer4_outputs(846) <= a and not b;
    layer4_outputs(847) <= not a;
    layer4_outputs(848) <= not a or b;
    layer4_outputs(849) <= not a or b;
    layer4_outputs(850) <= not a;
    layer4_outputs(851) <= not b or a;
    layer4_outputs(852) <= not b;
    layer4_outputs(853) <= a;
    layer4_outputs(854) <= a and b;
    layer4_outputs(855) <= not a;
    layer4_outputs(856) <= not a;
    layer4_outputs(857) <= a and not b;
    layer4_outputs(858) <= a xor b;
    layer4_outputs(859) <= not (a or b);
    layer4_outputs(860) <= not b;
    layer4_outputs(861) <= not b;
    layer4_outputs(862) <= a and not b;
    layer4_outputs(863) <= not (a and b);
    layer4_outputs(864) <= not b;
    layer4_outputs(865) <= b;
    layer4_outputs(866) <= not (a xor b);
    layer4_outputs(867) <= a;
    layer4_outputs(868) <= a;
    layer4_outputs(869) <= not a;
    layer4_outputs(870) <= b;
    layer4_outputs(871) <= not (a or b);
    layer4_outputs(872) <= not (a xor b);
    layer4_outputs(873) <= not b;
    layer4_outputs(874) <= not a;
    layer4_outputs(875) <= a;
    layer4_outputs(876) <= b;
    layer4_outputs(877) <= not a or b;
    layer4_outputs(878) <= b and not a;
    layer4_outputs(879) <= b;
    layer4_outputs(880) <= not (a or b);
    layer4_outputs(881) <= not (a or b);
    layer4_outputs(882) <= a xor b;
    layer4_outputs(883) <= a xor b;
    layer4_outputs(884) <= not (a or b);
    layer4_outputs(885) <= not b or a;
    layer4_outputs(886) <= '0';
    layer4_outputs(887) <= not b or a;
    layer4_outputs(888) <= a and b;
    layer4_outputs(889) <= a;
    layer4_outputs(890) <= not (a xor b);
    layer4_outputs(891) <= b and not a;
    layer4_outputs(892) <= not a;
    layer4_outputs(893) <= not (a or b);
    layer4_outputs(894) <= not b;
    layer4_outputs(895) <= '1';
    layer4_outputs(896) <= not b;
    layer4_outputs(897) <= not a;
    layer4_outputs(898) <= b;
    layer4_outputs(899) <= a or b;
    layer4_outputs(900) <= not (a and b);
    layer4_outputs(901) <= a;
    layer4_outputs(902) <= not b or a;
    layer4_outputs(903) <= a;
    layer4_outputs(904) <= a;
    layer4_outputs(905) <= not a or b;
    layer4_outputs(906) <= not a or b;
    layer4_outputs(907) <= '0';
    layer4_outputs(908) <= a xor b;
    layer4_outputs(909) <= not a or b;
    layer4_outputs(910) <= a xor b;
    layer4_outputs(911) <= b and not a;
    layer4_outputs(912) <= a;
    layer4_outputs(913) <= a xor b;
    layer4_outputs(914) <= not a;
    layer4_outputs(915) <= a and not b;
    layer4_outputs(916) <= not b;
    layer4_outputs(917) <= not (a or b);
    layer4_outputs(918) <= not a;
    layer4_outputs(919) <= '1';
    layer4_outputs(920) <= not a or b;
    layer4_outputs(921) <= not (a xor b);
    layer4_outputs(922) <= not b or a;
    layer4_outputs(923) <= a and not b;
    layer4_outputs(924) <= a and b;
    layer4_outputs(925) <= a or b;
    layer4_outputs(926) <= not b or a;
    layer4_outputs(927) <= b and not a;
    layer4_outputs(928) <= a or b;
    layer4_outputs(929) <= a and not b;
    layer4_outputs(930) <= a and b;
    layer4_outputs(931) <= not b;
    layer4_outputs(932) <= not (a and b);
    layer4_outputs(933) <= a and b;
    layer4_outputs(934) <= a and b;
    layer4_outputs(935) <= not (a xor b);
    layer4_outputs(936) <= b;
    layer4_outputs(937) <= a and b;
    layer4_outputs(938) <= not a;
    layer4_outputs(939) <= a xor b;
    layer4_outputs(940) <= b;
    layer4_outputs(941) <= not (a xor b);
    layer4_outputs(942) <= not (a and b);
    layer4_outputs(943) <= not a;
    layer4_outputs(944) <= not (a and b);
    layer4_outputs(945) <= not b;
    layer4_outputs(946) <= a and b;
    layer4_outputs(947) <= '1';
    layer4_outputs(948) <= b;
    layer4_outputs(949) <= not a or b;
    layer4_outputs(950) <= a or b;
    layer4_outputs(951) <= a and not b;
    layer4_outputs(952) <= a xor b;
    layer4_outputs(953) <= not b;
    layer4_outputs(954) <= a and b;
    layer4_outputs(955) <= not a;
    layer4_outputs(956) <= not (a or b);
    layer4_outputs(957) <= not a;
    layer4_outputs(958) <= not (a and b);
    layer4_outputs(959) <= not (a or b);
    layer4_outputs(960) <= a and b;
    layer4_outputs(961) <= not b or a;
    layer4_outputs(962) <= not b;
    layer4_outputs(963) <= a or b;
    layer4_outputs(964) <= not b;
    layer4_outputs(965) <= a;
    layer4_outputs(966) <= not (a or b);
    layer4_outputs(967) <= a and not b;
    layer4_outputs(968) <= not (a or b);
    layer4_outputs(969) <= '0';
    layer4_outputs(970) <= not a or b;
    layer4_outputs(971) <= '0';
    layer4_outputs(972) <= not b;
    layer4_outputs(973) <= b and not a;
    layer4_outputs(974) <= b and not a;
    layer4_outputs(975) <= b;
    layer4_outputs(976) <= not a or b;
    layer4_outputs(977) <= '0';
    layer4_outputs(978) <= not a;
    layer4_outputs(979) <= b;
    layer4_outputs(980) <= not a;
    layer4_outputs(981) <= b;
    layer4_outputs(982) <= b;
    layer4_outputs(983) <= a xor b;
    layer4_outputs(984) <= not a or b;
    layer4_outputs(985) <= a;
    layer4_outputs(986) <= not b;
    layer4_outputs(987) <= not a or b;
    layer4_outputs(988) <= a and b;
    layer4_outputs(989) <= not (a and b);
    layer4_outputs(990) <= not a;
    layer4_outputs(991) <= b;
    layer4_outputs(992) <= not b;
    layer4_outputs(993) <= b;
    layer4_outputs(994) <= a and not b;
    layer4_outputs(995) <= not b or a;
    layer4_outputs(996) <= not a;
    layer4_outputs(997) <= not b;
    layer4_outputs(998) <= a xor b;
    layer4_outputs(999) <= a;
    layer4_outputs(1000) <= a;
    layer4_outputs(1001) <= a;
    layer4_outputs(1002) <= b;
    layer4_outputs(1003) <= not b;
    layer4_outputs(1004) <= not a or b;
    layer4_outputs(1005) <= not a;
    layer4_outputs(1006) <= b;
    layer4_outputs(1007) <= not (a and b);
    layer4_outputs(1008) <= a xor b;
    layer4_outputs(1009) <= a and not b;
    layer4_outputs(1010) <= not a;
    layer4_outputs(1011) <= a;
    layer4_outputs(1012) <= not a;
    layer4_outputs(1013) <= not (a xor b);
    layer4_outputs(1014) <= a and not b;
    layer4_outputs(1015) <= b and not a;
    layer4_outputs(1016) <= b;
    layer4_outputs(1017) <= b;
    layer4_outputs(1018) <= not a or b;
    layer4_outputs(1019) <= b and not a;
    layer4_outputs(1020) <= not b;
    layer4_outputs(1021) <= not a;
    layer4_outputs(1022) <= a;
    layer4_outputs(1023) <= not b;
    layer4_outputs(1024) <= not a or b;
    layer4_outputs(1025) <= b;
    layer4_outputs(1026) <= not a;
    layer4_outputs(1027) <= b;
    layer4_outputs(1028) <= a and b;
    layer4_outputs(1029) <= not (a xor b);
    layer4_outputs(1030) <= not b;
    layer4_outputs(1031) <= a and b;
    layer4_outputs(1032) <= b;
    layer4_outputs(1033) <= a or b;
    layer4_outputs(1034) <= not (a or b);
    layer4_outputs(1035) <= '1';
    layer4_outputs(1036) <= a;
    layer4_outputs(1037) <= a;
    layer4_outputs(1038) <= a;
    layer4_outputs(1039) <= not b;
    layer4_outputs(1040) <= b and not a;
    layer4_outputs(1041) <= not b;
    layer4_outputs(1042) <= b;
    layer4_outputs(1043) <= a xor b;
    layer4_outputs(1044) <= not b;
    layer4_outputs(1045) <= not a or b;
    layer4_outputs(1046) <= a xor b;
    layer4_outputs(1047) <= not b or a;
    layer4_outputs(1048) <= a;
    layer4_outputs(1049) <= b and not a;
    layer4_outputs(1050) <= not (a and b);
    layer4_outputs(1051) <= not b;
    layer4_outputs(1052) <= a;
    layer4_outputs(1053) <= b;
    layer4_outputs(1054) <= a and not b;
    layer4_outputs(1055) <= not b;
    layer4_outputs(1056) <= a or b;
    layer4_outputs(1057) <= a;
    layer4_outputs(1058) <= b;
    layer4_outputs(1059) <= b and not a;
    layer4_outputs(1060) <= not b;
    layer4_outputs(1061) <= not b or a;
    layer4_outputs(1062) <= not (a or b);
    layer4_outputs(1063) <= not b;
    layer4_outputs(1064) <= not a or b;
    layer4_outputs(1065) <= not a or b;
    layer4_outputs(1066) <= not a;
    layer4_outputs(1067) <= not a;
    layer4_outputs(1068) <= not b;
    layer4_outputs(1069) <= a;
    layer4_outputs(1070) <= not b;
    layer4_outputs(1071) <= a;
    layer4_outputs(1072) <= '0';
    layer4_outputs(1073) <= not (a and b);
    layer4_outputs(1074) <= a and b;
    layer4_outputs(1075) <= a;
    layer4_outputs(1076) <= not (a or b);
    layer4_outputs(1077) <= a xor b;
    layer4_outputs(1078) <= not b or a;
    layer4_outputs(1079) <= not (a and b);
    layer4_outputs(1080) <= not (a and b);
    layer4_outputs(1081) <= not b;
    layer4_outputs(1082) <= not a or b;
    layer4_outputs(1083) <= a;
    layer4_outputs(1084) <= b;
    layer4_outputs(1085) <= not (a and b);
    layer4_outputs(1086) <= not b;
    layer4_outputs(1087) <= not a;
    layer4_outputs(1088) <= a or b;
    layer4_outputs(1089) <= a and not b;
    layer4_outputs(1090) <= not a;
    layer4_outputs(1091) <= b and not a;
    layer4_outputs(1092) <= not (a or b);
    layer4_outputs(1093) <= not b or a;
    layer4_outputs(1094) <= not b or a;
    layer4_outputs(1095) <= not b;
    layer4_outputs(1096) <= a or b;
    layer4_outputs(1097) <= a and not b;
    layer4_outputs(1098) <= not a;
    layer4_outputs(1099) <= a and not b;
    layer4_outputs(1100) <= b;
    layer4_outputs(1101) <= a;
    layer4_outputs(1102) <= '1';
    layer4_outputs(1103) <= not b;
    layer4_outputs(1104) <= not (a and b);
    layer4_outputs(1105) <= '0';
    layer4_outputs(1106) <= not a or b;
    layer4_outputs(1107) <= a or b;
    layer4_outputs(1108) <= a;
    layer4_outputs(1109) <= a;
    layer4_outputs(1110) <= not a;
    layer4_outputs(1111) <= a and b;
    layer4_outputs(1112) <= not (a and b);
    layer4_outputs(1113) <= a xor b;
    layer4_outputs(1114) <= a;
    layer4_outputs(1115) <= '1';
    layer4_outputs(1116) <= a xor b;
    layer4_outputs(1117) <= b;
    layer4_outputs(1118) <= a and not b;
    layer4_outputs(1119) <= a or b;
    layer4_outputs(1120) <= not b;
    layer4_outputs(1121) <= a and b;
    layer4_outputs(1122) <= a;
    layer4_outputs(1123) <= a;
    layer4_outputs(1124) <= not b;
    layer4_outputs(1125) <= a or b;
    layer4_outputs(1126) <= not (a or b);
    layer4_outputs(1127) <= a and not b;
    layer4_outputs(1128) <= b;
    layer4_outputs(1129) <= not (a or b);
    layer4_outputs(1130) <= not a;
    layer4_outputs(1131) <= b and not a;
    layer4_outputs(1132) <= b;
    layer4_outputs(1133) <= a xor b;
    layer4_outputs(1134) <= not (a or b);
    layer4_outputs(1135) <= not b or a;
    layer4_outputs(1136) <= not b;
    layer4_outputs(1137) <= not (a and b);
    layer4_outputs(1138) <= not b;
    layer4_outputs(1139) <= not a or b;
    layer4_outputs(1140) <= b;
    layer4_outputs(1141) <= a;
    layer4_outputs(1142) <= not (a and b);
    layer4_outputs(1143) <= not a;
    layer4_outputs(1144) <= a xor b;
    layer4_outputs(1145) <= b and not a;
    layer4_outputs(1146) <= not (a and b);
    layer4_outputs(1147) <= not a;
    layer4_outputs(1148) <= not a;
    layer4_outputs(1149) <= not a or b;
    layer4_outputs(1150) <= not b;
    layer4_outputs(1151) <= not b or a;
    layer4_outputs(1152) <= not a;
    layer4_outputs(1153) <= not b;
    layer4_outputs(1154) <= a;
    layer4_outputs(1155) <= b;
    layer4_outputs(1156) <= b;
    layer4_outputs(1157) <= not b;
    layer4_outputs(1158) <= a and b;
    layer4_outputs(1159) <= not a or b;
    layer4_outputs(1160) <= a and not b;
    layer4_outputs(1161) <= not a;
    layer4_outputs(1162) <= not a;
    layer4_outputs(1163) <= b;
    layer4_outputs(1164) <= '0';
    layer4_outputs(1165) <= a;
    layer4_outputs(1166) <= not (a xor b);
    layer4_outputs(1167) <= a and not b;
    layer4_outputs(1168) <= a;
    layer4_outputs(1169) <= not a;
    layer4_outputs(1170) <= not a;
    layer4_outputs(1171) <= not a;
    layer4_outputs(1172) <= b;
    layer4_outputs(1173) <= '0';
    layer4_outputs(1174) <= not b;
    layer4_outputs(1175) <= a;
    layer4_outputs(1176) <= not (a xor b);
    layer4_outputs(1177) <= not a;
    layer4_outputs(1178) <= '0';
    layer4_outputs(1179) <= not (a or b);
    layer4_outputs(1180) <= not (a xor b);
    layer4_outputs(1181) <= a;
    layer4_outputs(1182) <= '1';
    layer4_outputs(1183) <= b;
    layer4_outputs(1184) <= not (a or b);
    layer4_outputs(1185) <= a;
    layer4_outputs(1186) <= b and not a;
    layer4_outputs(1187) <= not a;
    layer4_outputs(1188) <= a and not b;
    layer4_outputs(1189) <= a;
    layer4_outputs(1190) <= not a or b;
    layer4_outputs(1191) <= not (a and b);
    layer4_outputs(1192) <= a and not b;
    layer4_outputs(1193) <= a and not b;
    layer4_outputs(1194) <= a;
    layer4_outputs(1195) <= not b;
    layer4_outputs(1196) <= a and not b;
    layer4_outputs(1197) <= not b or a;
    layer4_outputs(1198) <= a and b;
    layer4_outputs(1199) <= a and b;
    layer4_outputs(1200) <= not (a or b);
    layer4_outputs(1201) <= b;
    layer4_outputs(1202) <= a xor b;
    layer4_outputs(1203) <= b;
    layer4_outputs(1204) <= not b or a;
    layer4_outputs(1205) <= not b or a;
    layer4_outputs(1206) <= not (a and b);
    layer4_outputs(1207) <= not b or a;
    layer4_outputs(1208) <= not a or b;
    layer4_outputs(1209) <= b;
    layer4_outputs(1210) <= b;
    layer4_outputs(1211) <= not b;
    layer4_outputs(1212) <= a and not b;
    layer4_outputs(1213) <= not a or b;
    layer4_outputs(1214) <= a;
    layer4_outputs(1215) <= b;
    layer4_outputs(1216) <= a and b;
    layer4_outputs(1217) <= a and not b;
    layer4_outputs(1218) <= a;
    layer4_outputs(1219) <= a xor b;
    layer4_outputs(1220) <= not (a and b);
    layer4_outputs(1221) <= a;
    layer4_outputs(1222) <= '0';
    layer4_outputs(1223) <= not (a or b);
    layer4_outputs(1224) <= not a;
    layer4_outputs(1225) <= not (a and b);
    layer4_outputs(1226) <= not a;
    layer4_outputs(1227) <= a;
    layer4_outputs(1228) <= a;
    layer4_outputs(1229) <= a xor b;
    layer4_outputs(1230) <= a;
    layer4_outputs(1231) <= not (a xor b);
    layer4_outputs(1232) <= a;
    layer4_outputs(1233) <= not (a xor b);
    layer4_outputs(1234) <= a and not b;
    layer4_outputs(1235) <= a and b;
    layer4_outputs(1236) <= b;
    layer4_outputs(1237) <= b and not a;
    layer4_outputs(1238) <= not a;
    layer4_outputs(1239) <= a or b;
    layer4_outputs(1240) <= not b;
    layer4_outputs(1241) <= not a;
    layer4_outputs(1242) <= a and b;
    layer4_outputs(1243) <= not (a and b);
    layer4_outputs(1244) <= not a;
    layer4_outputs(1245) <= a;
    layer4_outputs(1246) <= '1';
    layer4_outputs(1247) <= a;
    layer4_outputs(1248) <= a or b;
    layer4_outputs(1249) <= not (a or b);
    layer4_outputs(1250) <= not a;
    layer4_outputs(1251) <= a xor b;
    layer4_outputs(1252) <= not a;
    layer4_outputs(1253) <= not (a or b);
    layer4_outputs(1254) <= a xor b;
    layer4_outputs(1255) <= a and b;
    layer4_outputs(1256) <= a and b;
    layer4_outputs(1257) <= not (a or b);
    layer4_outputs(1258) <= not (a and b);
    layer4_outputs(1259) <= not a;
    layer4_outputs(1260) <= b;
    layer4_outputs(1261) <= '0';
    layer4_outputs(1262) <= not (a and b);
    layer4_outputs(1263) <= not (a or b);
    layer4_outputs(1264) <= b;
    layer4_outputs(1265) <= '0';
    layer4_outputs(1266) <= not b or a;
    layer4_outputs(1267) <= b and not a;
    layer4_outputs(1268) <= a;
    layer4_outputs(1269) <= not (a and b);
    layer4_outputs(1270) <= not b;
    layer4_outputs(1271) <= not b;
    layer4_outputs(1272) <= not b;
    layer4_outputs(1273) <= not a or b;
    layer4_outputs(1274) <= a;
    layer4_outputs(1275) <= b and not a;
    layer4_outputs(1276) <= a and b;
    layer4_outputs(1277) <= a;
    layer4_outputs(1278) <= not (a and b);
    layer4_outputs(1279) <= not (a and b);
    layer4_outputs(1280) <= not (a and b);
    layer4_outputs(1281) <= not (a or b);
    layer4_outputs(1282) <= a;
    layer4_outputs(1283) <= b;
    layer4_outputs(1284) <= not (a or b);
    layer4_outputs(1285) <= a and b;
    layer4_outputs(1286) <= not b;
    layer4_outputs(1287) <= '1';
    layer4_outputs(1288) <= a or b;
    layer4_outputs(1289) <= a xor b;
    layer4_outputs(1290) <= a xor b;
    layer4_outputs(1291) <= a;
    layer4_outputs(1292) <= not b;
    layer4_outputs(1293) <= a or b;
    layer4_outputs(1294) <= a and not b;
    layer4_outputs(1295) <= a and not b;
    layer4_outputs(1296) <= b;
    layer4_outputs(1297) <= a and not b;
    layer4_outputs(1298) <= not (a or b);
    layer4_outputs(1299) <= a xor b;
    layer4_outputs(1300) <= b;
    layer4_outputs(1301) <= b and not a;
    layer4_outputs(1302) <= not b or a;
    layer4_outputs(1303) <= b;
    layer4_outputs(1304) <= not a;
    layer4_outputs(1305) <= b;
    layer4_outputs(1306) <= a;
    layer4_outputs(1307) <= not a or b;
    layer4_outputs(1308) <= b;
    layer4_outputs(1309) <= not (a or b);
    layer4_outputs(1310) <= not a;
    layer4_outputs(1311) <= '1';
    layer4_outputs(1312) <= b;
    layer4_outputs(1313) <= not b;
    layer4_outputs(1314) <= a and not b;
    layer4_outputs(1315) <= not b or a;
    layer4_outputs(1316) <= not a;
    layer4_outputs(1317) <= a and not b;
    layer4_outputs(1318) <= a;
    layer4_outputs(1319) <= a;
    layer4_outputs(1320) <= a and not b;
    layer4_outputs(1321) <= not b;
    layer4_outputs(1322) <= not a;
    layer4_outputs(1323) <= not a or b;
    layer4_outputs(1324) <= not a;
    layer4_outputs(1325) <= a and not b;
    layer4_outputs(1326) <= b and not a;
    layer4_outputs(1327) <= a or b;
    layer4_outputs(1328) <= a and b;
    layer4_outputs(1329) <= a or b;
    layer4_outputs(1330) <= not b;
    layer4_outputs(1331) <= not a or b;
    layer4_outputs(1332) <= '1';
    layer4_outputs(1333) <= a and b;
    layer4_outputs(1334) <= not b;
    layer4_outputs(1335) <= not a;
    layer4_outputs(1336) <= a xor b;
    layer4_outputs(1337) <= a or b;
    layer4_outputs(1338) <= not (a or b);
    layer4_outputs(1339) <= a;
    layer4_outputs(1340) <= not a or b;
    layer4_outputs(1341) <= b;
    layer4_outputs(1342) <= a or b;
    layer4_outputs(1343) <= a and not b;
    layer4_outputs(1344) <= not b or a;
    layer4_outputs(1345) <= not (a xor b);
    layer4_outputs(1346) <= b and not a;
    layer4_outputs(1347) <= not b;
    layer4_outputs(1348) <= not (a xor b);
    layer4_outputs(1349) <= a;
    layer4_outputs(1350) <= not b;
    layer4_outputs(1351) <= a and b;
    layer4_outputs(1352) <= not a;
    layer4_outputs(1353) <= not (a or b);
    layer4_outputs(1354) <= a or b;
    layer4_outputs(1355) <= b;
    layer4_outputs(1356) <= a xor b;
    layer4_outputs(1357) <= not (a or b);
    layer4_outputs(1358) <= a or b;
    layer4_outputs(1359) <= not a;
    layer4_outputs(1360) <= not b;
    layer4_outputs(1361) <= not (a xor b);
    layer4_outputs(1362) <= b;
    layer4_outputs(1363) <= a;
    layer4_outputs(1364) <= not a or b;
    layer4_outputs(1365) <= not b or a;
    layer4_outputs(1366) <= b;
    layer4_outputs(1367) <= a and not b;
    layer4_outputs(1368) <= b;
    layer4_outputs(1369) <= a;
    layer4_outputs(1370) <= a;
    layer4_outputs(1371) <= not (a and b);
    layer4_outputs(1372) <= a and not b;
    layer4_outputs(1373) <= '1';
    layer4_outputs(1374) <= a or b;
    layer4_outputs(1375) <= not b;
    layer4_outputs(1376) <= not (a xor b);
    layer4_outputs(1377) <= '0';
    layer4_outputs(1378) <= a or b;
    layer4_outputs(1379) <= a xor b;
    layer4_outputs(1380) <= a;
    layer4_outputs(1381) <= a and b;
    layer4_outputs(1382) <= b;
    layer4_outputs(1383) <= not a;
    layer4_outputs(1384) <= a;
    layer4_outputs(1385) <= a and b;
    layer4_outputs(1386) <= not (a or b);
    layer4_outputs(1387) <= b;
    layer4_outputs(1388) <= not a;
    layer4_outputs(1389) <= a or b;
    layer4_outputs(1390) <= not b or a;
    layer4_outputs(1391) <= a;
    layer4_outputs(1392) <= not a;
    layer4_outputs(1393) <= not b;
    layer4_outputs(1394) <= not (a and b);
    layer4_outputs(1395) <= a and not b;
    layer4_outputs(1396) <= a or b;
    layer4_outputs(1397) <= not (a or b);
    layer4_outputs(1398) <= b and not a;
    layer4_outputs(1399) <= not b;
    layer4_outputs(1400) <= a xor b;
    layer4_outputs(1401) <= a xor b;
    layer4_outputs(1402) <= a xor b;
    layer4_outputs(1403) <= a;
    layer4_outputs(1404) <= b and not a;
    layer4_outputs(1405) <= not b or a;
    layer4_outputs(1406) <= b;
    layer4_outputs(1407) <= not (a xor b);
    layer4_outputs(1408) <= a and b;
    layer4_outputs(1409) <= not (a or b);
    layer4_outputs(1410) <= b and not a;
    layer4_outputs(1411) <= a and b;
    layer4_outputs(1412) <= '1';
    layer4_outputs(1413) <= a;
    layer4_outputs(1414) <= not a;
    layer4_outputs(1415) <= a and not b;
    layer4_outputs(1416) <= not a;
    layer4_outputs(1417) <= not (a and b);
    layer4_outputs(1418) <= not (a and b);
    layer4_outputs(1419) <= a and b;
    layer4_outputs(1420) <= b and not a;
    layer4_outputs(1421) <= not a;
    layer4_outputs(1422) <= not a or b;
    layer4_outputs(1423) <= '1';
    layer4_outputs(1424) <= '1';
    layer4_outputs(1425) <= not (a or b);
    layer4_outputs(1426) <= not b;
    layer4_outputs(1427) <= '0';
    layer4_outputs(1428) <= b;
    layer4_outputs(1429) <= not (a and b);
    layer4_outputs(1430) <= a xor b;
    layer4_outputs(1431) <= a and not b;
    layer4_outputs(1432) <= not a;
    layer4_outputs(1433) <= a;
    layer4_outputs(1434) <= not a;
    layer4_outputs(1435) <= not b;
    layer4_outputs(1436) <= not (a and b);
    layer4_outputs(1437) <= b;
    layer4_outputs(1438) <= b and not a;
    layer4_outputs(1439) <= b;
    layer4_outputs(1440) <= b;
    layer4_outputs(1441) <= not a or b;
    layer4_outputs(1442) <= a and not b;
    layer4_outputs(1443) <= b;
    layer4_outputs(1444) <= b;
    layer4_outputs(1445) <= not a;
    layer4_outputs(1446) <= a and not b;
    layer4_outputs(1447) <= not a;
    layer4_outputs(1448) <= not b or a;
    layer4_outputs(1449) <= b;
    layer4_outputs(1450) <= b;
    layer4_outputs(1451) <= not (a xor b);
    layer4_outputs(1452) <= not a;
    layer4_outputs(1453) <= not b;
    layer4_outputs(1454) <= not a;
    layer4_outputs(1455) <= a and b;
    layer4_outputs(1456) <= '1';
    layer4_outputs(1457) <= a;
    layer4_outputs(1458) <= not (a or b);
    layer4_outputs(1459) <= a;
    layer4_outputs(1460) <= not a;
    layer4_outputs(1461) <= not (a and b);
    layer4_outputs(1462) <= a and not b;
    layer4_outputs(1463) <= '1';
    layer4_outputs(1464) <= not b or a;
    layer4_outputs(1465) <= b;
    layer4_outputs(1466) <= a or b;
    layer4_outputs(1467) <= not (a and b);
    layer4_outputs(1468) <= a xor b;
    layer4_outputs(1469) <= not b or a;
    layer4_outputs(1470) <= b and not a;
    layer4_outputs(1471) <= not b;
    layer4_outputs(1472) <= '0';
    layer4_outputs(1473) <= not (a or b);
    layer4_outputs(1474) <= not b or a;
    layer4_outputs(1475) <= not b;
    layer4_outputs(1476) <= not a;
    layer4_outputs(1477) <= a;
    layer4_outputs(1478) <= b;
    layer4_outputs(1479) <= not a;
    layer4_outputs(1480) <= a and not b;
    layer4_outputs(1481) <= a and not b;
    layer4_outputs(1482) <= b;
    layer4_outputs(1483) <= not a;
    layer4_outputs(1484) <= b and not a;
    layer4_outputs(1485) <= not a;
    layer4_outputs(1486) <= not a;
    layer4_outputs(1487) <= not b;
    layer4_outputs(1488) <= a;
    layer4_outputs(1489) <= not b;
    layer4_outputs(1490) <= b;
    layer4_outputs(1491) <= not a;
    layer4_outputs(1492) <= a and not b;
    layer4_outputs(1493) <= not (a xor b);
    layer4_outputs(1494) <= not (a and b);
    layer4_outputs(1495) <= a;
    layer4_outputs(1496) <= not (a xor b);
    layer4_outputs(1497) <= '0';
    layer4_outputs(1498) <= not b;
    layer4_outputs(1499) <= not b or a;
    layer4_outputs(1500) <= a or b;
    layer4_outputs(1501) <= a xor b;
    layer4_outputs(1502) <= '1';
    layer4_outputs(1503) <= b;
    layer4_outputs(1504) <= not (a or b);
    layer4_outputs(1505) <= not (a or b);
    layer4_outputs(1506) <= not a;
    layer4_outputs(1507) <= a and b;
    layer4_outputs(1508) <= a;
    layer4_outputs(1509) <= a and b;
    layer4_outputs(1510) <= a;
    layer4_outputs(1511) <= a xor b;
    layer4_outputs(1512) <= not a;
    layer4_outputs(1513) <= a or b;
    layer4_outputs(1514) <= not b;
    layer4_outputs(1515) <= not b;
    layer4_outputs(1516) <= a and b;
    layer4_outputs(1517) <= a or b;
    layer4_outputs(1518) <= '1';
    layer4_outputs(1519) <= a;
    layer4_outputs(1520) <= a and not b;
    layer4_outputs(1521) <= a;
    layer4_outputs(1522) <= '1';
    layer4_outputs(1523) <= a or b;
    layer4_outputs(1524) <= a and b;
    layer4_outputs(1525) <= a xor b;
    layer4_outputs(1526) <= not b;
    layer4_outputs(1527) <= a and not b;
    layer4_outputs(1528) <= a or b;
    layer4_outputs(1529) <= not b;
    layer4_outputs(1530) <= not a;
    layer4_outputs(1531) <= '1';
    layer4_outputs(1532) <= '1';
    layer4_outputs(1533) <= not a or b;
    layer4_outputs(1534) <= b;
    layer4_outputs(1535) <= a or b;
    layer4_outputs(1536) <= not (a xor b);
    layer4_outputs(1537) <= a and not b;
    layer4_outputs(1538) <= b;
    layer4_outputs(1539) <= not b;
    layer4_outputs(1540) <= a xor b;
    layer4_outputs(1541) <= a or b;
    layer4_outputs(1542) <= b and not a;
    layer4_outputs(1543) <= a and not b;
    layer4_outputs(1544) <= a;
    layer4_outputs(1545) <= a and b;
    layer4_outputs(1546) <= a and b;
    layer4_outputs(1547) <= not b;
    layer4_outputs(1548) <= b and not a;
    layer4_outputs(1549) <= '0';
    layer4_outputs(1550) <= '0';
    layer4_outputs(1551) <= not (a or b);
    layer4_outputs(1552) <= '1';
    layer4_outputs(1553) <= a;
    layer4_outputs(1554) <= b;
    layer4_outputs(1555) <= not a;
    layer4_outputs(1556) <= not b;
    layer4_outputs(1557) <= not b or a;
    layer4_outputs(1558) <= not b;
    layer4_outputs(1559) <= not a or b;
    layer4_outputs(1560) <= not a;
    layer4_outputs(1561) <= not (a and b);
    layer4_outputs(1562) <= not a;
    layer4_outputs(1563) <= a and not b;
    layer4_outputs(1564) <= not (a or b);
    layer4_outputs(1565) <= not a;
    layer4_outputs(1566) <= '0';
    layer4_outputs(1567) <= not (a or b);
    layer4_outputs(1568) <= not b;
    layer4_outputs(1569) <= not b;
    layer4_outputs(1570) <= a;
    layer4_outputs(1571) <= a and b;
    layer4_outputs(1572) <= not a or b;
    layer4_outputs(1573) <= a;
    layer4_outputs(1574) <= not a or b;
    layer4_outputs(1575) <= '0';
    layer4_outputs(1576) <= not a or b;
    layer4_outputs(1577) <= not a;
    layer4_outputs(1578) <= a;
    layer4_outputs(1579) <= not (a xor b);
    layer4_outputs(1580) <= a or b;
    layer4_outputs(1581) <= not a;
    layer4_outputs(1582) <= b;
    layer4_outputs(1583) <= not b or a;
    layer4_outputs(1584) <= not a;
    layer4_outputs(1585) <= b and not a;
    layer4_outputs(1586) <= not b or a;
    layer4_outputs(1587) <= a and not b;
    layer4_outputs(1588) <= not (a xor b);
    layer4_outputs(1589) <= '1';
    layer4_outputs(1590) <= a;
    layer4_outputs(1591) <= not a;
    layer4_outputs(1592) <= a and b;
    layer4_outputs(1593) <= not a;
    layer4_outputs(1594) <= not a;
    layer4_outputs(1595) <= b;
    layer4_outputs(1596) <= not a or b;
    layer4_outputs(1597) <= '1';
    layer4_outputs(1598) <= not (a xor b);
    layer4_outputs(1599) <= not a or b;
    layer4_outputs(1600) <= not b;
    layer4_outputs(1601) <= a and b;
    layer4_outputs(1602) <= a;
    layer4_outputs(1603) <= not b;
    layer4_outputs(1604) <= not (a or b);
    layer4_outputs(1605) <= not (a and b);
    layer4_outputs(1606) <= '1';
    layer4_outputs(1607) <= '0';
    layer4_outputs(1608) <= b;
    layer4_outputs(1609) <= not a;
    layer4_outputs(1610) <= b;
    layer4_outputs(1611) <= not a;
    layer4_outputs(1612) <= b and not a;
    layer4_outputs(1613) <= not (a and b);
    layer4_outputs(1614) <= not a;
    layer4_outputs(1615) <= not b;
    layer4_outputs(1616) <= b;
    layer4_outputs(1617) <= not a;
    layer4_outputs(1618) <= a;
    layer4_outputs(1619) <= not a;
    layer4_outputs(1620) <= not a;
    layer4_outputs(1621) <= a;
    layer4_outputs(1622) <= b;
    layer4_outputs(1623) <= not (a xor b);
    layer4_outputs(1624) <= b;
    layer4_outputs(1625) <= a;
    layer4_outputs(1626) <= a or b;
    layer4_outputs(1627) <= not (a and b);
    layer4_outputs(1628) <= not a;
    layer4_outputs(1629) <= a and not b;
    layer4_outputs(1630) <= not b;
    layer4_outputs(1631) <= not a;
    layer4_outputs(1632) <= b;
    layer4_outputs(1633) <= not b or a;
    layer4_outputs(1634) <= b;
    layer4_outputs(1635) <= '0';
    layer4_outputs(1636) <= not b;
    layer4_outputs(1637) <= not b or a;
    layer4_outputs(1638) <= not b;
    layer4_outputs(1639) <= a;
    layer4_outputs(1640) <= a or b;
    layer4_outputs(1641) <= b;
    layer4_outputs(1642) <= not a or b;
    layer4_outputs(1643) <= not b or a;
    layer4_outputs(1644) <= a or b;
    layer4_outputs(1645) <= not (a and b);
    layer4_outputs(1646) <= a xor b;
    layer4_outputs(1647) <= b;
    layer4_outputs(1648) <= not (a and b);
    layer4_outputs(1649) <= not a;
    layer4_outputs(1650) <= not b;
    layer4_outputs(1651) <= b;
    layer4_outputs(1652) <= not b or a;
    layer4_outputs(1653) <= b;
    layer4_outputs(1654) <= a and not b;
    layer4_outputs(1655) <= not (a xor b);
    layer4_outputs(1656) <= b;
    layer4_outputs(1657) <= not a;
    layer4_outputs(1658) <= not a;
    layer4_outputs(1659) <= not (a xor b);
    layer4_outputs(1660) <= not b;
    layer4_outputs(1661) <= a or b;
    layer4_outputs(1662) <= not b;
    layer4_outputs(1663) <= a;
    layer4_outputs(1664) <= not b;
    layer4_outputs(1665) <= '0';
    layer4_outputs(1666) <= b;
    layer4_outputs(1667) <= not a;
    layer4_outputs(1668) <= not (a or b);
    layer4_outputs(1669) <= a and b;
    layer4_outputs(1670) <= not a or b;
    layer4_outputs(1671) <= b;
    layer4_outputs(1672) <= a;
    layer4_outputs(1673) <= not (a and b);
    layer4_outputs(1674) <= not a;
    layer4_outputs(1675) <= a or b;
    layer4_outputs(1676) <= not a or b;
    layer4_outputs(1677) <= not a or b;
    layer4_outputs(1678) <= '1';
    layer4_outputs(1679) <= not a or b;
    layer4_outputs(1680) <= a;
    layer4_outputs(1681) <= b;
    layer4_outputs(1682) <= a;
    layer4_outputs(1683) <= a;
    layer4_outputs(1684) <= a;
    layer4_outputs(1685) <= not a or b;
    layer4_outputs(1686) <= not a;
    layer4_outputs(1687) <= not a;
    layer4_outputs(1688) <= a;
    layer4_outputs(1689) <= not a;
    layer4_outputs(1690) <= a and not b;
    layer4_outputs(1691) <= a and b;
    layer4_outputs(1692) <= not b;
    layer4_outputs(1693) <= b;
    layer4_outputs(1694) <= a and not b;
    layer4_outputs(1695) <= not (a and b);
    layer4_outputs(1696) <= b;
    layer4_outputs(1697) <= not b;
    layer4_outputs(1698) <= a and not b;
    layer4_outputs(1699) <= '1';
    layer4_outputs(1700) <= not a;
    layer4_outputs(1701) <= a xor b;
    layer4_outputs(1702) <= a;
    layer4_outputs(1703) <= not a or b;
    layer4_outputs(1704) <= not a;
    layer4_outputs(1705) <= b;
    layer4_outputs(1706) <= b and not a;
    layer4_outputs(1707) <= not a or b;
    layer4_outputs(1708) <= not b;
    layer4_outputs(1709) <= not b;
    layer4_outputs(1710) <= not (a xor b);
    layer4_outputs(1711) <= b;
    layer4_outputs(1712) <= not a or b;
    layer4_outputs(1713) <= not a;
    layer4_outputs(1714) <= not b or a;
    layer4_outputs(1715) <= a and not b;
    layer4_outputs(1716) <= b;
    layer4_outputs(1717) <= not b or a;
    layer4_outputs(1718) <= a or b;
    layer4_outputs(1719) <= not a;
    layer4_outputs(1720) <= b and not a;
    layer4_outputs(1721) <= not (a xor b);
    layer4_outputs(1722) <= a xor b;
    layer4_outputs(1723) <= not (a and b);
    layer4_outputs(1724) <= not (a or b);
    layer4_outputs(1725) <= '1';
    layer4_outputs(1726) <= a;
    layer4_outputs(1727) <= a;
    layer4_outputs(1728) <= b and not a;
    layer4_outputs(1729) <= not (a and b);
    layer4_outputs(1730) <= a;
    layer4_outputs(1731) <= not a;
    layer4_outputs(1732) <= not b;
    layer4_outputs(1733) <= not a;
    layer4_outputs(1734) <= a xor b;
    layer4_outputs(1735) <= a or b;
    layer4_outputs(1736) <= not a;
    layer4_outputs(1737) <= a or b;
    layer4_outputs(1738) <= not b or a;
    layer4_outputs(1739) <= b;
    layer4_outputs(1740) <= a xor b;
    layer4_outputs(1741) <= b;
    layer4_outputs(1742) <= not b or a;
    layer4_outputs(1743) <= a and b;
    layer4_outputs(1744) <= a xor b;
    layer4_outputs(1745) <= not (a xor b);
    layer4_outputs(1746) <= a and b;
    layer4_outputs(1747) <= a and b;
    layer4_outputs(1748) <= not b;
    layer4_outputs(1749) <= not (a or b);
    layer4_outputs(1750) <= not a or b;
    layer4_outputs(1751) <= not a;
    layer4_outputs(1752) <= not b;
    layer4_outputs(1753) <= a or b;
    layer4_outputs(1754) <= not a;
    layer4_outputs(1755) <= a xor b;
    layer4_outputs(1756) <= a or b;
    layer4_outputs(1757) <= a xor b;
    layer4_outputs(1758) <= b;
    layer4_outputs(1759) <= a and b;
    layer4_outputs(1760) <= a or b;
    layer4_outputs(1761) <= not b;
    layer4_outputs(1762) <= not b or a;
    layer4_outputs(1763) <= not (a or b);
    layer4_outputs(1764) <= b;
    layer4_outputs(1765) <= b;
    layer4_outputs(1766) <= not (a xor b);
    layer4_outputs(1767) <= not b;
    layer4_outputs(1768) <= not b;
    layer4_outputs(1769) <= not (a or b);
    layer4_outputs(1770) <= a and not b;
    layer4_outputs(1771) <= not a;
    layer4_outputs(1772) <= a or b;
    layer4_outputs(1773) <= a or b;
    layer4_outputs(1774) <= not (a xor b);
    layer4_outputs(1775) <= b and not a;
    layer4_outputs(1776) <= a and b;
    layer4_outputs(1777) <= not b or a;
    layer4_outputs(1778) <= a;
    layer4_outputs(1779) <= a;
    layer4_outputs(1780) <= not b or a;
    layer4_outputs(1781) <= b;
    layer4_outputs(1782) <= b and not a;
    layer4_outputs(1783) <= not (a or b);
    layer4_outputs(1784) <= b and not a;
    layer4_outputs(1785) <= a;
    layer4_outputs(1786) <= not b;
    layer4_outputs(1787) <= a and b;
    layer4_outputs(1788) <= b and not a;
    layer4_outputs(1789) <= not a or b;
    layer4_outputs(1790) <= a or b;
    layer4_outputs(1791) <= a;
    layer4_outputs(1792) <= not b;
    layer4_outputs(1793) <= not (a xor b);
    layer4_outputs(1794) <= not a;
    layer4_outputs(1795) <= a or b;
    layer4_outputs(1796) <= not a;
    layer4_outputs(1797) <= b and not a;
    layer4_outputs(1798) <= not b;
    layer4_outputs(1799) <= not b;
    layer4_outputs(1800) <= not (a xor b);
    layer4_outputs(1801) <= not a;
    layer4_outputs(1802) <= '1';
    layer4_outputs(1803) <= a and not b;
    layer4_outputs(1804) <= a and b;
    layer4_outputs(1805) <= not (a or b);
    layer4_outputs(1806) <= a xor b;
    layer4_outputs(1807) <= a and not b;
    layer4_outputs(1808) <= a and b;
    layer4_outputs(1809) <= a;
    layer4_outputs(1810) <= not b;
    layer4_outputs(1811) <= not b or a;
    layer4_outputs(1812) <= b and not a;
    layer4_outputs(1813) <= not a;
    layer4_outputs(1814) <= a and not b;
    layer4_outputs(1815) <= not a;
    layer4_outputs(1816) <= not a or b;
    layer4_outputs(1817) <= not b;
    layer4_outputs(1818) <= not b;
    layer4_outputs(1819) <= b;
    layer4_outputs(1820) <= not (a xor b);
    layer4_outputs(1821) <= b;
    layer4_outputs(1822) <= not (a or b);
    layer4_outputs(1823) <= not (a or b);
    layer4_outputs(1824) <= a;
    layer4_outputs(1825) <= not b;
    layer4_outputs(1826) <= not a or b;
    layer4_outputs(1827) <= b;
    layer4_outputs(1828) <= a xor b;
    layer4_outputs(1829) <= a;
    layer4_outputs(1830) <= a xor b;
    layer4_outputs(1831) <= a and b;
    layer4_outputs(1832) <= a;
    layer4_outputs(1833) <= a and not b;
    layer4_outputs(1834) <= b and not a;
    layer4_outputs(1835) <= not a;
    layer4_outputs(1836) <= not b;
    layer4_outputs(1837) <= not (a and b);
    layer4_outputs(1838) <= a;
    layer4_outputs(1839) <= not (a and b);
    layer4_outputs(1840) <= not (a and b);
    layer4_outputs(1841) <= b;
    layer4_outputs(1842) <= not b;
    layer4_outputs(1843) <= a;
    layer4_outputs(1844) <= not (a xor b);
    layer4_outputs(1845) <= not (a and b);
    layer4_outputs(1846) <= not a or b;
    layer4_outputs(1847) <= a xor b;
    layer4_outputs(1848) <= b and not a;
    layer4_outputs(1849) <= a and b;
    layer4_outputs(1850) <= not (a or b);
    layer4_outputs(1851) <= not b;
    layer4_outputs(1852) <= b and not a;
    layer4_outputs(1853) <= a and not b;
    layer4_outputs(1854) <= a and not b;
    layer4_outputs(1855) <= not a;
    layer4_outputs(1856) <= not a or b;
    layer4_outputs(1857) <= b and not a;
    layer4_outputs(1858) <= not (a and b);
    layer4_outputs(1859) <= a and b;
    layer4_outputs(1860) <= not b or a;
    layer4_outputs(1861) <= not b;
    layer4_outputs(1862) <= b;
    layer4_outputs(1863) <= a;
    layer4_outputs(1864) <= a and b;
    layer4_outputs(1865) <= a and not b;
    layer4_outputs(1866) <= not b;
    layer4_outputs(1867) <= a or b;
    layer4_outputs(1868) <= not b;
    layer4_outputs(1869) <= not a or b;
    layer4_outputs(1870) <= a;
    layer4_outputs(1871) <= a and b;
    layer4_outputs(1872) <= not b;
    layer4_outputs(1873) <= a and b;
    layer4_outputs(1874) <= b and not a;
    layer4_outputs(1875) <= not b;
    layer4_outputs(1876) <= not (a xor b);
    layer4_outputs(1877) <= not (a and b);
    layer4_outputs(1878) <= not a or b;
    layer4_outputs(1879) <= b;
    layer4_outputs(1880) <= not b;
    layer4_outputs(1881) <= a or b;
    layer4_outputs(1882) <= not b;
    layer4_outputs(1883) <= not a;
    layer4_outputs(1884) <= a;
    layer4_outputs(1885) <= not a or b;
    layer4_outputs(1886) <= b;
    layer4_outputs(1887) <= not (a and b);
    layer4_outputs(1888) <= a or b;
    layer4_outputs(1889) <= a xor b;
    layer4_outputs(1890) <= a and b;
    layer4_outputs(1891) <= a and b;
    layer4_outputs(1892) <= not a;
    layer4_outputs(1893) <= a and not b;
    layer4_outputs(1894) <= not a;
    layer4_outputs(1895) <= a and not b;
    layer4_outputs(1896) <= a;
    layer4_outputs(1897) <= not (a or b);
    layer4_outputs(1898) <= a or b;
    layer4_outputs(1899) <= a and b;
    layer4_outputs(1900) <= not b;
    layer4_outputs(1901) <= a xor b;
    layer4_outputs(1902) <= a and not b;
    layer4_outputs(1903) <= a;
    layer4_outputs(1904) <= not a;
    layer4_outputs(1905) <= b;
    layer4_outputs(1906) <= not b;
    layer4_outputs(1907) <= a and not b;
    layer4_outputs(1908) <= not b;
    layer4_outputs(1909) <= a;
    layer4_outputs(1910) <= a;
    layer4_outputs(1911) <= not a or b;
    layer4_outputs(1912) <= not b;
    layer4_outputs(1913) <= not a;
    layer4_outputs(1914) <= not b;
    layer4_outputs(1915) <= not (a or b);
    layer4_outputs(1916) <= a xor b;
    layer4_outputs(1917) <= a and b;
    layer4_outputs(1918) <= b;
    layer4_outputs(1919) <= b;
    layer4_outputs(1920) <= not b;
    layer4_outputs(1921) <= not b or a;
    layer4_outputs(1922) <= a xor b;
    layer4_outputs(1923) <= a and not b;
    layer4_outputs(1924) <= not b;
    layer4_outputs(1925) <= b;
    layer4_outputs(1926) <= b;
    layer4_outputs(1927) <= b and not a;
    layer4_outputs(1928) <= '0';
    layer4_outputs(1929) <= b;
    layer4_outputs(1930) <= not b;
    layer4_outputs(1931) <= b and not a;
    layer4_outputs(1932) <= b and not a;
    layer4_outputs(1933) <= b;
    layer4_outputs(1934) <= a and not b;
    layer4_outputs(1935) <= b;
    layer4_outputs(1936) <= not b;
    layer4_outputs(1937) <= not b;
    layer4_outputs(1938) <= a or b;
    layer4_outputs(1939) <= a or b;
    layer4_outputs(1940) <= a;
    layer4_outputs(1941) <= b;
    layer4_outputs(1942) <= '1';
    layer4_outputs(1943) <= not b or a;
    layer4_outputs(1944) <= not b or a;
    layer4_outputs(1945) <= not a or b;
    layer4_outputs(1946) <= a and not b;
    layer4_outputs(1947) <= b and not a;
    layer4_outputs(1948) <= a xor b;
    layer4_outputs(1949) <= b and not a;
    layer4_outputs(1950) <= a;
    layer4_outputs(1951) <= a and b;
    layer4_outputs(1952) <= a;
    layer4_outputs(1953) <= not b;
    layer4_outputs(1954) <= a xor b;
    layer4_outputs(1955) <= b and not a;
    layer4_outputs(1956) <= not (a xor b);
    layer4_outputs(1957) <= b;
    layer4_outputs(1958) <= b;
    layer4_outputs(1959) <= not (a and b);
    layer4_outputs(1960) <= a;
    layer4_outputs(1961) <= a and not b;
    layer4_outputs(1962) <= '0';
    layer4_outputs(1963) <= a xor b;
    layer4_outputs(1964) <= not b;
    layer4_outputs(1965) <= '0';
    layer4_outputs(1966) <= not a;
    layer4_outputs(1967) <= not b;
    layer4_outputs(1968) <= a and b;
    layer4_outputs(1969) <= '0';
    layer4_outputs(1970) <= a;
    layer4_outputs(1971) <= a;
    layer4_outputs(1972) <= not b;
    layer4_outputs(1973) <= not b;
    layer4_outputs(1974) <= b;
    layer4_outputs(1975) <= not b;
    layer4_outputs(1976) <= b;
    layer4_outputs(1977) <= '0';
    layer4_outputs(1978) <= not (a and b);
    layer4_outputs(1979) <= not (a or b);
    layer4_outputs(1980) <= not b;
    layer4_outputs(1981) <= a or b;
    layer4_outputs(1982) <= not b;
    layer4_outputs(1983) <= not b;
    layer4_outputs(1984) <= not (a and b);
    layer4_outputs(1985) <= not (a xor b);
    layer4_outputs(1986) <= not (a or b);
    layer4_outputs(1987) <= b;
    layer4_outputs(1988) <= not b;
    layer4_outputs(1989) <= not b or a;
    layer4_outputs(1990) <= not (a or b);
    layer4_outputs(1991) <= not a or b;
    layer4_outputs(1992) <= not a or b;
    layer4_outputs(1993) <= not a;
    layer4_outputs(1994) <= b and not a;
    layer4_outputs(1995) <= a and b;
    layer4_outputs(1996) <= b;
    layer4_outputs(1997) <= not b or a;
    layer4_outputs(1998) <= b and not a;
    layer4_outputs(1999) <= '1';
    layer4_outputs(2000) <= b and not a;
    layer4_outputs(2001) <= not b;
    layer4_outputs(2002) <= a xor b;
    layer4_outputs(2003) <= not b or a;
    layer4_outputs(2004) <= a;
    layer4_outputs(2005) <= a and b;
    layer4_outputs(2006) <= b;
    layer4_outputs(2007) <= a and not b;
    layer4_outputs(2008) <= not a or b;
    layer4_outputs(2009) <= a or b;
    layer4_outputs(2010) <= not a or b;
    layer4_outputs(2011) <= not a or b;
    layer4_outputs(2012) <= not b;
    layer4_outputs(2013) <= b;
    layer4_outputs(2014) <= b;
    layer4_outputs(2015) <= b;
    layer4_outputs(2016) <= b;
    layer4_outputs(2017) <= not b;
    layer4_outputs(2018) <= a or b;
    layer4_outputs(2019) <= a xor b;
    layer4_outputs(2020) <= a and b;
    layer4_outputs(2021) <= a and not b;
    layer4_outputs(2022) <= a and not b;
    layer4_outputs(2023) <= not a or b;
    layer4_outputs(2024) <= not (a or b);
    layer4_outputs(2025) <= b and not a;
    layer4_outputs(2026) <= a or b;
    layer4_outputs(2027) <= a and not b;
    layer4_outputs(2028) <= b and not a;
    layer4_outputs(2029) <= b;
    layer4_outputs(2030) <= b;
    layer4_outputs(2031) <= not b or a;
    layer4_outputs(2032) <= not b or a;
    layer4_outputs(2033) <= b;
    layer4_outputs(2034) <= a or b;
    layer4_outputs(2035) <= a or b;
    layer4_outputs(2036) <= not b or a;
    layer4_outputs(2037) <= '1';
    layer4_outputs(2038) <= b;
    layer4_outputs(2039) <= '0';
    layer4_outputs(2040) <= not (a or b);
    layer4_outputs(2041) <= '1';
    layer4_outputs(2042) <= not (a or b);
    layer4_outputs(2043) <= b;
    layer4_outputs(2044) <= not b or a;
    layer4_outputs(2045) <= not b or a;
    layer4_outputs(2046) <= b and not a;
    layer4_outputs(2047) <= a and b;
    layer4_outputs(2048) <= a and not b;
    layer4_outputs(2049) <= not (a xor b);
    layer4_outputs(2050) <= not a;
    layer4_outputs(2051) <= not (a xor b);
    layer4_outputs(2052) <= a and b;
    layer4_outputs(2053) <= not a;
    layer4_outputs(2054) <= a and b;
    layer4_outputs(2055) <= a or b;
    layer4_outputs(2056) <= a xor b;
    layer4_outputs(2057) <= not a;
    layer4_outputs(2058) <= b;
    layer4_outputs(2059) <= '0';
    layer4_outputs(2060) <= not a or b;
    layer4_outputs(2061) <= b;
    layer4_outputs(2062) <= b and not a;
    layer4_outputs(2063) <= b and not a;
    layer4_outputs(2064) <= not b or a;
    layer4_outputs(2065) <= a xor b;
    layer4_outputs(2066) <= a and not b;
    layer4_outputs(2067) <= not a;
    layer4_outputs(2068) <= '1';
    layer4_outputs(2069) <= '1';
    layer4_outputs(2070) <= not a;
    layer4_outputs(2071) <= a;
    layer4_outputs(2072) <= not b;
    layer4_outputs(2073) <= b and not a;
    layer4_outputs(2074) <= not a;
    layer4_outputs(2075) <= a;
    layer4_outputs(2076) <= not b;
    layer4_outputs(2077) <= not a;
    layer4_outputs(2078) <= a;
    layer4_outputs(2079) <= not a;
    layer4_outputs(2080) <= not (a xor b);
    layer4_outputs(2081) <= not a;
    layer4_outputs(2082) <= not b;
    layer4_outputs(2083) <= not (a and b);
    layer4_outputs(2084) <= not a;
    layer4_outputs(2085) <= not b or a;
    layer4_outputs(2086) <= b;
    layer4_outputs(2087) <= not b;
    layer4_outputs(2088) <= a and b;
    layer4_outputs(2089) <= '0';
    layer4_outputs(2090) <= a and b;
    layer4_outputs(2091) <= not (a and b);
    layer4_outputs(2092) <= a;
    layer4_outputs(2093) <= not a;
    layer4_outputs(2094) <= not a;
    layer4_outputs(2095) <= not (a and b);
    layer4_outputs(2096) <= a and b;
    layer4_outputs(2097) <= not a or b;
    layer4_outputs(2098) <= b;
    layer4_outputs(2099) <= not b or a;
    layer4_outputs(2100) <= a or b;
    layer4_outputs(2101) <= not a;
    layer4_outputs(2102) <= not (a and b);
    layer4_outputs(2103) <= not b or a;
    layer4_outputs(2104) <= not a;
    layer4_outputs(2105) <= '1';
    layer4_outputs(2106) <= a;
    layer4_outputs(2107) <= not (a or b);
    layer4_outputs(2108) <= '0';
    layer4_outputs(2109) <= '1';
    layer4_outputs(2110) <= not (a or b);
    layer4_outputs(2111) <= a and b;
    layer4_outputs(2112) <= b;
    layer4_outputs(2113) <= b;
    layer4_outputs(2114) <= b;
    layer4_outputs(2115) <= b;
    layer4_outputs(2116) <= a;
    layer4_outputs(2117) <= a and b;
    layer4_outputs(2118) <= not b;
    layer4_outputs(2119) <= b and not a;
    layer4_outputs(2120) <= a or b;
    layer4_outputs(2121) <= a and not b;
    layer4_outputs(2122) <= b;
    layer4_outputs(2123) <= b;
    layer4_outputs(2124) <= not a;
    layer4_outputs(2125) <= not a;
    layer4_outputs(2126) <= a or b;
    layer4_outputs(2127) <= b;
    layer4_outputs(2128) <= a or b;
    layer4_outputs(2129) <= not (a xor b);
    layer4_outputs(2130) <= '0';
    layer4_outputs(2131) <= not (a and b);
    layer4_outputs(2132) <= not (a or b);
    layer4_outputs(2133) <= not b;
    layer4_outputs(2134) <= '1';
    layer4_outputs(2135) <= not a or b;
    layer4_outputs(2136) <= a xor b;
    layer4_outputs(2137) <= b;
    layer4_outputs(2138) <= not a;
    layer4_outputs(2139) <= '1';
    layer4_outputs(2140) <= '0';
    layer4_outputs(2141) <= a and b;
    layer4_outputs(2142) <= b;
    layer4_outputs(2143) <= not (a or b);
    layer4_outputs(2144) <= not a;
    layer4_outputs(2145) <= not a or b;
    layer4_outputs(2146) <= '1';
    layer4_outputs(2147) <= not b;
    layer4_outputs(2148) <= a and not b;
    layer4_outputs(2149) <= not a;
    layer4_outputs(2150) <= not a;
    layer4_outputs(2151) <= '1';
    layer4_outputs(2152) <= a or b;
    layer4_outputs(2153) <= not (a and b);
    layer4_outputs(2154) <= not b;
    layer4_outputs(2155) <= not b;
    layer4_outputs(2156) <= a or b;
    layer4_outputs(2157) <= b;
    layer4_outputs(2158) <= not a or b;
    layer4_outputs(2159) <= a xor b;
    layer4_outputs(2160) <= b and not a;
    layer4_outputs(2161) <= not a;
    layer4_outputs(2162) <= a;
    layer4_outputs(2163) <= b;
    layer4_outputs(2164) <= b and not a;
    layer4_outputs(2165) <= not a;
    layer4_outputs(2166) <= b;
    layer4_outputs(2167) <= a or b;
    layer4_outputs(2168) <= not b or a;
    layer4_outputs(2169) <= a xor b;
    layer4_outputs(2170) <= '0';
    layer4_outputs(2171) <= not (a or b);
    layer4_outputs(2172) <= b;
    layer4_outputs(2173) <= not (a xor b);
    layer4_outputs(2174) <= not (a xor b);
    layer4_outputs(2175) <= a;
    layer4_outputs(2176) <= '0';
    layer4_outputs(2177) <= b;
    layer4_outputs(2178) <= not (a xor b);
    layer4_outputs(2179) <= a;
    layer4_outputs(2180) <= a or b;
    layer4_outputs(2181) <= a xor b;
    layer4_outputs(2182) <= b;
    layer4_outputs(2183) <= a xor b;
    layer4_outputs(2184) <= a and not b;
    layer4_outputs(2185) <= b;
    layer4_outputs(2186) <= a;
    layer4_outputs(2187) <= a;
    layer4_outputs(2188) <= a or b;
    layer4_outputs(2189) <= not (a or b);
    layer4_outputs(2190) <= a and not b;
    layer4_outputs(2191) <= b;
    layer4_outputs(2192) <= a and not b;
    layer4_outputs(2193) <= a and b;
    layer4_outputs(2194) <= a or b;
    layer4_outputs(2195) <= not b;
    layer4_outputs(2196) <= not (a or b);
    layer4_outputs(2197) <= not (a xor b);
    layer4_outputs(2198) <= not b or a;
    layer4_outputs(2199) <= a or b;
    layer4_outputs(2200) <= b;
    layer4_outputs(2201) <= a or b;
    layer4_outputs(2202) <= b;
    layer4_outputs(2203) <= a;
    layer4_outputs(2204) <= a;
    layer4_outputs(2205) <= b and not a;
    layer4_outputs(2206) <= not b;
    layer4_outputs(2207) <= not a or b;
    layer4_outputs(2208) <= not b;
    layer4_outputs(2209) <= a xor b;
    layer4_outputs(2210) <= not b;
    layer4_outputs(2211) <= a and b;
    layer4_outputs(2212) <= b;
    layer4_outputs(2213) <= b;
    layer4_outputs(2214) <= not b;
    layer4_outputs(2215) <= not a;
    layer4_outputs(2216) <= b;
    layer4_outputs(2217) <= b and not a;
    layer4_outputs(2218) <= not b or a;
    layer4_outputs(2219) <= a and b;
    layer4_outputs(2220) <= b;
    layer4_outputs(2221) <= not (a and b);
    layer4_outputs(2222) <= b;
    layer4_outputs(2223) <= not a or b;
    layer4_outputs(2224) <= not a;
    layer4_outputs(2225) <= '0';
    layer4_outputs(2226) <= not a;
    layer4_outputs(2227) <= b;
    layer4_outputs(2228) <= not b or a;
    layer4_outputs(2229) <= not (a xor b);
    layer4_outputs(2230) <= b;
    layer4_outputs(2231) <= b;
    layer4_outputs(2232) <= not (a or b);
    layer4_outputs(2233) <= a;
    layer4_outputs(2234) <= not b or a;
    layer4_outputs(2235) <= a and b;
    layer4_outputs(2236) <= a xor b;
    layer4_outputs(2237) <= a and b;
    layer4_outputs(2238) <= b;
    layer4_outputs(2239) <= a and not b;
    layer4_outputs(2240) <= not b or a;
    layer4_outputs(2241) <= not (a or b);
    layer4_outputs(2242) <= a and not b;
    layer4_outputs(2243) <= a;
    layer4_outputs(2244) <= b;
    layer4_outputs(2245) <= a xor b;
    layer4_outputs(2246) <= not (a or b);
    layer4_outputs(2247) <= '0';
    layer4_outputs(2248) <= not b;
    layer4_outputs(2249) <= '0';
    layer4_outputs(2250) <= '0';
    layer4_outputs(2251) <= a;
    layer4_outputs(2252) <= a and b;
    layer4_outputs(2253) <= a and not b;
    layer4_outputs(2254) <= b;
    layer4_outputs(2255) <= a xor b;
    layer4_outputs(2256) <= not a or b;
    layer4_outputs(2257) <= not (a or b);
    layer4_outputs(2258) <= not b or a;
    layer4_outputs(2259) <= a and not b;
    layer4_outputs(2260) <= a or b;
    layer4_outputs(2261) <= not a;
    layer4_outputs(2262) <= '0';
    layer4_outputs(2263) <= b and not a;
    layer4_outputs(2264) <= b and not a;
    layer4_outputs(2265) <= a;
    layer4_outputs(2266) <= b;
    layer4_outputs(2267) <= a and b;
    layer4_outputs(2268) <= not b;
    layer4_outputs(2269) <= a and b;
    layer4_outputs(2270) <= not b;
    layer4_outputs(2271) <= b and not a;
    layer4_outputs(2272) <= not b;
    layer4_outputs(2273) <= not (a or b);
    layer4_outputs(2274) <= b;
    layer4_outputs(2275) <= a and not b;
    layer4_outputs(2276) <= a and not b;
    layer4_outputs(2277) <= a;
    layer4_outputs(2278) <= not (a and b);
    layer4_outputs(2279) <= '0';
    layer4_outputs(2280) <= a and b;
    layer4_outputs(2281) <= not (a or b);
    layer4_outputs(2282) <= a;
    layer4_outputs(2283) <= not (a xor b);
    layer4_outputs(2284) <= a;
    layer4_outputs(2285) <= a xor b;
    layer4_outputs(2286) <= a or b;
    layer4_outputs(2287) <= b and not a;
    layer4_outputs(2288) <= not b or a;
    layer4_outputs(2289) <= a;
    layer4_outputs(2290) <= not (a and b);
    layer4_outputs(2291) <= not b;
    layer4_outputs(2292) <= not (a or b);
    layer4_outputs(2293) <= a and b;
    layer4_outputs(2294) <= b;
    layer4_outputs(2295) <= not b;
    layer4_outputs(2296) <= a or b;
    layer4_outputs(2297) <= not (a and b);
    layer4_outputs(2298) <= a;
    layer4_outputs(2299) <= not b or a;
    layer4_outputs(2300) <= a;
    layer4_outputs(2301) <= a;
    layer4_outputs(2302) <= a or b;
    layer4_outputs(2303) <= not b or a;
    layer4_outputs(2304) <= not b;
    layer4_outputs(2305) <= b;
    layer4_outputs(2306) <= not a or b;
    layer4_outputs(2307) <= not b or a;
    layer4_outputs(2308) <= a or b;
    layer4_outputs(2309) <= not (a and b);
    layer4_outputs(2310) <= b;
    layer4_outputs(2311) <= a xor b;
    layer4_outputs(2312) <= not b;
    layer4_outputs(2313) <= a;
    layer4_outputs(2314) <= not b;
    layer4_outputs(2315) <= not (a or b);
    layer4_outputs(2316) <= a and not b;
    layer4_outputs(2317) <= not (a or b);
    layer4_outputs(2318) <= not a or b;
    layer4_outputs(2319) <= a and b;
    layer4_outputs(2320) <= b and not a;
    layer4_outputs(2321) <= a and not b;
    layer4_outputs(2322) <= a xor b;
    layer4_outputs(2323) <= a xor b;
    layer4_outputs(2324) <= a xor b;
    layer4_outputs(2325) <= '1';
    layer4_outputs(2326) <= a;
    layer4_outputs(2327) <= not a;
    layer4_outputs(2328) <= a;
    layer4_outputs(2329) <= not (a and b);
    layer4_outputs(2330) <= not a;
    layer4_outputs(2331) <= not (a and b);
    layer4_outputs(2332) <= a and b;
    layer4_outputs(2333) <= not a;
    layer4_outputs(2334) <= not b;
    layer4_outputs(2335) <= not (a and b);
    layer4_outputs(2336) <= not a;
    layer4_outputs(2337) <= b;
    layer4_outputs(2338) <= a or b;
    layer4_outputs(2339) <= not b;
    layer4_outputs(2340) <= not a or b;
    layer4_outputs(2341) <= b;
    layer4_outputs(2342) <= not b;
    layer4_outputs(2343) <= a and b;
    layer4_outputs(2344) <= not b or a;
    layer4_outputs(2345) <= not (a and b);
    layer4_outputs(2346) <= a or b;
    layer4_outputs(2347) <= not a or b;
    layer4_outputs(2348) <= not b or a;
    layer4_outputs(2349) <= not (a xor b);
    layer4_outputs(2350) <= not b or a;
    layer4_outputs(2351) <= a or b;
    layer4_outputs(2352) <= not (a or b);
    layer4_outputs(2353) <= not (a xor b);
    layer4_outputs(2354) <= '0';
    layer4_outputs(2355) <= not b;
    layer4_outputs(2356) <= not b;
    layer4_outputs(2357) <= not a;
    layer4_outputs(2358) <= not b;
    layer4_outputs(2359) <= b and not a;
    layer4_outputs(2360) <= a and b;
    layer4_outputs(2361) <= not b;
    layer4_outputs(2362) <= a;
    layer4_outputs(2363) <= not b;
    layer4_outputs(2364) <= not a;
    layer4_outputs(2365) <= '0';
    layer4_outputs(2366) <= not a or b;
    layer4_outputs(2367) <= not b;
    layer4_outputs(2368) <= not (a and b);
    layer4_outputs(2369) <= not (a or b);
    layer4_outputs(2370) <= not b;
    layer4_outputs(2371) <= not b or a;
    layer4_outputs(2372) <= b;
    layer4_outputs(2373) <= not b or a;
    layer4_outputs(2374) <= a and not b;
    layer4_outputs(2375) <= a or b;
    layer4_outputs(2376) <= a;
    layer4_outputs(2377) <= not a or b;
    layer4_outputs(2378) <= not (a and b);
    layer4_outputs(2379) <= b;
    layer4_outputs(2380) <= a or b;
    layer4_outputs(2381) <= not a;
    layer4_outputs(2382) <= a xor b;
    layer4_outputs(2383) <= b;
    layer4_outputs(2384) <= not (a and b);
    layer4_outputs(2385) <= a xor b;
    layer4_outputs(2386) <= not a or b;
    layer4_outputs(2387) <= b and not a;
    layer4_outputs(2388) <= b and not a;
    layer4_outputs(2389) <= not a or b;
    layer4_outputs(2390) <= not a;
    layer4_outputs(2391) <= b and not a;
    layer4_outputs(2392) <= not a;
    layer4_outputs(2393) <= not a;
    layer4_outputs(2394) <= not b;
    layer4_outputs(2395) <= a and b;
    layer4_outputs(2396) <= not a;
    layer4_outputs(2397) <= not a;
    layer4_outputs(2398) <= '1';
    layer4_outputs(2399) <= not a;
    layer4_outputs(2400) <= not b;
    layer4_outputs(2401) <= b and not a;
    layer4_outputs(2402) <= not (a xor b);
    layer4_outputs(2403) <= not b;
    layer4_outputs(2404) <= not a;
    layer4_outputs(2405) <= '0';
    layer4_outputs(2406) <= b and not a;
    layer4_outputs(2407) <= not b;
    layer4_outputs(2408) <= b;
    layer4_outputs(2409) <= a and b;
    layer4_outputs(2410) <= not a;
    layer4_outputs(2411) <= not a;
    layer4_outputs(2412) <= not (a or b);
    layer4_outputs(2413) <= not b;
    layer4_outputs(2414) <= not b;
    layer4_outputs(2415) <= not (a xor b);
    layer4_outputs(2416) <= a or b;
    layer4_outputs(2417) <= not b;
    layer4_outputs(2418) <= a;
    layer4_outputs(2419) <= not a;
    layer4_outputs(2420) <= '1';
    layer4_outputs(2421) <= not a or b;
    layer4_outputs(2422) <= a;
    layer4_outputs(2423) <= not b or a;
    layer4_outputs(2424) <= a and not b;
    layer4_outputs(2425) <= a or b;
    layer4_outputs(2426) <= not a;
    layer4_outputs(2427) <= a xor b;
    layer4_outputs(2428) <= a;
    layer4_outputs(2429) <= a and b;
    layer4_outputs(2430) <= not b or a;
    layer4_outputs(2431) <= not a or b;
    layer4_outputs(2432) <= not (a xor b);
    layer4_outputs(2433) <= '0';
    layer4_outputs(2434) <= a;
    layer4_outputs(2435) <= not b or a;
    layer4_outputs(2436) <= not b;
    layer4_outputs(2437) <= not (a xor b);
    layer4_outputs(2438) <= a or b;
    layer4_outputs(2439) <= a or b;
    layer4_outputs(2440) <= a and not b;
    layer4_outputs(2441) <= not b;
    layer4_outputs(2442) <= b and not a;
    layer4_outputs(2443) <= b;
    layer4_outputs(2444) <= not a;
    layer4_outputs(2445) <= a xor b;
    layer4_outputs(2446) <= a or b;
    layer4_outputs(2447) <= a and b;
    layer4_outputs(2448) <= not b;
    layer4_outputs(2449) <= b and not a;
    layer4_outputs(2450) <= a;
    layer4_outputs(2451) <= a xor b;
    layer4_outputs(2452) <= not (a or b);
    layer4_outputs(2453) <= a or b;
    layer4_outputs(2454) <= a and b;
    layer4_outputs(2455) <= not a or b;
    layer4_outputs(2456) <= b;
    layer4_outputs(2457) <= not (a and b);
    layer4_outputs(2458) <= b and not a;
    layer4_outputs(2459) <= not b;
    layer4_outputs(2460) <= not a;
    layer4_outputs(2461) <= a or b;
    layer4_outputs(2462) <= a;
    layer4_outputs(2463) <= a;
    layer4_outputs(2464) <= b and not a;
    layer4_outputs(2465) <= a;
    layer4_outputs(2466) <= a xor b;
    layer4_outputs(2467) <= a;
    layer4_outputs(2468) <= not b;
    layer4_outputs(2469) <= not b;
    layer4_outputs(2470) <= a and b;
    layer4_outputs(2471) <= not (a and b);
    layer4_outputs(2472) <= b;
    layer4_outputs(2473) <= a;
    layer4_outputs(2474) <= b;
    layer4_outputs(2475) <= b and not a;
    layer4_outputs(2476) <= not (a xor b);
    layer4_outputs(2477) <= b and not a;
    layer4_outputs(2478) <= b and not a;
    layer4_outputs(2479) <= b;
    layer4_outputs(2480) <= not b or a;
    layer4_outputs(2481) <= a and b;
    layer4_outputs(2482) <= not (a and b);
    layer4_outputs(2483) <= not (a or b);
    layer4_outputs(2484) <= b;
    layer4_outputs(2485) <= not b;
    layer4_outputs(2486) <= a;
    layer4_outputs(2487) <= b and not a;
    layer4_outputs(2488) <= b;
    layer4_outputs(2489) <= b;
    layer4_outputs(2490) <= a or b;
    layer4_outputs(2491) <= not (a or b);
    layer4_outputs(2492) <= not a;
    layer4_outputs(2493) <= a and b;
    layer4_outputs(2494) <= not b;
    layer4_outputs(2495) <= not (a or b);
    layer4_outputs(2496) <= not (a xor b);
    layer4_outputs(2497) <= a xor b;
    layer4_outputs(2498) <= a and not b;
    layer4_outputs(2499) <= not (a or b);
    layer4_outputs(2500) <= not a;
    layer4_outputs(2501) <= not b;
    layer4_outputs(2502) <= a;
    layer4_outputs(2503) <= a or b;
    layer4_outputs(2504) <= not b;
    layer4_outputs(2505) <= b;
    layer4_outputs(2506) <= b;
    layer4_outputs(2507) <= b and not a;
    layer4_outputs(2508) <= b;
    layer4_outputs(2509) <= b;
    layer4_outputs(2510) <= not b;
    layer4_outputs(2511) <= b and not a;
    layer4_outputs(2512) <= not (a and b);
    layer4_outputs(2513) <= not a or b;
    layer4_outputs(2514) <= '0';
    layer4_outputs(2515) <= a;
    layer4_outputs(2516) <= a xor b;
    layer4_outputs(2517) <= a xor b;
    layer4_outputs(2518) <= a or b;
    layer4_outputs(2519) <= not a or b;
    layer4_outputs(2520) <= a or b;
    layer4_outputs(2521) <= not a or b;
    layer4_outputs(2522) <= b and not a;
    layer4_outputs(2523) <= a;
    layer4_outputs(2524) <= not (a xor b);
    layer4_outputs(2525) <= a;
    layer4_outputs(2526) <= b;
    layer4_outputs(2527) <= not (a and b);
    layer4_outputs(2528) <= not b;
    layer4_outputs(2529) <= a and b;
    layer4_outputs(2530) <= not a;
    layer4_outputs(2531) <= a and not b;
    layer4_outputs(2532) <= '0';
    layer4_outputs(2533) <= a xor b;
    layer4_outputs(2534) <= not b or a;
    layer4_outputs(2535) <= b and not a;
    layer4_outputs(2536) <= a xor b;
    layer4_outputs(2537) <= not (a and b);
    layer4_outputs(2538) <= a xor b;
    layer4_outputs(2539) <= not b or a;
    layer4_outputs(2540) <= '1';
    layer4_outputs(2541) <= a xor b;
    layer4_outputs(2542) <= a;
    layer4_outputs(2543) <= a and b;
    layer4_outputs(2544) <= not b or a;
    layer4_outputs(2545) <= b;
    layer4_outputs(2546) <= a;
    layer4_outputs(2547) <= not a or b;
    layer4_outputs(2548) <= not b;
    layer4_outputs(2549) <= b and not a;
    layer4_outputs(2550) <= not b or a;
    layer4_outputs(2551) <= not b;
    layer4_outputs(2552) <= not (a and b);
    layer4_outputs(2553) <= not (a xor b);
    layer4_outputs(2554) <= not a;
    layer4_outputs(2555) <= not (a xor b);
    layer4_outputs(2556) <= a and not b;
    layer4_outputs(2557) <= '0';
    layer4_outputs(2558) <= not a;
    layer4_outputs(2559) <= not (a and b);
    layer4_outputs(2560) <= not (a xor b);
    layer4_outputs(2561) <= a and not b;
    layer4_outputs(2562) <= a or b;
    layer4_outputs(2563) <= a;
    layer4_outputs(2564) <= not b or a;
    layer4_outputs(2565) <= not (a or b);
    layer4_outputs(2566) <= not b or a;
    layer4_outputs(2567) <= not a;
    layer4_outputs(2568) <= a;
    layer4_outputs(2569) <= b;
    layer4_outputs(2570) <= not (a xor b);
    layer4_outputs(2571) <= not (a xor b);
    layer4_outputs(2572) <= not b or a;
    layer4_outputs(2573) <= a;
    layer4_outputs(2574) <= not a;
    layer4_outputs(2575) <= not (a or b);
    layer4_outputs(2576) <= a and b;
    layer4_outputs(2577) <= a or b;
    layer4_outputs(2578) <= b;
    layer4_outputs(2579) <= a;
    layer4_outputs(2580) <= a and not b;
    layer4_outputs(2581) <= not b;
    layer4_outputs(2582) <= a or b;
    layer4_outputs(2583) <= not a;
    layer4_outputs(2584) <= not (a xor b);
    layer4_outputs(2585) <= not (a or b);
    layer4_outputs(2586) <= not a or b;
    layer4_outputs(2587) <= not a or b;
    layer4_outputs(2588) <= a and b;
    layer4_outputs(2589) <= a;
    layer4_outputs(2590) <= a;
    layer4_outputs(2591) <= not b;
    layer4_outputs(2592) <= not b;
    layer4_outputs(2593) <= '1';
    layer4_outputs(2594) <= b and not a;
    layer4_outputs(2595) <= not (a or b);
    layer4_outputs(2596) <= '0';
    layer4_outputs(2597) <= a and not b;
    layer4_outputs(2598) <= not (a or b);
    layer4_outputs(2599) <= b;
    layer4_outputs(2600) <= a xor b;
    layer4_outputs(2601) <= not a;
    layer4_outputs(2602) <= not (a xor b);
    layer4_outputs(2603) <= not b;
    layer4_outputs(2604) <= not b;
    layer4_outputs(2605) <= not a;
    layer4_outputs(2606) <= not b or a;
    layer4_outputs(2607) <= b;
    layer4_outputs(2608) <= a and not b;
    layer4_outputs(2609) <= not (a or b);
    layer4_outputs(2610) <= not b or a;
    layer4_outputs(2611) <= not (a and b);
    layer4_outputs(2612) <= not a;
    layer4_outputs(2613) <= a and not b;
    layer4_outputs(2614) <= a and not b;
    layer4_outputs(2615) <= a and b;
    layer4_outputs(2616) <= not a or b;
    layer4_outputs(2617) <= not b;
    layer4_outputs(2618) <= b and not a;
    layer4_outputs(2619) <= a and b;
    layer4_outputs(2620) <= not a;
    layer4_outputs(2621) <= a and b;
    layer4_outputs(2622) <= not a;
    layer4_outputs(2623) <= a and not b;
    layer4_outputs(2624) <= not b or a;
    layer4_outputs(2625) <= not b;
    layer4_outputs(2626) <= b and not a;
    layer4_outputs(2627) <= not (a and b);
    layer4_outputs(2628) <= '1';
    layer4_outputs(2629) <= not b;
    layer4_outputs(2630) <= a or b;
    layer4_outputs(2631) <= b and not a;
    layer4_outputs(2632) <= a;
    layer4_outputs(2633) <= a;
    layer4_outputs(2634) <= a;
    layer4_outputs(2635) <= not a;
    layer4_outputs(2636) <= a and not b;
    layer4_outputs(2637) <= '0';
    layer4_outputs(2638) <= a and not b;
    layer4_outputs(2639) <= not a;
    layer4_outputs(2640) <= '0';
    layer4_outputs(2641) <= a or b;
    layer4_outputs(2642) <= a and b;
    layer4_outputs(2643) <= b;
    layer4_outputs(2644) <= not b or a;
    layer4_outputs(2645) <= not a;
    layer4_outputs(2646) <= not (a or b);
    layer4_outputs(2647) <= not (a or b);
    layer4_outputs(2648) <= a and b;
    layer4_outputs(2649) <= a and not b;
    layer4_outputs(2650) <= not b;
    layer4_outputs(2651) <= a;
    layer4_outputs(2652) <= not (a and b);
    layer4_outputs(2653) <= a;
    layer4_outputs(2654) <= b;
    layer4_outputs(2655) <= not b;
    layer4_outputs(2656) <= b;
    layer4_outputs(2657) <= not b;
    layer4_outputs(2658) <= not b or a;
    layer4_outputs(2659) <= b;
    layer4_outputs(2660) <= not (a xor b);
    layer4_outputs(2661) <= a xor b;
    layer4_outputs(2662) <= not (a or b);
    layer4_outputs(2663) <= not (a or b);
    layer4_outputs(2664) <= not a;
    layer4_outputs(2665) <= a;
    layer4_outputs(2666) <= '0';
    layer4_outputs(2667) <= not b;
    layer4_outputs(2668) <= a and b;
    layer4_outputs(2669) <= not (a or b);
    layer4_outputs(2670) <= a;
    layer4_outputs(2671) <= not a;
    layer4_outputs(2672) <= not a;
    layer4_outputs(2673) <= not (a xor b);
    layer4_outputs(2674) <= not a;
    layer4_outputs(2675) <= a or b;
    layer4_outputs(2676) <= not (a and b);
    layer4_outputs(2677) <= not (a or b);
    layer4_outputs(2678) <= not b or a;
    layer4_outputs(2679) <= a xor b;
    layer4_outputs(2680) <= not a or b;
    layer4_outputs(2681) <= not a;
    layer4_outputs(2682) <= not a;
    layer4_outputs(2683) <= '0';
    layer4_outputs(2684) <= not b;
    layer4_outputs(2685) <= not a;
    layer4_outputs(2686) <= a and not b;
    layer4_outputs(2687) <= not a;
    layer4_outputs(2688) <= a and b;
    layer4_outputs(2689) <= a xor b;
    layer4_outputs(2690) <= not (a or b);
    layer4_outputs(2691) <= not a or b;
    layer4_outputs(2692) <= a or b;
    layer4_outputs(2693) <= not a;
    layer4_outputs(2694) <= a and not b;
    layer4_outputs(2695) <= a xor b;
    layer4_outputs(2696) <= not a;
    layer4_outputs(2697) <= b and not a;
    layer4_outputs(2698) <= not (a or b);
    layer4_outputs(2699) <= not a;
    layer4_outputs(2700) <= not (a or b);
    layer4_outputs(2701) <= not (a and b);
    layer4_outputs(2702) <= not (a and b);
    layer4_outputs(2703) <= a;
    layer4_outputs(2704) <= not (a or b);
    layer4_outputs(2705) <= not b;
    layer4_outputs(2706) <= b and not a;
    layer4_outputs(2707) <= not a or b;
    layer4_outputs(2708) <= not (a xor b);
    layer4_outputs(2709) <= not (a and b);
    layer4_outputs(2710) <= not b or a;
    layer4_outputs(2711) <= a xor b;
    layer4_outputs(2712) <= not b or a;
    layer4_outputs(2713) <= not a or b;
    layer4_outputs(2714) <= not (a xor b);
    layer4_outputs(2715) <= not (a or b);
    layer4_outputs(2716) <= not b;
    layer4_outputs(2717) <= b;
    layer4_outputs(2718) <= a and b;
    layer4_outputs(2719) <= a;
    layer4_outputs(2720) <= not b or a;
    layer4_outputs(2721) <= not (a or b);
    layer4_outputs(2722) <= not (a and b);
    layer4_outputs(2723) <= a and b;
    layer4_outputs(2724) <= not (a or b);
    layer4_outputs(2725) <= a and not b;
    layer4_outputs(2726) <= not a or b;
    layer4_outputs(2727) <= a;
    layer4_outputs(2728) <= not a;
    layer4_outputs(2729) <= not a;
    layer4_outputs(2730) <= '0';
    layer4_outputs(2731) <= not b;
    layer4_outputs(2732) <= b and not a;
    layer4_outputs(2733) <= not (a or b);
    layer4_outputs(2734) <= not a;
    layer4_outputs(2735) <= b;
    layer4_outputs(2736) <= a or b;
    layer4_outputs(2737) <= a or b;
    layer4_outputs(2738) <= b and not a;
    layer4_outputs(2739) <= not (a xor b);
    layer4_outputs(2740) <= not b;
    layer4_outputs(2741) <= not (a and b);
    layer4_outputs(2742) <= not (a xor b);
    layer4_outputs(2743) <= '0';
    layer4_outputs(2744) <= not (a and b);
    layer4_outputs(2745) <= not b;
    layer4_outputs(2746) <= a;
    layer4_outputs(2747) <= not (a xor b);
    layer4_outputs(2748) <= a and b;
    layer4_outputs(2749) <= not a;
    layer4_outputs(2750) <= '0';
    layer4_outputs(2751) <= a and b;
    layer4_outputs(2752) <= not b;
    layer4_outputs(2753) <= '1';
    layer4_outputs(2754) <= b;
    layer4_outputs(2755) <= '1';
    layer4_outputs(2756) <= a;
    layer4_outputs(2757) <= not a;
    layer4_outputs(2758) <= a and not b;
    layer4_outputs(2759) <= a;
    layer4_outputs(2760) <= not b;
    layer4_outputs(2761) <= not a;
    layer4_outputs(2762) <= a and not b;
    layer4_outputs(2763) <= not b;
    layer4_outputs(2764) <= '1';
    layer4_outputs(2765) <= not b;
    layer4_outputs(2766) <= '0';
    layer4_outputs(2767) <= b and not a;
    layer4_outputs(2768) <= b and not a;
    layer4_outputs(2769) <= not a or b;
    layer4_outputs(2770) <= a and b;
    layer4_outputs(2771) <= not a;
    layer4_outputs(2772) <= b;
    layer4_outputs(2773) <= a and b;
    layer4_outputs(2774) <= not (a or b);
    layer4_outputs(2775) <= not (a and b);
    layer4_outputs(2776) <= a and not b;
    layer4_outputs(2777) <= a and not b;
    layer4_outputs(2778) <= '0';
    layer4_outputs(2779) <= a;
    layer4_outputs(2780) <= not a;
    layer4_outputs(2781) <= a or b;
    layer4_outputs(2782) <= not b;
    layer4_outputs(2783) <= a or b;
    layer4_outputs(2784) <= not (a and b);
    layer4_outputs(2785) <= not a;
    layer4_outputs(2786) <= a;
    layer4_outputs(2787) <= '1';
    layer4_outputs(2788) <= '1';
    layer4_outputs(2789) <= not (a or b);
    layer4_outputs(2790) <= not (a or b);
    layer4_outputs(2791) <= a and b;
    layer4_outputs(2792) <= b;
    layer4_outputs(2793) <= a xor b;
    layer4_outputs(2794) <= not b or a;
    layer4_outputs(2795) <= b and not a;
    layer4_outputs(2796) <= not b;
    layer4_outputs(2797) <= not b;
    layer4_outputs(2798) <= b;
    layer4_outputs(2799) <= a xor b;
    layer4_outputs(2800) <= b;
    layer4_outputs(2801) <= a and not b;
    layer4_outputs(2802) <= not (a or b);
    layer4_outputs(2803) <= not (a xor b);
    layer4_outputs(2804) <= not b or a;
    layer4_outputs(2805) <= a and not b;
    layer4_outputs(2806) <= a or b;
    layer4_outputs(2807) <= b and not a;
    layer4_outputs(2808) <= a;
    layer4_outputs(2809) <= b and not a;
    layer4_outputs(2810) <= '0';
    layer4_outputs(2811) <= a xor b;
    layer4_outputs(2812) <= not a or b;
    layer4_outputs(2813) <= '0';
    layer4_outputs(2814) <= not a or b;
    layer4_outputs(2815) <= '0';
    layer4_outputs(2816) <= a or b;
    layer4_outputs(2817) <= a or b;
    layer4_outputs(2818) <= not (a or b);
    layer4_outputs(2819) <= not b;
    layer4_outputs(2820) <= not b or a;
    layer4_outputs(2821) <= not a or b;
    layer4_outputs(2822) <= not b;
    layer4_outputs(2823) <= not b or a;
    layer4_outputs(2824) <= not (a and b);
    layer4_outputs(2825) <= a or b;
    layer4_outputs(2826) <= b;
    layer4_outputs(2827) <= not (a or b);
    layer4_outputs(2828) <= not b;
    layer4_outputs(2829) <= not b;
    layer4_outputs(2830) <= not a;
    layer4_outputs(2831) <= not (a or b);
    layer4_outputs(2832) <= b and not a;
    layer4_outputs(2833) <= not b or a;
    layer4_outputs(2834) <= b and not a;
    layer4_outputs(2835) <= b;
    layer4_outputs(2836) <= a and not b;
    layer4_outputs(2837) <= not a;
    layer4_outputs(2838) <= b;
    layer4_outputs(2839) <= b;
    layer4_outputs(2840) <= a and b;
    layer4_outputs(2841) <= not a or b;
    layer4_outputs(2842) <= a and not b;
    layer4_outputs(2843) <= a and b;
    layer4_outputs(2844) <= b;
    layer4_outputs(2845) <= a and not b;
    layer4_outputs(2846) <= not (a and b);
    layer4_outputs(2847) <= a;
    layer4_outputs(2848) <= a and not b;
    layer4_outputs(2849) <= not b;
    layer4_outputs(2850) <= a xor b;
    layer4_outputs(2851) <= a and not b;
    layer4_outputs(2852) <= b;
    layer4_outputs(2853) <= not a or b;
    layer4_outputs(2854) <= not b;
    layer4_outputs(2855) <= b;
    layer4_outputs(2856) <= a or b;
    layer4_outputs(2857) <= a or b;
    layer4_outputs(2858) <= a or b;
    layer4_outputs(2859) <= not b;
    layer4_outputs(2860) <= not b;
    layer4_outputs(2861) <= b;
    layer4_outputs(2862) <= a and not b;
    layer4_outputs(2863) <= not a;
    layer4_outputs(2864) <= not (a xor b);
    layer4_outputs(2865) <= a or b;
    layer4_outputs(2866) <= not (a or b);
    layer4_outputs(2867) <= not (a or b);
    layer4_outputs(2868) <= '1';
    layer4_outputs(2869) <= not (a or b);
    layer4_outputs(2870) <= a and not b;
    layer4_outputs(2871) <= not b or a;
    layer4_outputs(2872) <= b;
    layer4_outputs(2873) <= not (a xor b);
    layer4_outputs(2874) <= not a;
    layer4_outputs(2875) <= not a;
    layer4_outputs(2876) <= a;
    layer4_outputs(2877) <= b;
    layer4_outputs(2878) <= not b;
    layer4_outputs(2879) <= not a or b;
    layer4_outputs(2880) <= not b or a;
    layer4_outputs(2881) <= b;
    layer4_outputs(2882) <= not (a or b);
    layer4_outputs(2883) <= '0';
    layer4_outputs(2884) <= not b;
    layer4_outputs(2885) <= b;
    layer4_outputs(2886) <= a or b;
    layer4_outputs(2887) <= b;
    layer4_outputs(2888) <= a or b;
    layer4_outputs(2889) <= a xor b;
    layer4_outputs(2890) <= a and b;
    layer4_outputs(2891) <= '0';
    layer4_outputs(2892) <= a;
    layer4_outputs(2893) <= not a;
    layer4_outputs(2894) <= b;
    layer4_outputs(2895) <= a or b;
    layer4_outputs(2896) <= not b;
    layer4_outputs(2897) <= not a;
    layer4_outputs(2898) <= a;
    layer4_outputs(2899) <= a and b;
    layer4_outputs(2900) <= not b;
    layer4_outputs(2901) <= b;
    layer4_outputs(2902) <= '0';
    layer4_outputs(2903) <= a xor b;
    layer4_outputs(2904) <= not a or b;
    layer4_outputs(2905) <= not a;
    layer4_outputs(2906) <= not a;
    layer4_outputs(2907) <= not b or a;
    layer4_outputs(2908) <= not b or a;
    layer4_outputs(2909) <= not b;
    layer4_outputs(2910) <= a or b;
    layer4_outputs(2911) <= a or b;
    layer4_outputs(2912) <= not (a or b);
    layer4_outputs(2913) <= not a or b;
    layer4_outputs(2914) <= a xor b;
    layer4_outputs(2915) <= not (a or b);
    layer4_outputs(2916) <= b and not a;
    layer4_outputs(2917) <= not a;
    layer4_outputs(2918) <= a and b;
    layer4_outputs(2919) <= not b;
    layer4_outputs(2920) <= not a or b;
    layer4_outputs(2921) <= not b or a;
    layer4_outputs(2922) <= not b or a;
    layer4_outputs(2923) <= not (a xor b);
    layer4_outputs(2924) <= not (a xor b);
    layer4_outputs(2925) <= not (a and b);
    layer4_outputs(2926) <= a and b;
    layer4_outputs(2927) <= a or b;
    layer4_outputs(2928) <= '0';
    layer4_outputs(2929) <= '1';
    layer4_outputs(2930) <= b and not a;
    layer4_outputs(2931) <= not a;
    layer4_outputs(2932) <= a;
    layer4_outputs(2933) <= not a;
    layer4_outputs(2934) <= not b;
    layer4_outputs(2935) <= not (a or b);
    layer4_outputs(2936) <= not b or a;
    layer4_outputs(2937) <= not b;
    layer4_outputs(2938) <= not a;
    layer4_outputs(2939) <= not a;
    layer4_outputs(2940) <= not (a xor b);
    layer4_outputs(2941) <= a;
    layer4_outputs(2942) <= a and b;
    layer4_outputs(2943) <= not b or a;
    layer4_outputs(2944) <= a or b;
    layer4_outputs(2945) <= a or b;
    layer4_outputs(2946) <= not a;
    layer4_outputs(2947) <= not a;
    layer4_outputs(2948) <= not b;
    layer4_outputs(2949) <= not b;
    layer4_outputs(2950) <= not (a and b);
    layer4_outputs(2951) <= not a;
    layer4_outputs(2952) <= not (a and b);
    layer4_outputs(2953) <= not a or b;
    layer4_outputs(2954) <= not b;
    layer4_outputs(2955) <= a;
    layer4_outputs(2956) <= a;
    layer4_outputs(2957) <= a;
    layer4_outputs(2958) <= a or b;
    layer4_outputs(2959) <= '0';
    layer4_outputs(2960) <= a or b;
    layer4_outputs(2961) <= not (a or b);
    layer4_outputs(2962) <= not a or b;
    layer4_outputs(2963) <= a and not b;
    layer4_outputs(2964) <= a xor b;
    layer4_outputs(2965) <= not b or a;
    layer4_outputs(2966) <= a;
    layer4_outputs(2967) <= a;
    layer4_outputs(2968) <= b and not a;
    layer4_outputs(2969) <= not a or b;
    layer4_outputs(2970) <= a;
    layer4_outputs(2971) <= not (a and b);
    layer4_outputs(2972) <= a and not b;
    layer4_outputs(2973) <= not (a xor b);
    layer4_outputs(2974) <= b;
    layer4_outputs(2975) <= a xor b;
    layer4_outputs(2976) <= not (a and b);
    layer4_outputs(2977) <= b and not a;
    layer4_outputs(2978) <= not a;
    layer4_outputs(2979) <= b;
    layer4_outputs(2980) <= b;
    layer4_outputs(2981) <= not b or a;
    layer4_outputs(2982) <= not a;
    layer4_outputs(2983) <= not (a and b);
    layer4_outputs(2984) <= a and b;
    layer4_outputs(2985) <= not a;
    layer4_outputs(2986) <= not (a and b);
    layer4_outputs(2987) <= a xor b;
    layer4_outputs(2988) <= a and b;
    layer4_outputs(2989) <= b;
    layer4_outputs(2990) <= not (a and b);
    layer4_outputs(2991) <= a or b;
    layer4_outputs(2992) <= '1';
    layer4_outputs(2993) <= not b;
    layer4_outputs(2994) <= not (a and b);
    layer4_outputs(2995) <= not b or a;
    layer4_outputs(2996) <= not a;
    layer4_outputs(2997) <= b and not a;
    layer4_outputs(2998) <= not b or a;
    layer4_outputs(2999) <= not a;
    layer4_outputs(3000) <= '0';
    layer4_outputs(3001) <= not a;
    layer4_outputs(3002) <= a or b;
    layer4_outputs(3003) <= not (a or b);
    layer4_outputs(3004) <= a and b;
    layer4_outputs(3005) <= a;
    layer4_outputs(3006) <= a and b;
    layer4_outputs(3007) <= a and b;
    layer4_outputs(3008) <= not b;
    layer4_outputs(3009) <= '0';
    layer4_outputs(3010) <= b;
    layer4_outputs(3011) <= not (a or b);
    layer4_outputs(3012) <= not b;
    layer4_outputs(3013) <= not (a xor b);
    layer4_outputs(3014) <= a and not b;
    layer4_outputs(3015) <= a;
    layer4_outputs(3016) <= a and b;
    layer4_outputs(3017) <= a and b;
    layer4_outputs(3018) <= not (a xor b);
    layer4_outputs(3019) <= b and not a;
    layer4_outputs(3020) <= b and not a;
    layer4_outputs(3021) <= not (a or b);
    layer4_outputs(3022) <= not a or b;
    layer4_outputs(3023) <= a;
    layer4_outputs(3024) <= not a;
    layer4_outputs(3025) <= not a or b;
    layer4_outputs(3026) <= a or b;
    layer4_outputs(3027) <= a;
    layer4_outputs(3028) <= a and b;
    layer4_outputs(3029) <= a;
    layer4_outputs(3030) <= b;
    layer4_outputs(3031) <= a;
    layer4_outputs(3032) <= not b;
    layer4_outputs(3033) <= not a;
    layer4_outputs(3034) <= b;
    layer4_outputs(3035) <= a and b;
    layer4_outputs(3036) <= not a;
    layer4_outputs(3037) <= a or b;
    layer4_outputs(3038) <= '1';
    layer4_outputs(3039) <= a xor b;
    layer4_outputs(3040) <= not a;
    layer4_outputs(3041) <= a and not b;
    layer4_outputs(3042) <= not a;
    layer4_outputs(3043) <= not (a or b);
    layer4_outputs(3044) <= not (a or b);
    layer4_outputs(3045) <= not a;
    layer4_outputs(3046) <= a;
    layer4_outputs(3047) <= a and not b;
    layer4_outputs(3048) <= a and not b;
    layer4_outputs(3049) <= a;
    layer4_outputs(3050) <= b;
    layer4_outputs(3051) <= not b or a;
    layer4_outputs(3052) <= not a;
    layer4_outputs(3053) <= not a;
    layer4_outputs(3054) <= b;
    layer4_outputs(3055) <= not a;
    layer4_outputs(3056) <= a;
    layer4_outputs(3057) <= a xor b;
    layer4_outputs(3058) <= b;
    layer4_outputs(3059) <= a;
    layer4_outputs(3060) <= a;
    layer4_outputs(3061) <= a and b;
    layer4_outputs(3062) <= not a;
    layer4_outputs(3063) <= not (a xor b);
    layer4_outputs(3064) <= not a;
    layer4_outputs(3065) <= not (a or b);
    layer4_outputs(3066) <= not (a xor b);
    layer4_outputs(3067) <= a and b;
    layer4_outputs(3068) <= not a;
    layer4_outputs(3069) <= not a;
    layer4_outputs(3070) <= b;
    layer4_outputs(3071) <= not (a and b);
    layer4_outputs(3072) <= not a;
    layer4_outputs(3073) <= not a;
    layer4_outputs(3074) <= not (a or b);
    layer4_outputs(3075) <= b;
    layer4_outputs(3076) <= b;
    layer4_outputs(3077) <= not b;
    layer4_outputs(3078) <= b and not a;
    layer4_outputs(3079) <= not (a and b);
    layer4_outputs(3080) <= not b;
    layer4_outputs(3081) <= a and not b;
    layer4_outputs(3082) <= b;
    layer4_outputs(3083) <= a;
    layer4_outputs(3084) <= not a or b;
    layer4_outputs(3085) <= b;
    layer4_outputs(3086) <= a;
    layer4_outputs(3087) <= not b;
    layer4_outputs(3088) <= not a;
    layer4_outputs(3089) <= a xor b;
    layer4_outputs(3090) <= not (a xor b);
    layer4_outputs(3091) <= a;
    layer4_outputs(3092) <= b and not a;
    layer4_outputs(3093) <= not (a and b);
    layer4_outputs(3094) <= a xor b;
    layer4_outputs(3095) <= a or b;
    layer4_outputs(3096) <= not b;
    layer4_outputs(3097) <= not (a and b);
    layer4_outputs(3098) <= b and not a;
    layer4_outputs(3099) <= a;
    layer4_outputs(3100) <= a xor b;
    layer4_outputs(3101) <= a or b;
    layer4_outputs(3102) <= not a;
    layer4_outputs(3103) <= '1';
    layer4_outputs(3104) <= a and b;
    layer4_outputs(3105) <= not (a and b);
    layer4_outputs(3106) <= not a or b;
    layer4_outputs(3107) <= not a;
    layer4_outputs(3108) <= a and b;
    layer4_outputs(3109) <= a and b;
    layer4_outputs(3110) <= a and not b;
    layer4_outputs(3111) <= not b;
    layer4_outputs(3112) <= a;
    layer4_outputs(3113) <= not b;
    layer4_outputs(3114) <= a or b;
    layer4_outputs(3115) <= not (a and b);
    layer4_outputs(3116) <= b;
    layer4_outputs(3117) <= a xor b;
    layer4_outputs(3118) <= not (a xor b);
    layer4_outputs(3119) <= '1';
    layer4_outputs(3120) <= not b;
    layer4_outputs(3121) <= not b or a;
    layer4_outputs(3122) <= not (a or b);
    layer4_outputs(3123) <= not (a or b);
    layer4_outputs(3124) <= not (a xor b);
    layer4_outputs(3125) <= a;
    layer4_outputs(3126) <= not a;
    layer4_outputs(3127) <= b;
    layer4_outputs(3128) <= '1';
    layer4_outputs(3129) <= a and not b;
    layer4_outputs(3130) <= a and b;
    layer4_outputs(3131) <= b;
    layer4_outputs(3132) <= a and b;
    layer4_outputs(3133) <= not b;
    layer4_outputs(3134) <= a and b;
    layer4_outputs(3135) <= b and not a;
    layer4_outputs(3136) <= not (a or b);
    layer4_outputs(3137) <= not a or b;
    layer4_outputs(3138) <= a;
    layer4_outputs(3139) <= not a;
    layer4_outputs(3140) <= not b or a;
    layer4_outputs(3141) <= not a or b;
    layer4_outputs(3142) <= not a;
    layer4_outputs(3143) <= not b;
    layer4_outputs(3144) <= not (a or b);
    layer4_outputs(3145) <= not (a and b);
    layer4_outputs(3146) <= a and b;
    layer4_outputs(3147) <= b;
    layer4_outputs(3148) <= not b or a;
    layer4_outputs(3149) <= a xor b;
    layer4_outputs(3150) <= not (a or b);
    layer4_outputs(3151) <= not a;
    layer4_outputs(3152) <= b;
    layer4_outputs(3153) <= not a;
    layer4_outputs(3154) <= '0';
    layer4_outputs(3155) <= a;
    layer4_outputs(3156) <= a xor b;
    layer4_outputs(3157) <= a and b;
    layer4_outputs(3158) <= a and b;
    layer4_outputs(3159) <= a;
    layer4_outputs(3160) <= b;
    layer4_outputs(3161) <= not b;
    layer4_outputs(3162) <= not b;
    layer4_outputs(3163) <= not (a xor b);
    layer4_outputs(3164) <= a;
    layer4_outputs(3165) <= a and not b;
    layer4_outputs(3166) <= not b;
    layer4_outputs(3167) <= not a;
    layer4_outputs(3168) <= not a or b;
    layer4_outputs(3169) <= b;
    layer4_outputs(3170) <= a xor b;
    layer4_outputs(3171) <= b;
    layer4_outputs(3172) <= a and not b;
    layer4_outputs(3173) <= not (a and b);
    layer4_outputs(3174) <= b;
    layer4_outputs(3175) <= '0';
    layer4_outputs(3176) <= '1';
    layer4_outputs(3177) <= b;
    layer4_outputs(3178) <= not a;
    layer4_outputs(3179) <= a;
    layer4_outputs(3180) <= not (a and b);
    layer4_outputs(3181) <= b and not a;
    layer4_outputs(3182) <= a;
    layer4_outputs(3183) <= a;
    layer4_outputs(3184) <= a and not b;
    layer4_outputs(3185) <= '0';
    layer4_outputs(3186) <= not a or b;
    layer4_outputs(3187) <= a and b;
    layer4_outputs(3188) <= a;
    layer4_outputs(3189) <= b and not a;
    layer4_outputs(3190) <= not a;
    layer4_outputs(3191) <= not (a or b);
    layer4_outputs(3192) <= b;
    layer4_outputs(3193) <= not a;
    layer4_outputs(3194) <= not (a and b);
    layer4_outputs(3195) <= not b or a;
    layer4_outputs(3196) <= b;
    layer4_outputs(3197) <= b;
    layer4_outputs(3198) <= not b or a;
    layer4_outputs(3199) <= a;
    layer4_outputs(3200) <= a;
    layer4_outputs(3201) <= b;
    layer4_outputs(3202) <= not a;
    layer4_outputs(3203) <= b and not a;
    layer4_outputs(3204) <= not b;
    layer4_outputs(3205) <= a;
    layer4_outputs(3206) <= a xor b;
    layer4_outputs(3207) <= not (a or b);
    layer4_outputs(3208) <= not a or b;
    layer4_outputs(3209) <= b and not a;
    layer4_outputs(3210) <= a;
    layer4_outputs(3211) <= a xor b;
    layer4_outputs(3212) <= b;
    layer4_outputs(3213) <= a or b;
    layer4_outputs(3214) <= a or b;
    layer4_outputs(3215) <= not b;
    layer4_outputs(3216) <= a and b;
    layer4_outputs(3217) <= not a;
    layer4_outputs(3218) <= not a;
    layer4_outputs(3219) <= b and not a;
    layer4_outputs(3220) <= not a or b;
    layer4_outputs(3221) <= a xor b;
    layer4_outputs(3222) <= b;
    layer4_outputs(3223) <= not b;
    layer4_outputs(3224) <= b and not a;
    layer4_outputs(3225) <= not b;
    layer4_outputs(3226) <= a and not b;
    layer4_outputs(3227) <= a or b;
    layer4_outputs(3228) <= not (a and b);
    layer4_outputs(3229) <= not (a xor b);
    layer4_outputs(3230) <= not (a xor b);
    layer4_outputs(3231) <= not a;
    layer4_outputs(3232) <= a;
    layer4_outputs(3233) <= not (a and b);
    layer4_outputs(3234) <= not b;
    layer4_outputs(3235) <= b and not a;
    layer4_outputs(3236) <= a and b;
    layer4_outputs(3237) <= a;
    layer4_outputs(3238) <= not a;
    layer4_outputs(3239) <= not b;
    layer4_outputs(3240) <= not a;
    layer4_outputs(3241) <= a and b;
    layer4_outputs(3242) <= not (a or b);
    layer4_outputs(3243) <= b;
    layer4_outputs(3244) <= not b;
    layer4_outputs(3245) <= not a or b;
    layer4_outputs(3246) <= not a;
    layer4_outputs(3247) <= a;
    layer4_outputs(3248) <= not (a or b);
    layer4_outputs(3249) <= not (a and b);
    layer4_outputs(3250) <= a or b;
    layer4_outputs(3251) <= a and b;
    layer4_outputs(3252) <= b;
    layer4_outputs(3253) <= not (a xor b);
    layer4_outputs(3254) <= not a;
    layer4_outputs(3255) <= b and not a;
    layer4_outputs(3256) <= not a or b;
    layer4_outputs(3257) <= not b;
    layer4_outputs(3258) <= a;
    layer4_outputs(3259) <= not (a or b);
    layer4_outputs(3260) <= b;
    layer4_outputs(3261) <= a and not b;
    layer4_outputs(3262) <= not b or a;
    layer4_outputs(3263) <= not a;
    layer4_outputs(3264) <= not b;
    layer4_outputs(3265) <= not (a or b);
    layer4_outputs(3266) <= not b;
    layer4_outputs(3267) <= not (a xor b);
    layer4_outputs(3268) <= not (a and b);
    layer4_outputs(3269) <= b;
    layer4_outputs(3270) <= not b or a;
    layer4_outputs(3271) <= not b;
    layer4_outputs(3272) <= not b;
    layer4_outputs(3273) <= b;
    layer4_outputs(3274) <= a;
    layer4_outputs(3275) <= not b;
    layer4_outputs(3276) <= not b;
    layer4_outputs(3277) <= a and not b;
    layer4_outputs(3278) <= a and not b;
    layer4_outputs(3279) <= '1';
    layer4_outputs(3280) <= not b;
    layer4_outputs(3281) <= b and not a;
    layer4_outputs(3282) <= a and b;
    layer4_outputs(3283) <= a xor b;
    layer4_outputs(3284) <= not a or b;
    layer4_outputs(3285) <= not (a xor b);
    layer4_outputs(3286) <= b and not a;
    layer4_outputs(3287) <= a;
    layer4_outputs(3288) <= a and not b;
    layer4_outputs(3289) <= not (a xor b);
    layer4_outputs(3290) <= not b or a;
    layer4_outputs(3291) <= b;
    layer4_outputs(3292) <= not b;
    layer4_outputs(3293) <= not b or a;
    layer4_outputs(3294) <= not a or b;
    layer4_outputs(3295) <= a;
    layer4_outputs(3296) <= b and not a;
    layer4_outputs(3297) <= b;
    layer4_outputs(3298) <= a and not b;
    layer4_outputs(3299) <= not (a and b);
    layer4_outputs(3300) <= not b;
    layer4_outputs(3301) <= '0';
    layer4_outputs(3302) <= not a or b;
    layer4_outputs(3303) <= b;
    layer4_outputs(3304) <= not a;
    layer4_outputs(3305) <= a or b;
    layer4_outputs(3306) <= not (a or b);
    layer4_outputs(3307) <= a or b;
    layer4_outputs(3308) <= a and b;
    layer4_outputs(3309) <= a or b;
    layer4_outputs(3310) <= not (a xor b);
    layer4_outputs(3311) <= not b;
    layer4_outputs(3312) <= a or b;
    layer4_outputs(3313) <= '0';
    layer4_outputs(3314) <= a;
    layer4_outputs(3315) <= a;
    layer4_outputs(3316) <= a or b;
    layer4_outputs(3317) <= b and not a;
    layer4_outputs(3318) <= a xor b;
    layer4_outputs(3319) <= not b;
    layer4_outputs(3320) <= not b;
    layer4_outputs(3321) <= not a;
    layer4_outputs(3322) <= a or b;
    layer4_outputs(3323) <= not (a and b);
    layer4_outputs(3324) <= not a or b;
    layer4_outputs(3325) <= not b;
    layer4_outputs(3326) <= '1';
    layer4_outputs(3327) <= not (a or b);
    layer4_outputs(3328) <= not a;
    layer4_outputs(3329) <= a and not b;
    layer4_outputs(3330) <= a xor b;
    layer4_outputs(3331) <= not a;
    layer4_outputs(3332) <= not b or a;
    layer4_outputs(3333) <= not a;
    layer4_outputs(3334) <= not a;
    layer4_outputs(3335) <= a and not b;
    layer4_outputs(3336) <= b and not a;
    layer4_outputs(3337) <= not (a xor b);
    layer4_outputs(3338) <= not b;
    layer4_outputs(3339) <= b;
    layer4_outputs(3340) <= not (a or b);
    layer4_outputs(3341) <= b;
    layer4_outputs(3342) <= not a;
    layer4_outputs(3343) <= not a;
    layer4_outputs(3344) <= a xor b;
    layer4_outputs(3345) <= b and not a;
    layer4_outputs(3346) <= '0';
    layer4_outputs(3347) <= not b;
    layer4_outputs(3348) <= not b;
    layer4_outputs(3349) <= not b;
    layer4_outputs(3350) <= a and b;
    layer4_outputs(3351) <= a and b;
    layer4_outputs(3352) <= not (a and b);
    layer4_outputs(3353) <= not a;
    layer4_outputs(3354) <= a;
    layer4_outputs(3355) <= a;
    layer4_outputs(3356) <= '0';
    layer4_outputs(3357) <= '1';
    layer4_outputs(3358) <= b;
    layer4_outputs(3359) <= not (a xor b);
    layer4_outputs(3360) <= a;
    layer4_outputs(3361) <= a or b;
    layer4_outputs(3362) <= a and b;
    layer4_outputs(3363) <= a;
    layer4_outputs(3364) <= a and b;
    layer4_outputs(3365) <= b and not a;
    layer4_outputs(3366) <= not b;
    layer4_outputs(3367) <= not b;
    layer4_outputs(3368) <= not b;
    layer4_outputs(3369) <= not a or b;
    layer4_outputs(3370) <= a and not b;
    layer4_outputs(3371) <= not a;
    layer4_outputs(3372) <= not b;
    layer4_outputs(3373) <= not a or b;
    layer4_outputs(3374) <= not (a or b);
    layer4_outputs(3375) <= a or b;
    layer4_outputs(3376) <= b and not a;
    layer4_outputs(3377) <= a and not b;
    layer4_outputs(3378) <= a;
    layer4_outputs(3379) <= not a or b;
    layer4_outputs(3380) <= b;
    layer4_outputs(3381) <= a;
    layer4_outputs(3382) <= a;
    layer4_outputs(3383) <= not b or a;
    layer4_outputs(3384) <= a or b;
    layer4_outputs(3385) <= a and not b;
    layer4_outputs(3386) <= a and not b;
    layer4_outputs(3387) <= not a;
    layer4_outputs(3388) <= '0';
    layer4_outputs(3389) <= b;
    layer4_outputs(3390) <= not (a and b);
    layer4_outputs(3391) <= b and not a;
    layer4_outputs(3392) <= not b or a;
    layer4_outputs(3393) <= not (a xor b);
    layer4_outputs(3394) <= not a or b;
    layer4_outputs(3395) <= not (a and b);
    layer4_outputs(3396) <= b;
    layer4_outputs(3397) <= a or b;
    layer4_outputs(3398) <= not a;
    layer4_outputs(3399) <= a;
    layer4_outputs(3400) <= not b or a;
    layer4_outputs(3401) <= not a;
    layer4_outputs(3402) <= not a;
    layer4_outputs(3403) <= not a;
    layer4_outputs(3404) <= a or b;
    layer4_outputs(3405) <= a and b;
    layer4_outputs(3406) <= a;
    layer4_outputs(3407) <= not (a or b);
    layer4_outputs(3408) <= a and b;
    layer4_outputs(3409) <= not b or a;
    layer4_outputs(3410) <= not b;
    layer4_outputs(3411) <= not b or a;
    layer4_outputs(3412) <= not b or a;
    layer4_outputs(3413) <= not (a or b);
    layer4_outputs(3414) <= b;
    layer4_outputs(3415) <= not a or b;
    layer4_outputs(3416) <= not a or b;
    layer4_outputs(3417) <= b;
    layer4_outputs(3418) <= '0';
    layer4_outputs(3419) <= '0';
    layer4_outputs(3420) <= not a;
    layer4_outputs(3421) <= not b or a;
    layer4_outputs(3422) <= a;
    layer4_outputs(3423) <= '1';
    layer4_outputs(3424) <= a;
    layer4_outputs(3425) <= not a;
    layer4_outputs(3426) <= a;
    layer4_outputs(3427) <= not (a and b);
    layer4_outputs(3428) <= b;
    layer4_outputs(3429) <= a xor b;
    layer4_outputs(3430) <= not b;
    layer4_outputs(3431) <= a;
    layer4_outputs(3432) <= a;
    layer4_outputs(3433) <= a;
    layer4_outputs(3434) <= not (a or b);
    layer4_outputs(3435) <= b;
    layer4_outputs(3436) <= a and b;
    layer4_outputs(3437) <= b;
    layer4_outputs(3438) <= a or b;
    layer4_outputs(3439) <= b and not a;
    layer4_outputs(3440) <= a and b;
    layer4_outputs(3441) <= a or b;
    layer4_outputs(3442) <= not a or b;
    layer4_outputs(3443) <= not (a or b);
    layer4_outputs(3444) <= not (a xor b);
    layer4_outputs(3445) <= a and b;
    layer4_outputs(3446) <= not b or a;
    layer4_outputs(3447) <= a or b;
    layer4_outputs(3448) <= not b or a;
    layer4_outputs(3449) <= not a;
    layer4_outputs(3450) <= not b or a;
    layer4_outputs(3451) <= not (a xor b);
    layer4_outputs(3452) <= not (a and b);
    layer4_outputs(3453) <= not a;
    layer4_outputs(3454) <= b;
    layer4_outputs(3455) <= not b or a;
    layer4_outputs(3456) <= not a;
    layer4_outputs(3457) <= not (a xor b);
    layer4_outputs(3458) <= a;
    layer4_outputs(3459) <= not b or a;
    layer4_outputs(3460) <= b;
    layer4_outputs(3461) <= not b;
    layer4_outputs(3462) <= b and not a;
    layer4_outputs(3463) <= b;
    layer4_outputs(3464) <= a;
    layer4_outputs(3465) <= not (a or b);
    layer4_outputs(3466) <= a and b;
    layer4_outputs(3467) <= a or b;
    layer4_outputs(3468) <= a and b;
    layer4_outputs(3469) <= not a;
    layer4_outputs(3470) <= '0';
    layer4_outputs(3471) <= a;
    layer4_outputs(3472) <= b;
    layer4_outputs(3473) <= '1';
    layer4_outputs(3474) <= '0';
    layer4_outputs(3475) <= a and b;
    layer4_outputs(3476) <= not b;
    layer4_outputs(3477) <= b;
    layer4_outputs(3478) <= not a;
    layer4_outputs(3479) <= not b;
    layer4_outputs(3480) <= a or b;
    layer4_outputs(3481) <= a and b;
    layer4_outputs(3482) <= b;
    layer4_outputs(3483) <= a;
    layer4_outputs(3484) <= not b;
    layer4_outputs(3485) <= not a or b;
    layer4_outputs(3486) <= not a;
    layer4_outputs(3487) <= b;
    layer4_outputs(3488) <= b and not a;
    layer4_outputs(3489) <= not (a and b);
    layer4_outputs(3490) <= b;
    layer4_outputs(3491) <= a and not b;
    layer4_outputs(3492) <= not (a or b);
    layer4_outputs(3493) <= b and not a;
    layer4_outputs(3494) <= not (a or b);
    layer4_outputs(3495) <= not b;
    layer4_outputs(3496) <= b and not a;
    layer4_outputs(3497) <= a or b;
    layer4_outputs(3498) <= a xor b;
    layer4_outputs(3499) <= a;
    layer4_outputs(3500) <= not b or a;
    layer4_outputs(3501) <= b;
    layer4_outputs(3502) <= not (a xor b);
    layer4_outputs(3503) <= not (a xor b);
    layer4_outputs(3504) <= '1';
    layer4_outputs(3505) <= not (a or b);
    layer4_outputs(3506) <= b;
    layer4_outputs(3507) <= b;
    layer4_outputs(3508) <= a xor b;
    layer4_outputs(3509) <= not (a or b);
    layer4_outputs(3510) <= b;
    layer4_outputs(3511) <= not a or b;
    layer4_outputs(3512) <= not a;
    layer4_outputs(3513) <= not (a and b);
    layer4_outputs(3514) <= a or b;
    layer4_outputs(3515) <= a and not b;
    layer4_outputs(3516) <= not a;
    layer4_outputs(3517) <= a or b;
    layer4_outputs(3518) <= not a;
    layer4_outputs(3519) <= a;
    layer4_outputs(3520) <= a and not b;
    layer4_outputs(3521) <= not a or b;
    layer4_outputs(3522) <= b and not a;
    layer4_outputs(3523) <= not a;
    layer4_outputs(3524) <= b;
    layer4_outputs(3525) <= a and not b;
    layer4_outputs(3526) <= a or b;
    layer4_outputs(3527) <= b;
    layer4_outputs(3528) <= not (a xor b);
    layer4_outputs(3529) <= not a;
    layer4_outputs(3530) <= a and not b;
    layer4_outputs(3531) <= a and not b;
    layer4_outputs(3532) <= not a;
    layer4_outputs(3533) <= not a or b;
    layer4_outputs(3534) <= b;
    layer4_outputs(3535) <= not (a xor b);
    layer4_outputs(3536) <= a;
    layer4_outputs(3537) <= a;
    layer4_outputs(3538) <= '1';
    layer4_outputs(3539) <= b;
    layer4_outputs(3540) <= a;
    layer4_outputs(3541) <= a xor b;
    layer4_outputs(3542) <= not (a or b);
    layer4_outputs(3543) <= a;
    layer4_outputs(3544) <= not b or a;
    layer4_outputs(3545) <= not (a or b);
    layer4_outputs(3546) <= a and b;
    layer4_outputs(3547) <= b and not a;
    layer4_outputs(3548) <= b;
    layer4_outputs(3549) <= not a;
    layer4_outputs(3550) <= b;
    layer4_outputs(3551) <= not b;
    layer4_outputs(3552) <= a and b;
    layer4_outputs(3553) <= a;
    layer4_outputs(3554) <= b;
    layer4_outputs(3555) <= a;
    layer4_outputs(3556) <= a and not b;
    layer4_outputs(3557) <= not (a or b);
    layer4_outputs(3558) <= not b or a;
    layer4_outputs(3559) <= not (a or b);
    layer4_outputs(3560) <= not b;
    layer4_outputs(3561) <= '0';
    layer4_outputs(3562) <= '0';
    layer4_outputs(3563) <= not b;
    layer4_outputs(3564) <= not (a and b);
    layer4_outputs(3565) <= not b;
    layer4_outputs(3566) <= not a;
    layer4_outputs(3567) <= a and b;
    layer4_outputs(3568) <= a and b;
    layer4_outputs(3569) <= a or b;
    layer4_outputs(3570) <= not b;
    layer4_outputs(3571) <= b and not a;
    layer4_outputs(3572) <= not b;
    layer4_outputs(3573) <= a xor b;
    layer4_outputs(3574) <= b;
    layer4_outputs(3575) <= a and b;
    layer4_outputs(3576) <= a and not b;
    layer4_outputs(3577) <= not a;
    layer4_outputs(3578) <= a and b;
    layer4_outputs(3579) <= not (a or b);
    layer4_outputs(3580) <= not a;
    layer4_outputs(3581) <= not (a xor b);
    layer4_outputs(3582) <= '0';
    layer4_outputs(3583) <= not a;
    layer4_outputs(3584) <= not b;
    layer4_outputs(3585) <= not a;
    layer4_outputs(3586) <= b;
    layer4_outputs(3587) <= '0';
    layer4_outputs(3588) <= not b or a;
    layer4_outputs(3589) <= a;
    layer4_outputs(3590) <= '0';
    layer4_outputs(3591) <= not (a or b);
    layer4_outputs(3592) <= not a;
    layer4_outputs(3593) <= '1';
    layer4_outputs(3594) <= '1';
    layer4_outputs(3595) <= not (a and b);
    layer4_outputs(3596) <= not b;
    layer4_outputs(3597) <= not a;
    layer4_outputs(3598) <= not a or b;
    layer4_outputs(3599) <= a and b;
    layer4_outputs(3600) <= not a;
    layer4_outputs(3601) <= '0';
    layer4_outputs(3602) <= not a;
    layer4_outputs(3603) <= not (a xor b);
    layer4_outputs(3604) <= not (a and b);
    layer4_outputs(3605) <= not (a and b);
    layer4_outputs(3606) <= a and b;
    layer4_outputs(3607) <= a;
    layer4_outputs(3608) <= b;
    layer4_outputs(3609) <= not b;
    layer4_outputs(3610) <= a;
    layer4_outputs(3611) <= not (a or b);
    layer4_outputs(3612) <= not (a and b);
    layer4_outputs(3613) <= not (a and b);
    layer4_outputs(3614) <= a and b;
    layer4_outputs(3615) <= a and b;
    layer4_outputs(3616) <= not (a and b);
    layer4_outputs(3617) <= not a;
    layer4_outputs(3618) <= b;
    layer4_outputs(3619) <= not a;
    layer4_outputs(3620) <= not b;
    layer4_outputs(3621) <= not a;
    layer4_outputs(3622) <= not a;
    layer4_outputs(3623) <= a;
    layer4_outputs(3624) <= a and not b;
    layer4_outputs(3625) <= b and not a;
    layer4_outputs(3626) <= not (a or b);
    layer4_outputs(3627) <= a;
    layer4_outputs(3628) <= not (a xor b);
    layer4_outputs(3629) <= '0';
    layer4_outputs(3630) <= not (a and b);
    layer4_outputs(3631) <= b;
    layer4_outputs(3632) <= not a;
    layer4_outputs(3633) <= a or b;
    layer4_outputs(3634) <= b and not a;
    layer4_outputs(3635) <= a or b;
    layer4_outputs(3636) <= not a;
    layer4_outputs(3637) <= a and not b;
    layer4_outputs(3638) <= a and not b;
    layer4_outputs(3639) <= not (a or b);
    layer4_outputs(3640) <= a;
    layer4_outputs(3641) <= a;
    layer4_outputs(3642) <= not b or a;
    layer4_outputs(3643) <= b;
    layer4_outputs(3644) <= not (a xor b);
    layer4_outputs(3645) <= b and not a;
    layer4_outputs(3646) <= a;
    layer4_outputs(3647) <= not a or b;
    layer4_outputs(3648) <= b;
    layer4_outputs(3649) <= a and b;
    layer4_outputs(3650) <= a;
    layer4_outputs(3651) <= a xor b;
    layer4_outputs(3652) <= not (a or b);
    layer4_outputs(3653) <= not (a and b);
    layer4_outputs(3654) <= not a;
    layer4_outputs(3655) <= not b;
    layer4_outputs(3656) <= not (a or b);
    layer4_outputs(3657) <= not (a or b);
    layer4_outputs(3658) <= not b or a;
    layer4_outputs(3659) <= b;
    layer4_outputs(3660) <= not b or a;
    layer4_outputs(3661) <= not b;
    layer4_outputs(3662) <= not b;
    layer4_outputs(3663) <= not b or a;
    layer4_outputs(3664) <= b;
    layer4_outputs(3665) <= a or b;
    layer4_outputs(3666) <= not a;
    layer4_outputs(3667) <= b;
    layer4_outputs(3668) <= not a;
    layer4_outputs(3669) <= a;
    layer4_outputs(3670) <= not b;
    layer4_outputs(3671) <= a and b;
    layer4_outputs(3672) <= b and not a;
    layer4_outputs(3673) <= a and not b;
    layer4_outputs(3674) <= a or b;
    layer4_outputs(3675) <= a;
    layer4_outputs(3676) <= a and b;
    layer4_outputs(3677) <= not b;
    layer4_outputs(3678) <= b and not a;
    layer4_outputs(3679) <= not (a or b);
    layer4_outputs(3680) <= not a;
    layer4_outputs(3681) <= not (a or b);
    layer4_outputs(3682) <= not (a and b);
    layer4_outputs(3683) <= a and b;
    layer4_outputs(3684) <= not b;
    layer4_outputs(3685) <= not (a xor b);
    layer4_outputs(3686) <= a and not b;
    layer4_outputs(3687) <= a and b;
    layer4_outputs(3688) <= not a or b;
    layer4_outputs(3689) <= not b;
    layer4_outputs(3690) <= not a;
    layer4_outputs(3691) <= a;
    layer4_outputs(3692) <= not (a or b);
    layer4_outputs(3693) <= b;
    layer4_outputs(3694) <= '0';
    layer4_outputs(3695) <= b;
    layer4_outputs(3696) <= not a;
    layer4_outputs(3697) <= not b;
    layer4_outputs(3698) <= b;
    layer4_outputs(3699) <= not (a and b);
    layer4_outputs(3700) <= a;
    layer4_outputs(3701) <= not a;
    layer4_outputs(3702) <= b;
    layer4_outputs(3703) <= a;
    layer4_outputs(3704) <= not (a and b);
    layer4_outputs(3705) <= not b;
    layer4_outputs(3706) <= a xor b;
    layer4_outputs(3707) <= not a;
    layer4_outputs(3708) <= a and not b;
    layer4_outputs(3709) <= b and not a;
    layer4_outputs(3710) <= not a;
    layer4_outputs(3711) <= not (a or b);
    layer4_outputs(3712) <= not a;
    layer4_outputs(3713) <= a or b;
    layer4_outputs(3714) <= not a;
    layer4_outputs(3715) <= not b;
    layer4_outputs(3716) <= a;
    layer4_outputs(3717) <= '0';
    layer4_outputs(3718) <= '1';
    layer4_outputs(3719) <= a xor b;
    layer4_outputs(3720) <= not (a and b);
    layer4_outputs(3721) <= a or b;
    layer4_outputs(3722) <= '0';
    layer4_outputs(3723) <= not a or b;
    layer4_outputs(3724) <= a and b;
    layer4_outputs(3725) <= a;
    layer4_outputs(3726) <= not b or a;
    layer4_outputs(3727) <= a or b;
    layer4_outputs(3728) <= not a;
    layer4_outputs(3729) <= b and not a;
    layer4_outputs(3730) <= a;
    layer4_outputs(3731) <= a and not b;
    layer4_outputs(3732) <= not a or b;
    layer4_outputs(3733) <= not b or a;
    layer4_outputs(3734) <= not b;
    layer4_outputs(3735) <= a and not b;
    layer4_outputs(3736) <= a;
    layer4_outputs(3737) <= not a;
    layer4_outputs(3738) <= not b or a;
    layer4_outputs(3739) <= not b or a;
    layer4_outputs(3740) <= not b;
    layer4_outputs(3741) <= not (a xor b);
    layer4_outputs(3742) <= not a;
    layer4_outputs(3743) <= a and not b;
    layer4_outputs(3744) <= not b;
    layer4_outputs(3745) <= not b or a;
    layer4_outputs(3746) <= not b;
    layer4_outputs(3747) <= not a;
    layer4_outputs(3748) <= a;
    layer4_outputs(3749) <= not (a xor b);
    layer4_outputs(3750) <= not (a or b);
    layer4_outputs(3751) <= not (a xor b);
    layer4_outputs(3752) <= b;
    layer4_outputs(3753) <= a or b;
    layer4_outputs(3754) <= a and not b;
    layer4_outputs(3755) <= a and not b;
    layer4_outputs(3756) <= a xor b;
    layer4_outputs(3757) <= b;
    layer4_outputs(3758) <= not (a and b);
    layer4_outputs(3759) <= not (a and b);
    layer4_outputs(3760) <= '1';
    layer4_outputs(3761) <= not b or a;
    layer4_outputs(3762) <= not a or b;
    layer4_outputs(3763) <= b;
    layer4_outputs(3764) <= b;
    layer4_outputs(3765) <= a and b;
    layer4_outputs(3766) <= not a or b;
    layer4_outputs(3767) <= b;
    layer4_outputs(3768) <= not b or a;
    layer4_outputs(3769) <= not (a or b);
    layer4_outputs(3770) <= b;
    layer4_outputs(3771) <= b;
    layer4_outputs(3772) <= not b;
    layer4_outputs(3773) <= not a or b;
    layer4_outputs(3774) <= a or b;
    layer4_outputs(3775) <= not a;
    layer4_outputs(3776) <= not a or b;
    layer4_outputs(3777) <= not b;
    layer4_outputs(3778) <= not a;
    layer4_outputs(3779) <= a;
    layer4_outputs(3780) <= a xor b;
    layer4_outputs(3781) <= not (a xor b);
    layer4_outputs(3782) <= '1';
    layer4_outputs(3783) <= b;
    layer4_outputs(3784) <= a;
    layer4_outputs(3785) <= not a or b;
    layer4_outputs(3786) <= not a;
    layer4_outputs(3787) <= not (a xor b);
    layer4_outputs(3788) <= not a;
    layer4_outputs(3789) <= '0';
    layer4_outputs(3790) <= b;
    layer4_outputs(3791) <= a and not b;
    layer4_outputs(3792) <= b;
    layer4_outputs(3793) <= not (a or b);
    layer4_outputs(3794) <= '1';
    layer4_outputs(3795) <= not b;
    layer4_outputs(3796) <= not b;
    layer4_outputs(3797) <= not (a or b);
    layer4_outputs(3798) <= a and not b;
    layer4_outputs(3799) <= not (a and b);
    layer4_outputs(3800) <= not (a xor b);
    layer4_outputs(3801) <= a;
    layer4_outputs(3802) <= not a;
    layer4_outputs(3803) <= not b;
    layer4_outputs(3804) <= not b;
    layer4_outputs(3805) <= not a or b;
    layer4_outputs(3806) <= a;
    layer4_outputs(3807) <= b and not a;
    layer4_outputs(3808) <= b;
    layer4_outputs(3809) <= b;
    layer4_outputs(3810) <= not (a and b);
    layer4_outputs(3811) <= not a;
    layer4_outputs(3812) <= a xor b;
    layer4_outputs(3813) <= a or b;
    layer4_outputs(3814) <= a;
    layer4_outputs(3815) <= not a or b;
    layer4_outputs(3816) <= b and not a;
    layer4_outputs(3817) <= '1';
    layer4_outputs(3818) <= '0';
    layer4_outputs(3819) <= not (a xor b);
    layer4_outputs(3820) <= a;
    layer4_outputs(3821) <= b;
    layer4_outputs(3822) <= a and b;
    layer4_outputs(3823) <= a;
    layer4_outputs(3824) <= a;
    layer4_outputs(3825) <= not a or b;
    layer4_outputs(3826) <= a;
    layer4_outputs(3827) <= not a or b;
    layer4_outputs(3828) <= not b or a;
    layer4_outputs(3829) <= a or b;
    layer4_outputs(3830) <= not (a and b);
    layer4_outputs(3831) <= b;
    layer4_outputs(3832) <= not (a xor b);
    layer4_outputs(3833) <= not b;
    layer4_outputs(3834) <= b;
    layer4_outputs(3835) <= a xor b;
    layer4_outputs(3836) <= not (a or b);
    layer4_outputs(3837) <= not a;
    layer4_outputs(3838) <= not b or a;
    layer4_outputs(3839) <= not (a or b);
    layer4_outputs(3840) <= not b;
    layer4_outputs(3841) <= '1';
    layer4_outputs(3842) <= not (a or b);
    layer4_outputs(3843) <= a and b;
    layer4_outputs(3844) <= not (a or b);
    layer4_outputs(3845) <= a or b;
    layer4_outputs(3846) <= not a;
    layer4_outputs(3847) <= '0';
    layer4_outputs(3848) <= not (a or b);
    layer4_outputs(3849) <= not (a or b);
    layer4_outputs(3850) <= not (a or b);
    layer4_outputs(3851) <= a or b;
    layer4_outputs(3852) <= b and not a;
    layer4_outputs(3853) <= not b;
    layer4_outputs(3854) <= '0';
    layer4_outputs(3855) <= '1';
    layer4_outputs(3856) <= not a;
    layer4_outputs(3857) <= a and not b;
    layer4_outputs(3858) <= not (a and b);
    layer4_outputs(3859) <= not a;
    layer4_outputs(3860) <= not (a and b);
    layer4_outputs(3861) <= not a or b;
    layer4_outputs(3862) <= not b;
    layer4_outputs(3863) <= a and b;
    layer4_outputs(3864) <= not b;
    layer4_outputs(3865) <= a xor b;
    layer4_outputs(3866) <= not a;
    layer4_outputs(3867) <= not b or a;
    layer4_outputs(3868) <= not a;
    layer4_outputs(3869) <= a or b;
    layer4_outputs(3870) <= a and not b;
    layer4_outputs(3871) <= a;
    layer4_outputs(3872) <= not a or b;
    layer4_outputs(3873) <= a;
    layer4_outputs(3874) <= not a;
    layer4_outputs(3875) <= not (a or b);
    layer4_outputs(3876) <= not (a or b);
    layer4_outputs(3877) <= a and b;
    layer4_outputs(3878) <= a;
    layer4_outputs(3879) <= a and not b;
    layer4_outputs(3880) <= a;
    layer4_outputs(3881) <= a and not b;
    layer4_outputs(3882) <= a or b;
    layer4_outputs(3883) <= b;
    layer4_outputs(3884) <= not (a or b);
    layer4_outputs(3885) <= b;
    layer4_outputs(3886) <= a and not b;
    layer4_outputs(3887) <= not b;
    layer4_outputs(3888) <= a;
    layer4_outputs(3889) <= b;
    layer4_outputs(3890) <= not (a and b);
    layer4_outputs(3891) <= not b;
    layer4_outputs(3892) <= not (a xor b);
    layer4_outputs(3893) <= b;
    layer4_outputs(3894) <= not (a or b);
    layer4_outputs(3895) <= b;
    layer4_outputs(3896) <= a and b;
    layer4_outputs(3897) <= '0';
    layer4_outputs(3898) <= not a;
    layer4_outputs(3899) <= not b;
    layer4_outputs(3900) <= not b;
    layer4_outputs(3901) <= not a or b;
    layer4_outputs(3902) <= a or b;
    layer4_outputs(3903) <= not a;
    layer4_outputs(3904) <= a;
    layer4_outputs(3905) <= not (a or b);
    layer4_outputs(3906) <= b and not a;
    layer4_outputs(3907) <= not b;
    layer4_outputs(3908) <= a;
    layer4_outputs(3909) <= not b;
    layer4_outputs(3910) <= b;
    layer4_outputs(3911) <= a;
    layer4_outputs(3912) <= not b or a;
    layer4_outputs(3913) <= b;
    layer4_outputs(3914) <= not a;
    layer4_outputs(3915) <= a;
    layer4_outputs(3916) <= b;
    layer4_outputs(3917) <= not (a xor b);
    layer4_outputs(3918) <= not (a and b);
    layer4_outputs(3919) <= not (a xor b);
    layer4_outputs(3920) <= a;
    layer4_outputs(3921) <= not (a and b);
    layer4_outputs(3922) <= not a;
    layer4_outputs(3923) <= a and b;
    layer4_outputs(3924) <= not (a and b);
    layer4_outputs(3925) <= '1';
    layer4_outputs(3926) <= b;
    layer4_outputs(3927) <= not a or b;
    layer4_outputs(3928) <= a and b;
    layer4_outputs(3929) <= a and not b;
    layer4_outputs(3930) <= a and b;
    layer4_outputs(3931) <= a and b;
    layer4_outputs(3932) <= not (a and b);
    layer4_outputs(3933) <= a and not b;
    layer4_outputs(3934) <= not (a and b);
    layer4_outputs(3935) <= b;
    layer4_outputs(3936) <= not (a and b);
    layer4_outputs(3937) <= not b;
    layer4_outputs(3938) <= not a;
    layer4_outputs(3939) <= not (a xor b);
    layer4_outputs(3940) <= a or b;
    layer4_outputs(3941) <= not b;
    layer4_outputs(3942) <= a;
    layer4_outputs(3943) <= not b;
    layer4_outputs(3944) <= a and not b;
    layer4_outputs(3945) <= b;
    layer4_outputs(3946) <= not a;
    layer4_outputs(3947) <= not b;
    layer4_outputs(3948) <= not b or a;
    layer4_outputs(3949) <= a;
    layer4_outputs(3950) <= not a;
    layer4_outputs(3951) <= a and b;
    layer4_outputs(3952) <= a;
    layer4_outputs(3953) <= b and not a;
    layer4_outputs(3954) <= not b;
    layer4_outputs(3955) <= not (a and b);
    layer4_outputs(3956) <= not (a and b);
    layer4_outputs(3957) <= b;
    layer4_outputs(3958) <= a xor b;
    layer4_outputs(3959) <= not (a xor b);
    layer4_outputs(3960) <= not (a or b);
    layer4_outputs(3961) <= not a;
    layer4_outputs(3962) <= a;
    layer4_outputs(3963) <= not b;
    layer4_outputs(3964) <= a or b;
    layer4_outputs(3965) <= a;
    layer4_outputs(3966) <= not b;
    layer4_outputs(3967) <= b;
    layer4_outputs(3968) <= not b or a;
    layer4_outputs(3969) <= b and not a;
    layer4_outputs(3970) <= a or b;
    layer4_outputs(3971) <= a;
    layer4_outputs(3972) <= not b;
    layer4_outputs(3973) <= not (a xor b);
    layer4_outputs(3974) <= not (a xor b);
    layer4_outputs(3975) <= not b or a;
    layer4_outputs(3976) <= a and not b;
    layer4_outputs(3977) <= a and not b;
    layer4_outputs(3978) <= a and not b;
    layer4_outputs(3979) <= a or b;
    layer4_outputs(3980) <= not b or a;
    layer4_outputs(3981) <= not a;
    layer4_outputs(3982) <= a;
    layer4_outputs(3983) <= not a;
    layer4_outputs(3984) <= a and b;
    layer4_outputs(3985) <= not b or a;
    layer4_outputs(3986) <= not a;
    layer4_outputs(3987) <= b;
    layer4_outputs(3988) <= not a;
    layer4_outputs(3989) <= a xor b;
    layer4_outputs(3990) <= not b;
    layer4_outputs(3991) <= not a;
    layer4_outputs(3992) <= not b;
    layer4_outputs(3993) <= a;
    layer4_outputs(3994) <= a;
    layer4_outputs(3995) <= a;
    layer4_outputs(3996) <= not b;
    layer4_outputs(3997) <= b and not a;
    layer4_outputs(3998) <= not b or a;
    layer4_outputs(3999) <= b and not a;
    layer4_outputs(4000) <= a;
    layer4_outputs(4001) <= '1';
    layer4_outputs(4002) <= a;
    layer4_outputs(4003) <= b;
    layer4_outputs(4004) <= a or b;
    layer4_outputs(4005) <= not b or a;
    layer4_outputs(4006) <= not (a and b);
    layer4_outputs(4007) <= '1';
    layer4_outputs(4008) <= a or b;
    layer4_outputs(4009) <= not a or b;
    layer4_outputs(4010) <= a and not b;
    layer4_outputs(4011) <= not b or a;
    layer4_outputs(4012) <= a or b;
    layer4_outputs(4013) <= a and not b;
    layer4_outputs(4014) <= not (a and b);
    layer4_outputs(4015) <= '0';
    layer4_outputs(4016) <= not b or a;
    layer4_outputs(4017) <= b;
    layer4_outputs(4018) <= not b;
    layer4_outputs(4019) <= not a or b;
    layer4_outputs(4020) <= not a;
    layer4_outputs(4021) <= a and b;
    layer4_outputs(4022) <= not (a and b);
    layer4_outputs(4023) <= b and not a;
    layer4_outputs(4024) <= not b;
    layer4_outputs(4025) <= not (a or b);
    layer4_outputs(4026) <= a;
    layer4_outputs(4027) <= b and not a;
    layer4_outputs(4028) <= a or b;
    layer4_outputs(4029) <= not a;
    layer4_outputs(4030) <= not (a or b);
    layer4_outputs(4031) <= not (a and b);
    layer4_outputs(4032) <= not (a or b);
    layer4_outputs(4033) <= not (a or b);
    layer4_outputs(4034) <= '1';
    layer4_outputs(4035) <= b;
    layer4_outputs(4036) <= not (a or b);
    layer4_outputs(4037) <= not (a xor b);
    layer4_outputs(4038) <= a xor b;
    layer4_outputs(4039) <= not a or b;
    layer4_outputs(4040) <= a and b;
    layer4_outputs(4041) <= not a or b;
    layer4_outputs(4042) <= b;
    layer4_outputs(4043) <= not b;
    layer4_outputs(4044) <= not (a or b);
    layer4_outputs(4045) <= a xor b;
    layer4_outputs(4046) <= not a or b;
    layer4_outputs(4047) <= not a;
    layer4_outputs(4048) <= not (a or b);
    layer4_outputs(4049) <= not b;
    layer4_outputs(4050) <= not b or a;
    layer4_outputs(4051) <= a or b;
    layer4_outputs(4052) <= b;
    layer4_outputs(4053) <= not (a or b);
    layer4_outputs(4054) <= not a or b;
    layer4_outputs(4055) <= a;
    layer4_outputs(4056) <= not b;
    layer4_outputs(4057) <= a or b;
    layer4_outputs(4058) <= b;
    layer4_outputs(4059) <= not b;
    layer4_outputs(4060) <= '0';
    layer4_outputs(4061) <= a;
    layer4_outputs(4062) <= a xor b;
    layer4_outputs(4063) <= a or b;
    layer4_outputs(4064) <= not (a and b);
    layer4_outputs(4065) <= not (a xor b);
    layer4_outputs(4066) <= not a or b;
    layer4_outputs(4067) <= not b;
    layer4_outputs(4068) <= not a;
    layer4_outputs(4069) <= not (a or b);
    layer4_outputs(4070) <= a and not b;
    layer4_outputs(4071) <= not b;
    layer4_outputs(4072) <= b;
    layer4_outputs(4073) <= not (a xor b);
    layer4_outputs(4074) <= not a;
    layer4_outputs(4075) <= b;
    layer4_outputs(4076) <= b;
    layer4_outputs(4077) <= not b;
    layer4_outputs(4078) <= b and not a;
    layer4_outputs(4079) <= not a;
    layer4_outputs(4080) <= not (a and b);
    layer4_outputs(4081) <= b;
    layer4_outputs(4082) <= not a or b;
    layer4_outputs(4083) <= not b or a;
    layer4_outputs(4084) <= not (a xor b);
    layer4_outputs(4085) <= a and b;
    layer4_outputs(4086) <= not b;
    layer4_outputs(4087) <= '0';
    layer4_outputs(4088) <= b and not a;
    layer4_outputs(4089) <= not (a xor b);
    layer4_outputs(4090) <= a;
    layer4_outputs(4091) <= '1';
    layer4_outputs(4092) <= not b;
    layer4_outputs(4093) <= not (a or b);
    layer4_outputs(4094) <= not b;
    layer4_outputs(4095) <= a and b;
    layer4_outputs(4096) <= not b;
    layer4_outputs(4097) <= a and not b;
    layer4_outputs(4098) <= a or b;
    layer4_outputs(4099) <= '1';
    layer4_outputs(4100) <= a and b;
    layer4_outputs(4101) <= not (a xor b);
    layer4_outputs(4102) <= not a or b;
    layer4_outputs(4103) <= a and b;
    layer4_outputs(4104) <= not (a and b);
    layer4_outputs(4105) <= a;
    layer4_outputs(4106) <= b;
    layer4_outputs(4107) <= b;
    layer4_outputs(4108) <= a and not b;
    layer4_outputs(4109) <= b and not a;
    layer4_outputs(4110) <= a and b;
    layer4_outputs(4111) <= '1';
    layer4_outputs(4112) <= a;
    layer4_outputs(4113) <= b and not a;
    layer4_outputs(4114) <= b and not a;
    layer4_outputs(4115) <= a;
    layer4_outputs(4116) <= not (a and b);
    layer4_outputs(4117) <= not a;
    layer4_outputs(4118) <= b and not a;
    layer4_outputs(4119) <= not a;
    layer4_outputs(4120) <= a;
    layer4_outputs(4121) <= a;
    layer4_outputs(4122) <= a and b;
    layer4_outputs(4123) <= not b;
    layer4_outputs(4124) <= not (a xor b);
    layer4_outputs(4125) <= not a or b;
    layer4_outputs(4126) <= a;
    layer4_outputs(4127) <= not (a or b);
    layer4_outputs(4128) <= not a;
    layer4_outputs(4129) <= b;
    layer4_outputs(4130) <= '1';
    layer4_outputs(4131) <= a and not b;
    layer4_outputs(4132) <= not a or b;
    layer4_outputs(4133) <= a and b;
    layer4_outputs(4134) <= not b or a;
    layer4_outputs(4135) <= not a or b;
    layer4_outputs(4136) <= a and not b;
    layer4_outputs(4137) <= not (a xor b);
    layer4_outputs(4138) <= b and not a;
    layer4_outputs(4139) <= not (a xor b);
    layer4_outputs(4140) <= not b;
    layer4_outputs(4141) <= not (a and b);
    layer4_outputs(4142) <= b;
    layer4_outputs(4143) <= a;
    layer4_outputs(4144) <= b;
    layer4_outputs(4145) <= a;
    layer4_outputs(4146) <= a;
    layer4_outputs(4147) <= not b or a;
    layer4_outputs(4148) <= b;
    layer4_outputs(4149) <= b and not a;
    layer4_outputs(4150) <= not a;
    layer4_outputs(4151) <= not a;
    layer4_outputs(4152) <= '1';
    layer4_outputs(4153) <= a;
    layer4_outputs(4154) <= '1';
    layer4_outputs(4155) <= b;
    layer4_outputs(4156) <= a;
    layer4_outputs(4157) <= a;
    layer4_outputs(4158) <= not a;
    layer4_outputs(4159) <= a and b;
    layer4_outputs(4160) <= not b;
    layer4_outputs(4161) <= not a or b;
    layer4_outputs(4162) <= not (a and b);
    layer4_outputs(4163) <= not b;
    layer4_outputs(4164) <= not b;
    layer4_outputs(4165) <= b;
    layer4_outputs(4166) <= a and b;
    layer4_outputs(4167) <= not a or b;
    layer4_outputs(4168) <= '0';
    layer4_outputs(4169) <= b;
    layer4_outputs(4170) <= not b;
    layer4_outputs(4171) <= b;
    layer4_outputs(4172) <= b and not a;
    layer4_outputs(4173) <= a;
    layer4_outputs(4174) <= a or b;
    layer4_outputs(4175) <= not b;
    layer4_outputs(4176) <= b and not a;
    layer4_outputs(4177) <= '1';
    layer4_outputs(4178) <= not b;
    layer4_outputs(4179) <= a and b;
    layer4_outputs(4180) <= b;
    layer4_outputs(4181) <= b;
    layer4_outputs(4182) <= a;
    layer4_outputs(4183) <= not a;
    layer4_outputs(4184) <= not (a or b);
    layer4_outputs(4185) <= not b;
    layer4_outputs(4186) <= a;
    layer4_outputs(4187) <= a or b;
    layer4_outputs(4188) <= a and b;
    layer4_outputs(4189) <= not b;
    layer4_outputs(4190) <= a and b;
    layer4_outputs(4191) <= '1';
    layer4_outputs(4192) <= a;
    layer4_outputs(4193) <= a;
    layer4_outputs(4194) <= a and not b;
    layer4_outputs(4195) <= not b;
    layer4_outputs(4196) <= not b;
    layer4_outputs(4197) <= a xor b;
    layer4_outputs(4198) <= a and b;
    layer4_outputs(4199) <= b;
    layer4_outputs(4200) <= a and b;
    layer4_outputs(4201) <= a;
    layer4_outputs(4202) <= not a or b;
    layer4_outputs(4203) <= b and not a;
    layer4_outputs(4204) <= a xor b;
    layer4_outputs(4205) <= b;
    layer4_outputs(4206) <= a;
    layer4_outputs(4207) <= not b or a;
    layer4_outputs(4208) <= a xor b;
    layer4_outputs(4209) <= not (a xor b);
    layer4_outputs(4210) <= a;
    layer4_outputs(4211) <= not b or a;
    layer4_outputs(4212) <= b and not a;
    layer4_outputs(4213) <= not a;
    layer4_outputs(4214) <= not a;
    layer4_outputs(4215) <= a and not b;
    layer4_outputs(4216) <= not a;
    layer4_outputs(4217) <= '1';
    layer4_outputs(4218) <= a xor b;
    layer4_outputs(4219) <= not b;
    layer4_outputs(4220) <= b;
    layer4_outputs(4221) <= b;
    layer4_outputs(4222) <= not b;
    layer4_outputs(4223) <= not b or a;
    layer4_outputs(4224) <= b and not a;
    layer4_outputs(4225) <= b and not a;
    layer4_outputs(4226) <= b;
    layer4_outputs(4227) <= '0';
    layer4_outputs(4228) <= a or b;
    layer4_outputs(4229) <= not b;
    layer4_outputs(4230) <= not b;
    layer4_outputs(4231) <= not (a or b);
    layer4_outputs(4232) <= b;
    layer4_outputs(4233) <= not (a xor b);
    layer4_outputs(4234) <= a;
    layer4_outputs(4235) <= b;
    layer4_outputs(4236) <= a and not b;
    layer4_outputs(4237) <= not a or b;
    layer4_outputs(4238) <= not (a or b);
    layer4_outputs(4239) <= b and not a;
    layer4_outputs(4240) <= b;
    layer4_outputs(4241) <= b;
    layer4_outputs(4242) <= a and not b;
    layer4_outputs(4243) <= not b;
    layer4_outputs(4244) <= a;
    layer4_outputs(4245) <= not a;
    layer4_outputs(4246) <= not (a and b);
    layer4_outputs(4247) <= not (a xor b);
    layer4_outputs(4248) <= a xor b;
    layer4_outputs(4249) <= a;
    layer4_outputs(4250) <= not (a or b);
    layer4_outputs(4251) <= a and b;
    layer4_outputs(4252) <= a;
    layer4_outputs(4253) <= not (a or b);
    layer4_outputs(4254) <= b and not a;
    layer4_outputs(4255) <= a or b;
    layer4_outputs(4256) <= a or b;
    layer4_outputs(4257) <= not b;
    layer4_outputs(4258) <= a or b;
    layer4_outputs(4259) <= not a;
    layer4_outputs(4260) <= not a;
    layer4_outputs(4261) <= a and not b;
    layer4_outputs(4262) <= a;
    layer4_outputs(4263) <= not (a xor b);
    layer4_outputs(4264) <= not a;
    layer4_outputs(4265) <= a and not b;
    layer4_outputs(4266) <= not a;
    layer4_outputs(4267) <= not b or a;
    layer4_outputs(4268) <= not b;
    layer4_outputs(4269) <= a;
    layer4_outputs(4270) <= not (a or b);
    layer4_outputs(4271) <= a and b;
    layer4_outputs(4272) <= b;
    layer4_outputs(4273) <= a and b;
    layer4_outputs(4274) <= a or b;
    layer4_outputs(4275) <= not a or b;
    layer4_outputs(4276) <= a xor b;
    layer4_outputs(4277) <= b;
    layer4_outputs(4278) <= a;
    layer4_outputs(4279) <= b and not a;
    layer4_outputs(4280) <= not a or b;
    layer4_outputs(4281) <= a;
    layer4_outputs(4282) <= '1';
    layer4_outputs(4283) <= not a or b;
    layer4_outputs(4284) <= '1';
    layer4_outputs(4285) <= a or b;
    layer4_outputs(4286) <= a;
    layer4_outputs(4287) <= b;
    layer4_outputs(4288) <= a;
    layer4_outputs(4289) <= a xor b;
    layer4_outputs(4290) <= a xor b;
    layer4_outputs(4291) <= a and b;
    layer4_outputs(4292) <= not (a and b);
    layer4_outputs(4293) <= not (a xor b);
    layer4_outputs(4294) <= b;
    layer4_outputs(4295) <= b and not a;
    layer4_outputs(4296) <= not (a and b);
    layer4_outputs(4297) <= a and b;
    layer4_outputs(4298) <= a;
    layer4_outputs(4299) <= not b;
    layer4_outputs(4300) <= not a;
    layer4_outputs(4301) <= a xor b;
    layer4_outputs(4302) <= a and not b;
    layer4_outputs(4303) <= a or b;
    layer4_outputs(4304) <= not b or a;
    layer4_outputs(4305) <= b and not a;
    layer4_outputs(4306) <= not a;
    layer4_outputs(4307) <= not a;
    layer4_outputs(4308) <= b and not a;
    layer4_outputs(4309) <= not a;
    layer4_outputs(4310) <= b;
    layer4_outputs(4311) <= b;
    layer4_outputs(4312) <= a and b;
    layer4_outputs(4313) <= a or b;
    layer4_outputs(4314) <= not b;
    layer4_outputs(4315) <= not a or b;
    layer4_outputs(4316) <= a and b;
    layer4_outputs(4317) <= a xor b;
    layer4_outputs(4318) <= not (a or b);
    layer4_outputs(4319) <= not b;
    layer4_outputs(4320) <= not a;
    layer4_outputs(4321) <= b;
    layer4_outputs(4322) <= not (a or b);
    layer4_outputs(4323) <= a or b;
    layer4_outputs(4324) <= a;
    layer4_outputs(4325) <= a or b;
    layer4_outputs(4326) <= a or b;
    layer4_outputs(4327) <= not a;
    layer4_outputs(4328) <= not b;
    layer4_outputs(4329) <= '1';
    layer4_outputs(4330) <= a;
    layer4_outputs(4331) <= not (a xor b);
    layer4_outputs(4332) <= not b;
    layer4_outputs(4333) <= b;
    layer4_outputs(4334) <= a and not b;
    layer4_outputs(4335) <= b;
    layer4_outputs(4336) <= not a;
    layer4_outputs(4337) <= not b;
    layer4_outputs(4338) <= b;
    layer4_outputs(4339) <= a or b;
    layer4_outputs(4340) <= a;
    layer4_outputs(4341) <= a and b;
    layer4_outputs(4342) <= not (a xor b);
    layer4_outputs(4343) <= a;
    layer4_outputs(4344) <= a and b;
    layer4_outputs(4345) <= not (a and b);
    layer4_outputs(4346) <= a and b;
    layer4_outputs(4347) <= b;
    layer4_outputs(4348) <= a xor b;
    layer4_outputs(4349) <= not b;
    layer4_outputs(4350) <= a;
    layer4_outputs(4351) <= not a;
    layer4_outputs(4352) <= not (a and b);
    layer4_outputs(4353) <= b;
    layer4_outputs(4354) <= not a;
    layer4_outputs(4355) <= not b or a;
    layer4_outputs(4356) <= b;
    layer4_outputs(4357) <= b;
    layer4_outputs(4358) <= a;
    layer4_outputs(4359) <= a or b;
    layer4_outputs(4360) <= not (a xor b);
    layer4_outputs(4361) <= a and b;
    layer4_outputs(4362) <= a;
    layer4_outputs(4363) <= a;
    layer4_outputs(4364) <= not b or a;
    layer4_outputs(4365) <= not (a xor b);
    layer4_outputs(4366) <= a;
    layer4_outputs(4367) <= '0';
    layer4_outputs(4368) <= a;
    layer4_outputs(4369) <= not b;
    layer4_outputs(4370) <= not a or b;
    layer4_outputs(4371) <= a xor b;
    layer4_outputs(4372) <= not (a or b);
    layer4_outputs(4373) <= not (a xor b);
    layer4_outputs(4374) <= a xor b;
    layer4_outputs(4375) <= not b or a;
    layer4_outputs(4376) <= not b;
    layer4_outputs(4377) <= b;
    layer4_outputs(4378) <= not a;
    layer4_outputs(4379) <= not b or a;
    layer4_outputs(4380) <= a;
    layer4_outputs(4381) <= a;
    layer4_outputs(4382) <= not a;
    layer4_outputs(4383) <= not a;
    layer4_outputs(4384) <= not b;
    layer4_outputs(4385) <= not a;
    layer4_outputs(4386) <= b and not a;
    layer4_outputs(4387) <= a and not b;
    layer4_outputs(4388) <= not (a and b);
    layer4_outputs(4389) <= a;
    layer4_outputs(4390) <= not b or a;
    layer4_outputs(4391) <= b;
    layer4_outputs(4392) <= not (a or b);
    layer4_outputs(4393) <= not b;
    layer4_outputs(4394) <= not (a or b);
    layer4_outputs(4395) <= a;
    layer4_outputs(4396) <= not (a and b);
    layer4_outputs(4397) <= '1';
    layer4_outputs(4398) <= not a;
    layer4_outputs(4399) <= not b or a;
    layer4_outputs(4400) <= a and not b;
    layer4_outputs(4401) <= not b or a;
    layer4_outputs(4402) <= not b;
    layer4_outputs(4403) <= b and not a;
    layer4_outputs(4404) <= a and not b;
    layer4_outputs(4405) <= not a;
    layer4_outputs(4406) <= not (a and b);
    layer4_outputs(4407) <= not (a and b);
    layer4_outputs(4408) <= not a or b;
    layer4_outputs(4409) <= a or b;
    layer4_outputs(4410) <= not (a and b);
    layer4_outputs(4411) <= not b;
    layer4_outputs(4412) <= a;
    layer4_outputs(4413) <= not b;
    layer4_outputs(4414) <= not a or b;
    layer4_outputs(4415) <= not (a and b);
    layer4_outputs(4416) <= b;
    layer4_outputs(4417) <= b;
    layer4_outputs(4418) <= not (a and b);
    layer4_outputs(4419) <= not b;
    layer4_outputs(4420) <= not b;
    layer4_outputs(4421) <= b;
    layer4_outputs(4422) <= a xor b;
    layer4_outputs(4423) <= not a;
    layer4_outputs(4424) <= a and b;
    layer4_outputs(4425) <= not b;
    layer4_outputs(4426) <= '1';
    layer4_outputs(4427) <= not b or a;
    layer4_outputs(4428) <= not (a or b);
    layer4_outputs(4429) <= not a;
    layer4_outputs(4430) <= b;
    layer4_outputs(4431) <= not a;
    layer4_outputs(4432) <= not a or b;
    layer4_outputs(4433) <= not (a and b);
    layer4_outputs(4434) <= a;
    layer4_outputs(4435) <= not b or a;
    layer4_outputs(4436) <= not (a and b);
    layer4_outputs(4437) <= a and b;
    layer4_outputs(4438) <= a;
    layer4_outputs(4439) <= a;
    layer4_outputs(4440) <= not (a xor b);
    layer4_outputs(4441) <= not a or b;
    layer4_outputs(4442) <= not b or a;
    layer4_outputs(4443) <= a;
    layer4_outputs(4444) <= b and not a;
    layer4_outputs(4445) <= not a;
    layer4_outputs(4446) <= '1';
    layer4_outputs(4447) <= not (a or b);
    layer4_outputs(4448) <= not a or b;
    layer4_outputs(4449) <= a and b;
    layer4_outputs(4450) <= not (a and b);
    layer4_outputs(4451) <= b;
    layer4_outputs(4452) <= not b or a;
    layer4_outputs(4453) <= a and b;
    layer4_outputs(4454) <= not b;
    layer4_outputs(4455) <= not a;
    layer4_outputs(4456) <= a;
    layer4_outputs(4457) <= a and not b;
    layer4_outputs(4458) <= not (a xor b);
    layer4_outputs(4459) <= not (a xor b);
    layer4_outputs(4460) <= b;
    layer4_outputs(4461) <= b and not a;
    layer4_outputs(4462) <= not (a xor b);
    layer4_outputs(4463) <= not a;
    layer4_outputs(4464) <= not b;
    layer4_outputs(4465) <= '1';
    layer4_outputs(4466) <= not (a and b);
    layer4_outputs(4467) <= not (a xor b);
    layer4_outputs(4468) <= a and b;
    layer4_outputs(4469) <= a and b;
    layer4_outputs(4470) <= not b;
    layer4_outputs(4471) <= not (a and b);
    layer4_outputs(4472) <= not (a and b);
    layer4_outputs(4473) <= not a or b;
    layer4_outputs(4474) <= not b or a;
    layer4_outputs(4475) <= a xor b;
    layer4_outputs(4476) <= a or b;
    layer4_outputs(4477) <= b and not a;
    layer4_outputs(4478) <= not a or b;
    layer4_outputs(4479) <= a and not b;
    layer4_outputs(4480) <= not b or a;
    layer4_outputs(4481) <= not (a and b);
    layer4_outputs(4482) <= a and not b;
    layer4_outputs(4483) <= not a;
    layer4_outputs(4484) <= a;
    layer4_outputs(4485) <= not (a and b);
    layer4_outputs(4486) <= '0';
    layer4_outputs(4487) <= a;
    layer4_outputs(4488) <= not (a xor b);
    layer4_outputs(4489) <= not b;
    layer4_outputs(4490) <= not a or b;
    layer4_outputs(4491) <= '1';
    layer4_outputs(4492) <= '0';
    layer4_outputs(4493) <= a and b;
    layer4_outputs(4494) <= '1';
    layer4_outputs(4495) <= a;
    layer4_outputs(4496) <= a or b;
    layer4_outputs(4497) <= '0';
    layer4_outputs(4498) <= b;
    layer4_outputs(4499) <= b;
    layer4_outputs(4500) <= b;
    layer4_outputs(4501) <= not a or b;
    layer4_outputs(4502) <= '0';
    layer4_outputs(4503) <= not b or a;
    layer4_outputs(4504) <= not a;
    layer4_outputs(4505) <= a and b;
    layer4_outputs(4506) <= not (a and b);
    layer4_outputs(4507) <= not (a xor b);
    layer4_outputs(4508) <= a and not b;
    layer4_outputs(4509) <= not a or b;
    layer4_outputs(4510) <= a and b;
    layer4_outputs(4511) <= not b or a;
    layer4_outputs(4512) <= a xor b;
    layer4_outputs(4513) <= b and not a;
    layer4_outputs(4514) <= not a or b;
    layer4_outputs(4515) <= a xor b;
    layer4_outputs(4516) <= not a;
    layer4_outputs(4517) <= a or b;
    layer4_outputs(4518) <= not b or a;
    layer4_outputs(4519) <= not a;
    layer4_outputs(4520) <= not b or a;
    layer4_outputs(4521) <= b;
    layer4_outputs(4522) <= not (a and b);
    layer4_outputs(4523) <= b;
    layer4_outputs(4524) <= '1';
    layer4_outputs(4525) <= a and not b;
    layer4_outputs(4526) <= a and b;
    layer4_outputs(4527) <= not b or a;
    layer4_outputs(4528) <= a xor b;
    layer4_outputs(4529) <= not (a xor b);
    layer4_outputs(4530) <= not a;
    layer4_outputs(4531) <= not (a and b);
    layer4_outputs(4532) <= a xor b;
    layer4_outputs(4533) <= a;
    layer4_outputs(4534) <= a;
    layer4_outputs(4535) <= not b;
    layer4_outputs(4536) <= b;
    layer4_outputs(4537) <= not a;
    layer4_outputs(4538) <= a or b;
    layer4_outputs(4539) <= not a;
    layer4_outputs(4540) <= not a or b;
    layer4_outputs(4541) <= b;
    layer4_outputs(4542) <= b;
    layer4_outputs(4543) <= not a;
    layer4_outputs(4544) <= b and not a;
    layer4_outputs(4545) <= '0';
    layer4_outputs(4546) <= not b or a;
    layer4_outputs(4547) <= b and not a;
    layer4_outputs(4548) <= not b or a;
    layer4_outputs(4549) <= not a;
    layer4_outputs(4550) <= b;
    layer4_outputs(4551) <= not (a or b);
    layer4_outputs(4552) <= a;
    layer4_outputs(4553) <= b;
    layer4_outputs(4554) <= a and b;
    layer4_outputs(4555) <= not (a xor b);
    layer4_outputs(4556) <= not b;
    layer4_outputs(4557) <= b;
    layer4_outputs(4558) <= not b or a;
    layer4_outputs(4559) <= not (a and b);
    layer4_outputs(4560) <= not (a and b);
    layer4_outputs(4561) <= '1';
    layer4_outputs(4562) <= a;
    layer4_outputs(4563) <= not (a xor b);
    layer4_outputs(4564) <= not b or a;
    layer4_outputs(4565) <= b and not a;
    layer4_outputs(4566) <= '0';
    layer4_outputs(4567) <= b and not a;
    layer4_outputs(4568) <= a and not b;
    layer4_outputs(4569) <= a and b;
    layer4_outputs(4570) <= b;
    layer4_outputs(4571) <= not b or a;
    layer4_outputs(4572) <= b;
    layer4_outputs(4573) <= not a;
    layer4_outputs(4574) <= not a or b;
    layer4_outputs(4575) <= not a or b;
    layer4_outputs(4576) <= a and not b;
    layer4_outputs(4577) <= a xor b;
    layer4_outputs(4578) <= not (a and b);
    layer4_outputs(4579) <= not b;
    layer4_outputs(4580) <= a and not b;
    layer4_outputs(4581) <= not a;
    layer4_outputs(4582) <= not (a or b);
    layer4_outputs(4583) <= a;
    layer4_outputs(4584) <= a;
    layer4_outputs(4585) <= not (a and b);
    layer4_outputs(4586) <= b;
    layer4_outputs(4587) <= a;
    layer4_outputs(4588) <= not a;
    layer4_outputs(4589) <= a;
    layer4_outputs(4590) <= not b;
    layer4_outputs(4591) <= not b;
    layer4_outputs(4592) <= not (a or b);
    layer4_outputs(4593) <= not (a and b);
    layer4_outputs(4594) <= a and b;
    layer4_outputs(4595) <= a and b;
    layer4_outputs(4596) <= b and not a;
    layer4_outputs(4597) <= not a or b;
    layer4_outputs(4598) <= not a;
    layer4_outputs(4599) <= not b;
    layer4_outputs(4600) <= a;
    layer4_outputs(4601) <= not b;
    layer4_outputs(4602) <= not a or b;
    layer4_outputs(4603) <= a;
    layer4_outputs(4604) <= not a;
    layer4_outputs(4605) <= a or b;
    layer4_outputs(4606) <= b;
    layer4_outputs(4607) <= b and not a;
    layer4_outputs(4608) <= not a or b;
    layer4_outputs(4609) <= a xor b;
    layer4_outputs(4610) <= not a;
    layer4_outputs(4611) <= b;
    layer4_outputs(4612) <= not b or a;
    layer4_outputs(4613) <= not (a xor b);
    layer4_outputs(4614) <= a and b;
    layer4_outputs(4615) <= not a;
    layer4_outputs(4616) <= not b or a;
    layer4_outputs(4617) <= '0';
    layer4_outputs(4618) <= b;
    layer4_outputs(4619) <= '1';
    layer4_outputs(4620) <= not a;
    layer4_outputs(4621) <= not (a xor b);
    layer4_outputs(4622) <= not b;
    layer4_outputs(4623) <= not (a or b);
    layer4_outputs(4624) <= a and b;
    layer4_outputs(4625) <= b;
    layer4_outputs(4626) <= not (a or b);
    layer4_outputs(4627) <= not (a and b);
    layer4_outputs(4628) <= not (a and b);
    layer4_outputs(4629) <= b and not a;
    layer4_outputs(4630) <= not (a or b);
    layer4_outputs(4631) <= not a;
    layer4_outputs(4632) <= b;
    layer4_outputs(4633) <= not a;
    layer4_outputs(4634) <= '1';
    layer4_outputs(4635) <= b;
    layer4_outputs(4636) <= b and not a;
    layer4_outputs(4637) <= b;
    layer4_outputs(4638) <= not b or a;
    layer4_outputs(4639) <= b and not a;
    layer4_outputs(4640) <= a or b;
    layer4_outputs(4641) <= not (a xor b);
    layer4_outputs(4642) <= not a;
    layer4_outputs(4643) <= b and not a;
    layer4_outputs(4644) <= b;
    layer4_outputs(4645) <= not b;
    layer4_outputs(4646) <= not (a xor b);
    layer4_outputs(4647) <= not a or b;
    layer4_outputs(4648) <= not a or b;
    layer4_outputs(4649) <= b;
    layer4_outputs(4650) <= b;
    layer4_outputs(4651) <= not (a or b);
    layer4_outputs(4652) <= not b;
    layer4_outputs(4653) <= not (a xor b);
    layer4_outputs(4654) <= not a;
    layer4_outputs(4655) <= not b or a;
    layer4_outputs(4656) <= not b;
    layer4_outputs(4657) <= not (a or b);
    layer4_outputs(4658) <= a xor b;
    layer4_outputs(4659) <= a or b;
    layer4_outputs(4660) <= not a;
    layer4_outputs(4661) <= a xor b;
    layer4_outputs(4662) <= not (a and b);
    layer4_outputs(4663) <= not a;
    layer4_outputs(4664) <= not b or a;
    layer4_outputs(4665) <= not (a or b);
    layer4_outputs(4666) <= not (a xor b);
    layer4_outputs(4667) <= not a or b;
    layer4_outputs(4668) <= not (a xor b);
    layer4_outputs(4669) <= not a;
    layer4_outputs(4670) <= '0';
    layer4_outputs(4671) <= not b;
    layer4_outputs(4672) <= b;
    layer4_outputs(4673) <= a;
    layer4_outputs(4674) <= a and not b;
    layer4_outputs(4675) <= not b or a;
    layer4_outputs(4676) <= '0';
    layer4_outputs(4677) <= a;
    layer4_outputs(4678) <= a xor b;
    layer4_outputs(4679) <= a and not b;
    layer4_outputs(4680) <= not a or b;
    layer4_outputs(4681) <= a and not b;
    layer4_outputs(4682) <= a or b;
    layer4_outputs(4683) <= not (a xor b);
    layer4_outputs(4684) <= a and b;
    layer4_outputs(4685) <= not a or b;
    layer4_outputs(4686) <= not b;
    layer4_outputs(4687) <= a or b;
    layer4_outputs(4688) <= not (a xor b);
    layer4_outputs(4689) <= not b;
    layer4_outputs(4690) <= b and not a;
    layer4_outputs(4691) <= b;
    layer4_outputs(4692) <= not b or a;
    layer4_outputs(4693) <= a and b;
    layer4_outputs(4694) <= not b;
    layer4_outputs(4695) <= b;
    layer4_outputs(4696) <= not (a xor b);
    layer4_outputs(4697) <= not b;
    layer4_outputs(4698) <= not (a xor b);
    layer4_outputs(4699) <= a;
    layer4_outputs(4700) <= not (a or b);
    layer4_outputs(4701) <= not a;
    layer4_outputs(4702) <= not b;
    layer4_outputs(4703) <= not (a xor b);
    layer4_outputs(4704) <= not a;
    layer4_outputs(4705) <= a xor b;
    layer4_outputs(4706) <= not b;
    layer4_outputs(4707) <= not (a xor b);
    layer4_outputs(4708) <= a and not b;
    layer4_outputs(4709) <= not (a and b);
    layer4_outputs(4710) <= b;
    layer4_outputs(4711) <= b;
    layer4_outputs(4712) <= b and not a;
    layer4_outputs(4713) <= not a;
    layer4_outputs(4714) <= not b or a;
    layer4_outputs(4715) <= a xor b;
    layer4_outputs(4716) <= a;
    layer4_outputs(4717) <= not a;
    layer4_outputs(4718) <= not (a xor b);
    layer4_outputs(4719) <= not b or a;
    layer4_outputs(4720) <= not a or b;
    layer4_outputs(4721) <= not (a or b);
    layer4_outputs(4722) <= not a;
    layer4_outputs(4723) <= b;
    layer4_outputs(4724) <= not (a xor b);
    layer4_outputs(4725) <= not b;
    layer4_outputs(4726) <= not (a and b);
    layer4_outputs(4727) <= a or b;
    layer4_outputs(4728) <= not b;
    layer4_outputs(4729) <= not (a or b);
    layer4_outputs(4730) <= not b;
    layer4_outputs(4731) <= a and not b;
    layer4_outputs(4732) <= a;
    layer4_outputs(4733) <= not a;
    layer4_outputs(4734) <= not a or b;
    layer4_outputs(4735) <= not (a or b);
    layer4_outputs(4736) <= a xor b;
    layer4_outputs(4737) <= not b;
    layer4_outputs(4738) <= a;
    layer4_outputs(4739) <= a;
    layer4_outputs(4740) <= b and not a;
    layer4_outputs(4741) <= b;
    layer4_outputs(4742) <= not b or a;
    layer4_outputs(4743) <= not b;
    layer4_outputs(4744) <= not a or b;
    layer4_outputs(4745) <= b;
    layer4_outputs(4746) <= not a;
    layer4_outputs(4747) <= b and not a;
    layer4_outputs(4748) <= b;
    layer4_outputs(4749) <= a;
    layer4_outputs(4750) <= not a;
    layer4_outputs(4751) <= not a;
    layer4_outputs(4752) <= a and not b;
    layer4_outputs(4753) <= not (a and b);
    layer4_outputs(4754) <= not a;
    layer4_outputs(4755) <= b and not a;
    layer4_outputs(4756) <= a and b;
    layer4_outputs(4757) <= not b;
    layer4_outputs(4758) <= not (a or b);
    layer4_outputs(4759) <= not a or b;
    layer4_outputs(4760) <= b;
    layer4_outputs(4761) <= a and b;
    layer4_outputs(4762) <= not a or b;
    layer4_outputs(4763) <= a xor b;
    layer4_outputs(4764) <= a xor b;
    layer4_outputs(4765) <= b;
    layer4_outputs(4766) <= a and not b;
    layer4_outputs(4767) <= not a;
    layer4_outputs(4768) <= not b;
    layer4_outputs(4769) <= not (a and b);
    layer4_outputs(4770) <= not (a and b);
    layer4_outputs(4771) <= a or b;
    layer4_outputs(4772) <= not (a and b);
    layer4_outputs(4773) <= not (a or b);
    layer4_outputs(4774) <= b and not a;
    layer4_outputs(4775) <= b;
    layer4_outputs(4776) <= not (a xor b);
    layer4_outputs(4777) <= not a;
    layer4_outputs(4778) <= b;
    layer4_outputs(4779) <= not (a xor b);
    layer4_outputs(4780) <= b;
    layer4_outputs(4781) <= b and not a;
    layer4_outputs(4782) <= not b;
    layer4_outputs(4783) <= not a;
    layer4_outputs(4784) <= a or b;
    layer4_outputs(4785) <= not (a or b);
    layer4_outputs(4786) <= a and b;
    layer4_outputs(4787) <= b and not a;
    layer4_outputs(4788) <= not (a and b);
    layer4_outputs(4789) <= not (a or b);
    layer4_outputs(4790) <= b;
    layer4_outputs(4791) <= a xor b;
    layer4_outputs(4792) <= not a;
    layer4_outputs(4793) <= b and not a;
    layer4_outputs(4794) <= a;
    layer4_outputs(4795) <= not (a or b);
    layer4_outputs(4796) <= b and not a;
    layer4_outputs(4797) <= a or b;
    layer4_outputs(4798) <= b;
    layer4_outputs(4799) <= b and not a;
    layer4_outputs(4800) <= not b;
    layer4_outputs(4801) <= not (a and b);
    layer4_outputs(4802) <= not (a xor b);
    layer4_outputs(4803) <= not a or b;
    layer4_outputs(4804) <= b and not a;
    layer4_outputs(4805) <= not a or b;
    layer4_outputs(4806) <= a and not b;
    layer4_outputs(4807) <= a xor b;
    layer4_outputs(4808) <= a;
    layer4_outputs(4809) <= a;
    layer4_outputs(4810) <= a;
    layer4_outputs(4811) <= '0';
    layer4_outputs(4812) <= not (a and b);
    layer4_outputs(4813) <= b;
    layer4_outputs(4814) <= not b;
    layer4_outputs(4815) <= not a or b;
    layer4_outputs(4816) <= '1';
    layer4_outputs(4817) <= not a or b;
    layer4_outputs(4818) <= b;
    layer4_outputs(4819) <= a and not b;
    layer4_outputs(4820) <= not a;
    layer4_outputs(4821) <= a;
    layer4_outputs(4822) <= not (a and b);
    layer4_outputs(4823) <= not b;
    layer4_outputs(4824) <= a xor b;
    layer4_outputs(4825) <= a and not b;
    layer4_outputs(4826) <= b and not a;
    layer4_outputs(4827) <= b;
    layer4_outputs(4828) <= a;
    layer4_outputs(4829) <= b;
    layer4_outputs(4830) <= a and not b;
    layer4_outputs(4831) <= not a;
    layer4_outputs(4832) <= not b;
    layer4_outputs(4833) <= a;
    layer4_outputs(4834) <= a and not b;
    layer4_outputs(4835) <= a and b;
    layer4_outputs(4836) <= not (a xor b);
    layer4_outputs(4837) <= a xor b;
    layer4_outputs(4838) <= '0';
    layer4_outputs(4839) <= a xor b;
    layer4_outputs(4840) <= b;
    layer4_outputs(4841) <= not b or a;
    layer4_outputs(4842) <= a;
    layer4_outputs(4843) <= not a or b;
    layer4_outputs(4844) <= a or b;
    layer4_outputs(4845) <= not (a xor b);
    layer4_outputs(4846) <= a or b;
    layer4_outputs(4847) <= not a;
    layer4_outputs(4848) <= not a or b;
    layer4_outputs(4849) <= not (a or b);
    layer4_outputs(4850) <= not (a or b);
    layer4_outputs(4851) <= a and b;
    layer4_outputs(4852) <= not b;
    layer4_outputs(4853) <= not a or b;
    layer4_outputs(4854) <= a;
    layer4_outputs(4855) <= a or b;
    layer4_outputs(4856) <= not a;
    layer4_outputs(4857) <= not (a and b);
    layer4_outputs(4858) <= a;
    layer4_outputs(4859) <= not b;
    layer4_outputs(4860) <= not (a or b);
    layer4_outputs(4861) <= not b;
    layer4_outputs(4862) <= a and not b;
    layer4_outputs(4863) <= '1';
    layer4_outputs(4864) <= not a;
    layer4_outputs(4865) <= not b or a;
    layer4_outputs(4866) <= a and b;
    layer4_outputs(4867) <= not b or a;
    layer4_outputs(4868) <= not b;
    layer4_outputs(4869) <= a;
    layer4_outputs(4870) <= not b;
    layer4_outputs(4871) <= not a;
    layer4_outputs(4872) <= a;
    layer4_outputs(4873) <= not b;
    layer4_outputs(4874) <= a or b;
    layer4_outputs(4875) <= not b;
    layer4_outputs(4876) <= not (a and b);
    layer4_outputs(4877) <= a;
    layer4_outputs(4878) <= not a or b;
    layer4_outputs(4879) <= not (a or b);
    layer4_outputs(4880) <= not a or b;
    layer4_outputs(4881) <= not (a and b);
    layer4_outputs(4882) <= not b;
    layer4_outputs(4883) <= b;
    layer4_outputs(4884) <= a;
    layer4_outputs(4885) <= b and not a;
    layer4_outputs(4886) <= a and b;
    layer4_outputs(4887) <= b;
    layer4_outputs(4888) <= a;
    layer4_outputs(4889) <= not (a and b);
    layer4_outputs(4890) <= a and b;
    layer4_outputs(4891) <= not b or a;
    layer4_outputs(4892) <= a and b;
    layer4_outputs(4893) <= not a;
    layer4_outputs(4894) <= a xor b;
    layer4_outputs(4895) <= not a;
    layer4_outputs(4896) <= a or b;
    layer4_outputs(4897) <= '1';
    layer4_outputs(4898) <= not (a and b);
    layer4_outputs(4899) <= b;
    layer4_outputs(4900) <= '0';
    layer4_outputs(4901) <= a or b;
    layer4_outputs(4902) <= not b;
    layer4_outputs(4903) <= a;
    layer4_outputs(4904) <= not (a and b);
    layer4_outputs(4905) <= not (a or b);
    layer4_outputs(4906) <= '0';
    layer4_outputs(4907) <= b;
    layer4_outputs(4908) <= not (a or b);
    layer4_outputs(4909) <= not b;
    layer4_outputs(4910) <= b;
    layer4_outputs(4911) <= a or b;
    layer4_outputs(4912) <= a and not b;
    layer4_outputs(4913) <= b;
    layer4_outputs(4914) <= a;
    layer4_outputs(4915) <= a and not b;
    layer4_outputs(4916) <= not (a or b);
    layer4_outputs(4917) <= not b;
    layer4_outputs(4918) <= a xor b;
    layer4_outputs(4919) <= a or b;
    layer4_outputs(4920) <= not a;
    layer4_outputs(4921) <= not b;
    layer4_outputs(4922) <= not (a xor b);
    layer4_outputs(4923) <= b and not a;
    layer4_outputs(4924) <= b;
    layer4_outputs(4925) <= not a or b;
    layer4_outputs(4926) <= b;
    layer4_outputs(4927) <= b and not a;
    layer4_outputs(4928) <= a xor b;
    layer4_outputs(4929) <= b;
    layer4_outputs(4930) <= not (a or b);
    layer4_outputs(4931) <= a or b;
    layer4_outputs(4932) <= not a;
    layer4_outputs(4933) <= not a or b;
    layer4_outputs(4934) <= not b;
    layer4_outputs(4935) <= a and b;
    layer4_outputs(4936) <= a or b;
    layer4_outputs(4937) <= not (a xor b);
    layer4_outputs(4938) <= not b or a;
    layer4_outputs(4939) <= a and not b;
    layer4_outputs(4940) <= b and not a;
    layer4_outputs(4941) <= not a or b;
    layer4_outputs(4942) <= not a;
    layer4_outputs(4943) <= not (a or b);
    layer4_outputs(4944) <= not b or a;
    layer4_outputs(4945) <= not (a xor b);
    layer4_outputs(4946) <= not (a or b);
    layer4_outputs(4947) <= a;
    layer4_outputs(4948) <= a and not b;
    layer4_outputs(4949) <= a or b;
    layer4_outputs(4950) <= a and not b;
    layer4_outputs(4951) <= not a;
    layer4_outputs(4952) <= not a;
    layer4_outputs(4953) <= '1';
    layer4_outputs(4954) <= b;
    layer4_outputs(4955) <= b and not a;
    layer4_outputs(4956) <= not (a or b);
    layer4_outputs(4957) <= a or b;
    layer4_outputs(4958) <= not b or a;
    layer4_outputs(4959) <= not b;
    layer4_outputs(4960) <= a and not b;
    layer4_outputs(4961) <= not a;
    layer4_outputs(4962) <= b;
    layer4_outputs(4963) <= b;
    layer4_outputs(4964) <= not b or a;
    layer4_outputs(4965) <= not (a or b);
    layer4_outputs(4966) <= not a or b;
    layer4_outputs(4967) <= not a;
    layer4_outputs(4968) <= b;
    layer4_outputs(4969) <= not (a and b);
    layer4_outputs(4970) <= b and not a;
    layer4_outputs(4971) <= not (a or b);
    layer4_outputs(4972) <= a and b;
    layer4_outputs(4973) <= a and b;
    layer4_outputs(4974) <= not (a or b);
    layer4_outputs(4975) <= a and b;
    layer4_outputs(4976) <= a xor b;
    layer4_outputs(4977) <= not a or b;
    layer4_outputs(4978) <= not b or a;
    layer4_outputs(4979) <= b and not a;
    layer4_outputs(4980) <= not b;
    layer4_outputs(4981) <= a or b;
    layer4_outputs(4982) <= '0';
    layer4_outputs(4983) <= a and b;
    layer4_outputs(4984) <= not a;
    layer4_outputs(4985) <= '0';
    layer4_outputs(4986) <= not (a and b);
    layer4_outputs(4987) <= b;
    layer4_outputs(4988) <= not b or a;
    layer4_outputs(4989) <= not b;
    layer4_outputs(4990) <= not a;
    layer4_outputs(4991) <= b;
    layer4_outputs(4992) <= not (a xor b);
    layer4_outputs(4993) <= not b;
    layer4_outputs(4994) <= b and not a;
    layer4_outputs(4995) <= a and not b;
    layer4_outputs(4996) <= not b or a;
    layer4_outputs(4997) <= not b or a;
    layer4_outputs(4998) <= a and not b;
    layer4_outputs(4999) <= a;
    layer4_outputs(5000) <= b and not a;
    layer4_outputs(5001) <= not a;
    layer4_outputs(5002) <= not (a and b);
    layer4_outputs(5003) <= b;
    layer4_outputs(5004) <= not a;
    layer4_outputs(5005) <= b and not a;
    layer4_outputs(5006) <= b;
    layer4_outputs(5007) <= a and not b;
    layer4_outputs(5008) <= b;
    layer4_outputs(5009) <= '1';
    layer4_outputs(5010) <= b;
    layer4_outputs(5011) <= '1';
    layer4_outputs(5012) <= not b;
    layer4_outputs(5013) <= not (a or b);
    layer4_outputs(5014) <= not b or a;
    layer4_outputs(5015) <= not b or a;
    layer4_outputs(5016) <= '1';
    layer4_outputs(5017) <= a xor b;
    layer4_outputs(5018) <= not b;
    layer4_outputs(5019) <= not a;
    layer4_outputs(5020) <= b;
    layer4_outputs(5021) <= a and b;
    layer4_outputs(5022) <= not b;
    layer4_outputs(5023) <= not a;
    layer4_outputs(5024) <= a and b;
    layer4_outputs(5025) <= a and not b;
    layer4_outputs(5026) <= a or b;
    layer4_outputs(5027) <= not a;
    layer4_outputs(5028) <= b;
    layer4_outputs(5029) <= not a or b;
    layer4_outputs(5030) <= not b;
    layer4_outputs(5031) <= a and b;
    layer4_outputs(5032) <= not (a and b);
    layer4_outputs(5033) <= not b;
    layer4_outputs(5034) <= a or b;
    layer4_outputs(5035) <= not (a or b);
    layer4_outputs(5036) <= not a;
    layer4_outputs(5037) <= not a;
    layer4_outputs(5038) <= '0';
    layer4_outputs(5039) <= '1';
    layer4_outputs(5040) <= a or b;
    layer4_outputs(5041) <= '1';
    layer4_outputs(5042) <= not b;
    layer4_outputs(5043) <= not (a xor b);
    layer4_outputs(5044) <= not a;
    layer4_outputs(5045) <= a and not b;
    layer4_outputs(5046) <= a;
    layer4_outputs(5047) <= b and not a;
    layer4_outputs(5048) <= a and not b;
    layer4_outputs(5049) <= not b;
    layer4_outputs(5050) <= not (a xor b);
    layer4_outputs(5051) <= not b;
    layer4_outputs(5052) <= b and not a;
    layer4_outputs(5053) <= a or b;
    layer4_outputs(5054) <= not (a and b);
    layer4_outputs(5055) <= b;
    layer4_outputs(5056) <= not a;
    layer4_outputs(5057) <= a;
    layer4_outputs(5058) <= a or b;
    layer4_outputs(5059) <= a;
    layer4_outputs(5060) <= not (a and b);
    layer4_outputs(5061) <= a;
    layer4_outputs(5062) <= b and not a;
    layer4_outputs(5063) <= a and not b;
    layer4_outputs(5064) <= b;
    layer4_outputs(5065) <= not a or b;
    layer4_outputs(5066) <= not a;
    layer4_outputs(5067) <= not (a and b);
    layer4_outputs(5068) <= not (a or b);
    layer4_outputs(5069) <= a and not b;
    layer4_outputs(5070) <= a;
    layer4_outputs(5071) <= not a;
    layer4_outputs(5072) <= not (a and b);
    layer4_outputs(5073) <= a xor b;
    layer4_outputs(5074) <= not (a or b);
    layer4_outputs(5075) <= '0';
    layer4_outputs(5076) <= not (a or b);
    layer4_outputs(5077) <= b;
    layer4_outputs(5078) <= a;
    layer4_outputs(5079) <= a;
    layer4_outputs(5080) <= a;
    layer4_outputs(5081) <= not (a or b);
    layer4_outputs(5082) <= not b;
    layer4_outputs(5083) <= not a or b;
    layer4_outputs(5084) <= b;
    layer4_outputs(5085) <= not b;
    layer4_outputs(5086) <= b;
    layer4_outputs(5087) <= not b or a;
    layer4_outputs(5088) <= not a;
    layer4_outputs(5089) <= b and not a;
    layer4_outputs(5090) <= not a;
    layer4_outputs(5091) <= b and not a;
    layer4_outputs(5092) <= not a;
    layer4_outputs(5093) <= b;
    layer4_outputs(5094) <= a and b;
    layer4_outputs(5095) <= not (a and b);
    layer4_outputs(5096) <= not (a or b);
    layer4_outputs(5097) <= not a;
    layer4_outputs(5098) <= not a;
    layer4_outputs(5099) <= b;
    layer4_outputs(5100) <= '1';
    layer4_outputs(5101) <= a and not b;
    layer4_outputs(5102) <= a or b;
    layer4_outputs(5103) <= not a;
    layer4_outputs(5104) <= not (a or b);
    layer4_outputs(5105) <= not b;
    layer4_outputs(5106) <= not a;
    layer4_outputs(5107) <= not a;
    layer4_outputs(5108) <= '0';
    layer4_outputs(5109) <= not (a xor b);
    layer4_outputs(5110) <= not a;
    layer4_outputs(5111) <= a and b;
    layer4_outputs(5112) <= a;
    layer4_outputs(5113) <= b and not a;
    layer4_outputs(5114) <= '1';
    layer4_outputs(5115) <= not a or b;
    layer4_outputs(5116) <= a and not b;
    layer4_outputs(5117) <= a and not b;
    layer4_outputs(5118) <= a and b;
    layer4_outputs(5119) <= not a or b;
    layer4_outputs(5120) <= a and not b;
    layer4_outputs(5121) <= not b;
    layer4_outputs(5122) <= a or b;
    layer4_outputs(5123) <= not a or b;
    layer4_outputs(5124) <= not b;
    layer4_outputs(5125) <= a;
    layer4_outputs(5126) <= b;
    layer4_outputs(5127) <= b;
    layer4_outputs(5128) <= a or b;
    layer4_outputs(5129) <= a;
    layer4_outputs(5130) <= not (a and b);
    layer4_outputs(5131) <= not b;
    layer4_outputs(5132) <= b;
    layer4_outputs(5133) <= not b;
    layer4_outputs(5134) <= a and not b;
    layer4_outputs(5135) <= a;
    layer4_outputs(5136) <= not (a or b);
    layer4_outputs(5137) <= a;
    layer4_outputs(5138) <= not b or a;
    layer4_outputs(5139) <= a;
    layer4_outputs(5140) <= b;
    layer4_outputs(5141) <= a xor b;
    layer4_outputs(5142) <= a and not b;
    layer4_outputs(5143) <= a or b;
    layer4_outputs(5144) <= b;
    layer4_outputs(5145) <= a and not b;
    layer4_outputs(5146) <= a and b;
    layer4_outputs(5147) <= not (a and b);
    layer4_outputs(5148) <= '1';
    layer4_outputs(5149) <= a or b;
    layer4_outputs(5150) <= b;
    layer4_outputs(5151) <= not b;
    layer4_outputs(5152) <= a and b;
    layer4_outputs(5153) <= not b or a;
    layer4_outputs(5154) <= not b;
    layer4_outputs(5155) <= a;
    layer4_outputs(5156) <= not (a or b);
    layer4_outputs(5157) <= not b;
    layer4_outputs(5158) <= a;
    layer4_outputs(5159) <= not (a or b);
    layer4_outputs(5160) <= a;
    layer4_outputs(5161) <= b and not a;
    layer4_outputs(5162) <= not (a or b);
    layer4_outputs(5163) <= a or b;
    layer4_outputs(5164) <= a;
    layer4_outputs(5165) <= not (a and b);
    layer4_outputs(5166) <= b;
    layer4_outputs(5167) <= not b;
    layer4_outputs(5168) <= b;
    layer4_outputs(5169) <= a;
    layer4_outputs(5170) <= not b;
    layer4_outputs(5171) <= not b;
    layer4_outputs(5172) <= b;
    layer4_outputs(5173) <= not (a xor b);
    layer4_outputs(5174) <= not a;
    layer4_outputs(5175) <= a and b;
    layer4_outputs(5176) <= not (a xor b);
    layer4_outputs(5177) <= not a;
    layer4_outputs(5178) <= b;
    layer4_outputs(5179) <= a;
    layer4_outputs(5180) <= a and b;
    layer4_outputs(5181) <= '1';
    layer4_outputs(5182) <= not (a and b);
    layer4_outputs(5183) <= not (a xor b);
    layer4_outputs(5184) <= not a or b;
    layer4_outputs(5185) <= not a;
    layer4_outputs(5186) <= not (a xor b);
    layer4_outputs(5187) <= b;
    layer4_outputs(5188) <= b and not a;
    layer4_outputs(5189) <= a or b;
    layer4_outputs(5190) <= a;
    layer4_outputs(5191) <= a;
    layer4_outputs(5192) <= not (a or b);
    layer4_outputs(5193) <= not b or a;
    layer4_outputs(5194) <= b;
    layer4_outputs(5195) <= b;
    layer4_outputs(5196) <= a and b;
    layer4_outputs(5197) <= a;
    layer4_outputs(5198) <= not (a or b);
    layer4_outputs(5199) <= not a;
    layer4_outputs(5200) <= b and not a;
    layer4_outputs(5201) <= not a;
    layer4_outputs(5202) <= a and not b;
    layer4_outputs(5203) <= not b;
    layer4_outputs(5204) <= not a;
    layer4_outputs(5205) <= not (a and b);
    layer4_outputs(5206) <= not b or a;
    layer4_outputs(5207) <= '1';
    layer4_outputs(5208) <= a;
    layer4_outputs(5209) <= not (a or b);
    layer4_outputs(5210) <= a;
    layer4_outputs(5211) <= a and b;
    layer4_outputs(5212) <= a and b;
    layer4_outputs(5213) <= '0';
    layer4_outputs(5214) <= not (a and b);
    layer4_outputs(5215) <= a and b;
    layer4_outputs(5216) <= b;
    layer4_outputs(5217) <= b;
    layer4_outputs(5218) <= not a or b;
    layer4_outputs(5219) <= a and b;
    layer4_outputs(5220) <= not b;
    layer4_outputs(5221) <= a and not b;
    layer4_outputs(5222) <= not a;
    layer4_outputs(5223) <= not b or a;
    layer4_outputs(5224) <= not a;
    layer4_outputs(5225) <= b and not a;
    layer4_outputs(5226) <= b;
    layer4_outputs(5227) <= a xor b;
    layer4_outputs(5228) <= not b or a;
    layer4_outputs(5229) <= not a or b;
    layer4_outputs(5230) <= a and b;
    layer4_outputs(5231) <= b;
    layer4_outputs(5232) <= not b;
    layer4_outputs(5233) <= not (a xor b);
    layer4_outputs(5234) <= not a or b;
    layer4_outputs(5235) <= not a;
    layer4_outputs(5236) <= b;
    layer4_outputs(5237) <= not (a xor b);
    layer4_outputs(5238) <= not b;
    layer4_outputs(5239) <= a;
    layer4_outputs(5240) <= a and b;
    layer4_outputs(5241) <= not a;
    layer4_outputs(5242) <= not (a and b);
    layer4_outputs(5243) <= b;
    layer4_outputs(5244) <= not b;
    layer4_outputs(5245) <= b and not a;
    layer4_outputs(5246) <= '0';
    layer4_outputs(5247) <= not a;
    layer4_outputs(5248) <= a and not b;
    layer4_outputs(5249) <= not a;
    layer4_outputs(5250) <= not b;
    layer4_outputs(5251) <= not b;
    layer4_outputs(5252) <= not (a and b);
    layer4_outputs(5253) <= b;
    layer4_outputs(5254) <= b;
    layer4_outputs(5255) <= a or b;
    layer4_outputs(5256) <= '0';
    layer4_outputs(5257) <= not b;
    layer4_outputs(5258) <= not b;
    layer4_outputs(5259) <= not a;
    layer4_outputs(5260) <= a and b;
    layer4_outputs(5261) <= not b;
    layer4_outputs(5262) <= not b;
    layer4_outputs(5263) <= a;
    layer4_outputs(5264) <= not b;
    layer4_outputs(5265) <= a and b;
    layer4_outputs(5266) <= not b;
    layer4_outputs(5267) <= not (a xor b);
    layer4_outputs(5268) <= not b;
    layer4_outputs(5269) <= not a or b;
    layer4_outputs(5270) <= a and not b;
    layer4_outputs(5271) <= a and b;
    layer4_outputs(5272) <= not a;
    layer4_outputs(5273) <= not b;
    layer4_outputs(5274) <= a;
    layer4_outputs(5275) <= not b;
    layer4_outputs(5276) <= b;
    layer4_outputs(5277) <= a;
    layer4_outputs(5278) <= a;
    layer4_outputs(5279) <= a and b;
    layer4_outputs(5280) <= not b;
    layer4_outputs(5281) <= not a or b;
    layer4_outputs(5282) <= not a;
    layer4_outputs(5283) <= a;
    layer4_outputs(5284) <= '0';
    layer4_outputs(5285) <= b;
    layer4_outputs(5286) <= a xor b;
    layer4_outputs(5287) <= not (a xor b);
    layer4_outputs(5288) <= a or b;
    layer4_outputs(5289) <= not (a or b);
    layer4_outputs(5290) <= b;
    layer4_outputs(5291) <= not a;
    layer4_outputs(5292) <= '1';
    layer4_outputs(5293) <= b and not a;
    layer4_outputs(5294) <= a and b;
    layer4_outputs(5295) <= a and b;
    layer4_outputs(5296) <= b and not a;
    layer4_outputs(5297) <= not b or a;
    layer4_outputs(5298) <= a;
    layer4_outputs(5299) <= a;
    layer4_outputs(5300) <= a and b;
    layer4_outputs(5301) <= not b;
    layer4_outputs(5302) <= not a;
    layer4_outputs(5303) <= a;
    layer4_outputs(5304) <= not (a and b);
    layer4_outputs(5305) <= not (a xor b);
    layer4_outputs(5306) <= a or b;
    layer4_outputs(5307) <= b;
    layer4_outputs(5308) <= b;
    layer4_outputs(5309) <= '1';
    layer4_outputs(5310) <= a and b;
    layer4_outputs(5311) <= a or b;
    layer4_outputs(5312) <= a xor b;
    layer4_outputs(5313) <= not (a or b);
    layer4_outputs(5314) <= a or b;
    layer4_outputs(5315) <= not (a and b);
    layer4_outputs(5316) <= not a or b;
    layer4_outputs(5317) <= not b;
    layer4_outputs(5318) <= b;
    layer4_outputs(5319) <= b and not a;
    layer4_outputs(5320) <= a;
    layer4_outputs(5321) <= not a;
    layer4_outputs(5322) <= not b or a;
    layer4_outputs(5323) <= a xor b;
    layer4_outputs(5324) <= not a;
    layer4_outputs(5325) <= not b or a;
    layer4_outputs(5326) <= b;
    layer4_outputs(5327) <= a or b;
    layer4_outputs(5328) <= not b or a;
    layer4_outputs(5329) <= not (a or b);
    layer4_outputs(5330) <= a and not b;
    layer4_outputs(5331) <= not (a or b);
    layer4_outputs(5332) <= not a or b;
    layer4_outputs(5333) <= not a;
    layer4_outputs(5334) <= a xor b;
    layer4_outputs(5335) <= not a;
    layer4_outputs(5336) <= a and b;
    layer4_outputs(5337) <= not a or b;
    layer4_outputs(5338) <= not (a or b);
    layer4_outputs(5339) <= a;
    layer4_outputs(5340) <= a;
    layer4_outputs(5341) <= not (a or b);
    layer4_outputs(5342) <= a xor b;
    layer4_outputs(5343) <= a or b;
    layer4_outputs(5344) <= a xor b;
    layer4_outputs(5345) <= not (a or b);
    layer4_outputs(5346) <= b and not a;
    layer4_outputs(5347) <= a;
    layer4_outputs(5348) <= not b or a;
    layer4_outputs(5349) <= not (a xor b);
    layer4_outputs(5350) <= b and not a;
    layer4_outputs(5351) <= b;
    layer4_outputs(5352) <= not a or b;
    layer4_outputs(5353) <= not (a or b);
    layer4_outputs(5354) <= not b;
    layer4_outputs(5355) <= '0';
    layer4_outputs(5356) <= a;
    layer4_outputs(5357) <= not a;
    layer4_outputs(5358) <= b and not a;
    layer4_outputs(5359) <= not a;
    layer4_outputs(5360) <= a or b;
    layer4_outputs(5361) <= a or b;
    layer4_outputs(5362) <= not (a and b);
    layer4_outputs(5363) <= '0';
    layer4_outputs(5364) <= not b;
    layer4_outputs(5365) <= not a;
    layer4_outputs(5366) <= not (a or b);
    layer4_outputs(5367) <= not b or a;
    layer4_outputs(5368) <= '0';
    layer4_outputs(5369) <= '0';
    layer4_outputs(5370) <= b and not a;
    layer4_outputs(5371) <= a and not b;
    layer4_outputs(5372) <= '0';
    layer4_outputs(5373) <= not a;
    layer4_outputs(5374) <= a and b;
    layer4_outputs(5375) <= a or b;
    layer4_outputs(5376) <= not b;
    layer4_outputs(5377) <= not a;
    layer4_outputs(5378) <= not a;
    layer4_outputs(5379) <= not b or a;
    layer4_outputs(5380) <= not a;
    layer4_outputs(5381) <= b;
    layer4_outputs(5382) <= not b;
    layer4_outputs(5383) <= a and b;
    layer4_outputs(5384) <= not a or b;
    layer4_outputs(5385) <= not b or a;
    layer4_outputs(5386) <= b and not a;
    layer4_outputs(5387) <= '0';
    layer4_outputs(5388) <= b;
    layer4_outputs(5389) <= not a;
    layer4_outputs(5390) <= not (a and b);
    layer4_outputs(5391) <= a and b;
    layer4_outputs(5392) <= not b;
    layer4_outputs(5393) <= not (a or b);
    layer4_outputs(5394) <= b;
    layer4_outputs(5395) <= not (a and b);
    layer4_outputs(5396) <= a xor b;
    layer4_outputs(5397) <= not b;
    layer4_outputs(5398) <= a;
    layer4_outputs(5399) <= a or b;
    layer4_outputs(5400) <= a and not b;
    layer4_outputs(5401) <= b;
    layer4_outputs(5402) <= not b or a;
    layer4_outputs(5403) <= a and not b;
    layer4_outputs(5404) <= a;
    layer4_outputs(5405) <= not a;
    layer4_outputs(5406) <= b;
    layer4_outputs(5407) <= a;
    layer4_outputs(5408) <= not b or a;
    layer4_outputs(5409) <= a and not b;
    layer4_outputs(5410) <= a and not b;
    layer4_outputs(5411) <= not a or b;
    layer4_outputs(5412) <= b;
    layer4_outputs(5413) <= b and not a;
    layer4_outputs(5414) <= a;
    layer4_outputs(5415) <= not a;
    layer4_outputs(5416) <= not a or b;
    layer4_outputs(5417) <= not b or a;
    layer4_outputs(5418) <= a;
    layer4_outputs(5419) <= a xor b;
    layer4_outputs(5420) <= not a;
    layer4_outputs(5421) <= not (a or b);
    layer4_outputs(5422) <= a or b;
    layer4_outputs(5423) <= not b;
    layer4_outputs(5424) <= a or b;
    layer4_outputs(5425) <= not b;
    layer4_outputs(5426) <= a or b;
    layer4_outputs(5427) <= not (a or b);
    layer4_outputs(5428) <= not b;
    layer4_outputs(5429) <= not (a and b);
    layer4_outputs(5430) <= a;
    layer4_outputs(5431) <= b and not a;
    layer4_outputs(5432) <= not a or b;
    layer4_outputs(5433) <= a;
    layer4_outputs(5434) <= not a;
    layer4_outputs(5435) <= b;
    layer4_outputs(5436) <= b and not a;
    layer4_outputs(5437) <= a and b;
    layer4_outputs(5438) <= b;
    layer4_outputs(5439) <= a;
    layer4_outputs(5440) <= not a;
    layer4_outputs(5441) <= a xor b;
    layer4_outputs(5442) <= a and b;
    layer4_outputs(5443) <= b and not a;
    layer4_outputs(5444) <= a;
    layer4_outputs(5445) <= not b or a;
    layer4_outputs(5446) <= not a;
    layer4_outputs(5447) <= not a;
    layer4_outputs(5448) <= not a or b;
    layer4_outputs(5449) <= '0';
    layer4_outputs(5450) <= a or b;
    layer4_outputs(5451) <= not (a and b);
    layer4_outputs(5452) <= a or b;
    layer4_outputs(5453) <= a or b;
    layer4_outputs(5454) <= a;
    layer4_outputs(5455) <= not b;
    layer4_outputs(5456) <= not b;
    layer4_outputs(5457) <= a xor b;
    layer4_outputs(5458) <= not (a xor b);
    layer4_outputs(5459) <= not a or b;
    layer4_outputs(5460) <= a and b;
    layer4_outputs(5461) <= a or b;
    layer4_outputs(5462) <= a and not b;
    layer4_outputs(5463) <= a or b;
    layer4_outputs(5464) <= not (a xor b);
    layer4_outputs(5465) <= a and b;
    layer4_outputs(5466) <= not a;
    layer4_outputs(5467) <= a and b;
    layer4_outputs(5468) <= a xor b;
    layer4_outputs(5469) <= a;
    layer4_outputs(5470) <= a xor b;
    layer4_outputs(5471) <= not a;
    layer4_outputs(5472) <= b;
    layer4_outputs(5473) <= not (a or b);
    layer4_outputs(5474) <= not b or a;
    layer4_outputs(5475) <= a or b;
    layer4_outputs(5476) <= not b;
    layer4_outputs(5477) <= a or b;
    layer4_outputs(5478) <= b and not a;
    layer4_outputs(5479) <= '1';
    layer4_outputs(5480) <= a xor b;
    layer4_outputs(5481) <= b;
    layer4_outputs(5482) <= a xor b;
    layer4_outputs(5483) <= not (a and b);
    layer4_outputs(5484) <= not a;
    layer4_outputs(5485) <= not b;
    layer4_outputs(5486) <= not b;
    layer4_outputs(5487) <= not b or a;
    layer4_outputs(5488) <= a xor b;
    layer4_outputs(5489) <= b;
    layer4_outputs(5490) <= a;
    layer4_outputs(5491) <= not (a xor b);
    layer4_outputs(5492) <= not a;
    layer4_outputs(5493) <= a and b;
    layer4_outputs(5494) <= not a;
    layer4_outputs(5495) <= not a;
    layer4_outputs(5496) <= not a;
    layer4_outputs(5497) <= not (a xor b);
    layer4_outputs(5498) <= b;
    layer4_outputs(5499) <= a or b;
    layer4_outputs(5500) <= not (a xor b);
    layer4_outputs(5501) <= a and not b;
    layer4_outputs(5502) <= a and not b;
    layer4_outputs(5503) <= not (a xor b);
    layer4_outputs(5504) <= not (a xor b);
    layer4_outputs(5505) <= a xor b;
    layer4_outputs(5506) <= a;
    layer4_outputs(5507) <= not b;
    layer4_outputs(5508) <= not (a xor b);
    layer4_outputs(5509) <= b;
    layer4_outputs(5510) <= a and b;
    layer4_outputs(5511) <= not (a xor b);
    layer4_outputs(5512) <= a and b;
    layer4_outputs(5513) <= not b;
    layer4_outputs(5514) <= a or b;
    layer4_outputs(5515) <= not (a or b);
    layer4_outputs(5516) <= not b;
    layer4_outputs(5517) <= not a;
    layer4_outputs(5518) <= b and not a;
    layer4_outputs(5519) <= b and not a;
    layer4_outputs(5520) <= a;
    layer4_outputs(5521) <= a;
    layer4_outputs(5522) <= not b;
    layer4_outputs(5523) <= a and b;
    layer4_outputs(5524) <= b;
    layer4_outputs(5525) <= b;
    layer4_outputs(5526) <= not a;
    layer4_outputs(5527) <= a;
    layer4_outputs(5528) <= not a;
    layer4_outputs(5529) <= not (a xor b);
    layer4_outputs(5530) <= a;
    layer4_outputs(5531) <= a xor b;
    layer4_outputs(5532) <= not (a xor b);
    layer4_outputs(5533) <= not a;
    layer4_outputs(5534) <= a and not b;
    layer4_outputs(5535) <= a xor b;
    layer4_outputs(5536) <= a and not b;
    layer4_outputs(5537) <= not (a or b);
    layer4_outputs(5538) <= not b or a;
    layer4_outputs(5539) <= not (a or b);
    layer4_outputs(5540) <= b and not a;
    layer4_outputs(5541) <= not b;
    layer4_outputs(5542) <= a or b;
    layer4_outputs(5543) <= not b or a;
    layer4_outputs(5544) <= a or b;
    layer4_outputs(5545) <= not a;
    layer4_outputs(5546) <= not a;
    layer4_outputs(5547) <= not a or b;
    layer4_outputs(5548) <= not (a xor b);
    layer4_outputs(5549) <= not a;
    layer4_outputs(5550) <= b and not a;
    layer4_outputs(5551) <= not b or a;
    layer4_outputs(5552) <= b and not a;
    layer4_outputs(5553) <= a;
    layer4_outputs(5554) <= not (a or b);
    layer4_outputs(5555) <= a;
    layer4_outputs(5556) <= b;
    layer4_outputs(5557) <= not b;
    layer4_outputs(5558) <= a or b;
    layer4_outputs(5559) <= '0';
    layer4_outputs(5560) <= not (a and b);
    layer4_outputs(5561) <= a xor b;
    layer4_outputs(5562) <= a and not b;
    layer4_outputs(5563) <= not b;
    layer4_outputs(5564) <= a or b;
    layer4_outputs(5565) <= not (a xor b);
    layer4_outputs(5566) <= not a;
    layer4_outputs(5567) <= not b;
    layer4_outputs(5568) <= not (a and b);
    layer4_outputs(5569) <= b and not a;
    layer4_outputs(5570) <= not a;
    layer4_outputs(5571) <= b;
    layer4_outputs(5572) <= not (a xor b);
    layer4_outputs(5573) <= b and not a;
    layer4_outputs(5574) <= a and b;
    layer4_outputs(5575) <= a and b;
    layer4_outputs(5576) <= not a or b;
    layer4_outputs(5577) <= a xor b;
    layer4_outputs(5578) <= a xor b;
    layer4_outputs(5579) <= b;
    layer4_outputs(5580) <= not (a xor b);
    layer4_outputs(5581) <= not a;
    layer4_outputs(5582) <= not a;
    layer4_outputs(5583) <= a or b;
    layer4_outputs(5584) <= b;
    layer4_outputs(5585) <= not b or a;
    layer4_outputs(5586) <= not (a and b);
    layer4_outputs(5587) <= not a;
    layer4_outputs(5588) <= not (a or b);
    layer4_outputs(5589) <= '1';
    layer4_outputs(5590) <= not a or b;
    layer4_outputs(5591) <= a;
    layer4_outputs(5592) <= not (a and b);
    layer4_outputs(5593) <= b;
    layer4_outputs(5594) <= a;
    layer4_outputs(5595) <= '0';
    layer4_outputs(5596) <= a and not b;
    layer4_outputs(5597) <= not b;
    layer4_outputs(5598) <= a xor b;
    layer4_outputs(5599) <= not b;
    layer4_outputs(5600) <= not a or b;
    layer4_outputs(5601) <= b;
    layer4_outputs(5602) <= not a;
    layer4_outputs(5603) <= a or b;
    layer4_outputs(5604) <= b;
    layer4_outputs(5605) <= '1';
    layer4_outputs(5606) <= not b;
    layer4_outputs(5607) <= a;
    layer4_outputs(5608) <= not a;
    layer4_outputs(5609) <= a and b;
    layer4_outputs(5610) <= a xor b;
    layer4_outputs(5611) <= b;
    layer4_outputs(5612) <= not b or a;
    layer4_outputs(5613) <= b;
    layer4_outputs(5614) <= b;
    layer4_outputs(5615) <= not b;
    layer4_outputs(5616) <= '0';
    layer4_outputs(5617) <= b;
    layer4_outputs(5618) <= not a;
    layer4_outputs(5619) <= a or b;
    layer4_outputs(5620) <= not (a xor b);
    layer4_outputs(5621) <= a;
    layer4_outputs(5622) <= not b;
    layer4_outputs(5623) <= not (a xor b);
    layer4_outputs(5624) <= not (a or b);
    layer4_outputs(5625) <= not (a or b);
    layer4_outputs(5626) <= not a;
    layer4_outputs(5627) <= a xor b;
    layer4_outputs(5628) <= not b or a;
    layer4_outputs(5629) <= not (a or b);
    layer4_outputs(5630) <= not (a and b);
    layer4_outputs(5631) <= not (a xor b);
    layer4_outputs(5632) <= not b;
    layer4_outputs(5633) <= b and not a;
    layer4_outputs(5634) <= not a;
    layer4_outputs(5635) <= not b or a;
    layer4_outputs(5636) <= a;
    layer4_outputs(5637) <= not b;
    layer4_outputs(5638) <= a and not b;
    layer4_outputs(5639) <= not (a xor b);
    layer4_outputs(5640) <= b;
    layer4_outputs(5641) <= b;
    layer4_outputs(5642) <= a or b;
    layer4_outputs(5643) <= not (a and b);
    layer4_outputs(5644) <= not (a xor b);
    layer4_outputs(5645) <= not (a or b);
    layer4_outputs(5646) <= a and not b;
    layer4_outputs(5647) <= a and not b;
    layer4_outputs(5648) <= a xor b;
    layer4_outputs(5649) <= a xor b;
    layer4_outputs(5650) <= not b;
    layer4_outputs(5651) <= not b;
    layer4_outputs(5652) <= a xor b;
    layer4_outputs(5653) <= a and b;
    layer4_outputs(5654) <= b and not a;
    layer4_outputs(5655) <= not a;
    layer4_outputs(5656) <= a and not b;
    layer4_outputs(5657) <= b;
    layer4_outputs(5658) <= not a or b;
    layer4_outputs(5659) <= not (a and b);
    layer4_outputs(5660) <= not a;
    layer4_outputs(5661) <= not b;
    layer4_outputs(5662) <= not b;
    layer4_outputs(5663) <= b;
    layer4_outputs(5664) <= not b or a;
    layer4_outputs(5665) <= a and not b;
    layer4_outputs(5666) <= a xor b;
    layer4_outputs(5667) <= a or b;
    layer4_outputs(5668) <= not (a and b);
    layer4_outputs(5669) <= a;
    layer4_outputs(5670) <= a and b;
    layer4_outputs(5671) <= '0';
    layer4_outputs(5672) <= b;
    layer4_outputs(5673) <= not a;
    layer4_outputs(5674) <= not b;
    layer4_outputs(5675) <= a;
    layer4_outputs(5676) <= a and not b;
    layer4_outputs(5677) <= not b;
    layer4_outputs(5678) <= not (a or b);
    layer4_outputs(5679) <= b;
    layer4_outputs(5680) <= not (a and b);
    layer4_outputs(5681) <= a and not b;
    layer4_outputs(5682) <= not a or b;
    layer4_outputs(5683) <= not b or a;
    layer4_outputs(5684) <= a and not b;
    layer4_outputs(5685) <= not b or a;
    layer4_outputs(5686) <= not (a and b);
    layer4_outputs(5687) <= not (a xor b);
    layer4_outputs(5688) <= a and b;
    layer4_outputs(5689) <= a;
    layer4_outputs(5690) <= not (a and b);
    layer4_outputs(5691) <= not a or b;
    layer4_outputs(5692) <= a xor b;
    layer4_outputs(5693) <= not b or a;
    layer4_outputs(5694) <= not b;
    layer4_outputs(5695) <= a and not b;
    layer4_outputs(5696) <= not (a and b);
    layer4_outputs(5697) <= a and not b;
    layer4_outputs(5698) <= a;
    layer4_outputs(5699) <= not b;
    layer4_outputs(5700) <= not (a and b);
    layer4_outputs(5701) <= not (a and b);
    layer4_outputs(5702) <= a and b;
    layer4_outputs(5703) <= not a;
    layer4_outputs(5704) <= a;
    layer4_outputs(5705) <= a;
    layer4_outputs(5706) <= a;
    layer4_outputs(5707) <= not b;
    layer4_outputs(5708) <= not (a or b);
    layer4_outputs(5709) <= not a;
    layer4_outputs(5710) <= not a;
    layer4_outputs(5711) <= '0';
    layer4_outputs(5712) <= b and not a;
    layer4_outputs(5713) <= a and not b;
    layer4_outputs(5714) <= a xor b;
    layer4_outputs(5715) <= a;
    layer4_outputs(5716) <= a;
    layer4_outputs(5717) <= b;
    layer4_outputs(5718) <= b and not a;
    layer4_outputs(5719) <= not (a and b);
    layer4_outputs(5720) <= not b;
    layer4_outputs(5721) <= a xor b;
    layer4_outputs(5722) <= not a;
    layer4_outputs(5723) <= a;
    layer4_outputs(5724) <= a and not b;
    layer4_outputs(5725) <= a and not b;
    layer4_outputs(5726) <= b;
    layer4_outputs(5727) <= not a;
    layer4_outputs(5728) <= a;
    layer4_outputs(5729) <= not a;
    layer4_outputs(5730) <= not (a xor b);
    layer4_outputs(5731) <= not a;
    layer4_outputs(5732) <= not (a and b);
    layer4_outputs(5733) <= a or b;
    layer4_outputs(5734) <= not b;
    layer4_outputs(5735) <= not b;
    layer4_outputs(5736) <= b;
    layer4_outputs(5737) <= a and not b;
    layer4_outputs(5738) <= a;
    layer4_outputs(5739) <= a and not b;
    layer4_outputs(5740) <= not b;
    layer4_outputs(5741) <= not (a or b);
    layer4_outputs(5742) <= a or b;
    layer4_outputs(5743) <= not a or b;
    layer4_outputs(5744) <= a and not b;
    layer4_outputs(5745) <= a;
    layer4_outputs(5746) <= b;
    layer4_outputs(5747) <= a xor b;
    layer4_outputs(5748) <= not (a or b);
    layer4_outputs(5749) <= not (a or b);
    layer4_outputs(5750) <= a and b;
    layer4_outputs(5751) <= b;
    layer4_outputs(5752) <= not a;
    layer4_outputs(5753) <= a;
    layer4_outputs(5754) <= a and b;
    layer4_outputs(5755) <= not a or b;
    layer4_outputs(5756) <= a or b;
    layer4_outputs(5757) <= not a;
    layer4_outputs(5758) <= b;
    layer4_outputs(5759) <= not (a and b);
    layer4_outputs(5760) <= not (a xor b);
    layer4_outputs(5761) <= a or b;
    layer4_outputs(5762) <= not b;
    layer4_outputs(5763) <= b;
    layer4_outputs(5764) <= not (a and b);
    layer4_outputs(5765) <= a xor b;
    layer4_outputs(5766) <= not (a xor b);
    layer4_outputs(5767) <= not a;
    layer4_outputs(5768) <= a or b;
    layer4_outputs(5769) <= not (a and b);
    layer4_outputs(5770) <= not (a and b);
    layer4_outputs(5771) <= a and not b;
    layer4_outputs(5772) <= not (a or b);
    layer4_outputs(5773) <= b;
    layer4_outputs(5774) <= b;
    layer4_outputs(5775) <= not (a xor b);
    layer4_outputs(5776) <= b;
    layer4_outputs(5777) <= b and not a;
    layer4_outputs(5778) <= a and not b;
    layer4_outputs(5779) <= not b;
    layer4_outputs(5780) <= not b or a;
    layer4_outputs(5781) <= a xor b;
    layer4_outputs(5782) <= not a;
    layer4_outputs(5783) <= a and b;
    layer4_outputs(5784) <= a and b;
    layer4_outputs(5785) <= not a;
    layer4_outputs(5786) <= a;
    layer4_outputs(5787) <= b and not a;
    layer4_outputs(5788) <= not (a and b);
    layer4_outputs(5789) <= a;
    layer4_outputs(5790) <= '1';
    layer4_outputs(5791) <= not b;
    layer4_outputs(5792) <= not b;
    layer4_outputs(5793) <= not (a xor b);
    layer4_outputs(5794) <= a and b;
    layer4_outputs(5795) <= not a;
    layer4_outputs(5796) <= a and not b;
    layer4_outputs(5797) <= not (a xor b);
    layer4_outputs(5798) <= not a;
    layer4_outputs(5799) <= a and not b;
    layer4_outputs(5800) <= '1';
    layer4_outputs(5801) <= a;
    layer4_outputs(5802) <= a and b;
    layer4_outputs(5803) <= '1';
    layer4_outputs(5804) <= not b;
    layer4_outputs(5805) <= b;
    layer4_outputs(5806) <= b;
    layer4_outputs(5807) <= a;
    layer4_outputs(5808) <= not a or b;
    layer4_outputs(5809) <= a and not b;
    layer4_outputs(5810) <= not (a or b);
    layer4_outputs(5811) <= not b;
    layer4_outputs(5812) <= '0';
    layer4_outputs(5813) <= b and not a;
    layer4_outputs(5814) <= not b;
    layer4_outputs(5815) <= not (a or b);
    layer4_outputs(5816) <= not a or b;
    layer4_outputs(5817) <= not a;
    layer4_outputs(5818) <= b;
    layer4_outputs(5819) <= a and b;
    layer4_outputs(5820) <= not b;
    layer4_outputs(5821) <= b;
    layer4_outputs(5822) <= b;
    layer4_outputs(5823) <= not b;
    layer4_outputs(5824) <= not (a and b);
    layer4_outputs(5825) <= a;
    layer4_outputs(5826) <= a and not b;
    layer4_outputs(5827) <= a xor b;
    layer4_outputs(5828) <= not (a xor b);
    layer4_outputs(5829) <= '1';
    layer4_outputs(5830) <= not (a and b);
    layer4_outputs(5831) <= a xor b;
    layer4_outputs(5832) <= a;
    layer4_outputs(5833) <= a or b;
    layer4_outputs(5834) <= b and not a;
    layer4_outputs(5835) <= not b;
    layer4_outputs(5836) <= a or b;
    layer4_outputs(5837) <= a and b;
    layer4_outputs(5838) <= a and not b;
    layer4_outputs(5839) <= a;
    layer4_outputs(5840) <= a;
    layer4_outputs(5841) <= not (a xor b);
    layer4_outputs(5842) <= b and not a;
    layer4_outputs(5843) <= b;
    layer4_outputs(5844) <= b;
    layer4_outputs(5845) <= '1';
    layer4_outputs(5846) <= not a or b;
    layer4_outputs(5847) <= b;
    layer4_outputs(5848) <= not (a xor b);
    layer4_outputs(5849) <= not a;
    layer4_outputs(5850) <= not b;
    layer4_outputs(5851) <= a or b;
    layer4_outputs(5852) <= not b;
    layer4_outputs(5853) <= not (a and b);
    layer4_outputs(5854) <= a and not b;
    layer4_outputs(5855) <= b and not a;
    layer4_outputs(5856) <= a and b;
    layer4_outputs(5857) <= not a;
    layer4_outputs(5858) <= a and not b;
    layer4_outputs(5859) <= a or b;
    layer4_outputs(5860) <= not a;
    layer4_outputs(5861) <= not a or b;
    layer4_outputs(5862) <= not a or b;
    layer4_outputs(5863) <= not (a or b);
    layer4_outputs(5864) <= not (a and b);
    layer4_outputs(5865) <= not a;
    layer4_outputs(5866) <= b and not a;
    layer4_outputs(5867) <= a and b;
    layer4_outputs(5868) <= not (a or b);
    layer4_outputs(5869) <= not (a and b);
    layer4_outputs(5870) <= not a;
    layer4_outputs(5871) <= b and not a;
    layer4_outputs(5872) <= a or b;
    layer4_outputs(5873) <= a and not b;
    layer4_outputs(5874) <= not (a or b);
    layer4_outputs(5875) <= b;
    layer4_outputs(5876) <= a or b;
    layer4_outputs(5877) <= not a;
    layer4_outputs(5878) <= a and not b;
    layer4_outputs(5879) <= not a;
    layer4_outputs(5880) <= a;
    layer4_outputs(5881) <= a and b;
    layer4_outputs(5882) <= b and not a;
    layer4_outputs(5883) <= a and not b;
    layer4_outputs(5884) <= a and not b;
    layer4_outputs(5885) <= not (a or b);
    layer4_outputs(5886) <= not a or b;
    layer4_outputs(5887) <= a xor b;
    layer4_outputs(5888) <= not (a and b);
    layer4_outputs(5889) <= '1';
    layer4_outputs(5890) <= a and b;
    layer4_outputs(5891) <= not b or a;
    layer4_outputs(5892) <= not b or a;
    layer4_outputs(5893) <= b;
    layer4_outputs(5894) <= b;
    layer4_outputs(5895) <= a;
    layer4_outputs(5896) <= not b;
    layer4_outputs(5897) <= a;
    layer4_outputs(5898) <= a;
    layer4_outputs(5899) <= '0';
    layer4_outputs(5900) <= b;
    layer4_outputs(5901) <= a;
    layer4_outputs(5902) <= b;
    layer4_outputs(5903) <= b;
    layer4_outputs(5904) <= a xor b;
    layer4_outputs(5905) <= b and not a;
    layer4_outputs(5906) <= not b;
    layer4_outputs(5907) <= b;
    layer4_outputs(5908) <= b;
    layer4_outputs(5909) <= b and not a;
    layer4_outputs(5910) <= b;
    layer4_outputs(5911) <= a or b;
    layer4_outputs(5912) <= a;
    layer4_outputs(5913) <= not (a xor b);
    layer4_outputs(5914) <= a xor b;
    layer4_outputs(5915) <= a;
    layer4_outputs(5916) <= not (a and b);
    layer4_outputs(5917) <= '0';
    layer4_outputs(5918) <= b;
    layer4_outputs(5919) <= not a or b;
    layer4_outputs(5920) <= a and not b;
    layer4_outputs(5921) <= a or b;
    layer4_outputs(5922) <= not b;
    layer4_outputs(5923) <= not b or a;
    layer4_outputs(5924) <= not a;
    layer4_outputs(5925) <= a;
    layer4_outputs(5926) <= b and not a;
    layer4_outputs(5927) <= a;
    layer4_outputs(5928) <= b;
    layer4_outputs(5929) <= b and not a;
    layer4_outputs(5930) <= a or b;
    layer4_outputs(5931) <= '0';
    layer4_outputs(5932) <= b;
    layer4_outputs(5933) <= b;
    layer4_outputs(5934) <= a;
    layer4_outputs(5935) <= not (a or b);
    layer4_outputs(5936) <= not (a xor b);
    layer4_outputs(5937) <= not (a xor b);
    layer4_outputs(5938) <= b;
    layer4_outputs(5939) <= not b or a;
    layer4_outputs(5940) <= not b;
    layer4_outputs(5941) <= a xor b;
    layer4_outputs(5942) <= a and not b;
    layer4_outputs(5943) <= a;
    layer4_outputs(5944) <= a;
    layer4_outputs(5945) <= not (a xor b);
    layer4_outputs(5946) <= not b;
    layer4_outputs(5947) <= a and b;
    layer4_outputs(5948) <= not b;
    layer4_outputs(5949) <= b;
    layer4_outputs(5950) <= not (a xor b);
    layer4_outputs(5951) <= b;
    layer4_outputs(5952) <= not a;
    layer4_outputs(5953) <= a or b;
    layer4_outputs(5954) <= a;
    layer4_outputs(5955) <= not a or b;
    layer4_outputs(5956) <= not a;
    layer4_outputs(5957) <= not (a or b);
    layer4_outputs(5958) <= b;
    layer4_outputs(5959) <= not a or b;
    layer4_outputs(5960) <= a;
    layer4_outputs(5961) <= not b or a;
    layer4_outputs(5962) <= not a;
    layer4_outputs(5963) <= not a;
    layer4_outputs(5964) <= not (a or b);
    layer4_outputs(5965) <= not (a and b);
    layer4_outputs(5966) <= not b;
    layer4_outputs(5967) <= not a or b;
    layer4_outputs(5968) <= not (a and b);
    layer4_outputs(5969) <= b and not a;
    layer4_outputs(5970) <= not b or a;
    layer4_outputs(5971) <= not a or b;
    layer4_outputs(5972) <= not b;
    layer4_outputs(5973) <= a;
    layer4_outputs(5974) <= not b;
    layer4_outputs(5975) <= '1';
    layer4_outputs(5976) <= b;
    layer4_outputs(5977) <= b and not a;
    layer4_outputs(5978) <= a and not b;
    layer4_outputs(5979) <= b;
    layer4_outputs(5980) <= b and not a;
    layer4_outputs(5981) <= b and not a;
    layer4_outputs(5982) <= a or b;
    layer4_outputs(5983) <= a and b;
    layer4_outputs(5984) <= a and not b;
    layer4_outputs(5985) <= not (a xor b);
    layer4_outputs(5986) <= not a;
    layer4_outputs(5987) <= not b;
    layer4_outputs(5988) <= a or b;
    layer4_outputs(5989) <= a;
    layer4_outputs(5990) <= a;
    layer4_outputs(5991) <= a and not b;
    layer4_outputs(5992) <= b;
    layer4_outputs(5993) <= not b;
    layer4_outputs(5994) <= a and not b;
    layer4_outputs(5995) <= a and b;
    layer4_outputs(5996) <= b;
    layer4_outputs(5997) <= a;
    layer4_outputs(5998) <= '1';
    layer4_outputs(5999) <= a and b;
    layer4_outputs(6000) <= a;
    layer4_outputs(6001) <= b and not a;
    layer4_outputs(6002) <= a;
    layer4_outputs(6003) <= a and not b;
    layer4_outputs(6004) <= not (a xor b);
    layer4_outputs(6005) <= not (a or b);
    layer4_outputs(6006) <= b;
    layer4_outputs(6007) <= not b;
    layer4_outputs(6008) <= not (a or b);
    layer4_outputs(6009) <= not (a and b);
    layer4_outputs(6010) <= not b or a;
    layer4_outputs(6011) <= not a;
    layer4_outputs(6012) <= a and b;
    layer4_outputs(6013) <= a and b;
    layer4_outputs(6014) <= a and b;
    layer4_outputs(6015) <= not a;
    layer4_outputs(6016) <= '1';
    layer4_outputs(6017) <= b;
    layer4_outputs(6018) <= a or b;
    layer4_outputs(6019) <= a and not b;
    layer4_outputs(6020) <= a and b;
    layer4_outputs(6021) <= '0';
    layer4_outputs(6022) <= a;
    layer4_outputs(6023) <= a and not b;
    layer4_outputs(6024) <= b and not a;
    layer4_outputs(6025) <= a xor b;
    layer4_outputs(6026) <= not a or b;
    layer4_outputs(6027) <= not (a xor b);
    layer4_outputs(6028) <= not (a xor b);
    layer4_outputs(6029) <= not (a or b);
    layer4_outputs(6030) <= not (a and b);
    layer4_outputs(6031) <= a and not b;
    layer4_outputs(6032) <= not a;
    layer4_outputs(6033) <= not a;
    layer4_outputs(6034) <= b and not a;
    layer4_outputs(6035) <= b and not a;
    layer4_outputs(6036) <= b and not a;
    layer4_outputs(6037) <= b;
    layer4_outputs(6038) <= not b;
    layer4_outputs(6039) <= a and not b;
    layer4_outputs(6040) <= not (a and b);
    layer4_outputs(6041) <= '1';
    layer4_outputs(6042) <= a;
    layer4_outputs(6043) <= not a or b;
    layer4_outputs(6044) <= a and b;
    layer4_outputs(6045) <= a or b;
    layer4_outputs(6046) <= not a;
    layer4_outputs(6047) <= not b;
    layer4_outputs(6048) <= not a;
    layer4_outputs(6049) <= a and b;
    layer4_outputs(6050) <= not a;
    layer4_outputs(6051) <= a and not b;
    layer4_outputs(6052) <= not a;
    layer4_outputs(6053) <= b;
    layer4_outputs(6054) <= not a;
    layer4_outputs(6055) <= not (a and b);
    layer4_outputs(6056) <= not a;
    layer4_outputs(6057) <= not b;
    layer4_outputs(6058) <= b;
    layer4_outputs(6059) <= not b;
    layer4_outputs(6060) <= a and b;
    layer4_outputs(6061) <= not (a xor b);
    layer4_outputs(6062) <= not (a or b);
    layer4_outputs(6063) <= not b;
    layer4_outputs(6064) <= a or b;
    layer4_outputs(6065) <= b and not a;
    layer4_outputs(6066) <= not a or b;
    layer4_outputs(6067) <= b;
    layer4_outputs(6068) <= not b;
    layer4_outputs(6069) <= b;
    layer4_outputs(6070) <= not a;
    layer4_outputs(6071) <= not a;
    layer4_outputs(6072) <= a xor b;
    layer4_outputs(6073) <= not b;
    layer4_outputs(6074) <= not a;
    layer4_outputs(6075) <= b and not a;
    layer4_outputs(6076) <= a;
    layer4_outputs(6077) <= b and not a;
    layer4_outputs(6078) <= not a or b;
    layer4_outputs(6079) <= a xor b;
    layer4_outputs(6080) <= a and b;
    layer4_outputs(6081) <= not b or a;
    layer4_outputs(6082) <= '1';
    layer4_outputs(6083) <= not b;
    layer4_outputs(6084) <= not a or b;
    layer4_outputs(6085) <= b and not a;
    layer4_outputs(6086) <= not (a or b);
    layer4_outputs(6087) <= b;
    layer4_outputs(6088) <= not a;
    layer4_outputs(6089) <= not (a or b);
    layer4_outputs(6090) <= not a;
    layer4_outputs(6091) <= not (a xor b);
    layer4_outputs(6092) <= '1';
    layer4_outputs(6093) <= a;
    layer4_outputs(6094) <= a;
    layer4_outputs(6095) <= not (a and b);
    layer4_outputs(6096) <= not a;
    layer4_outputs(6097) <= not (a or b);
    layer4_outputs(6098) <= a;
    layer4_outputs(6099) <= b;
    layer4_outputs(6100) <= not (a or b);
    layer4_outputs(6101) <= not b;
    layer4_outputs(6102) <= not (a xor b);
    layer4_outputs(6103) <= a xor b;
    layer4_outputs(6104) <= not (a xor b);
    layer4_outputs(6105) <= a xor b;
    layer4_outputs(6106) <= not b or a;
    layer4_outputs(6107) <= not b or a;
    layer4_outputs(6108) <= not b;
    layer4_outputs(6109) <= a xor b;
    layer4_outputs(6110) <= a and not b;
    layer4_outputs(6111) <= a and b;
    layer4_outputs(6112) <= b;
    layer4_outputs(6113) <= not (a or b);
    layer4_outputs(6114) <= a or b;
    layer4_outputs(6115) <= b and not a;
    layer4_outputs(6116) <= a or b;
    layer4_outputs(6117) <= a;
    layer4_outputs(6118) <= a;
    layer4_outputs(6119) <= a or b;
    layer4_outputs(6120) <= not (a and b);
    layer4_outputs(6121) <= a and not b;
    layer4_outputs(6122) <= a;
    layer4_outputs(6123) <= not (a xor b);
    layer4_outputs(6124) <= b;
    layer4_outputs(6125) <= not a;
    layer4_outputs(6126) <= a xor b;
    layer4_outputs(6127) <= a or b;
    layer4_outputs(6128) <= not a;
    layer4_outputs(6129) <= not b or a;
    layer4_outputs(6130) <= not a or b;
    layer4_outputs(6131) <= a or b;
    layer4_outputs(6132) <= a and not b;
    layer4_outputs(6133) <= b;
    layer4_outputs(6134) <= a;
    layer4_outputs(6135) <= a;
    layer4_outputs(6136) <= not b or a;
    layer4_outputs(6137) <= b and not a;
    layer4_outputs(6138) <= a;
    layer4_outputs(6139) <= not b or a;
    layer4_outputs(6140) <= not (a and b);
    layer4_outputs(6141) <= b;
    layer4_outputs(6142) <= not b or a;
    layer4_outputs(6143) <= not a;
    layer4_outputs(6144) <= a xor b;
    layer4_outputs(6145) <= not b or a;
    layer4_outputs(6146) <= not a;
    layer4_outputs(6147) <= a;
    layer4_outputs(6148) <= not (a or b);
    layer4_outputs(6149) <= '1';
    layer4_outputs(6150) <= not (a and b);
    layer4_outputs(6151) <= b and not a;
    layer4_outputs(6152) <= not b;
    layer4_outputs(6153) <= not a or b;
    layer4_outputs(6154) <= not b or a;
    layer4_outputs(6155) <= a or b;
    layer4_outputs(6156) <= not a;
    layer4_outputs(6157) <= a and not b;
    layer4_outputs(6158) <= not (a and b);
    layer4_outputs(6159) <= a and b;
    layer4_outputs(6160) <= a xor b;
    layer4_outputs(6161) <= a or b;
    layer4_outputs(6162) <= not (a and b);
    layer4_outputs(6163) <= not (a or b);
    layer4_outputs(6164) <= not b;
    layer4_outputs(6165) <= a and b;
    layer4_outputs(6166) <= not b or a;
    layer4_outputs(6167) <= a and b;
    layer4_outputs(6168) <= not b or a;
    layer4_outputs(6169) <= not (a xor b);
    layer4_outputs(6170) <= not (a or b);
    layer4_outputs(6171) <= not (a xor b);
    layer4_outputs(6172) <= b;
    layer4_outputs(6173) <= not (a and b);
    layer4_outputs(6174) <= b;
    layer4_outputs(6175) <= a;
    layer4_outputs(6176) <= not (a or b);
    layer4_outputs(6177) <= not (a xor b);
    layer4_outputs(6178) <= a xor b;
    layer4_outputs(6179) <= not b;
    layer4_outputs(6180) <= not b or a;
    layer4_outputs(6181) <= not b;
    layer4_outputs(6182) <= b;
    layer4_outputs(6183) <= a and not b;
    layer4_outputs(6184) <= not (a and b);
    layer4_outputs(6185) <= not a;
    layer4_outputs(6186) <= b;
    layer4_outputs(6187) <= not (a or b);
    layer4_outputs(6188) <= b;
    layer4_outputs(6189) <= not a;
    layer4_outputs(6190) <= not a;
    layer4_outputs(6191) <= not b or a;
    layer4_outputs(6192) <= not (a or b);
    layer4_outputs(6193) <= not b;
    layer4_outputs(6194) <= b and not a;
    layer4_outputs(6195) <= a and b;
    layer4_outputs(6196) <= b and not a;
    layer4_outputs(6197) <= not a;
    layer4_outputs(6198) <= not a;
    layer4_outputs(6199) <= not a;
    layer4_outputs(6200) <= not (a or b);
    layer4_outputs(6201) <= not a;
    layer4_outputs(6202) <= not b;
    layer4_outputs(6203) <= a and not b;
    layer4_outputs(6204) <= not a;
    layer4_outputs(6205) <= a;
    layer4_outputs(6206) <= '1';
    layer4_outputs(6207) <= b and not a;
    layer4_outputs(6208) <= not b;
    layer4_outputs(6209) <= b and not a;
    layer4_outputs(6210) <= '1';
    layer4_outputs(6211) <= not a;
    layer4_outputs(6212) <= b and not a;
    layer4_outputs(6213) <= not a;
    layer4_outputs(6214) <= not (a and b);
    layer4_outputs(6215) <= a or b;
    layer4_outputs(6216) <= a and not b;
    layer4_outputs(6217) <= not b;
    layer4_outputs(6218) <= not a;
    layer4_outputs(6219) <= not (a and b);
    layer4_outputs(6220) <= not a or b;
    layer4_outputs(6221) <= b;
    layer4_outputs(6222) <= a or b;
    layer4_outputs(6223) <= not a or b;
    layer4_outputs(6224) <= a and b;
    layer4_outputs(6225) <= a or b;
    layer4_outputs(6226) <= a and not b;
    layer4_outputs(6227) <= '0';
    layer4_outputs(6228) <= not (a or b);
    layer4_outputs(6229) <= b;
    layer4_outputs(6230) <= a;
    layer4_outputs(6231) <= a and not b;
    layer4_outputs(6232) <= not b or a;
    layer4_outputs(6233) <= not a or b;
    layer4_outputs(6234) <= a;
    layer4_outputs(6235) <= not a or b;
    layer4_outputs(6236) <= a and not b;
    layer4_outputs(6237) <= not a;
    layer4_outputs(6238) <= not b;
    layer4_outputs(6239) <= not b;
    layer4_outputs(6240) <= not (a or b);
    layer4_outputs(6241) <= not a;
    layer4_outputs(6242) <= not b or a;
    layer4_outputs(6243) <= not a;
    layer4_outputs(6244) <= not (a xor b);
    layer4_outputs(6245) <= not b or a;
    layer4_outputs(6246) <= not a;
    layer4_outputs(6247) <= a;
    layer4_outputs(6248) <= not (a or b);
    layer4_outputs(6249) <= b and not a;
    layer4_outputs(6250) <= a xor b;
    layer4_outputs(6251) <= not b;
    layer4_outputs(6252) <= b and not a;
    layer4_outputs(6253) <= not b;
    layer4_outputs(6254) <= a xor b;
    layer4_outputs(6255) <= a;
    layer4_outputs(6256) <= not b;
    layer4_outputs(6257) <= a xor b;
    layer4_outputs(6258) <= not b;
    layer4_outputs(6259) <= a and b;
    layer4_outputs(6260) <= not a;
    layer4_outputs(6261) <= b;
    layer4_outputs(6262) <= '0';
    layer4_outputs(6263) <= '0';
    layer4_outputs(6264) <= a;
    layer4_outputs(6265) <= not (a xor b);
    layer4_outputs(6266) <= not a;
    layer4_outputs(6267) <= not a;
    layer4_outputs(6268) <= b and not a;
    layer4_outputs(6269) <= a or b;
    layer4_outputs(6270) <= not b;
    layer4_outputs(6271) <= b and not a;
    layer4_outputs(6272) <= a or b;
    layer4_outputs(6273) <= a and not b;
    layer4_outputs(6274) <= a;
    layer4_outputs(6275) <= a and not b;
    layer4_outputs(6276) <= a and b;
    layer4_outputs(6277) <= a xor b;
    layer4_outputs(6278) <= not (a xor b);
    layer4_outputs(6279) <= not a or b;
    layer4_outputs(6280) <= not b;
    layer4_outputs(6281) <= '0';
    layer4_outputs(6282) <= not (a or b);
    layer4_outputs(6283) <= b and not a;
    layer4_outputs(6284) <= b;
    layer4_outputs(6285) <= not b;
    layer4_outputs(6286) <= b;
    layer4_outputs(6287) <= a or b;
    layer4_outputs(6288) <= not (a or b);
    layer4_outputs(6289) <= not a;
    layer4_outputs(6290) <= b;
    layer4_outputs(6291) <= a or b;
    layer4_outputs(6292) <= a xor b;
    layer4_outputs(6293) <= not a;
    layer4_outputs(6294) <= not a or b;
    layer4_outputs(6295) <= a;
    layer4_outputs(6296) <= a;
    layer4_outputs(6297) <= '0';
    layer4_outputs(6298) <= not a;
    layer4_outputs(6299) <= not (a or b);
    layer4_outputs(6300) <= not (a or b);
    layer4_outputs(6301) <= b;
    layer4_outputs(6302) <= a;
    layer4_outputs(6303) <= not a;
    layer4_outputs(6304) <= a and b;
    layer4_outputs(6305) <= a;
    layer4_outputs(6306) <= b;
    layer4_outputs(6307) <= '0';
    layer4_outputs(6308) <= not a;
    layer4_outputs(6309) <= not b;
    layer4_outputs(6310) <= not a;
    layer4_outputs(6311) <= '0';
    layer4_outputs(6312) <= a and not b;
    layer4_outputs(6313) <= not b;
    layer4_outputs(6314) <= a or b;
    layer4_outputs(6315) <= a or b;
    layer4_outputs(6316) <= '0';
    layer4_outputs(6317) <= not (a or b);
    layer4_outputs(6318) <= b;
    layer4_outputs(6319) <= a and not b;
    layer4_outputs(6320) <= not (a and b);
    layer4_outputs(6321) <= b;
    layer4_outputs(6322) <= a;
    layer4_outputs(6323) <= a;
    layer4_outputs(6324) <= not a or b;
    layer4_outputs(6325) <= not (a or b);
    layer4_outputs(6326) <= not b;
    layer4_outputs(6327) <= not (a and b);
    layer4_outputs(6328) <= not b;
    layer4_outputs(6329) <= b and not a;
    layer4_outputs(6330) <= not a;
    layer4_outputs(6331) <= b;
    layer4_outputs(6332) <= b;
    layer4_outputs(6333) <= a and not b;
    layer4_outputs(6334) <= b;
    layer4_outputs(6335) <= a and not b;
    layer4_outputs(6336) <= not a;
    layer4_outputs(6337) <= not (a and b);
    layer4_outputs(6338) <= b;
    layer4_outputs(6339) <= b;
    layer4_outputs(6340) <= not (a and b);
    layer4_outputs(6341) <= not (a and b);
    layer4_outputs(6342) <= b;
    layer4_outputs(6343) <= not a;
    layer4_outputs(6344) <= not b;
    layer4_outputs(6345) <= b and not a;
    layer4_outputs(6346) <= not b or a;
    layer4_outputs(6347) <= a xor b;
    layer4_outputs(6348) <= not b;
    layer4_outputs(6349) <= a and b;
    layer4_outputs(6350) <= not b or a;
    layer4_outputs(6351) <= b;
    layer4_outputs(6352) <= b;
    layer4_outputs(6353) <= not (a or b);
    layer4_outputs(6354) <= a or b;
    layer4_outputs(6355) <= a xor b;
    layer4_outputs(6356) <= not a or b;
    layer4_outputs(6357) <= b;
    layer4_outputs(6358) <= a xor b;
    layer4_outputs(6359) <= a;
    layer4_outputs(6360) <= b and not a;
    layer4_outputs(6361) <= a;
    layer4_outputs(6362) <= a or b;
    layer4_outputs(6363) <= '0';
    layer4_outputs(6364) <= b;
    layer4_outputs(6365) <= not a;
    layer4_outputs(6366) <= not (a xor b);
    layer4_outputs(6367) <= not a or b;
    layer4_outputs(6368) <= not a;
    layer4_outputs(6369) <= b;
    layer4_outputs(6370) <= not b or a;
    layer4_outputs(6371) <= b;
    layer4_outputs(6372) <= b;
    layer4_outputs(6373) <= a xor b;
    layer4_outputs(6374) <= a xor b;
    layer4_outputs(6375) <= not b or a;
    layer4_outputs(6376) <= not a;
    layer4_outputs(6377) <= a or b;
    layer4_outputs(6378) <= b and not a;
    layer4_outputs(6379) <= not b;
    layer4_outputs(6380) <= b;
    layer4_outputs(6381) <= not a;
    layer4_outputs(6382) <= b;
    layer4_outputs(6383) <= a xor b;
    layer4_outputs(6384) <= b;
    layer4_outputs(6385) <= a xor b;
    layer4_outputs(6386) <= not (a xor b);
    layer4_outputs(6387) <= not (a and b);
    layer4_outputs(6388) <= not b;
    layer4_outputs(6389) <= b;
    layer4_outputs(6390) <= a;
    layer4_outputs(6391) <= b;
    layer4_outputs(6392) <= not (a and b);
    layer4_outputs(6393) <= not a;
    layer4_outputs(6394) <= not (a and b);
    layer4_outputs(6395) <= b;
    layer4_outputs(6396) <= not b;
    layer4_outputs(6397) <= not a;
    layer4_outputs(6398) <= not a;
    layer4_outputs(6399) <= not (a or b);
    layer4_outputs(6400) <= not a;
    layer4_outputs(6401) <= not b;
    layer4_outputs(6402) <= not a;
    layer4_outputs(6403) <= a;
    layer4_outputs(6404) <= not b or a;
    layer4_outputs(6405) <= b and not a;
    layer4_outputs(6406) <= not b or a;
    layer4_outputs(6407) <= not b or a;
    layer4_outputs(6408) <= '1';
    layer4_outputs(6409) <= a;
    layer4_outputs(6410) <= a;
    layer4_outputs(6411) <= a;
    layer4_outputs(6412) <= not b;
    layer4_outputs(6413) <= not b or a;
    layer4_outputs(6414) <= not a;
    layer4_outputs(6415) <= not b or a;
    layer4_outputs(6416) <= not a or b;
    layer4_outputs(6417) <= a xor b;
    layer4_outputs(6418) <= not a;
    layer4_outputs(6419) <= a and b;
    layer4_outputs(6420) <= b and not a;
    layer4_outputs(6421) <= a;
    layer4_outputs(6422) <= a and not b;
    layer4_outputs(6423) <= a or b;
    layer4_outputs(6424) <= not (a and b);
    layer4_outputs(6425) <= b and not a;
    layer4_outputs(6426) <= a xor b;
    layer4_outputs(6427) <= not a;
    layer4_outputs(6428) <= b;
    layer4_outputs(6429) <= not (a or b);
    layer4_outputs(6430) <= b;
    layer4_outputs(6431) <= a;
    layer4_outputs(6432) <= a and not b;
    layer4_outputs(6433) <= a;
    layer4_outputs(6434) <= not a;
    layer4_outputs(6435) <= a or b;
    layer4_outputs(6436) <= a;
    layer4_outputs(6437) <= not a;
    layer4_outputs(6438) <= a;
    layer4_outputs(6439) <= not (a and b);
    layer4_outputs(6440) <= a;
    layer4_outputs(6441) <= b;
    layer4_outputs(6442) <= a;
    layer4_outputs(6443) <= a and not b;
    layer4_outputs(6444) <= '0';
    layer4_outputs(6445) <= not (a xor b);
    layer4_outputs(6446) <= not a;
    layer4_outputs(6447) <= a and b;
    layer4_outputs(6448) <= not (a and b);
    layer4_outputs(6449) <= not a or b;
    layer4_outputs(6450) <= not a;
    layer4_outputs(6451) <= b;
    layer4_outputs(6452) <= not b;
    layer4_outputs(6453) <= a;
    layer4_outputs(6454) <= b and not a;
    layer4_outputs(6455) <= a;
    layer4_outputs(6456) <= not (a and b);
    layer4_outputs(6457) <= not (a xor b);
    layer4_outputs(6458) <= b and not a;
    layer4_outputs(6459) <= not b;
    layer4_outputs(6460) <= not a;
    layer4_outputs(6461) <= not b;
    layer4_outputs(6462) <= not b or a;
    layer4_outputs(6463) <= not a or b;
    layer4_outputs(6464) <= not a or b;
    layer4_outputs(6465) <= not (a and b);
    layer4_outputs(6466) <= b;
    layer4_outputs(6467) <= not b;
    layer4_outputs(6468) <= not b;
    layer4_outputs(6469) <= not a;
    layer4_outputs(6470) <= a and not b;
    layer4_outputs(6471) <= not a;
    layer4_outputs(6472) <= a;
    layer4_outputs(6473) <= a and b;
    layer4_outputs(6474) <= not b;
    layer4_outputs(6475) <= not (a and b);
    layer4_outputs(6476) <= a or b;
    layer4_outputs(6477) <= not a or b;
    layer4_outputs(6478) <= b;
    layer4_outputs(6479) <= not (a xor b);
    layer4_outputs(6480) <= b;
    layer4_outputs(6481) <= not b;
    layer4_outputs(6482) <= not (a xor b);
    layer4_outputs(6483) <= a;
    layer4_outputs(6484) <= a;
    layer4_outputs(6485) <= a and b;
    layer4_outputs(6486) <= not (a xor b);
    layer4_outputs(6487) <= b;
    layer4_outputs(6488) <= not b;
    layer4_outputs(6489) <= not a or b;
    layer4_outputs(6490) <= not b;
    layer4_outputs(6491) <= a and b;
    layer4_outputs(6492) <= not a;
    layer4_outputs(6493) <= not a;
    layer4_outputs(6494) <= not a;
    layer4_outputs(6495) <= a;
    layer4_outputs(6496) <= not a or b;
    layer4_outputs(6497) <= a;
    layer4_outputs(6498) <= not b;
    layer4_outputs(6499) <= not (a xor b);
    layer4_outputs(6500) <= a and not b;
    layer4_outputs(6501) <= a and b;
    layer4_outputs(6502) <= not b;
    layer4_outputs(6503) <= a and b;
    layer4_outputs(6504) <= a xor b;
    layer4_outputs(6505) <= b;
    layer4_outputs(6506) <= not a or b;
    layer4_outputs(6507) <= not b;
    layer4_outputs(6508) <= not a;
    layer4_outputs(6509) <= a or b;
    layer4_outputs(6510) <= not b or a;
    layer4_outputs(6511) <= not a;
    layer4_outputs(6512) <= not (a or b);
    layer4_outputs(6513) <= '1';
    layer4_outputs(6514) <= not b or a;
    layer4_outputs(6515) <= not (a and b);
    layer4_outputs(6516) <= '0';
    layer4_outputs(6517) <= b and not a;
    layer4_outputs(6518) <= not a;
    layer4_outputs(6519) <= not b or a;
    layer4_outputs(6520) <= b and not a;
    layer4_outputs(6521) <= not (a or b);
    layer4_outputs(6522) <= a and b;
    layer4_outputs(6523) <= not (a and b);
    layer4_outputs(6524) <= not a or b;
    layer4_outputs(6525) <= b;
    layer4_outputs(6526) <= not (a or b);
    layer4_outputs(6527) <= not b or a;
    layer4_outputs(6528) <= not b;
    layer4_outputs(6529) <= not a;
    layer4_outputs(6530) <= '0';
    layer4_outputs(6531) <= not b;
    layer4_outputs(6532) <= '0';
    layer4_outputs(6533) <= not a or b;
    layer4_outputs(6534) <= b and not a;
    layer4_outputs(6535) <= b and not a;
    layer4_outputs(6536) <= '1';
    layer4_outputs(6537) <= b;
    layer4_outputs(6538) <= b;
    layer4_outputs(6539) <= '0';
    layer4_outputs(6540) <= not (a xor b);
    layer4_outputs(6541) <= a and not b;
    layer4_outputs(6542) <= not (a or b);
    layer4_outputs(6543) <= a or b;
    layer4_outputs(6544) <= not a or b;
    layer4_outputs(6545) <= a and not b;
    layer4_outputs(6546) <= not a;
    layer4_outputs(6547) <= a;
    layer4_outputs(6548) <= b;
    layer4_outputs(6549) <= '0';
    layer4_outputs(6550) <= a and not b;
    layer4_outputs(6551) <= a;
    layer4_outputs(6552) <= '0';
    layer4_outputs(6553) <= a;
    layer4_outputs(6554) <= b;
    layer4_outputs(6555) <= not (a and b);
    layer4_outputs(6556) <= a;
    layer4_outputs(6557) <= a and not b;
    layer4_outputs(6558) <= b and not a;
    layer4_outputs(6559) <= a and not b;
    layer4_outputs(6560) <= not (a or b);
    layer4_outputs(6561) <= a or b;
    layer4_outputs(6562) <= not a;
    layer4_outputs(6563) <= a and not b;
    layer4_outputs(6564) <= '1';
    layer4_outputs(6565) <= not b;
    layer4_outputs(6566) <= a and b;
    layer4_outputs(6567) <= a;
    layer4_outputs(6568) <= b;
    layer4_outputs(6569) <= a xor b;
    layer4_outputs(6570) <= '1';
    layer4_outputs(6571) <= not b or a;
    layer4_outputs(6572) <= not (a or b);
    layer4_outputs(6573) <= not (a xor b);
    layer4_outputs(6574) <= a or b;
    layer4_outputs(6575) <= not b or a;
    layer4_outputs(6576) <= not b or a;
    layer4_outputs(6577) <= b;
    layer4_outputs(6578) <= not a or b;
    layer4_outputs(6579) <= a;
    layer4_outputs(6580) <= not a;
    layer4_outputs(6581) <= not b;
    layer4_outputs(6582) <= b;
    layer4_outputs(6583) <= not (a or b);
    layer4_outputs(6584) <= a and b;
    layer4_outputs(6585) <= not (a and b);
    layer4_outputs(6586) <= not b;
    layer4_outputs(6587) <= not a or b;
    layer4_outputs(6588) <= a;
    layer4_outputs(6589) <= not b;
    layer4_outputs(6590) <= b and not a;
    layer4_outputs(6591) <= not a;
    layer4_outputs(6592) <= not b;
    layer4_outputs(6593) <= not (a and b);
    layer4_outputs(6594) <= not (a xor b);
    layer4_outputs(6595) <= not (a and b);
    layer4_outputs(6596) <= b;
    layer4_outputs(6597) <= a;
    layer4_outputs(6598) <= not a or b;
    layer4_outputs(6599) <= not b;
    layer4_outputs(6600) <= not a;
    layer4_outputs(6601) <= a or b;
    layer4_outputs(6602) <= b and not a;
    layer4_outputs(6603) <= not (a or b);
    layer4_outputs(6604) <= not b or a;
    layer4_outputs(6605) <= a xor b;
    layer4_outputs(6606) <= a xor b;
    layer4_outputs(6607) <= a or b;
    layer4_outputs(6608) <= not b;
    layer4_outputs(6609) <= not (a and b);
    layer4_outputs(6610) <= a xor b;
    layer4_outputs(6611) <= not (a or b);
    layer4_outputs(6612) <= not a;
    layer4_outputs(6613) <= not (a and b);
    layer4_outputs(6614) <= not (a and b);
    layer4_outputs(6615) <= b;
    layer4_outputs(6616) <= not a;
    layer4_outputs(6617) <= a;
    layer4_outputs(6618) <= not a;
    layer4_outputs(6619) <= a;
    layer4_outputs(6620) <= not a;
    layer4_outputs(6621) <= not (a and b);
    layer4_outputs(6622) <= a or b;
    layer4_outputs(6623) <= b;
    layer4_outputs(6624) <= a and not b;
    layer4_outputs(6625) <= not (a and b);
    layer4_outputs(6626) <= b and not a;
    layer4_outputs(6627) <= not a;
    layer4_outputs(6628) <= b;
    layer4_outputs(6629) <= b;
    layer4_outputs(6630) <= not a;
    layer4_outputs(6631) <= not b;
    layer4_outputs(6632) <= not a or b;
    layer4_outputs(6633) <= not a;
    layer4_outputs(6634) <= a and b;
    layer4_outputs(6635) <= not a or b;
    layer4_outputs(6636) <= not b;
    layer4_outputs(6637) <= a;
    layer4_outputs(6638) <= b and not a;
    layer4_outputs(6639) <= not (a or b);
    layer4_outputs(6640) <= not (a or b);
    layer4_outputs(6641) <= '0';
    layer4_outputs(6642) <= '0';
    layer4_outputs(6643) <= not b or a;
    layer4_outputs(6644) <= not (a and b);
    layer4_outputs(6645) <= not (a or b);
    layer4_outputs(6646) <= a;
    layer4_outputs(6647) <= '0';
    layer4_outputs(6648) <= a and b;
    layer4_outputs(6649) <= b;
    layer4_outputs(6650) <= a and not b;
    layer4_outputs(6651) <= a xor b;
    layer4_outputs(6652) <= a and not b;
    layer4_outputs(6653) <= not a;
    layer4_outputs(6654) <= not a or b;
    layer4_outputs(6655) <= b and not a;
    layer4_outputs(6656) <= b and not a;
    layer4_outputs(6657) <= not a;
    layer4_outputs(6658) <= a xor b;
    layer4_outputs(6659) <= a and b;
    layer4_outputs(6660) <= b and not a;
    layer4_outputs(6661) <= not b or a;
    layer4_outputs(6662) <= not a or b;
    layer4_outputs(6663) <= a or b;
    layer4_outputs(6664) <= not a or b;
    layer4_outputs(6665) <= a and not b;
    layer4_outputs(6666) <= not b;
    layer4_outputs(6667) <= not b;
    layer4_outputs(6668) <= b and not a;
    layer4_outputs(6669) <= a and b;
    layer4_outputs(6670) <= not a;
    layer4_outputs(6671) <= b;
    layer4_outputs(6672) <= b;
    layer4_outputs(6673) <= a and not b;
    layer4_outputs(6674) <= not b or a;
    layer4_outputs(6675) <= b and not a;
    layer4_outputs(6676) <= a or b;
    layer4_outputs(6677) <= not (a xor b);
    layer4_outputs(6678) <= a;
    layer4_outputs(6679) <= a xor b;
    layer4_outputs(6680) <= not a;
    layer4_outputs(6681) <= not (a and b);
    layer4_outputs(6682) <= '0';
    layer4_outputs(6683) <= not (a or b);
    layer4_outputs(6684) <= a;
    layer4_outputs(6685) <= not b or a;
    layer4_outputs(6686) <= not b or a;
    layer4_outputs(6687) <= a xor b;
    layer4_outputs(6688) <= b;
    layer4_outputs(6689) <= b;
    layer4_outputs(6690) <= not a;
    layer4_outputs(6691) <= '1';
    layer4_outputs(6692) <= not b;
    layer4_outputs(6693) <= not b;
    layer4_outputs(6694) <= a;
    layer4_outputs(6695) <= a;
    layer4_outputs(6696) <= not (a xor b);
    layer4_outputs(6697) <= b;
    layer4_outputs(6698) <= a xor b;
    layer4_outputs(6699) <= not a or b;
    layer4_outputs(6700) <= b and not a;
    layer4_outputs(6701) <= not b;
    layer4_outputs(6702) <= not (a xor b);
    layer4_outputs(6703) <= '0';
    layer4_outputs(6704) <= b;
    layer4_outputs(6705) <= not (a and b);
    layer4_outputs(6706) <= not (a or b);
    layer4_outputs(6707) <= not a;
    layer4_outputs(6708) <= not (a xor b);
    layer4_outputs(6709) <= b;
    layer4_outputs(6710) <= a;
    layer4_outputs(6711) <= not a or b;
    layer4_outputs(6712) <= b and not a;
    layer4_outputs(6713) <= a xor b;
    layer4_outputs(6714) <= b;
    layer4_outputs(6715) <= not (a xor b);
    layer4_outputs(6716) <= a or b;
    layer4_outputs(6717) <= a and not b;
    layer4_outputs(6718) <= not b or a;
    layer4_outputs(6719) <= a or b;
    layer4_outputs(6720) <= b;
    layer4_outputs(6721) <= not (a and b);
    layer4_outputs(6722) <= a and b;
    layer4_outputs(6723) <= b;
    layer4_outputs(6724) <= b and not a;
    layer4_outputs(6725) <= not (a xor b);
    layer4_outputs(6726) <= not (a or b);
    layer4_outputs(6727) <= a;
    layer4_outputs(6728) <= '1';
    layer4_outputs(6729) <= not b;
    layer4_outputs(6730) <= not b or a;
    layer4_outputs(6731) <= not (a or b);
    layer4_outputs(6732) <= a and not b;
    layer4_outputs(6733) <= '1';
    layer4_outputs(6734) <= not b;
    layer4_outputs(6735) <= not (a or b);
    layer4_outputs(6736) <= not a;
    layer4_outputs(6737) <= b;
    layer4_outputs(6738) <= '0';
    layer4_outputs(6739) <= a and b;
    layer4_outputs(6740) <= not (a or b);
    layer4_outputs(6741) <= a or b;
    layer4_outputs(6742) <= not (a and b);
    layer4_outputs(6743) <= a and not b;
    layer4_outputs(6744) <= a or b;
    layer4_outputs(6745) <= a and b;
    layer4_outputs(6746) <= a and b;
    layer4_outputs(6747) <= a;
    layer4_outputs(6748) <= not (a xor b);
    layer4_outputs(6749) <= a and b;
    layer4_outputs(6750) <= a or b;
    layer4_outputs(6751) <= not b;
    layer4_outputs(6752) <= a and b;
    layer4_outputs(6753) <= not b or a;
    layer4_outputs(6754) <= a xor b;
    layer4_outputs(6755) <= not b;
    layer4_outputs(6756) <= a and b;
    layer4_outputs(6757) <= not a or b;
    layer4_outputs(6758) <= not (a or b);
    layer4_outputs(6759) <= b and not a;
    layer4_outputs(6760) <= not b or a;
    layer4_outputs(6761) <= b;
    layer4_outputs(6762) <= a;
    layer4_outputs(6763) <= not b;
    layer4_outputs(6764) <= not (a xor b);
    layer4_outputs(6765) <= a and b;
    layer4_outputs(6766) <= not (a or b);
    layer4_outputs(6767) <= '1';
    layer4_outputs(6768) <= a and b;
    layer4_outputs(6769) <= '0';
    layer4_outputs(6770) <= not a;
    layer4_outputs(6771) <= a and not b;
    layer4_outputs(6772) <= not (a xor b);
    layer4_outputs(6773) <= b;
    layer4_outputs(6774) <= not (a xor b);
    layer4_outputs(6775) <= not b;
    layer4_outputs(6776) <= not a;
    layer4_outputs(6777) <= a and not b;
    layer4_outputs(6778) <= b and not a;
    layer4_outputs(6779) <= not b or a;
    layer4_outputs(6780) <= a and not b;
    layer4_outputs(6781) <= a and not b;
    layer4_outputs(6782) <= not (a xor b);
    layer4_outputs(6783) <= a or b;
    layer4_outputs(6784) <= b and not a;
    layer4_outputs(6785) <= not (a xor b);
    layer4_outputs(6786) <= not a;
    layer4_outputs(6787) <= not (a and b);
    layer4_outputs(6788) <= a xor b;
    layer4_outputs(6789) <= b;
    layer4_outputs(6790) <= not (a or b);
    layer4_outputs(6791) <= not (a or b);
    layer4_outputs(6792) <= not b;
    layer4_outputs(6793) <= a or b;
    layer4_outputs(6794) <= not (a xor b);
    layer4_outputs(6795) <= not a;
    layer4_outputs(6796) <= not b;
    layer4_outputs(6797) <= not a;
    layer4_outputs(6798) <= not a;
    layer4_outputs(6799) <= not b or a;
    layer4_outputs(6800) <= a;
    layer4_outputs(6801) <= a or b;
    layer4_outputs(6802) <= '0';
    layer4_outputs(6803) <= not a or b;
    layer4_outputs(6804) <= not b or a;
    layer4_outputs(6805) <= not b;
    layer4_outputs(6806) <= '0';
    layer4_outputs(6807) <= a;
    layer4_outputs(6808) <= a or b;
    layer4_outputs(6809) <= not a;
    layer4_outputs(6810) <= not (a xor b);
    layer4_outputs(6811) <= a;
    layer4_outputs(6812) <= a xor b;
    layer4_outputs(6813) <= a;
    layer4_outputs(6814) <= a;
    layer4_outputs(6815) <= a or b;
    layer4_outputs(6816) <= a;
    layer4_outputs(6817) <= not b;
    layer4_outputs(6818) <= not b;
    layer4_outputs(6819) <= '0';
    layer4_outputs(6820) <= not a;
    layer4_outputs(6821) <= a or b;
    layer4_outputs(6822) <= b;
    layer4_outputs(6823) <= b;
    layer4_outputs(6824) <= a or b;
    layer4_outputs(6825) <= '1';
    layer4_outputs(6826) <= not (a xor b);
    layer4_outputs(6827) <= not b;
    layer4_outputs(6828) <= b and not a;
    layer4_outputs(6829) <= not b;
    layer4_outputs(6830) <= a;
    layer4_outputs(6831) <= not b;
    layer4_outputs(6832) <= a and not b;
    layer4_outputs(6833) <= a;
    layer4_outputs(6834) <= b and not a;
    layer4_outputs(6835) <= '1';
    layer4_outputs(6836) <= b;
    layer4_outputs(6837) <= a and not b;
    layer4_outputs(6838) <= not a or b;
    layer4_outputs(6839) <= a;
    layer4_outputs(6840) <= not a;
    layer4_outputs(6841) <= not (a or b);
    layer4_outputs(6842) <= not a or b;
    layer4_outputs(6843) <= not a or b;
    layer4_outputs(6844) <= a and not b;
    layer4_outputs(6845) <= not b;
    layer4_outputs(6846) <= b;
    layer4_outputs(6847) <= not a or b;
    layer4_outputs(6848) <= '1';
    layer4_outputs(6849) <= b;
    layer4_outputs(6850) <= a and not b;
    layer4_outputs(6851) <= a and not b;
    layer4_outputs(6852) <= not b or a;
    layer4_outputs(6853) <= a and b;
    layer4_outputs(6854) <= not a;
    layer4_outputs(6855) <= a;
    layer4_outputs(6856) <= '0';
    layer4_outputs(6857) <= not b or a;
    layer4_outputs(6858) <= b and not a;
    layer4_outputs(6859) <= b and not a;
    layer4_outputs(6860) <= not b;
    layer4_outputs(6861) <= not a or b;
    layer4_outputs(6862) <= not b;
    layer4_outputs(6863) <= a and not b;
    layer4_outputs(6864) <= b;
    layer4_outputs(6865) <= '1';
    layer4_outputs(6866) <= not a or b;
    layer4_outputs(6867) <= not a;
    layer4_outputs(6868) <= a;
    layer4_outputs(6869) <= a;
    layer4_outputs(6870) <= not b;
    layer4_outputs(6871) <= a xor b;
    layer4_outputs(6872) <= not (a or b);
    layer4_outputs(6873) <= a xor b;
    layer4_outputs(6874) <= a;
    layer4_outputs(6875) <= a and not b;
    layer4_outputs(6876) <= a;
    layer4_outputs(6877) <= not a;
    layer4_outputs(6878) <= not a;
    layer4_outputs(6879) <= not a;
    layer4_outputs(6880) <= a xor b;
    layer4_outputs(6881) <= a and not b;
    layer4_outputs(6882) <= not b;
    layer4_outputs(6883) <= b;
    layer4_outputs(6884) <= a;
    layer4_outputs(6885) <= not (a and b);
    layer4_outputs(6886) <= '1';
    layer4_outputs(6887) <= '0';
    layer4_outputs(6888) <= a;
    layer4_outputs(6889) <= not a or b;
    layer4_outputs(6890) <= not (a and b);
    layer4_outputs(6891) <= a;
    layer4_outputs(6892) <= a xor b;
    layer4_outputs(6893) <= not a;
    layer4_outputs(6894) <= a and not b;
    layer4_outputs(6895) <= b;
    layer4_outputs(6896) <= a and b;
    layer4_outputs(6897) <= b;
    layer4_outputs(6898) <= a;
    layer4_outputs(6899) <= not (a xor b);
    layer4_outputs(6900) <= not (a or b);
    layer4_outputs(6901) <= a and not b;
    layer4_outputs(6902) <= a xor b;
    layer4_outputs(6903) <= a xor b;
    layer4_outputs(6904) <= not a;
    layer4_outputs(6905) <= not b or a;
    layer4_outputs(6906) <= a and not b;
    layer4_outputs(6907) <= b;
    layer4_outputs(6908) <= not a;
    layer4_outputs(6909) <= not b;
    layer4_outputs(6910) <= a;
    layer4_outputs(6911) <= b and not a;
    layer4_outputs(6912) <= a and not b;
    layer4_outputs(6913) <= a and not b;
    layer4_outputs(6914) <= not a or b;
    layer4_outputs(6915) <= not b or a;
    layer4_outputs(6916) <= not (a or b);
    layer4_outputs(6917) <= a;
    layer4_outputs(6918) <= a and b;
    layer4_outputs(6919) <= not b;
    layer4_outputs(6920) <= b;
    layer4_outputs(6921) <= not b or a;
    layer4_outputs(6922) <= a and not b;
    layer4_outputs(6923) <= a;
    layer4_outputs(6924) <= not a or b;
    layer4_outputs(6925) <= a and not b;
    layer4_outputs(6926) <= b;
    layer4_outputs(6927) <= b and not a;
    layer4_outputs(6928) <= a and b;
    layer4_outputs(6929) <= not a;
    layer4_outputs(6930) <= b;
    layer4_outputs(6931) <= not (a and b);
    layer4_outputs(6932) <= not (a xor b);
    layer4_outputs(6933) <= b;
    layer4_outputs(6934) <= not a;
    layer4_outputs(6935) <= not b or a;
    layer4_outputs(6936) <= a or b;
    layer4_outputs(6937) <= b;
    layer4_outputs(6938) <= b;
    layer4_outputs(6939) <= not (a or b);
    layer4_outputs(6940) <= not (a xor b);
    layer4_outputs(6941) <= a;
    layer4_outputs(6942) <= a;
    layer4_outputs(6943) <= not a;
    layer4_outputs(6944) <= not (a and b);
    layer4_outputs(6945) <= not (a and b);
    layer4_outputs(6946) <= not (a and b);
    layer4_outputs(6947) <= not (a xor b);
    layer4_outputs(6948) <= b;
    layer4_outputs(6949) <= b;
    layer4_outputs(6950) <= not b or a;
    layer4_outputs(6951) <= a;
    layer4_outputs(6952) <= not a;
    layer4_outputs(6953) <= not (a or b);
    layer4_outputs(6954) <= a xor b;
    layer4_outputs(6955) <= a xor b;
    layer4_outputs(6956) <= not b;
    layer4_outputs(6957) <= a;
    layer4_outputs(6958) <= '0';
    layer4_outputs(6959) <= a and not b;
    layer4_outputs(6960) <= a;
    layer4_outputs(6961) <= a;
    layer4_outputs(6962) <= not b;
    layer4_outputs(6963) <= not b or a;
    layer4_outputs(6964) <= not a or b;
    layer4_outputs(6965) <= not (a or b);
    layer4_outputs(6966) <= a or b;
    layer4_outputs(6967) <= not (a xor b);
    layer4_outputs(6968) <= '0';
    layer4_outputs(6969) <= a xor b;
    layer4_outputs(6970) <= not b or a;
    layer4_outputs(6971) <= a and b;
    layer4_outputs(6972) <= not b or a;
    layer4_outputs(6973) <= b and not a;
    layer4_outputs(6974) <= not b or a;
    layer4_outputs(6975) <= a;
    layer4_outputs(6976) <= not b;
    layer4_outputs(6977) <= a xor b;
    layer4_outputs(6978) <= not (a xor b);
    layer4_outputs(6979) <= a;
    layer4_outputs(6980) <= not (a and b);
    layer4_outputs(6981) <= a and b;
    layer4_outputs(6982) <= b and not a;
    layer4_outputs(6983) <= not (a or b);
    layer4_outputs(6984) <= a and b;
    layer4_outputs(6985) <= a xor b;
    layer4_outputs(6986) <= not a;
    layer4_outputs(6987) <= not a or b;
    layer4_outputs(6988) <= not a or b;
    layer4_outputs(6989) <= not (a and b);
    layer4_outputs(6990) <= b and not a;
    layer4_outputs(6991) <= '0';
    layer4_outputs(6992) <= not a or b;
    layer4_outputs(6993) <= not b;
    layer4_outputs(6994) <= '0';
    layer4_outputs(6995) <= b and not a;
    layer4_outputs(6996) <= a xor b;
    layer4_outputs(6997) <= b;
    layer4_outputs(6998) <= b and not a;
    layer4_outputs(6999) <= a;
    layer4_outputs(7000) <= not (a xor b);
    layer4_outputs(7001) <= not b or a;
    layer4_outputs(7002) <= not b or a;
    layer4_outputs(7003) <= a or b;
    layer4_outputs(7004) <= '1';
    layer4_outputs(7005) <= not b;
    layer4_outputs(7006) <= a and b;
    layer4_outputs(7007) <= a xor b;
    layer4_outputs(7008) <= not (a xor b);
    layer4_outputs(7009) <= not b;
    layer4_outputs(7010) <= not b;
    layer4_outputs(7011) <= b and not a;
    layer4_outputs(7012) <= a and b;
    layer4_outputs(7013) <= a;
    layer4_outputs(7014) <= not (a or b);
    layer4_outputs(7015) <= not b;
    layer4_outputs(7016) <= not (a and b);
    layer4_outputs(7017) <= not a or b;
    layer4_outputs(7018) <= not a or b;
    layer4_outputs(7019) <= not b;
    layer4_outputs(7020) <= not a;
    layer4_outputs(7021) <= a or b;
    layer4_outputs(7022) <= not b;
    layer4_outputs(7023) <= not (a or b);
    layer4_outputs(7024) <= a;
    layer4_outputs(7025) <= not b;
    layer4_outputs(7026) <= b;
    layer4_outputs(7027) <= not b;
    layer4_outputs(7028) <= not (a xor b);
    layer4_outputs(7029) <= '1';
    layer4_outputs(7030) <= a;
    layer4_outputs(7031) <= b;
    layer4_outputs(7032) <= not (a xor b);
    layer4_outputs(7033) <= not (a and b);
    layer4_outputs(7034) <= b;
    layer4_outputs(7035) <= a xor b;
    layer4_outputs(7036) <= not (a and b);
    layer4_outputs(7037) <= a xor b;
    layer4_outputs(7038) <= not b;
    layer4_outputs(7039) <= not (a or b);
    layer4_outputs(7040) <= a xor b;
    layer4_outputs(7041) <= not a or b;
    layer4_outputs(7042) <= a or b;
    layer4_outputs(7043) <= a;
    layer4_outputs(7044) <= a;
    layer4_outputs(7045) <= not a;
    layer4_outputs(7046) <= not b;
    layer4_outputs(7047) <= not a;
    layer4_outputs(7048) <= a and b;
    layer4_outputs(7049) <= not (a or b);
    layer4_outputs(7050) <= not (a or b);
    layer4_outputs(7051) <= not b or a;
    layer4_outputs(7052) <= a and b;
    layer4_outputs(7053) <= not (a or b);
    layer4_outputs(7054) <= not a;
    layer4_outputs(7055) <= not b or a;
    layer4_outputs(7056) <= a;
    layer4_outputs(7057) <= b;
    layer4_outputs(7058) <= a xor b;
    layer4_outputs(7059) <= not b or a;
    layer4_outputs(7060) <= a and b;
    layer4_outputs(7061) <= a;
    layer4_outputs(7062) <= a;
    layer4_outputs(7063) <= a xor b;
    layer4_outputs(7064) <= not a;
    layer4_outputs(7065) <= b and not a;
    layer4_outputs(7066) <= a and not b;
    layer4_outputs(7067) <= not b or a;
    layer4_outputs(7068) <= a and not b;
    layer4_outputs(7069) <= '1';
    layer4_outputs(7070) <= a and b;
    layer4_outputs(7071) <= a xor b;
    layer4_outputs(7072) <= not (a xor b);
    layer4_outputs(7073) <= not a or b;
    layer4_outputs(7074) <= not (a xor b);
    layer4_outputs(7075) <= a or b;
    layer4_outputs(7076) <= not b or a;
    layer4_outputs(7077) <= b;
    layer4_outputs(7078) <= not a or b;
    layer4_outputs(7079) <= not b;
    layer4_outputs(7080) <= b;
    layer4_outputs(7081) <= not (a and b);
    layer4_outputs(7082) <= not b;
    layer4_outputs(7083) <= not a or b;
    layer4_outputs(7084) <= a or b;
    layer4_outputs(7085) <= not (a and b);
    layer4_outputs(7086) <= a or b;
    layer4_outputs(7087) <= a xor b;
    layer4_outputs(7088) <= a;
    layer4_outputs(7089) <= not b;
    layer4_outputs(7090) <= a and b;
    layer4_outputs(7091) <= a;
    layer4_outputs(7092) <= b and not a;
    layer4_outputs(7093) <= not a;
    layer4_outputs(7094) <= not (a xor b);
    layer4_outputs(7095) <= '0';
    layer4_outputs(7096) <= a or b;
    layer4_outputs(7097) <= a;
    layer4_outputs(7098) <= not (a and b);
    layer4_outputs(7099) <= not a;
    layer4_outputs(7100) <= not (a and b);
    layer4_outputs(7101) <= not b or a;
    layer4_outputs(7102) <= not b or a;
    layer4_outputs(7103) <= b;
    layer4_outputs(7104) <= not a;
    layer4_outputs(7105) <= not (a xor b);
    layer4_outputs(7106) <= not (a or b);
    layer4_outputs(7107) <= not (a xor b);
    layer4_outputs(7108) <= '0';
    layer4_outputs(7109) <= b and not a;
    layer4_outputs(7110) <= not b;
    layer4_outputs(7111) <= a xor b;
    layer4_outputs(7112) <= not a or b;
    layer4_outputs(7113) <= not (a or b);
    layer4_outputs(7114) <= a or b;
    layer4_outputs(7115) <= not b or a;
    layer4_outputs(7116) <= not a;
    layer4_outputs(7117) <= not a or b;
    layer4_outputs(7118) <= a;
    layer4_outputs(7119) <= not (a xor b);
    layer4_outputs(7120) <= b;
    layer4_outputs(7121) <= not b;
    layer4_outputs(7122) <= not (a xor b);
    layer4_outputs(7123) <= not b;
    layer4_outputs(7124) <= not (a and b);
    layer4_outputs(7125) <= not (a and b);
    layer4_outputs(7126) <= b;
    layer4_outputs(7127) <= b;
    layer4_outputs(7128) <= a and not b;
    layer4_outputs(7129) <= a or b;
    layer4_outputs(7130) <= not a;
    layer4_outputs(7131) <= not b or a;
    layer4_outputs(7132) <= b;
    layer4_outputs(7133) <= '1';
    layer4_outputs(7134) <= not (a or b);
    layer4_outputs(7135) <= '0';
    layer4_outputs(7136) <= not a;
    layer4_outputs(7137) <= a and not b;
    layer4_outputs(7138) <= not a or b;
    layer4_outputs(7139) <= a;
    layer4_outputs(7140) <= not b;
    layer4_outputs(7141) <= a and not b;
    layer4_outputs(7142) <= not a or b;
    layer4_outputs(7143) <= a;
    layer4_outputs(7144) <= not b;
    layer4_outputs(7145) <= a xor b;
    layer4_outputs(7146) <= not a;
    layer4_outputs(7147) <= not (a and b);
    layer4_outputs(7148) <= a or b;
    layer4_outputs(7149) <= a and b;
    layer4_outputs(7150) <= b and not a;
    layer4_outputs(7151) <= not (a xor b);
    layer4_outputs(7152) <= a;
    layer4_outputs(7153) <= not b or a;
    layer4_outputs(7154) <= not a or b;
    layer4_outputs(7155) <= a;
    layer4_outputs(7156) <= not b;
    layer4_outputs(7157) <= not (a and b);
    layer4_outputs(7158) <= not b;
    layer4_outputs(7159) <= not b or a;
    layer4_outputs(7160) <= not (a and b);
    layer4_outputs(7161) <= '1';
    layer4_outputs(7162) <= not b or a;
    layer4_outputs(7163) <= not a;
    layer4_outputs(7164) <= a xor b;
    layer4_outputs(7165) <= a xor b;
    layer4_outputs(7166) <= not b or a;
    layer4_outputs(7167) <= '0';
    layer4_outputs(7168) <= not (a and b);
    layer4_outputs(7169) <= not a or b;
    layer4_outputs(7170) <= a and b;
    layer4_outputs(7171) <= b;
    layer4_outputs(7172) <= a;
    layer4_outputs(7173) <= a and not b;
    layer4_outputs(7174) <= b and not a;
    layer4_outputs(7175) <= not (a and b);
    layer4_outputs(7176) <= not a or b;
    layer4_outputs(7177) <= not a or b;
    layer4_outputs(7178) <= a;
    layer4_outputs(7179) <= '0';
    layer4_outputs(7180) <= b;
    layer4_outputs(7181) <= a or b;
    layer4_outputs(7182) <= not a;
    layer4_outputs(7183) <= not (a or b);
    layer4_outputs(7184) <= a;
    layer4_outputs(7185) <= b;
    layer4_outputs(7186) <= not (a or b);
    layer4_outputs(7187) <= not (a and b);
    layer4_outputs(7188) <= b and not a;
    layer4_outputs(7189) <= not (a and b);
    layer4_outputs(7190) <= a xor b;
    layer4_outputs(7191) <= b and not a;
    layer4_outputs(7192) <= a or b;
    layer4_outputs(7193) <= '0';
    layer4_outputs(7194) <= a or b;
    layer4_outputs(7195) <= a;
    layer4_outputs(7196) <= b and not a;
    layer4_outputs(7197) <= not (a xor b);
    layer4_outputs(7198) <= not a or b;
    layer4_outputs(7199) <= a;
    layer4_outputs(7200) <= not a;
    layer4_outputs(7201) <= a;
    layer4_outputs(7202) <= b and not a;
    layer4_outputs(7203) <= b and not a;
    layer4_outputs(7204) <= not (a xor b);
    layer4_outputs(7205) <= not b;
    layer4_outputs(7206) <= a;
    layer4_outputs(7207) <= a;
    layer4_outputs(7208) <= a and not b;
    layer4_outputs(7209) <= not (a xor b);
    layer4_outputs(7210) <= b;
    layer4_outputs(7211) <= not (a and b);
    layer4_outputs(7212) <= not a;
    layer4_outputs(7213) <= not a or b;
    layer4_outputs(7214) <= a;
    layer4_outputs(7215) <= a xor b;
    layer4_outputs(7216) <= b and not a;
    layer4_outputs(7217) <= a and b;
    layer4_outputs(7218) <= not (a and b);
    layer4_outputs(7219) <= a and not b;
    layer4_outputs(7220) <= b and not a;
    layer4_outputs(7221) <= a;
    layer4_outputs(7222) <= a or b;
    layer4_outputs(7223) <= b;
    layer4_outputs(7224) <= a or b;
    layer4_outputs(7225) <= not (a or b);
    layer4_outputs(7226) <= a or b;
    layer4_outputs(7227) <= not a;
    layer4_outputs(7228) <= a;
    layer4_outputs(7229) <= not a;
    layer4_outputs(7230) <= not (a or b);
    layer4_outputs(7231) <= not a or b;
    layer4_outputs(7232) <= a xor b;
    layer4_outputs(7233) <= a and not b;
    layer4_outputs(7234) <= not b or a;
    layer4_outputs(7235) <= not (a or b);
    layer4_outputs(7236) <= not a or b;
    layer4_outputs(7237) <= a or b;
    layer4_outputs(7238) <= a;
    layer4_outputs(7239) <= a;
    layer4_outputs(7240) <= not a;
    layer4_outputs(7241) <= not b or a;
    layer4_outputs(7242) <= a xor b;
    layer4_outputs(7243) <= a xor b;
    layer4_outputs(7244) <= a and b;
    layer4_outputs(7245) <= b;
    layer4_outputs(7246) <= not a or b;
    layer4_outputs(7247) <= not (a and b);
    layer4_outputs(7248) <= not a or b;
    layer4_outputs(7249) <= not b or a;
    layer4_outputs(7250) <= not (a and b);
    layer4_outputs(7251) <= not b;
    layer4_outputs(7252) <= a and not b;
    layer4_outputs(7253) <= a and b;
    layer4_outputs(7254) <= a;
    layer4_outputs(7255) <= not a or b;
    layer4_outputs(7256) <= a;
    layer4_outputs(7257) <= not (a and b);
    layer4_outputs(7258) <= a;
    layer4_outputs(7259) <= not a;
    layer4_outputs(7260) <= not b;
    layer4_outputs(7261) <= b and not a;
    layer4_outputs(7262) <= not b;
    layer4_outputs(7263) <= a;
    layer4_outputs(7264) <= not (a or b);
    layer4_outputs(7265) <= b;
    layer4_outputs(7266) <= not a;
    layer4_outputs(7267) <= not a or b;
    layer4_outputs(7268) <= not a;
    layer4_outputs(7269) <= not (a or b);
    layer4_outputs(7270) <= '0';
    layer4_outputs(7271) <= a;
    layer4_outputs(7272) <= a or b;
    layer4_outputs(7273) <= b;
    layer4_outputs(7274) <= a xor b;
    layer4_outputs(7275) <= not a;
    layer4_outputs(7276) <= not (a or b);
    layer4_outputs(7277) <= a and b;
    layer4_outputs(7278) <= not b;
    layer4_outputs(7279) <= b;
    layer4_outputs(7280) <= a and not b;
    layer4_outputs(7281) <= a and not b;
    layer4_outputs(7282) <= not a;
    layer4_outputs(7283) <= '0';
    layer4_outputs(7284) <= a xor b;
    layer4_outputs(7285) <= not a or b;
    layer4_outputs(7286) <= a;
    layer4_outputs(7287) <= not a or b;
    layer4_outputs(7288) <= not a;
    layer4_outputs(7289) <= a and not b;
    layer4_outputs(7290) <= '1';
    layer4_outputs(7291) <= not a;
    layer4_outputs(7292) <= not a or b;
    layer4_outputs(7293) <= a;
    layer4_outputs(7294) <= a and b;
    layer4_outputs(7295) <= a;
    layer4_outputs(7296) <= not (a and b);
    layer4_outputs(7297) <= a and not b;
    layer4_outputs(7298) <= not b;
    layer4_outputs(7299) <= a;
    layer4_outputs(7300) <= a xor b;
    layer4_outputs(7301) <= b;
    layer4_outputs(7302) <= not b or a;
    layer4_outputs(7303) <= a and not b;
    layer4_outputs(7304) <= a and not b;
    layer4_outputs(7305) <= not a;
    layer4_outputs(7306) <= not (a or b);
    layer4_outputs(7307) <= b;
    layer4_outputs(7308) <= not a or b;
    layer4_outputs(7309) <= not a;
    layer4_outputs(7310) <= not b;
    layer4_outputs(7311) <= '0';
    layer4_outputs(7312) <= not a or b;
    layer4_outputs(7313) <= not (a or b);
    layer4_outputs(7314) <= not (a or b);
    layer4_outputs(7315) <= not b or a;
    layer4_outputs(7316) <= a xor b;
    layer4_outputs(7317) <= not (a and b);
    layer4_outputs(7318) <= a and not b;
    layer4_outputs(7319) <= not a or b;
    layer4_outputs(7320) <= not (a xor b);
    layer4_outputs(7321) <= b;
    layer4_outputs(7322) <= not b;
    layer4_outputs(7323) <= not (a xor b);
    layer4_outputs(7324) <= not a or b;
    layer4_outputs(7325) <= not (a or b);
    layer4_outputs(7326) <= a and b;
    layer4_outputs(7327) <= a or b;
    layer4_outputs(7328) <= b and not a;
    layer4_outputs(7329) <= not (a or b);
    layer4_outputs(7330) <= b;
    layer4_outputs(7331) <= not a or b;
    layer4_outputs(7332) <= b and not a;
    layer4_outputs(7333) <= not b;
    layer4_outputs(7334) <= a and not b;
    layer4_outputs(7335) <= b and not a;
    layer4_outputs(7336) <= not b;
    layer4_outputs(7337) <= not (a and b);
    layer4_outputs(7338) <= not b;
    layer4_outputs(7339) <= b and not a;
    layer4_outputs(7340) <= not b or a;
    layer4_outputs(7341) <= not b or a;
    layer4_outputs(7342) <= a and not b;
    layer4_outputs(7343) <= a or b;
    layer4_outputs(7344) <= not (a xor b);
    layer4_outputs(7345) <= a;
    layer4_outputs(7346) <= not b or a;
    layer4_outputs(7347) <= not a or b;
    layer4_outputs(7348) <= b;
    layer4_outputs(7349) <= not a;
    layer4_outputs(7350) <= not b;
    layer4_outputs(7351) <= not (a xor b);
    layer4_outputs(7352) <= not (a and b);
    layer4_outputs(7353) <= not b;
    layer4_outputs(7354) <= '0';
    layer4_outputs(7355) <= not b;
    layer4_outputs(7356) <= not b;
    layer4_outputs(7357) <= a and b;
    layer4_outputs(7358) <= not b or a;
    layer4_outputs(7359) <= not b;
    layer4_outputs(7360) <= b;
    layer4_outputs(7361) <= a xor b;
    layer4_outputs(7362) <= b;
    layer4_outputs(7363) <= not a;
    layer4_outputs(7364) <= not a or b;
    layer4_outputs(7365) <= b;
    layer4_outputs(7366) <= not a or b;
    layer4_outputs(7367) <= not (a xor b);
    layer4_outputs(7368) <= not a or b;
    layer4_outputs(7369) <= not a or b;
    layer4_outputs(7370) <= a and b;
    layer4_outputs(7371) <= b;
    layer4_outputs(7372) <= b;
    layer4_outputs(7373) <= not b;
    layer4_outputs(7374) <= a;
    layer4_outputs(7375) <= not (a xor b);
    layer4_outputs(7376) <= not a;
    layer4_outputs(7377) <= not (a and b);
    layer4_outputs(7378) <= not a or b;
    layer4_outputs(7379) <= a and not b;
    layer4_outputs(7380) <= not a or b;
    layer4_outputs(7381) <= not (a xor b);
    layer4_outputs(7382) <= a xor b;
    layer4_outputs(7383) <= not b;
    layer4_outputs(7384) <= not (a or b);
    layer4_outputs(7385) <= '1';
    layer4_outputs(7386) <= '0';
    layer4_outputs(7387) <= b and not a;
    layer4_outputs(7388) <= not (a xor b);
    layer4_outputs(7389) <= a or b;
    layer4_outputs(7390) <= not a or b;
    layer4_outputs(7391) <= not b;
    layer4_outputs(7392) <= b and not a;
    layer4_outputs(7393) <= b;
    layer4_outputs(7394) <= not (a or b);
    layer4_outputs(7395) <= not b;
    layer4_outputs(7396) <= not a;
    layer4_outputs(7397) <= not b or a;
    layer4_outputs(7398) <= a;
    layer4_outputs(7399) <= not (a or b);
    layer4_outputs(7400) <= not b or a;
    layer4_outputs(7401) <= a and b;
    layer4_outputs(7402) <= not (a and b);
    layer4_outputs(7403) <= not a or b;
    layer4_outputs(7404) <= a or b;
    layer4_outputs(7405) <= b;
    layer4_outputs(7406) <= a and b;
    layer4_outputs(7407) <= not (a xor b);
    layer4_outputs(7408) <= not b;
    layer4_outputs(7409) <= not (a and b);
    layer4_outputs(7410) <= not a or b;
    layer4_outputs(7411) <= b and not a;
    layer4_outputs(7412) <= b;
    layer4_outputs(7413) <= not (a or b);
    layer4_outputs(7414) <= not a;
    layer4_outputs(7415) <= not (a xor b);
    layer4_outputs(7416) <= not (a and b);
    layer4_outputs(7417) <= a;
    layer4_outputs(7418) <= not (a or b);
    layer4_outputs(7419) <= a;
    layer4_outputs(7420) <= '0';
    layer4_outputs(7421) <= a xor b;
    layer4_outputs(7422) <= not a or b;
    layer4_outputs(7423) <= a or b;
    layer4_outputs(7424) <= not a;
    layer4_outputs(7425) <= a or b;
    layer4_outputs(7426) <= not (a or b);
    layer4_outputs(7427) <= a or b;
    layer4_outputs(7428) <= b and not a;
    layer4_outputs(7429) <= b and not a;
    layer4_outputs(7430) <= not b;
    layer4_outputs(7431) <= a and not b;
    layer4_outputs(7432) <= not b;
    layer4_outputs(7433) <= not b or a;
    layer4_outputs(7434) <= a;
    layer4_outputs(7435) <= not a or b;
    layer4_outputs(7436) <= a;
    layer4_outputs(7437) <= not a;
    layer4_outputs(7438) <= not b;
    layer4_outputs(7439) <= not a or b;
    layer4_outputs(7440) <= not (a and b);
    layer4_outputs(7441) <= a or b;
    layer4_outputs(7442) <= not (a xor b);
    layer4_outputs(7443) <= not a;
    layer4_outputs(7444) <= not b;
    layer4_outputs(7445) <= not a or b;
    layer4_outputs(7446) <= not a;
    layer4_outputs(7447) <= not (a and b);
    layer4_outputs(7448) <= not a;
    layer4_outputs(7449) <= a and b;
    layer4_outputs(7450) <= a;
    layer4_outputs(7451) <= not a;
    layer4_outputs(7452) <= not (a xor b);
    layer4_outputs(7453) <= not (a or b);
    layer4_outputs(7454) <= not (a xor b);
    layer4_outputs(7455) <= b and not a;
    layer4_outputs(7456) <= a or b;
    layer4_outputs(7457) <= a and b;
    layer4_outputs(7458) <= a;
    layer4_outputs(7459) <= not (a and b);
    layer4_outputs(7460) <= not b or a;
    layer4_outputs(7461) <= not a;
    layer4_outputs(7462) <= not (a or b);
    layer4_outputs(7463) <= a and not b;
    layer4_outputs(7464) <= not a;
    layer4_outputs(7465) <= not a;
    layer4_outputs(7466) <= not b;
    layer4_outputs(7467) <= not b;
    layer4_outputs(7468) <= not (a xor b);
    layer4_outputs(7469) <= a and not b;
    layer4_outputs(7470) <= b and not a;
    layer4_outputs(7471) <= a xor b;
    layer4_outputs(7472) <= a and not b;
    layer4_outputs(7473) <= not b or a;
    layer4_outputs(7474) <= a;
    layer4_outputs(7475) <= b;
    layer4_outputs(7476) <= b;
    layer4_outputs(7477) <= not a or b;
    layer4_outputs(7478) <= not a;
    layer4_outputs(7479) <= a;
    layer4_outputs(7480) <= a xor b;
    layer4_outputs(7481) <= not b or a;
    layer4_outputs(7482) <= b;
    layer4_outputs(7483) <= not b or a;
    layer4_outputs(7484) <= a;
    layer4_outputs(7485) <= b;
    layer4_outputs(7486) <= a and not b;
    layer4_outputs(7487) <= not a;
    layer4_outputs(7488) <= b and not a;
    layer4_outputs(7489) <= a and not b;
    layer4_outputs(7490) <= not (a and b);
    layer4_outputs(7491) <= a or b;
    layer4_outputs(7492) <= a xor b;
    layer4_outputs(7493) <= not (a or b);
    layer4_outputs(7494) <= not (a and b);
    layer4_outputs(7495) <= not a;
    layer4_outputs(7496) <= not a;
    layer4_outputs(7497) <= a;
    layer4_outputs(7498) <= a and b;
    layer4_outputs(7499) <= not b;
    layer4_outputs(7500) <= a or b;
    layer4_outputs(7501) <= a;
    layer4_outputs(7502) <= not (a and b);
    layer4_outputs(7503) <= b and not a;
    layer4_outputs(7504) <= b;
    layer4_outputs(7505) <= not (a or b);
    layer4_outputs(7506) <= not a or b;
    layer4_outputs(7507) <= a and b;
    layer4_outputs(7508) <= not a;
    layer4_outputs(7509) <= b;
    layer4_outputs(7510) <= not a;
    layer4_outputs(7511) <= not (a or b);
    layer4_outputs(7512) <= not (a and b);
    layer4_outputs(7513) <= a xor b;
    layer4_outputs(7514) <= b and not a;
    layer4_outputs(7515) <= not a or b;
    layer4_outputs(7516) <= not (a and b);
    layer4_outputs(7517) <= not (a or b);
    layer4_outputs(7518) <= not a;
    layer4_outputs(7519) <= a xor b;
    layer4_outputs(7520) <= not b;
    layer4_outputs(7521) <= not (a or b);
    layer4_outputs(7522) <= not a;
    layer4_outputs(7523) <= b and not a;
    layer4_outputs(7524) <= a;
    layer4_outputs(7525) <= not (a or b);
    layer4_outputs(7526) <= a;
    layer4_outputs(7527) <= not a;
    layer4_outputs(7528) <= not b or a;
    layer4_outputs(7529) <= not (a and b);
    layer4_outputs(7530) <= not b;
    layer4_outputs(7531) <= a;
    layer4_outputs(7532) <= a and b;
    layer4_outputs(7533) <= b and not a;
    layer4_outputs(7534) <= a or b;
    layer4_outputs(7535) <= a or b;
    layer4_outputs(7536) <= a;
    layer4_outputs(7537) <= not a or b;
    layer4_outputs(7538) <= not b;
    layer4_outputs(7539) <= a;
    layer4_outputs(7540) <= not a;
    layer4_outputs(7541) <= not b;
    layer4_outputs(7542) <= a xor b;
    layer4_outputs(7543) <= '0';
    layer4_outputs(7544) <= a and not b;
    layer4_outputs(7545) <= '1';
    layer4_outputs(7546) <= not a;
    layer4_outputs(7547) <= b;
    layer4_outputs(7548) <= a;
    layer4_outputs(7549) <= b;
    layer4_outputs(7550) <= not b;
    layer4_outputs(7551) <= a and b;
    layer4_outputs(7552) <= '1';
    layer4_outputs(7553) <= b;
    layer4_outputs(7554) <= a;
    layer4_outputs(7555) <= not (a and b);
    layer4_outputs(7556) <= a or b;
    layer4_outputs(7557) <= b and not a;
    layer4_outputs(7558) <= not b;
    layer4_outputs(7559) <= '0';
    layer4_outputs(7560) <= not (a or b);
    layer4_outputs(7561) <= not (a and b);
    layer4_outputs(7562) <= not a;
    layer4_outputs(7563) <= a or b;
    layer4_outputs(7564) <= not b or a;
    layer4_outputs(7565) <= '1';
    layer4_outputs(7566) <= '1';
    layer4_outputs(7567) <= not a;
    layer4_outputs(7568) <= b and not a;
    layer4_outputs(7569) <= '1';
    layer4_outputs(7570) <= a and not b;
    layer4_outputs(7571) <= not a or b;
    layer4_outputs(7572) <= a or b;
    layer4_outputs(7573) <= not (a and b);
    layer4_outputs(7574) <= not a;
    layer4_outputs(7575) <= b and not a;
    layer4_outputs(7576) <= b and not a;
    layer4_outputs(7577) <= not (a or b);
    layer4_outputs(7578) <= not (a and b);
    layer4_outputs(7579) <= a and b;
    layer4_outputs(7580) <= a and b;
    layer4_outputs(7581) <= a or b;
    layer4_outputs(7582) <= not b;
    layer4_outputs(7583) <= a xor b;
    layer4_outputs(7584) <= a and b;
    layer4_outputs(7585) <= not (a or b);
    layer4_outputs(7586) <= '1';
    layer4_outputs(7587) <= a xor b;
    layer4_outputs(7588) <= not (a and b);
    layer4_outputs(7589) <= b;
    layer4_outputs(7590) <= not b;
    layer4_outputs(7591) <= a;
    layer4_outputs(7592) <= b and not a;
    layer4_outputs(7593) <= a or b;
    layer4_outputs(7594) <= b;
    layer4_outputs(7595) <= a;
    layer4_outputs(7596) <= a and b;
    layer4_outputs(7597) <= not b;
    layer4_outputs(7598) <= b;
    layer4_outputs(7599) <= '1';
    layer4_outputs(7600) <= a;
    layer4_outputs(7601) <= not (a xor b);
    layer4_outputs(7602) <= a or b;
    layer4_outputs(7603) <= a and b;
    layer4_outputs(7604) <= '1';
    layer4_outputs(7605) <= '1';
    layer4_outputs(7606) <= a xor b;
    layer4_outputs(7607) <= not a or b;
    layer4_outputs(7608) <= not a or b;
    layer4_outputs(7609) <= not (a and b);
    layer4_outputs(7610) <= '0';
    layer4_outputs(7611) <= a xor b;
    layer4_outputs(7612) <= a and not b;
    layer4_outputs(7613) <= a or b;
    layer4_outputs(7614) <= not (a or b);
    layer4_outputs(7615) <= a xor b;
    layer4_outputs(7616) <= b;
    layer4_outputs(7617) <= a and not b;
    layer4_outputs(7618) <= a and not b;
    layer4_outputs(7619) <= not b or a;
    layer4_outputs(7620) <= a xor b;
    layer4_outputs(7621) <= a or b;
    layer4_outputs(7622) <= not a or b;
    layer4_outputs(7623) <= b and not a;
    layer4_outputs(7624) <= not a;
    layer4_outputs(7625) <= not b;
    layer4_outputs(7626) <= not b or a;
    layer4_outputs(7627) <= '0';
    layer4_outputs(7628) <= a xor b;
    layer4_outputs(7629) <= not b;
    layer4_outputs(7630) <= b;
    layer4_outputs(7631) <= not b;
    layer4_outputs(7632) <= b;
    layer4_outputs(7633) <= a and not b;
    layer4_outputs(7634) <= not b or a;
    layer4_outputs(7635) <= not a;
    layer4_outputs(7636) <= not b;
    layer4_outputs(7637) <= a and not b;
    layer4_outputs(7638) <= a or b;
    layer4_outputs(7639) <= b and not a;
    layer4_outputs(7640) <= a;
    layer4_outputs(7641) <= not b or a;
    layer4_outputs(7642) <= a and b;
    layer4_outputs(7643) <= not a;
    layer4_outputs(7644) <= not a;
    layer4_outputs(7645) <= not a;
    layer4_outputs(7646) <= a;
    layer4_outputs(7647) <= not b or a;
    layer4_outputs(7648) <= not b;
    layer4_outputs(7649) <= not a;
    layer4_outputs(7650) <= b and not a;
    layer4_outputs(7651) <= not (a or b);
    layer4_outputs(7652) <= a and not b;
    layer4_outputs(7653) <= b;
    layer4_outputs(7654) <= b and not a;
    layer4_outputs(7655) <= not a;
    layer4_outputs(7656) <= b;
    layer4_outputs(7657) <= b;
    layer4_outputs(7658) <= not (a or b);
    layer4_outputs(7659) <= a or b;
    layer4_outputs(7660) <= a xor b;
    layer4_outputs(7661) <= not a or b;
    layer4_outputs(7662) <= b;
    layer4_outputs(7663) <= not a or b;
    layer4_outputs(7664) <= not (a or b);
    layer4_outputs(7665) <= a and b;
    layer4_outputs(7666) <= a or b;
    layer4_outputs(7667) <= a and b;
    layer4_outputs(7668) <= not a;
    layer4_outputs(7669) <= '0';
    layer4_outputs(7670) <= not a or b;
    layer4_outputs(7671) <= b and not a;
    layer4_outputs(7672) <= a;
    layer4_outputs(7673) <= a;
    layer4_outputs(7674) <= a and b;
    layer4_outputs(7675) <= a xor b;
    layer4_outputs(7676) <= a;
    layer4_outputs(7677) <= a and b;
    layer4_outputs(7678) <= not (a or b);
    layer4_outputs(7679) <= not b;
    layer4_outputs(7680) <= not b;
    layer4_outputs(7681) <= b;
    layer4_outputs(7682) <= a and b;
    layer4_outputs(7683) <= a or b;
    layer4_outputs(7684) <= not a or b;
    layer4_outputs(7685) <= not (a or b);
    layer4_outputs(7686) <= not (a and b);
    layer4_outputs(7687) <= b;
    layer4_outputs(7688) <= not a;
    layer4_outputs(7689) <= a;
    layer4_outputs(7690) <= a or b;
    layer4_outputs(7691) <= b;
    layer4_outputs(7692) <= not a;
    layer4_outputs(7693) <= b;
    layer4_outputs(7694) <= not a or b;
    layer4_outputs(7695) <= not a;
    layer4_outputs(7696) <= not b or a;
    layer4_outputs(7697) <= '1';
    layer4_outputs(7698) <= a and b;
    layer4_outputs(7699) <= a and b;
    layer4_outputs(7700) <= a;
    layer4_outputs(7701) <= not (a or b);
    layer4_outputs(7702) <= not b;
    layer4_outputs(7703) <= not b or a;
    layer4_outputs(7704) <= not a;
    layer4_outputs(7705) <= a and not b;
    layer4_outputs(7706) <= not a;
    layer4_outputs(7707) <= a and b;
    layer4_outputs(7708) <= b and not a;
    layer4_outputs(7709) <= a and b;
    layer4_outputs(7710) <= not (a and b);
    layer4_outputs(7711) <= not (a xor b);
    layer4_outputs(7712) <= not (a xor b);
    layer4_outputs(7713) <= b;
    layer4_outputs(7714) <= a;
    layer4_outputs(7715) <= a;
    layer4_outputs(7716) <= not (a and b);
    layer4_outputs(7717) <= '0';
    layer4_outputs(7718) <= not (a and b);
    layer4_outputs(7719) <= a;
    layer4_outputs(7720) <= not a;
    layer4_outputs(7721) <= not a;
    layer4_outputs(7722) <= a;
    layer4_outputs(7723) <= a;
    layer4_outputs(7724) <= b;
    layer4_outputs(7725) <= not (a and b);
    layer4_outputs(7726) <= not a or b;
    layer4_outputs(7727) <= a and b;
    layer4_outputs(7728) <= not b;
    layer4_outputs(7729) <= not (a xor b);
    layer4_outputs(7730) <= not b;
    layer4_outputs(7731) <= a and not b;
    layer4_outputs(7732) <= not a or b;
    layer4_outputs(7733) <= not b or a;
    layer4_outputs(7734) <= not b or a;
    layer4_outputs(7735) <= not b;
    layer4_outputs(7736) <= a or b;
    layer4_outputs(7737) <= a or b;
    layer4_outputs(7738) <= a and b;
    layer4_outputs(7739) <= b and not a;
    layer4_outputs(7740) <= b;
    layer4_outputs(7741) <= not (a xor b);
    layer4_outputs(7742) <= a or b;
    layer4_outputs(7743) <= not a;
    layer4_outputs(7744) <= not a;
    layer4_outputs(7745) <= a xor b;
    layer4_outputs(7746) <= a;
    layer4_outputs(7747) <= not b;
    layer4_outputs(7748) <= not (a or b);
    layer4_outputs(7749) <= b;
    layer4_outputs(7750) <= a xor b;
    layer4_outputs(7751) <= '0';
    layer4_outputs(7752) <= a;
    layer4_outputs(7753) <= not (a or b);
    layer4_outputs(7754) <= b;
    layer4_outputs(7755) <= not b;
    layer4_outputs(7756) <= a or b;
    layer4_outputs(7757) <= not (a xor b);
    layer4_outputs(7758) <= a and b;
    layer4_outputs(7759) <= b and not a;
    layer4_outputs(7760) <= '1';
    layer4_outputs(7761) <= not (a or b);
    layer4_outputs(7762) <= b and not a;
    layer4_outputs(7763) <= not b;
    layer4_outputs(7764) <= a or b;
    layer4_outputs(7765) <= not (a xor b);
    layer4_outputs(7766) <= not (a xor b);
    layer4_outputs(7767) <= a or b;
    layer4_outputs(7768) <= not a or b;
    layer4_outputs(7769) <= not b or a;
    layer4_outputs(7770) <= a;
    layer4_outputs(7771) <= a xor b;
    layer4_outputs(7772) <= not a or b;
    layer4_outputs(7773) <= not (a or b);
    layer4_outputs(7774) <= not a or b;
    layer4_outputs(7775) <= a or b;
    layer4_outputs(7776) <= b and not a;
    layer4_outputs(7777) <= not b;
    layer4_outputs(7778) <= a and not b;
    layer4_outputs(7779) <= not b;
    layer4_outputs(7780) <= a or b;
    layer4_outputs(7781) <= not b or a;
    layer4_outputs(7782) <= not (a and b);
    layer4_outputs(7783) <= b;
    layer4_outputs(7784) <= not (a and b);
    layer4_outputs(7785) <= not a;
    layer4_outputs(7786) <= not b;
    layer4_outputs(7787) <= a or b;
    layer4_outputs(7788) <= a and b;
    layer4_outputs(7789) <= not b;
    layer4_outputs(7790) <= a xor b;
    layer4_outputs(7791) <= not a;
    layer4_outputs(7792) <= not a;
    layer4_outputs(7793) <= b and not a;
    layer4_outputs(7794) <= b and not a;
    layer4_outputs(7795) <= '1';
    layer4_outputs(7796) <= a or b;
    layer4_outputs(7797) <= not b;
    layer4_outputs(7798) <= not (a or b);
    layer4_outputs(7799) <= b;
    layer4_outputs(7800) <= '0';
    layer4_outputs(7801) <= a;
    layer4_outputs(7802) <= b;
    layer4_outputs(7803) <= not (a and b);
    layer4_outputs(7804) <= a;
    layer4_outputs(7805) <= not (a or b);
    layer4_outputs(7806) <= a or b;
    layer4_outputs(7807) <= not (a or b);
    layer4_outputs(7808) <= not a or b;
    layer4_outputs(7809) <= not (a xor b);
    layer4_outputs(7810) <= not (a or b);
    layer4_outputs(7811) <= a and not b;
    layer4_outputs(7812) <= a xor b;
    layer4_outputs(7813) <= not (a or b);
    layer4_outputs(7814) <= a xor b;
    layer4_outputs(7815) <= a and b;
    layer4_outputs(7816) <= b and not a;
    layer4_outputs(7817) <= not b;
    layer4_outputs(7818) <= not a or b;
    layer4_outputs(7819) <= not a;
    layer4_outputs(7820) <= a xor b;
    layer4_outputs(7821) <= a;
    layer4_outputs(7822) <= not a or b;
    layer4_outputs(7823) <= not a;
    layer4_outputs(7824) <= b and not a;
    layer4_outputs(7825) <= a or b;
    layer4_outputs(7826) <= a or b;
    layer4_outputs(7827) <= not b or a;
    layer4_outputs(7828) <= a xor b;
    layer4_outputs(7829) <= not a or b;
    layer4_outputs(7830) <= a and not b;
    layer4_outputs(7831) <= not (a or b);
    layer4_outputs(7832) <= not b;
    layer4_outputs(7833) <= not a;
    layer4_outputs(7834) <= a xor b;
    layer4_outputs(7835) <= b and not a;
    layer4_outputs(7836) <= a or b;
    layer4_outputs(7837) <= b;
    layer4_outputs(7838) <= a and b;
    layer4_outputs(7839) <= not a;
    layer4_outputs(7840) <= not b;
    layer4_outputs(7841) <= not b or a;
    layer4_outputs(7842) <= a or b;
    layer4_outputs(7843) <= not (a xor b);
    layer4_outputs(7844) <= not b;
    layer4_outputs(7845) <= a xor b;
    layer4_outputs(7846) <= '1';
    layer4_outputs(7847) <= a;
    layer4_outputs(7848) <= a and not b;
    layer4_outputs(7849) <= a and b;
    layer4_outputs(7850) <= not b;
    layer4_outputs(7851) <= not (a and b);
    layer4_outputs(7852) <= a and b;
    layer4_outputs(7853) <= not (a xor b);
    layer4_outputs(7854) <= not a;
    layer4_outputs(7855) <= a xor b;
    layer4_outputs(7856) <= b;
    layer4_outputs(7857) <= not (a or b);
    layer4_outputs(7858) <= not a;
    layer4_outputs(7859) <= a;
    layer4_outputs(7860) <= not a or b;
    layer4_outputs(7861) <= a and b;
    layer4_outputs(7862) <= '1';
    layer4_outputs(7863) <= not b;
    layer4_outputs(7864) <= not (a and b);
    layer4_outputs(7865) <= a or b;
    layer4_outputs(7866) <= a;
    layer4_outputs(7867) <= not a;
    layer4_outputs(7868) <= b and not a;
    layer4_outputs(7869) <= b and not a;
    layer4_outputs(7870) <= a xor b;
    layer4_outputs(7871) <= not (a and b);
    layer4_outputs(7872) <= b;
    layer4_outputs(7873) <= a and not b;
    layer4_outputs(7874) <= b and not a;
    layer4_outputs(7875) <= not b;
    layer4_outputs(7876) <= not b;
    layer4_outputs(7877) <= not (a or b);
    layer4_outputs(7878) <= a;
    layer4_outputs(7879) <= b;
    layer4_outputs(7880) <= not (a or b);
    layer4_outputs(7881) <= not (a xor b);
    layer4_outputs(7882) <= not b;
    layer4_outputs(7883) <= not b;
    layer4_outputs(7884) <= not a;
    layer4_outputs(7885) <= not b;
    layer4_outputs(7886) <= not b;
    layer4_outputs(7887) <= not (a and b);
    layer4_outputs(7888) <= not a or b;
    layer4_outputs(7889) <= not b or a;
    layer4_outputs(7890) <= not (a xor b);
    layer4_outputs(7891) <= a or b;
    layer4_outputs(7892) <= not a;
    layer4_outputs(7893) <= '0';
    layer4_outputs(7894) <= not a or b;
    layer4_outputs(7895) <= not b;
    layer4_outputs(7896) <= not (a or b);
    layer4_outputs(7897) <= a or b;
    layer4_outputs(7898) <= a;
    layer4_outputs(7899) <= a;
    layer4_outputs(7900) <= a xor b;
    layer4_outputs(7901) <= not (a or b);
    layer4_outputs(7902) <= a and not b;
    layer4_outputs(7903) <= not b;
    layer4_outputs(7904) <= a or b;
    layer4_outputs(7905) <= not a;
    layer4_outputs(7906) <= a or b;
    layer4_outputs(7907) <= b;
    layer4_outputs(7908) <= b and not a;
    layer4_outputs(7909) <= not (a xor b);
    layer4_outputs(7910) <= not b or a;
    layer4_outputs(7911) <= a or b;
    layer4_outputs(7912) <= a or b;
    layer4_outputs(7913) <= a xor b;
    layer4_outputs(7914) <= '1';
    layer4_outputs(7915) <= not (a and b);
    layer4_outputs(7916) <= not b or a;
    layer4_outputs(7917) <= a or b;
    layer4_outputs(7918) <= not b;
    layer4_outputs(7919) <= a;
    layer4_outputs(7920) <= not b;
    layer4_outputs(7921) <= b;
    layer4_outputs(7922) <= a;
    layer4_outputs(7923) <= a and not b;
    layer4_outputs(7924) <= not (a xor b);
    layer4_outputs(7925) <= '1';
    layer4_outputs(7926) <= b;
    layer4_outputs(7927) <= a xor b;
    layer4_outputs(7928) <= b;
    layer4_outputs(7929) <= a and not b;
    layer4_outputs(7930) <= '0';
    layer4_outputs(7931) <= a;
    layer4_outputs(7932) <= not a;
    layer4_outputs(7933) <= not b or a;
    layer4_outputs(7934) <= a xor b;
    layer4_outputs(7935) <= a;
    layer4_outputs(7936) <= a;
    layer4_outputs(7937) <= a;
    layer4_outputs(7938) <= a and not b;
    layer4_outputs(7939) <= not (a and b);
    layer4_outputs(7940) <= a xor b;
    layer4_outputs(7941) <= a;
    layer4_outputs(7942) <= a and b;
    layer4_outputs(7943) <= a and not b;
    layer4_outputs(7944) <= a xor b;
    layer4_outputs(7945) <= not b;
    layer4_outputs(7946) <= not a;
    layer4_outputs(7947) <= a and b;
    layer4_outputs(7948) <= a and not b;
    layer4_outputs(7949) <= b;
    layer4_outputs(7950) <= a xor b;
    layer4_outputs(7951) <= not (a or b);
    layer4_outputs(7952) <= not a or b;
    layer4_outputs(7953) <= b and not a;
    layer4_outputs(7954) <= a or b;
    layer4_outputs(7955) <= b and not a;
    layer4_outputs(7956) <= a;
    layer4_outputs(7957) <= not a or b;
    layer4_outputs(7958) <= not b or a;
    layer4_outputs(7959) <= a;
    layer4_outputs(7960) <= not a;
    layer4_outputs(7961) <= a or b;
    layer4_outputs(7962) <= a and not b;
    layer4_outputs(7963) <= a and not b;
    layer4_outputs(7964) <= a;
    layer4_outputs(7965) <= not b or a;
    layer4_outputs(7966) <= a and b;
    layer4_outputs(7967) <= not b;
    layer4_outputs(7968) <= a;
    layer4_outputs(7969) <= not (a and b);
    layer4_outputs(7970) <= a;
    layer4_outputs(7971) <= b;
    layer4_outputs(7972) <= a xor b;
    layer4_outputs(7973) <= b;
    layer4_outputs(7974) <= b;
    layer4_outputs(7975) <= not a;
    layer4_outputs(7976) <= not a or b;
    layer4_outputs(7977) <= not b;
    layer4_outputs(7978) <= not a or b;
    layer4_outputs(7979) <= not a or b;
    layer4_outputs(7980) <= b;
    layer4_outputs(7981) <= not (a and b);
    layer4_outputs(7982) <= not (a or b);
    layer4_outputs(7983) <= not (a and b);
    layer4_outputs(7984) <= b and not a;
    layer4_outputs(7985) <= a;
    layer4_outputs(7986) <= b;
    layer4_outputs(7987) <= not b or a;
    layer4_outputs(7988) <= not (a and b);
    layer4_outputs(7989) <= a and b;
    layer4_outputs(7990) <= b;
    layer4_outputs(7991) <= not b or a;
    layer4_outputs(7992) <= a;
    layer4_outputs(7993) <= b;
    layer4_outputs(7994) <= not a;
    layer4_outputs(7995) <= a or b;
    layer4_outputs(7996) <= not b;
    layer4_outputs(7997) <= not (a xor b);
    layer4_outputs(7998) <= a;
    layer4_outputs(7999) <= not b or a;
    layer4_outputs(8000) <= b;
    layer4_outputs(8001) <= not b;
    layer4_outputs(8002) <= not (a xor b);
    layer4_outputs(8003) <= not (a or b);
    layer4_outputs(8004) <= a xor b;
    layer4_outputs(8005) <= not a;
    layer4_outputs(8006) <= a and not b;
    layer4_outputs(8007) <= b;
    layer4_outputs(8008) <= a xor b;
    layer4_outputs(8009) <= a or b;
    layer4_outputs(8010) <= b;
    layer4_outputs(8011) <= a and b;
    layer4_outputs(8012) <= not a;
    layer4_outputs(8013) <= b;
    layer4_outputs(8014) <= not b or a;
    layer4_outputs(8015) <= a xor b;
    layer4_outputs(8016) <= a and b;
    layer4_outputs(8017) <= b and not a;
    layer4_outputs(8018) <= a and b;
    layer4_outputs(8019) <= not b or a;
    layer4_outputs(8020) <= b and not a;
    layer4_outputs(8021) <= '0';
    layer4_outputs(8022) <= a and b;
    layer4_outputs(8023) <= not a;
    layer4_outputs(8024) <= b;
    layer4_outputs(8025) <= a xor b;
    layer4_outputs(8026) <= not (a or b);
    layer4_outputs(8027) <= a;
    layer4_outputs(8028) <= not b or a;
    layer4_outputs(8029) <= b;
    layer4_outputs(8030) <= a or b;
    layer4_outputs(8031) <= not (a or b);
    layer4_outputs(8032) <= not b;
    layer4_outputs(8033) <= not b;
    layer4_outputs(8034) <= not (a and b);
    layer4_outputs(8035) <= not a or b;
    layer4_outputs(8036) <= not a;
    layer4_outputs(8037) <= a and not b;
    layer4_outputs(8038) <= a xor b;
    layer4_outputs(8039) <= b;
    layer4_outputs(8040) <= not b or a;
    layer4_outputs(8041) <= a and b;
    layer4_outputs(8042) <= not a or b;
    layer4_outputs(8043) <= not a;
    layer4_outputs(8044) <= b and not a;
    layer4_outputs(8045) <= not a or b;
    layer4_outputs(8046) <= a or b;
    layer4_outputs(8047) <= b and not a;
    layer4_outputs(8048) <= a;
    layer4_outputs(8049) <= not (a or b);
    layer4_outputs(8050) <= not (a xor b);
    layer4_outputs(8051) <= a;
    layer4_outputs(8052) <= a xor b;
    layer4_outputs(8053) <= b and not a;
    layer4_outputs(8054) <= not b;
    layer4_outputs(8055) <= not a;
    layer4_outputs(8056) <= a or b;
    layer4_outputs(8057) <= not a;
    layer4_outputs(8058) <= a;
    layer4_outputs(8059) <= a;
    layer4_outputs(8060) <= not b or a;
    layer4_outputs(8061) <= b;
    layer4_outputs(8062) <= a xor b;
    layer4_outputs(8063) <= not a;
    layer4_outputs(8064) <= a and b;
    layer4_outputs(8065) <= not a;
    layer4_outputs(8066) <= a or b;
    layer4_outputs(8067) <= a xor b;
    layer4_outputs(8068) <= b;
    layer4_outputs(8069) <= b and not a;
    layer4_outputs(8070) <= b;
    layer4_outputs(8071) <= b;
    layer4_outputs(8072) <= a;
    layer4_outputs(8073) <= not a;
    layer4_outputs(8074) <= b;
    layer4_outputs(8075) <= a or b;
    layer4_outputs(8076) <= not a or b;
    layer4_outputs(8077) <= a or b;
    layer4_outputs(8078) <= a or b;
    layer4_outputs(8079) <= a and b;
    layer4_outputs(8080) <= b;
    layer4_outputs(8081) <= a xor b;
    layer4_outputs(8082) <= not (a xor b);
    layer4_outputs(8083) <= b;
    layer4_outputs(8084) <= a;
    layer4_outputs(8085) <= a or b;
    layer4_outputs(8086) <= not b;
    layer4_outputs(8087) <= a xor b;
    layer4_outputs(8088) <= not a;
    layer4_outputs(8089) <= a;
    layer4_outputs(8090) <= b;
    layer4_outputs(8091) <= not (a xor b);
    layer4_outputs(8092) <= not (a xor b);
    layer4_outputs(8093) <= a and b;
    layer4_outputs(8094) <= a or b;
    layer4_outputs(8095) <= b;
    layer4_outputs(8096) <= b;
    layer4_outputs(8097) <= b;
    layer4_outputs(8098) <= not b;
    layer4_outputs(8099) <= not a or b;
    layer4_outputs(8100) <= a;
    layer4_outputs(8101) <= not (a and b);
    layer4_outputs(8102) <= b;
    layer4_outputs(8103) <= a or b;
    layer4_outputs(8104) <= a and not b;
    layer4_outputs(8105) <= not (a xor b);
    layer4_outputs(8106) <= b and not a;
    layer4_outputs(8107) <= not b or a;
    layer4_outputs(8108) <= a xor b;
    layer4_outputs(8109) <= not b;
    layer4_outputs(8110) <= a xor b;
    layer4_outputs(8111) <= not (a and b);
    layer4_outputs(8112) <= '1';
    layer4_outputs(8113) <= b;
    layer4_outputs(8114) <= b;
    layer4_outputs(8115) <= not b;
    layer4_outputs(8116) <= not a or b;
    layer4_outputs(8117) <= not a;
    layer4_outputs(8118) <= not a;
    layer4_outputs(8119) <= not (a or b);
    layer4_outputs(8120) <= a;
    layer4_outputs(8121) <= not a;
    layer4_outputs(8122) <= not a;
    layer4_outputs(8123) <= not (a and b);
    layer4_outputs(8124) <= not a or b;
    layer4_outputs(8125) <= b;
    layer4_outputs(8126) <= not a or b;
    layer4_outputs(8127) <= '0';
    layer4_outputs(8128) <= not (a and b);
    layer4_outputs(8129) <= not (a xor b);
    layer4_outputs(8130) <= b;
    layer4_outputs(8131) <= b and not a;
    layer4_outputs(8132) <= not (a xor b);
    layer4_outputs(8133) <= not (a or b);
    layer4_outputs(8134) <= not b;
    layer4_outputs(8135) <= a or b;
    layer4_outputs(8136) <= not a;
    layer4_outputs(8137) <= a and not b;
    layer4_outputs(8138) <= a and b;
    layer4_outputs(8139) <= not b;
    layer4_outputs(8140) <= a and not b;
    layer4_outputs(8141) <= a and not b;
    layer4_outputs(8142) <= '0';
    layer4_outputs(8143) <= a or b;
    layer4_outputs(8144) <= not (a or b);
    layer4_outputs(8145) <= not (a xor b);
    layer4_outputs(8146) <= not a or b;
    layer4_outputs(8147) <= a and b;
    layer4_outputs(8148) <= not b;
    layer4_outputs(8149) <= a xor b;
    layer4_outputs(8150) <= a xor b;
    layer4_outputs(8151) <= a and not b;
    layer4_outputs(8152) <= not b or a;
    layer4_outputs(8153) <= b;
    layer4_outputs(8154) <= not b or a;
    layer4_outputs(8155) <= a and not b;
    layer4_outputs(8156) <= a and b;
    layer4_outputs(8157) <= not b or a;
    layer4_outputs(8158) <= not (a and b);
    layer4_outputs(8159) <= not (a xor b);
    layer4_outputs(8160) <= b;
    layer4_outputs(8161) <= not (a and b);
    layer4_outputs(8162) <= not a or b;
    layer4_outputs(8163) <= not a;
    layer4_outputs(8164) <= not b;
    layer4_outputs(8165) <= not a;
    layer4_outputs(8166) <= not a;
    layer4_outputs(8167) <= a and b;
    layer4_outputs(8168) <= a xor b;
    layer4_outputs(8169) <= a or b;
    layer4_outputs(8170) <= b and not a;
    layer4_outputs(8171) <= a;
    layer4_outputs(8172) <= not b;
    layer4_outputs(8173) <= a and b;
    layer4_outputs(8174) <= not a;
    layer4_outputs(8175) <= not a;
    layer4_outputs(8176) <= a and not b;
    layer4_outputs(8177) <= b and not a;
    layer4_outputs(8178) <= not (a and b);
    layer4_outputs(8179) <= not a;
    layer4_outputs(8180) <= a and not b;
    layer4_outputs(8181) <= not a;
    layer4_outputs(8182) <= a and b;
    layer4_outputs(8183) <= not (a xor b);
    layer4_outputs(8184) <= b;
    layer4_outputs(8185) <= not a or b;
    layer4_outputs(8186) <= a and not b;
    layer4_outputs(8187) <= b and not a;
    layer4_outputs(8188) <= '0';
    layer4_outputs(8189) <= b;
    layer4_outputs(8190) <= not b;
    layer4_outputs(8191) <= '0';
    layer4_outputs(8192) <= '1';
    layer4_outputs(8193) <= not a;
    layer4_outputs(8194) <= a or b;
    layer4_outputs(8195) <= a xor b;
    layer4_outputs(8196) <= a or b;
    layer4_outputs(8197) <= not a;
    layer4_outputs(8198) <= not a;
    layer4_outputs(8199) <= not (a or b);
    layer4_outputs(8200) <= a;
    layer4_outputs(8201) <= a;
    layer4_outputs(8202) <= a or b;
    layer4_outputs(8203) <= not a or b;
    layer4_outputs(8204) <= not (a and b);
    layer4_outputs(8205) <= not a;
    layer4_outputs(8206) <= not a;
    layer4_outputs(8207) <= a or b;
    layer4_outputs(8208) <= not (a or b);
    layer4_outputs(8209) <= '1';
    layer4_outputs(8210) <= not (a and b);
    layer4_outputs(8211) <= a;
    layer4_outputs(8212) <= not a;
    layer4_outputs(8213) <= b;
    layer4_outputs(8214) <= a;
    layer4_outputs(8215) <= not a or b;
    layer4_outputs(8216) <= not (a and b);
    layer4_outputs(8217) <= b;
    layer4_outputs(8218) <= not (a xor b);
    layer4_outputs(8219) <= a and b;
    layer4_outputs(8220) <= not (a and b);
    layer4_outputs(8221) <= not a;
    layer4_outputs(8222) <= not (a and b);
    layer4_outputs(8223) <= a xor b;
    layer4_outputs(8224) <= not b;
    layer4_outputs(8225) <= '1';
    layer4_outputs(8226) <= not (a xor b);
    layer4_outputs(8227) <= a or b;
    layer4_outputs(8228) <= not (a xor b);
    layer4_outputs(8229) <= not (a and b);
    layer4_outputs(8230) <= b;
    layer4_outputs(8231) <= not (a or b);
    layer4_outputs(8232) <= not b or a;
    layer4_outputs(8233) <= not b;
    layer4_outputs(8234) <= '0';
    layer4_outputs(8235) <= a or b;
    layer4_outputs(8236) <= not b;
    layer4_outputs(8237) <= a;
    layer4_outputs(8238) <= not b;
    layer4_outputs(8239) <= b and not a;
    layer4_outputs(8240) <= not b or a;
    layer4_outputs(8241) <= not (a xor b);
    layer4_outputs(8242) <= not (a and b);
    layer4_outputs(8243) <= b and not a;
    layer4_outputs(8244) <= '0';
    layer4_outputs(8245) <= b;
    layer4_outputs(8246) <= not (a or b);
    layer4_outputs(8247) <= b;
    layer4_outputs(8248) <= b and not a;
    layer4_outputs(8249) <= not (a or b);
    layer4_outputs(8250) <= '1';
    layer4_outputs(8251) <= not (a and b);
    layer4_outputs(8252) <= a;
    layer4_outputs(8253) <= a and b;
    layer4_outputs(8254) <= a or b;
    layer4_outputs(8255) <= not (a or b);
    layer4_outputs(8256) <= not (a and b);
    layer4_outputs(8257) <= not b;
    layer4_outputs(8258) <= b and not a;
    layer4_outputs(8259) <= not a or b;
    layer4_outputs(8260) <= b and not a;
    layer4_outputs(8261) <= a;
    layer4_outputs(8262) <= not a;
    layer4_outputs(8263) <= a or b;
    layer4_outputs(8264) <= not (a or b);
    layer4_outputs(8265) <= not b;
    layer4_outputs(8266) <= a and not b;
    layer4_outputs(8267) <= a;
    layer4_outputs(8268) <= not a;
    layer4_outputs(8269) <= not a;
    layer4_outputs(8270) <= a xor b;
    layer4_outputs(8271) <= not (a xor b);
    layer4_outputs(8272) <= not (a or b);
    layer4_outputs(8273) <= a and b;
    layer4_outputs(8274) <= not (a and b);
    layer4_outputs(8275) <= not (a or b);
    layer4_outputs(8276) <= not (a or b);
    layer4_outputs(8277) <= not b or a;
    layer4_outputs(8278) <= not (a xor b);
    layer4_outputs(8279) <= not a or b;
    layer4_outputs(8280) <= not a;
    layer4_outputs(8281) <= a and b;
    layer4_outputs(8282) <= not b;
    layer4_outputs(8283) <= b;
    layer4_outputs(8284) <= not (a xor b);
    layer4_outputs(8285) <= not b or a;
    layer4_outputs(8286) <= a and b;
    layer4_outputs(8287) <= b;
    layer4_outputs(8288) <= not (a xor b);
    layer4_outputs(8289) <= not b;
    layer4_outputs(8290) <= a or b;
    layer4_outputs(8291) <= not b or a;
    layer4_outputs(8292) <= not a or b;
    layer4_outputs(8293) <= a;
    layer4_outputs(8294) <= not a or b;
    layer4_outputs(8295) <= not a;
    layer4_outputs(8296) <= a and not b;
    layer4_outputs(8297) <= not (a and b);
    layer4_outputs(8298) <= a or b;
    layer4_outputs(8299) <= a or b;
    layer4_outputs(8300) <= not a;
    layer4_outputs(8301) <= a;
    layer4_outputs(8302) <= a and not b;
    layer4_outputs(8303) <= not (a or b);
    layer4_outputs(8304) <= a and not b;
    layer4_outputs(8305) <= not (a and b);
    layer4_outputs(8306) <= a and not b;
    layer4_outputs(8307) <= b;
    layer4_outputs(8308) <= a xor b;
    layer4_outputs(8309) <= not a;
    layer4_outputs(8310) <= not a;
    layer4_outputs(8311) <= a;
    layer4_outputs(8312) <= not (a and b);
    layer4_outputs(8313) <= not (a or b);
    layer4_outputs(8314) <= a and not b;
    layer4_outputs(8315) <= not (a or b);
    layer4_outputs(8316) <= a or b;
    layer4_outputs(8317) <= not b or a;
    layer4_outputs(8318) <= not b;
    layer4_outputs(8319) <= not b or a;
    layer4_outputs(8320) <= a;
    layer4_outputs(8321) <= not a;
    layer4_outputs(8322) <= not a or b;
    layer4_outputs(8323) <= not a;
    layer4_outputs(8324) <= not b;
    layer4_outputs(8325) <= not (a or b);
    layer4_outputs(8326) <= a and not b;
    layer4_outputs(8327) <= not (a or b);
    layer4_outputs(8328) <= not b;
    layer4_outputs(8329) <= '0';
    layer4_outputs(8330) <= '0';
    layer4_outputs(8331) <= not a;
    layer4_outputs(8332) <= a and b;
    layer4_outputs(8333) <= b;
    layer4_outputs(8334) <= '1';
    layer4_outputs(8335) <= a xor b;
    layer4_outputs(8336) <= a;
    layer4_outputs(8337) <= not b or a;
    layer4_outputs(8338) <= a;
    layer4_outputs(8339) <= not b;
    layer4_outputs(8340) <= a;
    layer4_outputs(8341) <= not (a or b);
    layer4_outputs(8342) <= not a or b;
    layer4_outputs(8343) <= not a or b;
    layer4_outputs(8344) <= not b;
    layer4_outputs(8345) <= not (a or b);
    layer4_outputs(8346) <= not b;
    layer4_outputs(8347) <= a;
    layer4_outputs(8348) <= b and not a;
    layer4_outputs(8349) <= a xor b;
    layer4_outputs(8350) <= a and b;
    layer4_outputs(8351) <= b;
    layer4_outputs(8352) <= b;
    layer4_outputs(8353) <= not (a and b);
    layer4_outputs(8354) <= not (a and b);
    layer4_outputs(8355) <= a or b;
    layer4_outputs(8356) <= not b or a;
    layer4_outputs(8357) <= a xor b;
    layer4_outputs(8358) <= a xor b;
    layer4_outputs(8359) <= a and not b;
    layer4_outputs(8360) <= not (a and b);
    layer4_outputs(8361) <= not b;
    layer4_outputs(8362) <= a and not b;
    layer4_outputs(8363) <= not b;
    layer4_outputs(8364) <= not b;
    layer4_outputs(8365) <= b;
    layer4_outputs(8366) <= a and b;
    layer4_outputs(8367) <= a xor b;
    layer4_outputs(8368) <= not b;
    layer4_outputs(8369) <= a and b;
    layer4_outputs(8370) <= '1';
    layer4_outputs(8371) <= a or b;
    layer4_outputs(8372) <= b;
    layer4_outputs(8373) <= not b;
    layer4_outputs(8374) <= a;
    layer4_outputs(8375) <= a or b;
    layer4_outputs(8376) <= not a;
    layer4_outputs(8377) <= not (a or b);
    layer4_outputs(8378) <= not a;
    layer4_outputs(8379) <= not (a or b);
    layer4_outputs(8380) <= not a;
    layer4_outputs(8381) <= not a or b;
    layer4_outputs(8382) <= a;
    layer4_outputs(8383) <= '1';
    layer4_outputs(8384) <= a;
    layer4_outputs(8385) <= not (a and b);
    layer4_outputs(8386) <= a or b;
    layer4_outputs(8387) <= not (a and b);
    layer4_outputs(8388) <= a or b;
    layer4_outputs(8389) <= not a or b;
    layer4_outputs(8390) <= a and not b;
    layer4_outputs(8391) <= a;
    layer4_outputs(8392) <= a or b;
    layer4_outputs(8393) <= not b;
    layer4_outputs(8394) <= not b;
    layer4_outputs(8395) <= a xor b;
    layer4_outputs(8396) <= not (a or b);
    layer4_outputs(8397) <= a and b;
    layer4_outputs(8398) <= '0';
    layer4_outputs(8399) <= b;
    layer4_outputs(8400) <= a xor b;
    layer4_outputs(8401) <= a;
    layer4_outputs(8402) <= not a;
    layer4_outputs(8403) <= b;
    layer4_outputs(8404) <= a and b;
    layer4_outputs(8405) <= a xor b;
    layer4_outputs(8406) <= a;
    layer4_outputs(8407) <= not a;
    layer4_outputs(8408) <= not (a or b);
    layer4_outputs(8409) <= a;
    layer4_outputs(8410) <= not b;
    layer4_outputs(8411) <= not a;
    layer4_outputs(8412) <= a and b;
    layer4_outputs(8413) <= not a or b;
    layer4_outputs(8414) <= not (a and b);
    layer4_outputs(8415) <= not (a and b);
    layer4_outputs(8416) <= a;
    layer4_outputs(8417) <= not b;
    layer4_outputs(8418) <= not (a or b);
    layer4_outputs(8419) <= not b;
    layer4_outputs(8420) <= not (a xor b);
    layer4_outputs(8421) <= a and b;
    layer4_outputs(8422) <= not (a or b);
    layer4_outputs(8423) <= b and not a;
    layer4_outputs(8424) <= not (a and b);
    layer4_outputs(8425) <= a and not b;
    layer4_outputs(8426) <= not a or b;
    layer4_outputs(8427) <= not b;
    layer4_outputs(8428) <= '0';
    layer4_outputs(8429) <= not (a and b);
    layer4_outputs(8430) <= b and not a;
    layer4_outputs(8431) <= not b;
    layer4_outputs(8432) <= a and not b;
    layer4_outputs(8433) <= a or b;
    layer4_outputs(8434) <= a or b;
    layer4_outputs(8435) <= not b;
    layer4_outputs(8436) <= b and not a;
    layer4_outputs(8437) <= not (a or b);
    layer4_outputs(8438) <= not (a and b);
    layer4_outputs(8439) <= a xor b;
    layer4_outputs(8440) <= b;
    layer4_outputs(8441) <= a or b;
    layer4_outputs(8442) <= not (a xor b);
    layer4_outputs(8443) <= b;
    layer4_outputs(8444) <= a;
    layer4_outputs(8445) <= a and not b;
    layer4_outputs(8446) <= a or b;
    layer4_outputs(8447) <= b and not a;
    layer4_outputs(8448) <= not a;
    layer4_outputs(8449) <= b;
    layer4_outputs(8450) <= not a or b;
    layer4_outputs(8451) <= not a;
    layer4_outputs(8452) <= a xor b;
    layer4_outputs(8453) <= a;
    layer4_outputs(8454) <= b;
    layer4_outputs(8455) <= b;
    layer4_outputs(8456) <= a;
    layer4_outputs(8457) <= b and not a;
    layer4_outputs(8458) <= not b or a;
    layer4_outputs(8459) <= not (a xor b);
    layer4_outputs(8460) <= a and b;
    layer4_outputs(8461) <= not b;
    layer4_outputs(8462) <= not a;
    layer4_outputs(8463) <= not (a and b);
    layer4_outputs(8464) <= not (a or b);
    layer4_outputs(8465) <= b and not a;
    layer4_outputs(8466) <= not a;
    layer4_outputs(8467) <= '0';
    layer4_outputs(8468) <= not a;
    layer4_outputs(8469) <= not (a and b);
    layer4_outputs(8470) <= not b;
    layer4_outputs(8471) <= b;
    layer4_outputs(8472) <= b;
    layer4_outputs(8473) <= '0';
    layer4_outputs(8474) <= not (a or b);
    layer4_outputs(8475) <= b and not a;
    layer4_outputs(8476) <= b;
    layer4_outputs(8477) <= not (a and b);
    layer4_outputs(8478) <= b;
    layer4_outputs(8479) <= a;
    layer4_outputs(8480) <= not (a or b);
    layer4_outputs(8481) <= not b;
    layer4_outputs(8482) <= b;
    layer4_outputs(8483) <= not (a and b);
    layer4_outputs(8484) <= not (a and b);
    layer4_outputs(8485) <= not (a xor b);
    layer4_outputs(8486) <= not (a xor b);
    layer4_outputs(8487) <= a and b;
    layer4_outputs(8488) <= not (a and b);
    layer4_outputs(8489) <= b;
    layer4_outputs(8490) <= b;
    layer4_outputs(8491) <= a and not b;
    layer4_outputs(8492) <= a;
    layer4_outputs(8493) <= not (a xor b);
    layer4_outputs(8494) <= not a;
    layer4_outputs(8495) <= not (a or b);
    layer4_outputs(8496) <= b;
    layer4_outputs(8497) <= not b;
    layer4_outputs(8498) <= a;
    layer4_outputs(8499) <= not a;
    layer4_outputs(8500) <= a;
    layer4_outputs(8501) <= a or b;
    layer4_outputs(8502) <= a;
    layer4_outputs(8503) <= not (a xor b);
    layer4_outputs(8504) <= b;
    layer4_outputs(8505) <= not a;
    layer4_outputs(8506) <= not (a or b);
    layer4_outputs(8507) <= b;
    layer4_outputs(8508) <= b and not a;
    layer4_outputs(8509) <= a and b;
    layer4_outputs(8510) <= b and not a;
    layer4_outputs(8511) <= a xor b;
    layer4_outputs(8512) <= b;
    layer4_outputs(8513) <= a;
    layer4_outputs(8514) <= not a;
    layer4_outputs(8515) <= not b or a;
    layer4_outputs(8516) <= a or b;
    layer4_outputs(8517) <= not a or b;
    layer4_outputs(8518) <= not a;
    layer4_outputs(8519) <= not b or a;
    layer4_outputs(8520) <= b and not a;
    layer4_outputs(8521) <= not b;
    layer4_outputs(8522) <= a or b;
    layer4_outputs(8523) <= a xor b;
    layer4_outputs(8524) <= a;
    layer4_outputs(8525) <= b;
    layer4_outputs(8526) <= not b;
    layer4_outputs(8527) <= b;
    layer4_outputs(8528) <= not (a or b);
    layer4_outputs(8529) <= a;
    layer4_outputs(8530) <= not (a xor b);
    layer4_outputs(8531) <= not a or b;
    layer4_outputs(8532) <= not b;
    layer4_outputs(8533) <= not a or b;
    layer4_outputs(8534) <= not a;
    layer4_outputs(8535) <= not (a and b);
    layer4_outputs(8536) <= a and not b;
    layer4_outputs(8537) <= not a or b;
    layer4_outputs(8538) <= not (a and b);
    layer4_outputs(8539) <= a and b;
    layer4_outputs(8540) <= a or b;
    layer4_outputs(8541) <= a and not b;
    layer4_outputs(8542) <= a or b;
    layer4_outputs(8543) <= not (a or b);
    layer4_outputs(8544) <= b and not a;
    layer4_outputs(8545) <= a;
    layer4_outputs(8546) <= a;
    layer4_outputs(8547) <= not b or a;
    layer4_outputs(8548) <= b;
    layer4_outputs(8549) <= not a or b;
    layer4_outputs(8550) <= not a;
    layer4_outputs(8551) <= not a or b;
    layer4_outputs(8552) <= not b or a;
    layer4_outputs(8553) <= not b or a;
    layer4_outputs(8554) <= b and not a;
    layer4_outputs(8555) <= not a;
    layer4_outputs(8556) <= not a;
    layer4_outputs(8557) <= a;
    layer4_outputs(8558) <= not a;
    layer4_outputs(8559) <= not a;
    layer4_outputs(8560) <= not b;
    layer4_outputs(8561) <= b;
    layer4_outputs(8562) <= a xor b;
    layer4_outputs(8563) <= a;
    layer4_outputs(8564) <= not a;
    layer4_outputs(8565) <= a xor b;
    layer4_outputs(8566) <= b;
    layer4_outputs(8567) <= b;
    layer4_outputs(8568) <= b;
    layer4_outputs(8569) <= a and not b;
    layer4_outputs(8570) <= b and not a;
    layer4_outputs(8571) <= not b;
    layer4_outputs(8572) <= a;
    layer4_outputs(8573) <= a and not b;
    layer4_outputs(8574) <= not a or b;
    layer4_outputs(8575) <= not a;
    layer4_outputs(8576) <= b;
    layer4_outputs(8577) <= a and b;
    layer4_outputs(8578) <= not b;
    layer4_outputs(8579) <= b and not a;
    layer4_outputs(8580) <= not a;
    layer4_outputs(8581) <= not a or b;
    layer4_outputs(8582) <= not a or b;
    layer4_outputs(8583) <= a and b;
    layer4_outputs(8584) <= a or b;
    layer4_outputs(8585) <= b;
    layer4_outputs(8586) <= b;
    layer4_outputs(8587) <= not b;
    layer4_outputs(8588) <= a and b;
    layer4_outputs(8589) <= a xor b;
    layer4_outputs(8590) <= b;
    layer4_outputs(8591) <= not a;
    layer4_outputs(8592) <= not (a or b);
    layer4_outputs(8593) <= not (a or b);
    layer4_outputs(8594) <= not a;
    layer4_outputs(8595) <= '1';
    layer4_outputs(8596) <= not a;
    layer4_outputs(8597) <= not a or b;
    layer4_outputs(8598) <= a or b;
    layer4_outputs(8599) <= not a;
    layer4_outputs(8600) <= not b or a;
    layer4_outputs(8601) <= '0';
    layer4_outputs(8602) <= a and b;
    layer4_outputs(8603) <= not b;
    layer4_outputs(8604) <= not a;
    layer4_outputs(8605) <= a;
    layer4_outputs(8606) <= a;
    layer4_outputs(8607) <= b;
    layer4_outputs(8608) <= a;
    layer4_outputs(8609) <= not (a or b);
    layer4_outputs(8610) <= a xor b;
    layer4_outputs(8611) <= not b or a;
    layer4_outputs(8612) <= b and not a;
    layer4_outputs(8613) <= not a;
    layer4_outputs(8614) <= b;
    layer4_outputs(8615) <= a and not b;
    layer4_outputs(8616) <= a xor b;
    layer4_outputs(8617) <= not b;
    layer4_outputs(8618) <= not a or b;
    layer4_outputs(8619) <= not (a xor b);
    layer4_outputs(8620) <= not (a xor b);
    layer4_outputs(8621) <= '1';
    layer4_outputs(8622) <= not a or b;
    layer4_outputs(8623) <= not (a or b);
    layer4_outputs(8624) <= not b or a;
    layer4_outputs(8625) <= not b or a;
    layer4_outputs(8626) <= a and not b;
    layer4_outputs(8627) <= a and b;
    layer4_outputs(8628) <= not (a and b);
    layer4_outputs(8629) <= a;
    layer4_outputs(8630) <= a;
    layer4_outputs(8631) <= a and b;
    layer4_outputs(8632) <= a and b;
    layer4_outputs(8633) <= not (a or b);
    layer4_outputs(8634) <= not a;
    layer4_outputs(8635) <= a;
    layer4_outputs(8636) <= a;
    layer4_outputs(8637) <= not b;
    layer4_outputs(8638) <= b;
    layer4_outputs(8639) <= b;
    layer4_outputs(8640) <= a;
    layer4_outputs(8641) <= not a or b;
    layer4_outputs(8642) <= b;
    layer4_outputs(8643) <= a and b;
    layer4_outputs(8644) <= a and b;
    layer4_outputs(8645) <= '0';
    layer4_outputs(8646) <= not (a or b);
    layer4_outputs(8647) <= not b;
    layer4_outputs(8648) <= not (a or b);
    layer4_outputs(8649) <= a or b;
    layer4_outputs(8650) <= a xor b;
    layer4_outputs(8651) <= a xor b;
    layer4_outputs(8652) <= a xor b;
    layer4_outputs(8653) <= a or b;
    layer4_outputs(8654) <= a and b;
    layer4_outputs(8655) <= a or b;
    layer4_outputs(8656) <= b;
    layer4_outputs(8657) <= b and not a;
    layer4_outputs(8658) <= a and not b;
    layer4_outputs(8659) <= a xor b;
    layer4_outputs(8660) <= not (a or b);
    layer4_outputs(8661) <= not b;
    layer4_outputs(8662) <= a xor b;
    layer4_outputs(8663) <= not b;
    layer4_outputs(8664) <= not (a xor b);
    layer4_outputs(8665) <= not a;
    layer4_outputs(8666) <= a or b;
    layer4_outputs(8667) <= not a;
    layer4_outputs(8668) <= a and not b;
    layer4_outputs(8669) <= a or b;
    layer4_outputs(8670) <= not a;
    layer4_outputs(8671) <= a;
    layer4_outputs(8672) <= a xor b;
    layer4_outputs(8673) <= a and not b;
    layer4_outputs(8674) <= not a;
    layer4_outputs(8675) <= a and not b;
    layer4_outputs(8676) <= not (a and b);
    layer4_outputs(8677) <= b;
    layer4_outputs(8678) <= not (a or b);
    layer4_outputs(8679) <= a or b;
    layer4_outputs(8680) <= a and b;
    layer4_outputs(8681) <= b;
    layer4_outputs(8682) <= a;
    layer4_outputs(8683) <= a;
    layer4_outputs(8684) <= a xor b;
    layer4_outputs(8685) <= a xor b;
    layer4_outputs(8686) <= not (a or b);
    layer4_outputs(8687) <= a and b;
    layer4_outputs(8688) <= not (a xor b);
    layer4_outputs(8689) <= not b;
    layer4_outputs(8690) <= b and not a;
    layer4_outputs(8691) <= a and not b;
    layer4_outputs(8692) <= b and not a;
    layer4_outputs(8693) <= not b;
    layer4_outputs(8694) <= b;
    layer4_outputs(8695) <= not b or a;
    layer4_outputs(8696) <= not b;
    layer4_outputs(8697) <= a;
    layer4_outputs(8698) <= not a or b;
    layer4_outputs(8699) <= a;
    layer4_outputs(8700) <= a;
    layer4_outputs(8701) <= a;
    layer4_outputs(8702) <= not b or a;
    layer4_outputs(8703) <= '1';
    layer4_outputs(8704) <= a and b;
    layer4_outputs(8705) <= not (a or b);
    layer4_outputs(8706) <= b;
    layer4_outputs(8707) <= not (a and b);
    layer4_outputs(8708) <= a or b;
    layer4_outputs(8709) <= not b;
    layer4_outputs(8710) <= not (a xor b);
    layer4_outputs(8711) <= not a;
    layer4_outputs(8712) <= a and not b;
    layer4_outputs(8713) <= not b;
    layer4_outputs(8714) <= '1';
    layer4_outputs(8715) <= not a;
    layer4_outputs(8716) <= not (a xor b);
    layer4_outputs(8717) <= not a;
    layer4_outputs(8718) <= a and not b;
    layer4_outputs(8719) <= not b or a;
    layer4_outputs(8720) <= not (a or b);
    layer4_outputs(8721) <= a or b;
    layer4_outputs(8722) <= not a;
    layer4_outputs(8723) <= a;
    layer4_outputs(8724) <= b;
    layer4_outputs(8725) <= not (a xor b);
    layer4_outputs(8726) <= not b;
    layer4_outputs(8727) <= a xor b;
    layer4_outputs(8728) <= b;
    layer4_outputs(8729) <= not b;
    layer4_outputs(8730) <= not b;
    layer4_outputs(8731) <= not a;
    layer4_outputs(8732) <= '1';
    layer4_outputs(8733) <= '1';
    layer4_outputs(8734) <= not a;
    layer4_outputs(8735) <= a;
    layer4_outputs(8736) <= not (a or b);
    layer4_outputs(8737) <= not a;
    layer4_outputs(8738) <= not (a and b);
    layer4_outputs(8739) <= b;
    layer4_outputs(8740) <= not a or b;
    layer4_outputs(8741) <= not (a or b);
    layer4_outputs(8742) <= a and not b;
    layer4_outputs(8743) <= not b or a;
    layer4_outputs(8744) <= not (a or b);
    layer4_outputs(8745) <= a or b;
    layer4_outputs(8746) <= not (a and b);
    layer4_outputs(8747) <= a;
    layer4_outputs(8748) <= a xor b;
    layer4_outputs(8749) <= a xor b;
    layer4_outputs(8750) <= '1';
    layer4_outputs(8751) <= not a;
    layer4_outputs(8752) <= not (a and b);
    layer4_outputs(8753) <= not b;
    layer4_outputs(8754) <= a or b;
    layer4_outputs(8755) <= not b or a;
    layer4_outputs(8756) <= a and b;
    layer4_outputs(8757) <= a;
    layer4_outputs(8758) <= not a;
    layer4_outputs(8759) <= not (a xor b);
    layer4_outputs(8760) <= a and b;
    layer4_outputs(8761) <= a xor b;
    layer4_outputs(8762) <= a xor b;
    layer4_outputs(8763) <= not b;
    layer4_outputs(8764) <= b and not a;
    layer4_outputs(8765) <= a or b;
    layer4_outputs(8766) <= not b;
    layer4_outputs(8767) <= not a;
    layer4_outputs(8768) <= a or b;
    layer4_outputs(8769) <= '0';
    layer4_outputs(8770) <= a;
    layer4_outputs(8771) <= a or b;
    layer4_outputs(8772) <= not (a and b);
    layer4_outputs(8773) <= not (a and b);
    layer4_outputs(8774) <= not b;
    layer4_outputs(8775) <= not b or a;
    layer4_outputs(8776) <= b and not a;
    layer4_outputs(8777) <= not b or a;
    layer4_outputs(8778) <= b;
    layer4_outputs(8779) <= b and not a;
    layer4_outputs(8780) <= a and b;
    layer4_outputs(8781) <= a or b;
    layer4_outputs(8782) <= b and not a;
    layer4_outputs(8783) <= not a or b;
    layer4_outputs(8784) <= not a;
    layer4_outputs(8785) <= a xor b;
    layer4_outputs(8786) <= not (a and b);
    layer4_outputs(8787) <= '0';
    layer4_outputs(8788) <= '1';
    layer4_outputs(8789) <= not a;
    layer4_outputs(8790) <= b;
    layer4_outputs(8791) <= a or b;
    layer4_outputs(8792) <= a;
    layer4_outputs(8793) <= a;
    layer4_outputs(8794) <= not (a xor b);
    layer4_outputs(8795) <= a xor b;
    layer4_outputs(8796) <= a and not b;
    layer4_outputs(8797) <= a and b;
    layer4_outputs(8798) <= not (a or b);
    layer4_outputs(8799) <= '0';
    layer4_outputs(8800) <= not a;
    layer4_outputs(8801) <= not a;
    layer4_outputs(8802) <= a and not b;
    layer4_outputs(8803) <= b;
    layer4_outputs(8804) <= not b;
    layer4_outputs(8805) <= not b;
    layer4_outputs(8806) <= '1';
    layer4_outputs(8807) <= '1';
    layer4_outputs(8808) <= not a;
    layer4_outputs(8809) <= b;
    layer4_outputs(8810) <= not a or b;
    layer4_outputs(8811) <= not a;
    layer4_outputs(8812) <= not (a or b);
    layer4_outputs(8813) <= not a;
    layer4_outputs(8814) <= not (a and b);
    layer4_outputs(8815) <= a;
    layer4_outputs(8816) <= a and b;
    layer4_outputs(8817) <= a and not b;
    layer4_outputs(8818) <= b and not a;
    layer4_outputs(8819) <= not b;
    layer4_outputs(8820) <= b;
    layer4_outputs(8821) <= not a;
    layer4_outputs(8822) <= not b;
    layer4_outputs(8823) <= not a or b;
    layer4_outputs(8824) <= a and not b;
    layer4_outputs(8825) <= a and b;
    layer4_outputs(8826) <= b;
    layer4_outputs(8827) <= not b or a;
    layer4_outputs(8828) <= '0';
    layer4_outputs(8829) <= not (a xor b);
    layer4_outputs(8830) <= a and not b;
    layer4_outputs(8831) <= not b or a;
    layer4_outputs(8832) <= a;
    layer4_outputs(8833) <= b and not a;
    layer4_outputs(8834) <= a and b;
    layer4_outputs(8835) <= a xor b;
    layer4_outputs(8836) <= not (a or b);
    layer4_outputs(8837) <= not b or a;
    layer4_outputs(8838) <= b and not a;
    layer4_outputs(8839) <= a and not b;
    layer4_outputs(8840) <= a;
    layer4_outputs(8841) <= not a;
    layer4_outputs(8842) <= a;
    layer4_outputs(8843) <= not b;
    layer4_outputs(8844) <= '0';
    layer4_outputs(8845) <= not (a xor b);
    layer4_outputs(8846) <= not b;
    layer4_outputs(8847) <= b and not a;
    layer4_outputs(8848) <= a and b;
    layer4_outputs(8849) <= not (a or b);
    layer4_outputs(8850) <= a and not b;
    layer4_outputs(8851) <= not b;
    layer4_outputs(8852) <= not (a and b);
    layer4_outputs(8853) <= a and not b;
    layer4_outputs(8854) <= not a;
    layer4_outputs(8855) <= a;
    layer4_outputs(8856) <= a and b;
    layer4_outputs(8857) <= not a or b;
    layer4_outputs(8858) <= a;
    layer4_outputs(8859) <= not (a and b);
    layer4_outputs(8860) <= not a;
    layer4_outputs(8861) <= a and not b;
    layer4_outputs(8862) <= b;
    layer4_outputs(8863) <= b;
    layer4_outputs(8864) <= not b;
    layer4_outputs(8865) <= not a;
    layer4_outputs(8866) <= a or b;
    layer4_outputs(8867) <= not b or a;
    layer4_outputs(8868) <= not (a xor b);
    layer4_outputs(8869) <= a and not b;
    layer4_outputs(8870) <= not a;
    layer4_outputs(8871) <= a;
    layer4_outputs(8872) <= b;
    layer4_outputs(8873) <= a and not b;
    layer4_outputs(8874) <= not b;
    layer4_outputs(8875) <= not b;
    layer4_outputs(8876) <= a;
    layer4_outputs(8877) <= a xor b;
    layer4_outputs(8878) <= not a;
    layer4_outputs(8879) <= not (a and b);
    layer4_outputs(8880) <= b;
    layer4_outputs(8881) <= '0';
    layer4_outputs(8882) <= not a or b;
    layer4_outputs(8883) <= not (a and b);
    layer4_outputs(8884) <= a or b;
    layer4_outputs(8885) <= not (a or b);
    layer4_outputs(8886) <= a;
    layer4_outputs(8887) <= a or b;
    layer4_outputs(8888) <= b;
    layer4_outputs(8889) <= a or b;
    layer4_outputs(8890) <= not b;
    layer4_outputs(8891) <= a;
    layer4_outputs(8892) <= a and not b;
    layer4_outputs(8893) <= a;
    layer4_outputs(8894) <= not b or a;
    layer4_outputs(8895) <= a;
    layer4_outputs(8896) <= not a;
    layer4_outputs(8897) <= not a;
    layer4_outputs(8898) <= not a;
    layer4_outputs(8899) <= not b;
    layer4_outputs(8900) <= b;
    layer4_outputs(8901) <= not (a or b);
    layer4_outputs(8902) <= a and not b;
    layer4_outputs(8903) <= b and not a;
    layer4_outputs(8904) <= not a or b;
    layer4_outputs(8905) <= not b or a;
    layer4_outputs(8906) <= not b or a;
    layer4_outputs(8907) <= not a;
    layer4_outputs(8908) <= not b or a;
    layer4_outputs(8909) <= b and not a;
    layer4_outputs(8910) <= not b or a;
    layer4_outputs(8911) <= not a;
    layer4_outputs(8912) <= a;
    layer4_outputs(8913) <= a xor b;
    layer4_outputs(8914) <= b and not a;
    layer4_outputs(8915) <= a or b;
    layer4_outputs(8916) <= a and not b;
    layer4_outputs(8917) <= not a;
    layer4_outputs(8918) <= not a or b;
    layer4_outputs(8919) <= '1';
    layer4_outputs(8920) <= a and b;
    layer4_outputs(8921) <= not b or a;
    layer4_outputs(8922) <= not (a xor b);
    layer4_outputs(8923) <= not (a and b);
    layer4_outputs(8924) <= not a;
    layer4_outputs(8925) <= not (a and b);
    layer4_outputs(8926) <= not (a and b);
    layer4_outputs(8927) <= a xor b;
    layer4_outputs(8928) <= a xor b;
    layer4_outputs(8929) <= '0';
    layer4_outputs(8930) <= not (a or b);
    layer4_outputs(8931) <= not a;
    layer4_outputs(8932) <= not a;
    layer4_outputs(8933) <= '0';
    layer4_outputs(8934) <= a;
    layer4_outputs(8935) <= b;
    layer4_outputs(8936) <= '0';
    layer4_outputs(8937) <= a;
    layer4_outputs(8938) <= not (a or b);
    layer4_outputs(8939) <= not (a or b);
    layer4_outputs(8940) <= a and b;
    layer4_outputs(8941) <= '1';
    layer4_outputs(8942) <= not a or b;
    layer4_outputs(8943) <= '0';
    layer4_outputs(8944) <= a;
    layer4_outputs(8945) <= a or b;
    layer4_outputs(8946) <= b;
    layer4_outputs(8947) <= not b or a;
    layer4_outputs(8948) <= not (a or b);
    layer4_outputs(8949) <= a and not b;
    layer4_outputs(8950) <= a and not b;
    layer4_outputs(8951) <= not b;
    layer4_outputs(8952) <= a and not b;
    layer4_outputs(8953) <= not (a and b);
    layer4_outputs(8954) <= b and not a;
    layer4_outputs(8955) <= '1';
    layer4_outputs(8956) <= b;
    layer4_outputs(8957) <= not (a xor b);
    layer4_outputs(8958) <= b;
    layer4_outputs(8959) <= a and b;
    layer4_outputs(8960) <= not (a and b);
    layer4_outputs(8961) <= a and b;
    layer4_outputs(8962) <= a;
    layer4_outputs(8963) <= a and not b;
    layer4_outputs(8964) <= a or b;
    layer4_outputs(8965) <= not a or b;
    layer4_outputs(8966) <= a or b;
    layer4_outputs(8967) <= not b or a;
    layer4_outputs(8968) <= not a;
    layer4_outputs(8969) <= not a;
    layer4_outputs(8970) <= b and not a;
    layer4_outputs(8971) <= b;
    layer4_outputs(8972) <= not b;
    layer4_outputs(8973) <= a or b;
    layer4_outputs(8974) <= b;
    layer4_outputs(8975) <= a;
    layer4_outputs(8976) <= not (a or b);
    layer4_outputs(8977) <= not b or a;
    layer4_outputs(8978) <= not (a and b);
    layer4_outputs(8979) <= '1';
    layer4_outputs(8980) <= not a;
    layer4_outputs(8981) <= a and b;
    layer4_outputs(8982) <= b and not a;
    layer4_outputs(8983) <= b and not a;
    layer4_outputs(8984) <= b;
    layer4_outputs(8985) <= a;
    layer4_outputs(8986) <= not b;
    layer4_outputs(8987) <= b;
    layer4_outputs(8988) <= b;
    layer4_outputs(8989) <= not (a or b);
    layer4_outputs(8990) <= b and not a;
    layer4_outputs(8991) <= not b or a;
    layer4_outputs(8992) <= not b;
    layer4_outputs(8993) <= not a;
    layer4_outputs(8994) <= not b or a;
    layer4_outputs(8995) <= not a;
    layer4_outputs(8996) <= not b or a;
    layer4_outputs(8997) <= not b;
    layer4_outputs(8998) <= a xor b;
    layer4_outputs(8999) <= not (a xor b);
    layer4_outputs(9000) <= a or b;
    layer4_outputs(9001) <= not a or b;
    layer4_outputs(9002) <= not a or b;
    layer4_outputs(9003) <= not a or b;
    layer4_outputs(9004) <= b;
    layer4_outputs(9005) <= not b;
    layer4_outputs(9006) <= a;
    layer4_outputs(9007) <= not (a or b);
    layer4_outputs(9008) <= a or b;
    layer4_outputs(9009) <= a;
    layer4_outputs(9010) <= not a;
    layer4_outputs(9011) <= not a;
    layer4_outputs(9012) <= a xor b;
    layer4_outputs(9013) <= not b;
    layer4_outputs(9014) <= a;
    layer4_outputs(9015) <= b and not a;
    layer4_outputs(9016) <= a;
    layer4_outputs(9017) <= a;
    layer4_outputs(9018) <= not a;
    layer4_outputs(9019) <= a and not b;
    layer4_outputs(9020) <= not b;
    layer4_outputs(9021) <= a and b;
    layer4_outputs(9022) <= b;
    layer4_outputs(9023) <= not a or b;
    layer4_outputs(9024) <= a;
    layer4_outputs(9025) <= a;
    layer4_outputs(9026) <= not (a or b);
    layer4_outputs(9027) <= not (a or b);
    layer4_outputs(9028) <= not (a and b);
    layer4_outputs(9029) <= a;
    layer4_outputs(9030) <= not a or b;
    layer4_outputs(9031) <= not a;
    layer4_outputs(9032) <= b;
    layer4_outputs(9033) <= not b or a;
    layer4_outputs(9034) <= a;
    layer4_outputs(9035) <= not a;
    layer4_outputs(9036) <= a and b;
    layer4_outputs(9037) <= not a;
    layer4_outputs(9038) <= not (a or b);
    layer4_outputs(9039) <= b;
    layer4_outputs(9040) <= not b;
    layer4_outputs(9041) <= not (a or b);
    layer4_outputs(9042) <= a and not b;
    layer4_outputs(9043) <= a xor b;
    layer4_outputs(9044) <= not (a or b);
    layer4_outputs(9045) <= not (a and b);
    layer4_outputs(9046) <= not (a and b);
    layer4_outputs(9047) <= not b;
    layer4_outputs(9048) <= a;
    layer4_outputs(9049) <= a xor b;
    layer4_outputs(9050) <= a;
    layer4_outputs(9051) <= a or b;
    layer4_outputs(9052) <= a;
    layer4_outputs(9053) <= not a or b;
    layer4_outputs(9054) <= not b;
    layer4_outputs(9055) <= not a or b;
    layer4_outputs(9056) <= a;
    layer4_outputs(9057) <= b;
    layer4_outputs(9058) <= a;
    layer4_outputs(9059) <= a or b;
    layer4_outputs(9060) <= '1';
    layer4_outputs(9061) <= not (a xor b);
    layer4_outputs(9062) <= a and b;
    layer4_outputs(9063) <= not a or b;
    layer4_outputs(9064) <= b and not a;
    layer4_outputs(9065) <= not b or a;
    layer4_outputs(9066) <= a;
    layer4_outputs(9067) <= not b;
    layer4_outputs(9068) <= not (a or b);
    layer4_outputs(9069) <= not a;
    layer4_outputs(9070) <= not b;
    layer4_outputs(9071) <= a or b;
    layer4_outputs(9072) <= not b or a;
    layer4_outputs(9073) <= a and b;
    layer4_outputs(9074) <= b;
    layer4_outputs(9075) <= a or b;
    layer4_outputs(9076) <= a and not b;
    layer4_outputs(9077) <= not (a and b);
    layer4_outputs(9078) <= not (a xor b);
    layer4_outputs(9079) <= a xor b;
    layer4_outputs(9080) <= not a;
    layer4_outputs(9081) <= not (a and b);
    layer4_outputs(9082) <= not a or b;
    layer4_outputs(9083) <= '0';
    layer4_outputs(9084) <= a;
    layer4_outputs(9085) <= not (a or b);
    layer4_outputs(9086) <= a and b;
    layer4_outputs(9087) <= a;
    layer4_outputs(9088) <= not b;
    layer4_outputs(9089) <= a;
    layer4_outputs(9090) <= not b or a;
    layer4_outputs(9091) <= a and not b;
    layer4_outputs(9092) <= not b or a;
    layer4_outputs(9093) <= not b;
    layer4_outputs(9094) <= a and b;
    layer4_outputs(9095) <= a xor b;
    layer4_outputs(9096) <= a or b;
    layer4_outputs(9097) <= not (a and b);
    layer4_outputs(9098) <= b;
    layer4_outputs(9099) <= not a or b;
    layer4_outputs(9100) <= not a or b;
    layer4_outputs(9101) <= not (a and b);
    layer4_outputs(9102) <= a;
    layer4_outputs(9103) <= not a or b;
    layer4_outputs(9104) <= not a or b;
    layer4_outputs(9105) <= b;
    layer4_outputs(9106) <= not b;
    layer4_outputs(9107) <= not (a and b);
    layer4_outputs(9108) <= b;
    layer4_outputs(9109) <= '0';
    layer4_outputs(9110) <= a and b;
    layer4_outputs(9111) <= a;
    layer4_outputs(9112) <= not a or b;
    layer4_outputs(9113) <= not (a or b);
    layer4_outputs(9114) <= '1';
    layer4_outputs(9115) <= b and not a;
    layer4_outputs(9116) <= b;
    layer4_outputs(9117) <= '1';
    layer4_outputs(9118) <= b and not a;
    layer4_outputs(9119) <= not a;
    layer4_outputs(9120) <= not b or a;
    layer4_outputs(9121) <= a or b;
    layer4_outputs(9122) <= '1';
    layer4_outputs(9123) <= not (a and b);
    layer4_outputs(9124) <= not a or b;
    layer4_outputs(9125) <= not b or a;
    layer4_outputs(9126) <= b and not a;
    layer4_outputs(9127) <= b;
    layer4_outputs(9128) <= not b;
    layer4_outputs(9129) <= a and not b;
    layer4_outputs(9130) <= a;
    layer4_outputs(9131) <= b;
    layer4_outputs(9132) <= b;
    layer4_outputs(9133) <= a;
    layer4_outputs(9134) <= not (a or b);
    layer4_outputs(9135) <= a;
    layer4_outputs(9136) <= b;
    layer4_outputs(9137) <= a and not b;
    layer4_outputs(9138) <= not b;
    layer4_outputs(9139) <= a and not b;
    layer4_outputs(9140) <= not a or b;
    layer4_outputs(9141) <= not a;
    layer4_outputs(9142) <= a and not b;
    layer4_outputs(9143) <= '1';
    layer4_outputs(9144) <= not b;
    layer4_outputs(9145) <= a xor b;
    layer4_outputs(9146) <= not b;
    layer4_outputs(9147) <= not a or b;
    layer4_outputs(9148) <= not b;
    layer4_outputs(9149) <= a;
    layer4_outputs(9150) <= not a;
    layer4_outputs(9151) <= not a or b;
    layer4_outputs(9152) <= not b;
    layer4_outputs(9153) <= not b;
    layer4_outputs(9154) <= a or b;
    layer4_outputs(9155) <= a xor b;
    layer4_outputs(9156) <= b;
    layer4_outputs(9157) <= not a or b;
    layer4_outputs(9158) <= b;
    layer4_outputs(9159) <= not (a xor b);
    layer4_outputs(9160) <= a;
    layer4_outputs(9161) <= not a;
    layer4_outputs(9162) <= not (a or b);
    layer4_outputs(9163) <= not (a xor b);
    layer4_outputs(9164) <= '0';
    layer4_outputs(9165) <= a and b;
    layer4_outputs(9166) <= not b;
    layer4_outputs(9167) <= a or b;
    layer4_outputs(9168) <= not a;
    layer4_outputs(9169) <= not a;
    layer4_outputs(9170) <= '0';
    layer4_outputs(9171) <= a or b;
    layer4_outputs(9172) <= a and not b;
    layer4_outputs(9173) <= a and b;
    layer4_outputs(9174) <= '0';
    layer4_outputs(9175) <= b;
    layer4_outputs(9176) <= a;
    layer4_outputs(9177) <= a or b;
    layer4_outputs(9178) <= b;
    layer4_outputs(9179) <= a;
    layer4_outputs(9180) <= a;
    layer4_outputs(9181) <= a and not b;
    layer4_outputs(9182) <= not b or a;
    layer4_outputs(9183) <= b;
    layer4_outputs(9184) <= not b or a;
    layer4_outputs(9185) <= not a or b;
    layer4_outputs(9186) <= a or b;
    layer4_outputs(9187) <= not (a or b);
    layer4_outputs(9188) <= a and b;
    layer4_outputs(9189) <= not a;
    layer4_outputs(9190) <= not a;
    layer4_outputs(9191) <= not a or b;
    layer4_outputs(9192) <= a and not b;
    layer4_outputs(9193) <= a or b;
    layer4_outputs(9194) <= b and not a;
    layer4_outputs(9195) <= a or b;
    layer4_outputs(9196) <= b;
    layer4_outputs(9197) <= a;
    layer4_outputs(9198) <= a or b;
    layer4_outputs(9199) <= not b;
    layer4_outputs(9200) <= b;
    layer4_outputs(9201) <= b and not a;
    layer4_outputs(9202) <= a;
    layer4_outputs(9203) <= not a;
    layer4_outputs(9204) <= b;
    layer4_outputs(9205) <= not a;
    layer4_outputs(9206) <= not b;
    layer4_outputs(9207) <= b and not a;
    layer4_outputs(9208) <= not a;
    layer4_outputs(9209) <= not b;
    layer4_outputs(9210) <= b and not a;
    layer4_outputs(9211) <= not a or b;
    layer4_outputs(9212) <= not a;
    layer4_outputs(9213) <= b and not a;
    layer4_outputs(9214) <= not b;
    layer4_outputs(9215) <= a;
    layer4_outputs(9216) <= not (a xor b);
    layer4_outputs(9217) <= a;
    layer4_outputs(9218) <= b and not a;
    layer4_outputs(9219) <= a and b;
    layer4_outputs(9220) <= b;
    layer4_outputs(9221) <= not b;
    layer4_outputs(9222) <= a xor b;
    layer4_outputs(9223) <= not (a or b);
    layer4_outputs(9224) <= '1';
    layer4_outputs(9225) <= b and not a;
    layer4_outputs(9226) <= not b;
    layer4_outputs(9227) <= not a;
    layer4_outputs(9228) <= a and b;
    layer4_outputs(9229) <= b;
    layer4_outputs(9230) <= b and not a;
    layer4_outputs(9231) <= not a;
    layer4_outputs(9232) <= b;
    layer4_outputs(9233) <= b;
    layer4_outputs(9234) <= b and not a;
    layer4_outputs(9235) <= not b;
    layer4_outputs(9236) <= not b;
    layer4_outputs(9237) <= b;
    layer4_outputs(9238) <= b;
    layer4_outputs(9239) <= not a or b;
    layer4_outputs(9240) <= a xor b;
    layer4_outputs(9241) <= not b;
    layer4_outputs(9242) <= not a or b;
    layer4_outputs(9243) <= a;
    layer4_outputs(9244) <= a;
    layer4_outputs(9245) <= not b;
    layer4_outputs(9246) <= not (a and b);
    layer4_outputs(9247) <= b;
    layer4_outputs(9248) <= not a;
    layer4_outputs(9249) <= a and b;
    layer4_outputs(9250) <= not a or b;
    layer4_outputs(9251) <= not b or a;
    layer4_outputs(9252) <= not b or a;
    layer4_outputs(9253) <= b and not a;
    layer4_outputs(9254) <= a or b;
    layer4_outputs(9255) <= a and not b;
    layer4_outputs(9256) <= a xor b;
    layer4_outputs(9257) <= not a;
    layer4_outputs(9258) <= '0';
    layer4_outputs(9259) <= not b;
    layer4_outputs(9260) <= a or b;
    layer4_outputs(9261) <= not a;
    layer4_outputs(9262) <= not b or a;
    layer4_outputs(9263) <= not b;
    layer4_outputs(9264) <= '0';
    layer4_outputs(9265) <= b;
    layer4_outputs(9266) <= '0';
    layer4_outputs(9267) <= a and not b;
    layer4_outputs(9268) <= not a or b;
    layer4_outputs(9269) <= a;
    layer4_outputs(9270) <= a;
    layer4_outputs(9271) <= a;
    layer4_outputs(9272) <= a and b;
    layer4_outputs(9273) <= not (a or b);
    layer4_outputs(9274) <= b;
    layer4_outputs(9275) <= a and b;
    layer4_outputs(9276) <= not (a xor b);
    layer4_outputs(9277) <= a and b;
    layer4_outputs(9278) <= not a;
    layer4_outputs(9279) <= not a or b;
    layer4_outputs(9280) <= a;
    layer4_outputs(9281) <= a;
    layer4_outputs(9282) <= a xor b;
    layer4_outputs(9283) <= not b or a;
    layer4_outputs(9284) <= not a or b;
    layer4_outputs(9285) <= not b or a;
    layer4_outputs(9286) <= not (a or b);
    layer4_outputs(9287) <= not a or b;
    layer4_outputs(9288) <= b and not a;
    layer4_outputs(9289) <= not (a or b);
    layer4_outputs(9290) <= not (a and b);
    layer4_outputs(9291) <= a or b;
    layer4_outputs(9292) <= not b;
    layer4_outputs(9293) <= b and not a;
    layer4_outputs(9294) <= b and not a;
    layer4_outputs(9295) <= a or b;
    layer4_outputs(9296) <= not b;
    layer4_outputs(9297) <= not b or a;
    layer4_outputs(9298) <= not b;
    layer4_outputs(9299) <= not (a or b);
    layer4_outputs(9300) <= not b;
    layer4_outputs(9301) <= b;
    layer4_outputs(9302) <= not a;
    layer4_outputs(9303) <= b and not a;
    layer4_outputs(9304) <= not b;
    layer4_outputs(9305) <= not b or a;
    layer4_outputs(9306) <= not a or b;
    layer4_outputs(9307) <= a and not b;
    layer4_outputs(9308) <= b;
    layer4_outputs(9309) <= not (a and b);
    layer4_outputs(9310) <= b and not a;
    layer4_outputs(9311) <= a;
    layer4_outputs(9312) <= not (a and b);
    layer4_outputs(9313) <= b and not a;
    layer4_outputs(9314) <= not b;
    layer4_outputs(9315) <= a;
    layer4_outputs(9316) <= a;
    layer4_outputs(9317) <= not (a xor b);
    layer4_outputs(9318) <= a or b;
    layer4_outputs(9319) <= a or b;
    layer4_outputs(9320) <= a and b;
    layer4_outputs(9321) <= b and not a;
    layer4_outputs(9322) <= not b;
    layer4_outputs(9323) <= not (a xor b);
    layer4_outputs(9324) <= '0';
    layer4_outputs(9325) <= a xor b;
    layer4_outputs(9326) <= not b;
    layer4_outputs(9327) <= b;
    layer4_outputs(9328) <= a and not b;
    layer4_outputs(9329) <= not b;
    layer4_outputs(9330) <= not (a or b);
    layer4_outputs(9331) <= a;
    layer4_outputs(9332) <= b;
    layer4_outputs(9333) <= not b;
    layer4_outputs(9334) <= not b;
    layer4_outputs(9335) <= b;
    layer4_outputs(9336) <= a or b;
    layer4_outputs(9337) <= b and not a;
    layer4_outputs(9338) <= a;
    layer4_outputs(9339) <= b;
    layer4_outputs(9340) <= not a;
    layer4_outputs(9341) <= not a or b;
    layer4_outputs(9342) <= not (a and b);
    layer4_outputs(9343) <= a;
    layer4_outputs(9344) <= not (a xor b);
    layer4_outputs(9345) <= b;
    layer4_outputs(9346) <= a or b;
    layer4_outputs(9347) <= not b;
    layer4_outputs(9348) <= not a or b;
    layer4_outputs(9349) <= not b;
    layer4_outputs(9350) <= not b or a;
    layer4_outputs(9351) <= not a;
    layer4_outputs(9352) <= not b or a;
    layer4_outputs(9353) <= not b;
    layer4_outputs(9354) <= not a;
    layer4_outputs(9355) <= b;
    layer4_outputs(9356) <= a and not b;
    layer4_outputs(9357) <= b;
    layer4_outputs(9358) <= a xor b;
    layer4_outputs(9359) <= a;
    layer4_outputs(9360) <= a and b;
    layer4_outputs(9361) <= '0';
    layer4_outputs(9362) <= a and b;
    layer4_outputs(9363) <= not b;
    layer4_outputs(9364) <= a and b;
    layer4_outputs(9365) <= not a or b;
    layer4_outputs(9366) <= not a;
    layer4_outputs(9367) <= not (a or b);
    layer4_outputs(9368) <= '1';
    layer4_outputs(9369) <= not a;
    layer4_outputs(9370) <= not b or a;
    layer4_outputs(9371) <= not b or a;
    layer4_outputs(9372) <= a;
    layer4_outputs(9373) <= '0';
    layer4_outputs(9374) <= a and not b;
    layer4_outputs(9375) <= a and b;
    layer4_outputs(9376) <= a and not b;
    layer4_outputs(9377) <= a;
    layer4_outputs(9378) <= not b or a;
    layer4_outputs(9379) <= not b;
    layer4_outputs(9380) <= not b;
    layer4_outputs(9381) <= not (a or b);
    layer4_outputs(9382) <= not b;
    layer4_outputs(9383) <= '1';
    layer4_outputs(9384) <= '1';
    layer4_outputs(9385) <= a and b;
    layer4_outputs(9386) <= not (a xor b);
    layer4_outputs(9387) <= a;
    layer4_outputs(9388) <= b;
    layer4_outputs(9389) <= not (a xor b);
    layer4_outputs(9390) <= not b;
    layer4_outputs(9391) <= b;
    layer4_outputs(9392) <= a and not b;
    layer4_outputs(9393) <= not b or a;
    layer4_outputs(9394) <= b;
    layer4_outputs(9395) <= a or b;
    layer4_outputs(9396) <= b;
    layer4_outputs(9397) <= a;
    layer4_outputs(9398) <= '1';
    layer4_outputs(9399) <= not a;
    layer4_outputs(9400) <= not a;
    layer4_outputs(9401) <= b;
    layer4_outputs(9402) <= a or b;
    layer4_outputs(9403) <= not (a and b);
    layer4_outputs(9404) <= not (a and b);
    layer4_outputs(9405) <= a;
    layer4_outputs(9406) <= not (a or b);
    layer4_outputs(9407) <= b and not a;
    layer4_outputs(9408) <= not a;
    layer4_outputs(9409) <= not a;
    layer4_outputs(9410) <= not (a and b);
    layer4_outputs(9411) <= a xor b;
    layer4_outputs(9412) <= a and b;
    layer4_outputs(9413) <= a;
    layer4_outputs(9414) <= a;
    layer4_outputs(9415) <= a;
    layer4_outputs(9416) <= not a or b;
    layer4_outputs(9417) <= not a;
    layer4_outputs(9418) <= b;
    layer4_outputs(9419) <= not (a or b);
    layer4_outputs(9420) <= not a or b;
    layer4_outputs(9421) <= not b;
    layer4_outputs(9422) <= a and not b;
    layer4_outputs(9423) <= not (a and b);
    layer4_outputs(9424) <= b;
    layer4_outputs(9425) <= not a;
    layer4_outputs(9426) <= not a;
    layer4_outputs(9427) <= b;
    layer4_outputs(9428) <= a xor b;
    layer4_outputs(9429) <= b and not a;
    layer4_outputs(9430) <= b;
    layer4_outputs(9431) <= not b;
    layer4_outputs(9432) <= not a;
    layer4_outputs(9433) <= a and b;
    layer4_outputs(9434) <= a or b;
    layer4_outputs(9435) <= b and not a;
    layer4_outputs(9436) <= a;
    layer4_outputs(9437) <= a and b;
    layer4_outputs(9438) <= not (a or b);
    layer4_outputs(9439) <= not b;
    layer4_outputs(9440) <= not (a xor b);
    layer4_outputs(9441) <= not b;
    layer4_outputs(9442) <= b;
    layer4_outputs(9443) <= not b;
    layer4_outputs(9444) <= not b;
    layer4_outputs(9445) <= b;
    layer4_outputs(9446) <= a;
    layer4_outputs(9447) <= a;
    layer4_outputs(9448) <= b;
    layer4_outputs(9449) <= not a or b;
    layer4_outputs(9450) <= a or b;
    layer4_outputs(9451) <= not a;
    layer4_outputs(9452) <= b;
    layer4_outputs(9453) <= a and b;
    layer4_outputs(9454) <= a and b;
    layer4_outputs(9455) <= not b;
    layer4_outputs(9456) <= not (a and b);
    layer4_outputs(9457) <= not b;
    layer4_outputs(9458) <= '1';
    layer4_outputs(9459) <= a and not b;
    layer4_outputs(9460) <= a or b;
    layer4_outputs(9461) <= a xor b;
    layer4_outputs(9462) <= not a;
    layer4_outputs(9463) <= not b;
    layer4_outputs(9464) <= not a or b;
    layer4_outputs(9465) <= not a or b;
    layer4_outputs(9466) <= not b;
    layer4_outputs(9467) <= not b;
    layer4_outputs(9468) <= not a;
    layer4_outputs(9469) <= not (a or b);
    layer4_outputs(9470) <= a;
    layer4_outputs(9471) <= not b or a;
    layer4_outputs(9472) <= not a or b;
    layer4_outputs(9473) <= '1';
    layer4_outputs(9474) <= not (a and b);
    layer4_outputs(9475) <= a;
    layer4_outputs(9476) <= not (a xor b);
    layer4_outputs(9477) <= not a or b;
    layer4_outputs(9478) <= not a;
    layer4_outputs(9479) <= b and not a;
    layer4_outputs(9480) <= b;
    layer4_outputs(9481) <= not a;
    layer4_outputs(9482) <= not b;
    layer4_outputs(9483) <= not a or b;
    layer4_outputs(9484) <= b;
    layer4_outputs(9485) <= not b;
    layer4_outputs(9486) <= a xor b;
    layer4_outputs(9487) <= a xor b;
    layer4_outputs(9488) <= a xor b;
    layer4_outputs(9489) <= b and not a;
    layer4_outputs(9490) <= not b;
    layer4_outputs(9491) <= not b;
    layer4_outputs(9492) <= not a;
    layer4_outputs(9493) <= b and not a;
    layer4_outputs(9494) <= not b;
    layer4_outputs(9495) <= a or b;
    layer4_outputs(9496) <= not a or b;
    layer4_outputs(9497) <= not (a xor b);
    layer4_outputs(9498) <= not (a and b);
    layer4_outputs(9499) <= a or b;
    layer4_outputs(9500) <= not a or b;
    layer4_outputs(9501) <= b;
    layer4_outputs(9502) <= not (a or b);
    layer4_outputs(9503) <= b;
    layer4_outputs(9504) <= not (a or b);
    layer4_outputs(9505) <= b;
    layer4_outputs(9506) <= b and not a;
    layer4_outputs(9507) <= a or b;
    layer4_outputs(9508) <= a;
    layer4_outputs(9509) <= not a;
    layer4_outputs(9510) <= not a or b;
    layer4_outputs(9511) <= not (a or b);
    layer4_outputs(9512) <= not b or a;
    layer4_outputs(9513) <= not (a xor b);
    layer4_outputs(9514) <= a and not b;
    layer4_outputs(9515) <= not a;
    layer4_outputs(9516) <= not (a xor b);
    layer4_outputs(9517) <= not b;
    layer4_outputs(9518) <= a or b;
    layer4_outputs(9519) <= a and not b;
    layer4_outputs(9520) <= '0';
    layer4_outputs(9521) <= '1';
    layer4_outputs(9522) <= not a or b;
    layer4_outputs(9523) <= '1';
    layer4_outputs(9524) <= b;
    layer4_outputs(9525) <= not b or a;
    layer4_outputs(9526) <= not a or b;
    layer4_outputs(9527) <= a and b;
    layer4_outputs(9528) <= b;
    layer4_outputs(9529) <= b;
    layer4_outputs(9530) <= b;
    layer4_outputs(9531) <= not a or b;
    layer4_outputs(9532) <= not (a or b);
    layer4_outputs(9533) <= b;
    layer4_outputs(9534) <= not (a xor b);
    layer4_outputs(9535) <= b;
    layer4_outputs(9536) <= not b or a;
    layer4_outputs(9537) <= not b;
    layer4_outputs(9538) <= not (a or b);
    layer4_outputs(9539) <= b;
    layer4_outputs(9540) <= b and not a;
    layer4_outputs(9541) <= a and b;
    layer4_outputs(9542) <= not a;
    layer4_outputs(9543) <= a and not b;
    layer4_outputs(9544) <= '1';
    layer4_outputs(9545) <= not b;
    layer4_outputs(9546) <= a and b;
    layer4_outputs(9547) <= b;
    layer4_outputs(9548) <= not (a and b);
    layer4_outputs(9549) <= a xor b;
    layer4_outputs(9550) <= not a;
    layer4_outputs(9551) <= not b;
    layer4_outputs(9552) <= not b or a;
    layer4_outputs(9553) <= not a;
    layer4_outputs(9554) <= a and not b;
    layer4_outputs(9555) <= a;
    layer4_outputs(9556) <= '1';
    layer4_outputs(9557) <= a xor b;
    layer4_outputs(9558) <= not (a xor b);
    layer4_outputs(9559) <= not b;
    layer4_outputs(9560) <= not (a and b);
    layer4_outputs(9561) <= a;
    layer4_outputs(9562) <= a xor b;
    layer4_outputs(9563) <= b;
    layer4_outputs(9564) <= not a;
    layer4_outputs(9565) <= a;
    layer4_outputs(9566) <= a and b;
    layer4_outputs(9567) <= not (a and b);
    layer4_outputs(9568) <= '1';
    layer4_outputs(9569) <= not a;
    layer4_outputs(9570) <= a and not b;
    layer4_outputs(9571) <= not b;
    layer4_outputs(9572) <= '1';
    layer4_outputs(9573) <= a;
    layer4_outputs(9574) <= a and not b;
    layer4_outputs(9575) <= a;
    layer4_outputs(9576) <= a or b;
    layer4_outputs(9577) <= a xor b;
    layer4_outputs(9578) <= b and not a;
    layer4_outputs(9579) <= not (a or b);
    layer4_outputs(9580) <= not (a or b);
    layer4_outputs(9581) <= not a;
    layer4_outputs(9582) <= not a;
    layer4_outputs(9583) <= a and b;
    layer4_outputs(9584) <= not a;
    layer4_outputs(9585) <= not b;
    layer4_outputs(9586) <= a or b;
    layer4_outputs(9587) <= not a or b;
    layer4_outputs(9588) <= not a;
    layer4_outputs(9589) <= not a or b;
    layer4_outputs(9590) <= a;
    layer4_outputs(9591) <= b;
    layer4_outputs(9592) <= not b;
    layer4_outputs(9593) <= '0';
    layer4_outputs(9594) <= not a;
    layer4_outputs(9595) <= not b or a;
    layer4_outputs(9596) <= a xor b;
    layer4_outputs(9597) <= a;
    layer4_outputs(9598) <= not b or a;
    layer4_outputs(9599) <= b and not a;
    layer4_outputs(9600) <= '0';
    layer4_outputs(9601) <= not b;
    layer4_outputs(9602) <= not b;
    layer4_outputs(9603) <= not b;
    layer4_outputs(9604) <= a and b;
    layer4_outputs(9605) <= b and not a;
    layer4_outputs(9606) <= '1';
    layer4_outputs(9607) <= a;
    layer4_outputs(9608) <= a and b;
    layer4_outputs(9609) <= not b or a;
    layer4_outputs(9610) <= '0';
    layer4_outputs(9611) <= not (a xor b);
    layer4_outputs(9612) <= not (a xor b);
    layer4_outputs(9613) <= not a;
    layer4_outputs(9614) <= a and not b;
    layer4_outputs(9615) <= b and not a;
    layer4_outputs(9616) <= not (a or b);
    layer4_outputs(9617) <= b and not a;
    layer4_outputs(9618) <= not (a or b);
    layer4_outputs(9619) <= not (a or b);
    layer4_outputs(9620) <= not (a xor b);
    layer4_outputs(9621) <= a or b;
    layer4_outputs(9622) <= not a or b;
    layer4_outputs(9623) <= a xor b;
    layer4_outputs(9624) <= not a;
    layer4_outputs(9625) <= b;
    layer4_outputs(9626) <= not b;
    layer4_outputs(9627) <= a and b;
    layer4_outputs(9628) <= not a;
    layer4_outputs(9629) <= a;
    layer4_outputs(9630) <= not (a or b);
    layer4_outputs(9631) <= not a;
    layer4_outputs(9632) <= a;
    layer4_outputs(9633) <= not a;
    layer4_outputs(9634) <= not b;
    layer4_outputs(9635) <= not (a or b);
    layer4_outputs(9636) <= '1';
    layer4_outputs(9637) <= not b;
    layer4_outputs(9638) <= a;
    layer4_outputs(9639) <= not b;
    layer4_outputs(9640) <= not b;
    layer4_outputs(9641) <= not (a and b);
    layer4_outputs(9642) <= '0';
    layer4_outputs(9643) <= not b;
    layer4_outputs(9644) <= '1';
    layer4_outputs(9645) <= '1';
    layer4_outputs(9646) <= a or b;
    layer4_outputs(9647) <= not a or b;
    layer4_outputs(9648) <= a and b;
    layer4_outputs(9649) <= a xor b;
    layer4_outputs(9650) <= not (a and b);
    layer4_outputs(9651) <= not (a or b);
    layer4_outputs(9652) <= not b;
    layer4_outputs(9653) <= b;
    layer4_outputs(9654) <= not b;
    layer4_outputs(9655) <= a or b;
    layer4_outputs(9656) <= '1';
    layer4_outputs(9657) <= not a;
    layer4_outputs(9658) <= a;
    layer4_outputs(9659) <= not (a xor b);
    layer4_outputs(9660) <= not a or b;
    layer4_outputs(9661) <= '0';
    layer4_outputs(9662) <= a and not b;
    layer4_outputs(9663) <= b;
    layer4_outputs(9664) <= not b;
    layer4_outputs(9665) <= not a or b;
    layer4_outputs(9666) <= b and not a;
    layer4_outputs(9667) <= '0';
    layer4_outputs(9668) <= not (a xor b);
    layer4_outputs(9669) <= a xor b;
    layer4_outputs(9670) <= b and not a;
    layer4_outputs(9671) <= not (a and b);
    layer4_outputs(9672) <= b;
    layer4_outputs(9673) <= not (a or b);
    layer4_outputs(9674) <= b;
    layer4_outputs(9675) <= b and not a;
    layer4_outputs(9676) <= not a;
    layer4_outputs(9677) <= not b;
    layer4_outputs(9678) <= a or b;
    layer4_outputs(9679) <= b;
    layer4_outputs(9680) <= not a;
    layer4_outputs(9681) <= b;
    layer4_outputs(9682) <= not (a xor b);
    layer4_outputs(9683) <= a and b;
    layer4_outputs(9684) <= b;
    layer4_outputs(9685) <= a and not b;
    layer4_outputs(9686) <= b;
    layer4_outputs(9687) <= not (a or b);
    layer4_outputs(9688) <= not a or b;
    layer4_outputs(9689) <= not b or a;
    layer4_outputs(9690) <= b;
    layer4_outputs(9691) <= not b or a;
    layer4_outputs(9692) <= b;
    layer4_outputs(9693) <= a or b;
    layer4_outputs(9694) <= a and not b;
    layer4_outputs(9695) <= b and not a;
    layer4_outputs(9696) <= not (a or b);
    layer4_outputs(9697) <= not a;
    layer4_outputs(9698) <= not b;
    layer4_outputs(9699) <= a or b;
    layer4_outputs(9700) <= a and b;
    layer4_outputs(9701) <= a;
    layer4_outputs(9702) <= a and b;
    layer4_outputs(9703) <= b and not a;
    layer4_outputs(9704) <= '0';
    layer4_outputs(9705) <= a xor b;
    layer4_outputs(9706) <= a xor b;
    layer4_outputs(9707) <= '0';
    layer4_outputs(9708) <= not (a xor b);
    layer4_outputs(9709) <= a and not b;
    layer4_outputs(9710) <= a;
    layer4_outputs(9711) <= b;
    layer4_outputs(9712) <= a;
    layer4_outputs(9713) <= a;
    layer4_outputs(9714) <= a xor b;
    layer4_outputs(9715) <= '1';
    layer4_outputs(9716) <= b and not a;
    layer4_outputs(9717) <= '1';
    layer4_outputs(9718) <= not (a or b);
    layer4_outputs(9719) <= not b;
    layer4_outputs(9720) <= b;
    layer4_outputs(9721) <= not b;
    layer4_outputs(9722) <= b;
    layer4_outputs(9723) <= b and not a;
    layer4_outputs(9724) <= b;
    layer4_outputs(9725) <= b;
    layer4_outputs(9726) <= not (a or b);
    layer4_outputs(9727) <= a xor b;
    layer4_outputs(9728) <= not b or a;
    layer4_outputs(9729) <= not b or a;
    layer4_outputs(9730) <= '0';
    layer4_outputs(9731) <= a and not b;
    layer4_outputs(9732) <= not a or b;
    layer4_outputs(9733) <= a xor b;
    layer4_outputs(9734) <= not (a and b);
    layer4_outputs(9735) <= not (a xor b);
    layer4_outputs(9736) <= not b;
    layer4_outputs(9737) <= b and not a;
    layer4_outputs(9738) <= a and not b;
    layer4_outputs(9739) <= not (a and b);
    layer4_outputs(9740) <= a and not b;
    layer4_outputs(9741) <= a;
    layer4_outputs(9742) <= a and not b;
    layer4_outputs(9743) <= not b;
    layer4_outputs(9744) <= b;
    layer4_outputs(9745) <= b and not a;
    layer4_outputs(9746) <= a;
    layer4_outputs(9747) <= b and not a;
    layer4_outputs(9748) <= not (a or b);
    layer4_outputs(9749) <= a;
    layer4_outputs(9750) <= not a;
    layer4_outputs(9751) <= b;
    layer4_outputs(9752) <= not b;
    layer4_outputs(9753) <= b;
    layer4_outputs(9754) <= a or b;
    layer4_outputs(9755) <= not (a xor b);
    layer4_outputs(9756) <= a and b;
    layer4_outputs(9757) <= a;
    layer4_outputs(9758) <= not (a and b);
    layer4_outputs(9759) <= a xor b;
    layer4_outputs(9760) <= not b;
    layer4_outputs(9761) <= not (a xor b);
    layer4_outputs(9762) <= a and b;
    layer4_outputs(9763) <= b;
    layer4_outputs(9764) <= a or b;
    layer4_outputs(9765) <= a;
    layer4_outputs(9766) <= b and not a;
    layer4_outputs(9767) <= not (a xor b);
    layer4_outputs(9768) <= a and not b;
    layer4_outputs(9769) <= a and not b;
    layer4_outputs(9770) <= not b or a;
    layer4_outputs(9771) <= not (a and b);
    layer4_outputs(9772) <= not a or b;
    layer4_outputs(9773) <= a and not b;
    layer4_outputs(9774) <= not (a and b);
    layer4_outputs(9775) <= a and not b;
    layer4_outputs(9776) <= '1';
    layer4_outputs(9777) <= not (a and b);
    layer4_outputs(9778) <= b and not a;
    layer4_outputs(9779) <= b;
    layer4_outputs(9780) <= not a or b;
    layer4_outputs(9781) <= not a;
    layer4_outputs(9782) <= a;
    layer4_outputs(9783) <= not a or b;
    layer4_outputs(9784) <= not a;
    layer4_outputs(9785) <= b and not a;
    layer4_outputs(9786) <= a;
    layer4_outputs(9787) <= not (a or b);
    layer4_outputs(9788) <= not b;
    layer4_outputs(9789) <= not (a and b);
    layer4_outputs(9790) <= a or b;
    layer4_outputs(9791) <= not a;
    layer4_outputs(9792) <= not b or a;
    layer4_outputs(9793) <= a;
    layer4_outputs(9794) <= b and not a;
    layer4_outputs(9795) <= a or b;
    layer4_outputs(9796) <= b;
    layer4_outputs(9797) <= b and not a;
    layer4_outputs(9798) <= not a or b;
    layer4_outputs(9799) <= not a;
    layer4_outputs(9800) <= not a;
    layer4_outputs(9801) <= b;
    layer4_outputs(9802) <= not a or b;
    layer4_outputs(9803) <= not b or a;
    layer4_outputs(9804) <= not a;
    layer4_outputs(9805) <= not b;
    layer4_outputs(9806) <= b;
    layer4_outputs(9807) <= a;
    layer4_outputs(9808) <= not (a and b);
    layer4_outputs(9809) <= b;
    layer4_outputs(9810) <= a and not b;
    layer4_outputs(9811) <= a;
    layer4_outputs(9812) <= b and not a;
    layer4_outputs(9813) <= not (a or b);
    layer4_outputs(9814) <= not b;
    layer4_outputs(9815) <= a and b;
    layer4_outputs(9816) <= not b or a;
    layer4_outputs(9817) <= a or b;
    layer4_outputs(9818) <= a;
    layer4_outputs(9819) <= a;
    layer4_outputs(9820) <= not a;
    layer4_outputs(9821) <= not a or b;
    layer4_outputs(9822) <= not (a and b);
    layer4_outputs(9823) <= not b;
    layer4_outputs(9824) <= a and b;
    layer4_outputs(9825) <= '1';
    layer4_outputs(9826) <= a xor b;
    layer4_outputs(9827) <= not a;
    layer4_outputs(9828) <= not b or a;
    layer4_outputs(9829) <= a or b;
    layer4_outputs(9830) <= b and not a;
    layer4_outputs(9831) <= not b;
    layer4_outputs(9832) <= b and not a;
    layer4_outputs(9833) <= not b or a;
    layer4_outputs(9834) <= '1';
    layer4_outputs(9835) <= a;
    layer4_outputs(9836) <= not b;
    layer4_outputs(9837) <= a and not b;
    layer4_outputs(9838) <= b;
    layer4_outputs(9839) <= not a;
    layer4_outputs(9840) <= b and not a;
    layer4_outputs(9841) <= a or b;
    layer4_outputs(9842) <= not a;
    layer4_outputs(9843) <= a xor b;
    layer4_outputs(9844) <= a;
    layer4_outputs(9845) <= not (a xor b);
    layer4_outputs(9846) <= not a;
    layer4_outputs(9847) <= b and not a;
    layer4_outputs(9848) <= not b;
    layer4_outputs(9849) <= not a;
    layer4_outputs(9850) <= a;
    layer4_outputs(9851) <= a;
    layer4_outputs(9852) <= not a;
    layer4_outputs(9853) <= not a;
    layer4_outputs(9854) <= not b;
    layer4_outputs(9855) <= not a;
    layer4_outputs(9856) <= not b or a;
    layer4_outputs(9857) <= b;
    layer4_outputs(9858) <= a and not b;
    layer4_outputs(9859) <= b and not a;
    layer4_outputs(9860) <= a or b;
    layer4_outputs(9861) <= not a;
    layer4_outputs(9862) <= a and not b;
    layer4_outputs(9863) <= b;
    layer4_outputs(9864) <= not b or a;
    layer4_outputs(9865) <= not b;
    layer4_outputs(9866) <= a and not b;
    layer4_outputs(9867) <= not b;
    layer4_outputs(9868) <= not b;
    layer4_outputs(9869) <= not b;
    layer4_outputs(9870) <= b;
    layer4_outputs(9871) <= not (a and b);
    layer4_outputs(9872) <= not b;
    layer4_outputs(9873) <= not a;
    layer4_outputs(9874) <= not (a or b);
    layer4_outputs(9875) <= b and not a;
    layer4_outputs(9876) <= a and not b;
    layer4_outputs(9877) <= '1';
    layer4_outputs(9878) <= not b;
    layer4_outputs(9879) <= b and not a;
    layer4_outputs(9880) <= not (a or b);
    layer4_outputs(9881) <= b and not a;
    layer4_outputs(9882) <= not b or a;
    layer4_outputs(9883) <= a;
    layer4_outputs(9884) <= not b or a;
    layer4_outputs(9885) <= not (a and b);
    layer4_outputs(9886) <= a or b;
    layer4_outputs(9887) <= not (a xor b);
    layer4_outputs(9888) <= not b;
    layer4_outputs(9889) <= a and b;
    layer4_outputs(9890) <= not a or b;
    layer4_outputs(9891) <= a xor b;
    layer4_outputs(9892) <= b and not a;
    layer4_outputs(9893) <= a or b;
    layer4_outputs(9894) <= b;
    layer4_outputs(9895) <= not b or a;
    layer4_outputs(9896) <= not (a and b);
    layer4_outputs(9897) <= a xor b;
    layer4_outputs(9898) <= not a;
    layer4_outputs(9899) <= a and not b;
    layer4_outputs(9900) <= a;
    layer4_outputs(9901) <= a;
    layer4_outputs(9902) <= not (a or b);
    layer4_outputs(9903) <= not (a and b);
    layer4_outputs(9904) <= '0';
    layer4_outputs(9905) <= a;
    layer4_outputs(9906) <= a xor b;
    layer4_outputs(9907) <= b;
    layer4_outputs(9908) <= not (a and b);
    layer4_outputs(9909) <= a and b;
    layer4_outputs(9910) <= not b;
    layer4_outputs(9911) <= a;
    layer4_outputs(9912) <= a or b;
    layer4_outputs(9913) <= not a;
    layer4_outputs(9914) <= not (a xor b);
    layer4_outputs(9915) <= not (a and b);
    layer4_outputs(9916) <= b and not a;
    layer4_outputs(9917) <= a and not b;
    layer4_outputs(9918) <= not (a xor b);
    layer4_outputs(9919) <= a and not b;
    layer4_outputs(9920) <= not b;
    layer4_outputs(9921) <= a and b;
    layer4_outputs(9922) <= b;
    layer4_outputs(9923) <= a and b;
    layer4_outputs(9924) <= not (a and b);
    layer4_outputs(9925) <= not b or a;
    layer4_outputs(9926) <= a;
    layer4_outputs(9927) <= b and not a;
    layer4_outputs(9928) <= b and not a;
    layer4_outputs(9929) <= a or b;
    layer4_outputs(9930) <= b and not a;
    layer4_outputs(9931) <= b;
    layer4_outputs(9932) <= a and b;
    layer4_outputs(9933) <= b;
    layer4_outputs(9934) <= not (a and b);
    layer4_outputs(9935) <= a or b;
    layer4_outputs(9936) <= a and not b;
    layer4_outputs(9937) <= a and not b;
    layer4_outputs(9938) <= b and not a;
    layer4_outputs(9939) <= b and not a;
    layer4_outputs(9940) <= a and b;
    layer4_outputs(9941) <= a;
    layer4_outputs(9942) <= not (a xor b);
    layer4_outputs(9943) <= a xor b;
    layer4_outputs(9944) <= b and not a;
    layer4_outputs(9945) <= not b;
    layer4_outputs(9946) <= a or b;
    layer4_outputs(9947) <= not a or b;
    layer4_outputs(9948) <= a and b;
    layer4_outputs(9949) <= b;
    layer4_outputs(9950) <= not b;
    layer4_outputs(9951) <= a or b;
    layer4_outputs(9952) <= not b;
    layer4_outputs(9953) <= a or b;
    layer4_outputs(9954) <= not b;
    layer4_outputs(9955) <= b and not a;
    layer4_outputs(9956) <= a;
    layer4_outputs(9957) <= b and not a;
    layer4_outputs(9958) <= '1';
    layer4_outputs(9959) <= a;
    layer4_outputs(9960) <= not (a or b);
    layer4_outputs(9961) <= a or b;
    layer4_outputs(9962) <= a and not b;
    layer4_outputs(9963) <= a xor b;
    layer4_outputs(9964) <= not a;
    layer4_outputs(9965) <= a and b;
    layer4_outputs(9966) <= not b;
    layer4_outputs(9967) <= not b;
    layer4_outputs(9968) <= '0';
    layer4_outputs(9969) <= a and b;
    layer4_outputs(9970) <= not a;
    layer4_outputs(9971) <= a;
    layer4_outputs(9972) <= not b;
    layer4_outputs(9973) <= not a;
    layer4_outputs(9974) <= not (a or b);
    layer4_outputs(9975) <= a;
    layer4_outputs(9976) <= a xor b;
    layer4_outputs(9977) <= a;
    layer4_outputs(9978) <= not a;
    layer4_outputs(9979) <= '0';
    layer4_outputs(9980) <= a and b;
    layer4_outputs(9981) <= not b;
    layer4_outputs(9982) <= '1';
    layer4_outputs(9983) <= a and not b;
    layer4_outputs(9984) <= not b;
    layer4_outputs(9985) <= b;
    layer4_outputs(9986) <= not b;
    layer4_outputs(9987) <= not (a or b);
    layer4_outputs(9988) <= not a or b;
    layer4_outputs(9989) <= not (a and b);
    layer4_outputs(9990) <= not b or a;
    layer4_outputs(9991) <= a;
    layer4_outputs(9992) <= b;
    layer4_outputs(9993) <= not b or a;
    layer4_outputs(9994) <= a;
    layer4_outputs(9995) <= not a or b;
    layer4_outputs(9996) <= not b;
    layer4_outputs(9997) <= not (a and b);
    layer4_outputs(9998) <= not b;
    layer4_outputs(9999) <= a;
    layer4_outputs(10000) <= a xor b;
    layer4_outputs(10001) <= not (a and b);
    layer4_outputs(10002) <= a;
    layer4_outputs(10003) <= not a or b;
    layer4_outputs(10004) <= a and b;
    layer4_outputs(10005) <= not (a and b);
    layer4_outputs(10006) <= a xor b;
    layer4_outputs(10007) <= not a;
    layer4_outputs(10008) <= not (a xor b);
    layer4_outputs(10009) <= not a;
    layer4_outputs(10010) <= '0';
    layer4_outputs(10011) <= not (a and b);
    layer4_outputs(10012) <= b and not a;
    layer4_outputs(10013) <= not (a and b);
    layer4_outputs(10014) <= not a;
    layer4_outputs(10015) <= a or b;
    layer4_outputs(10016) <= not b;
    layer4_outputs(10017) <= not (a xor b);
    layer4_outputs(10018) <= not b;
    layer4_outputs(10019) <= not (a and b);
    layer4_outputs(10020) <= b;
    layer4_outputs(10021) <= not (a xor b);
    layer4_outputs(10022) <= a and b;
    layer4_outputs(10023) <= not a or b;
    layer4_outputs(10024) <= a and not b;
    layer4_outputs(10025) <= a xor b;
    layer4_outputs(10026) <= not (a and b);
    layer4_outputs(10027) <= not a or b;
    layer4_outputs(10028) <= a and b;
    layer4_outputs(10029) <= a and b;
    layer4_outputs(10030) <= not a;
    layer4_outputs(10031) <= a or b;
    layer4_outputs(10032) <= a;
    layer4_outputs(10033) <= not b;
    layer4_outputs(10034) <= not b;
    layer4_outputs(10035) <= a and b;
    layer4_outputs(10036) <= a;
    layer4_outputs(10037) <= not a;
    layer4_outputs(10038) <= a or b;
    layer4_outputs(10039) <= '1';
    layer4_outputs(10040) <= a and not b;
    layer4_outputs(10041) <= not (a xor b);
    layer4_outputs(10042) <= not a or b;
    layer4_outputs(10043) <= not a;
    layer4_outputs(10044) <= a or b;
    layer4_outputs(10045) <= a;
    layer4_outputs(10046) <= not a;
    layer4_outputs(10047) <= a or b;
    layer4_outputs(10048) <= a and b;
    layer4_outputs(10049) <= not b or a;
    layer4_outputs(10050) <= a xor b;
    layer4_outputs(10051) <= not b;
    layer4_outputs(10052) <= not a;
    layer4_outputs(10053) <= a xor b;
    layer4_outputs(10054) <= a;
    layer4_outputs(10055) <= not b;
    layer4_outputs(10056) <= not b;
    layer4_outputs(10057) <= '0';
    layer4_outputs(10058) <= a and b;
    layer4_outputs(10059) <= not (a or b);
    layer4_outputs(10060) <= a;
    layer4_outputs(10061) <= b;
    layer4_outputs(10062) <= a and b;
    layer4_outputs(10063) <= a or b;
    layer4_outputs(10064) <= not b or a;
    layer4_outputs(10065) <= not a or b;
    layer4_outputs(10066) <= not (a and b);
    layer4_outputs(10067) <= not b or a;
    layer4_outputs(10068) <= not a or b;
    layer4_outputs(10069) <= not a;
    layer4_outputs(10070) <= a xor b;
    layer4_outputs(10071) <= not a or b;
    layer4_outputs(10072) <= not a or b;
    layer4_outputs(10073) <= a or b;
    layer4_outputs(10074) <= a or b;
    layer4_outputs(10075) <= b and not a;
    layer4_outputs(10076) <= a or b;
    layer4_outputs(10077) <= b and not a;
    layer4_outputs(10078) <= not b;
    layer4_outputs(10079) <= a and b;
    layer4_outputs(10080) <= not a;
    layer4_outputs(10081) <= a and b;
    layer4_outputs(10082) <= a or b;
    layer4_outputs(10083) <= b;
    layer4_outputs(10084) <= a and b;
    layer4_outputs(10085) <= b and not a;
    layer4_outputs(10086) <= not (a xor b);
    layer4_outputs(10087) <= not a;
    layer4_outputs(10088) <= not a;
    layer4_outputs(10089) <= a and not b;
    layer4_outputs(10090) <= not b or a;
    layer4_outputs(10091) <= b;
    layer4_outputs(10092) <= not a;
    layer4_outputs(10093) <= not a or b;
    layer4_outputs(10094) <= a or b;
    layer4_outputs(10095) <= not b or a;
    layer4_outputs(10096) <= a xor b;
    layer4_outputs(10097) <= a xor b;
    layer4_outputs(10098) <= not b or a;
    layer4_outputs(10099) <= not (a and b);
    layer4_outputs(10100) <= '1';
    layer4_outputs(10101) <= not a;
    layer4_outputs(10102) <= a;
    layer4_outputs(10103) <= a or b;
    layer4_outputs(10104) <= a;
    layer4_outputs(10105) <= a or b;
    layer4_outputs(10106) <= a or b;
    layer4_outputs(10107) <= not (a or b);
    layer4_outputs(10108) <= not a or b;
    layer4_outputs(10109) <= a;
    layer4_outputs(10110) <= not b;
    layer4_outputs(10111) <= not b or a;
    layer4_outputs(10112) <= not b or a;
    layer4_outputs(10113) <= '0';
    layer4_outputs(10114) <= a or b;
    layer4_outputs(10115) <= '1';
    layer4_outputs(10116) <= a and not b;
    layer4_outputs(10117) <= not (a or b);
    layer4_outputs(10118) <= '0';
    layer4_outputs(10119) <= not b;
    layer4_outputs(10120) <= a;
    layer4_outputs(10121) <= not (a xor b);
    layer4_outputs(10122) <= b;
    layer4_outputs(10123) <= a;
    layer4_outputs(10124) <= not a or b;
    layer4_outputs(10125) <= not b or a;
    layer4_outputs(10126) <= not b or a;
    layer4_outputs(10127) <= a and b;
    layer4_outputs(10128) <= not b;
    layer4_outputs(10129) <= not (a or b);
    layer4_outputs(10130) <= a;
    layer4_outputs(10131) <= not (a or b);
    layer4_outputs(10132) <= a xor b;
    layer4_outputs(10133) <= a;
    layer4_outputs(10134) <= not (a or b);
    layer4_outputs(10135) <= not (a or b);
    layer4_outputs(10136) <= b;
    layer4_outputs(10137) <= a;
    layer4_outputs(10138) <= not a or b;
    layer4_outputs(10139) <= not a or b;
    layer4_outputs(10140) <= not a or b;
    layer4_outputs(10141) <= a and b;
    layer4_outputs(10142) <= not (a xor b);
    layer4_outputs(10143) <= not a;
    layer4_outputs(10144) <= not (a or b);
    layer4_outputs(10145) <= not b;
    layer4_outputs(10146) <= b;
    layer4_outputs(10147) <= not a or b;
    layer4_outputs(10148) <= not a;
    layer4_outputs(10149) <= not b or a;
    layer4_outputs(10150) <= b;
    layer4_outputs(10151) <= not b or a;
    layer4_outputs(10152) <= not a or b;
    layer4_outputs(10153) <= b;
    layer4_outputs(10154) <= not (a or b);
    layer4_outputs(10155) <= a and b;
    layer4_outputs(10156) <= not b;
    layer4_outputs(10157) <= a and not b;
    layer4_outputs(10158) <= b;
    layer4_outputs(10159) <= not a;
    layer4_outputs(10160) <= not b;
    layer4_outputs(10161) <= not b;
    layer4_outputs(10162) <= a and not b;
    layer4_outputs(10163) <= '1';
    layer4_outputs(10164) <= not a;
    layer4_outputs(10165) <= not (a or b);
    layer4_outputs(10166) <= a xor b;
    layer4_outputs(10167) <= a and not b;
    layer4_outputs(10168) <= a or b;
    layer4_outputs(10169) <= b and not a;
    layer4_outputs(10170) <= b and not a;
    layer4_outputs(10171) <= not (a or b);
    layer4_outputs(10172) <= not a;
    layer4_outputs(10173) <= not a or b;
    layer4_outputs(10174) <= a or b;
    layer4_outputs(10175) <= a xor b;
    layer4_outputs(10176) <= not a;
    layer4_outputs(10177) <= not (a or b);
    layer4_outputs(10178) <= not a;
    layer4_outputs(10179) <= not a;
    layer4_outputs(10180) <= b;
    layer4_outputs(10181) <= not b;
    layer4_outputs(10182) <= a and not b;
    layer4_outputs(10183) <= not (a and b);
    layer4_outputs(10184) <= not a or b;
    layer4_outputs(10185) <= b;
    layer4_outputs(10186) <= not a or b;
    layer4_outputs(10187) <= a and b;
    layer4_outputs(10188) <= a or b;
    layer4_outputs(10189) <= a and b;
    layer4_outputs(10190) <= b;
    layer4_outputs(10191) <= a;
    layer4_outputs(10192) <= a;
    layer4_outputs(10193) <= not b or a;
    layer4_outputs(10194) <= a xor b;
    layer4_outputs(10195) <= b and not a;
    layer4_outputs(10196) <= not a;
    layer4_outputs(10197) <= not b;
    layer4_outputs(10198) <= a;
    layer4_outputs(10199) <= b;
    layer4_outputs(10200) <= not (a or b);
    layer4_outputs(10201) <= '1';
    layer4_outputs(10202) <= not a;
    layer4_outputs(10203) <= not b;
    layer4_outputs(10204) <= a and not b;
    layer4_outputs(10205) <= a;
    layer4_outputs(10206) <= not b or a;
    layer4_outputs(10207) <= not b;
    layer4_outputs(10208) <= not b;
    layer4_outputs(10209) <= not a or b;
    layer4_outputs(10210) <= b;
    layer4_outputs(10211) <= '0';
    layer4_outputs(10212) <= not a;
    layer4_outputs(10213) <= not b;
    layer4_outputs(10214) <= not b;
    layer4_outputs(10215) <= a;
    layer4_outputs(10216) <= not a;
    layer4_outputs(10217) <= a xor b;
    layer4_outputs(10218) <= not (a xor b);
    layer4_outputs(10219) <= not (a or b);
    layer4_outputs(10220) <= b and not a;
    layer4_outputs(10221) <= a and b;
    layer4_outputs(10222) <= not a;
    layer4_outputs(10223) <= '0';
    layer4_outputs(10224) <= not (a xor b);
    layer4_outputs(10225) <= a and b;
    layer4_outputs(10226) <= b;
    layer4_outputs(10227) <= b and not a;
    layer4_outputs(10228) <= not b or a;
    layer4_outputs(10229) <= not (a and b);
    layer4_outputs(10230) <= not (a and b);
    layer4_outputs(10231) <= not a or b;
    layer4_outputs(10232) <= b and not a;
    layer4_outputs(10233) <= a and not b;
    layer4_outputs(10234) <= not (a or b);
    layer4_outputs(10235) <= a or b;
    layer4_outputs(10236) <= not b;
    layer4_outputs(10237) <= b;
    layer4_outputs(10238) <= not b;
    layer4_outputs(10239) <= a and not b;
    layer5_outputs(0) <= not a;
    layer5_outputs(1) <= not b;
    layer5_outputs(2) <= not (a or b);
    layer5_outputs(3) <= a and not b;
    layer5_outputs(4) <= b and not a;
    layer5_outputs(5) <= not b;
    layer5_outputs(6) <= b;
    layer5_outputs(7) <= a xor b;
    layer5_outputs(8) <= not b;
    layer5_outputs(9) <= not (a xor b);
    layer5_outputs(10) <= a;
    layer5_outputs(11) <= a;
    layer5_outputs(12) <= not a;
    layer5_outputs(13) <= not b;
    layer5_outputs(14) <= a and b;
    layer5_outputs(15) <= not a;
    layer5_outputs(16) <= a;
    layer5_outputs(17) <= a;
    layer5_outputs(18) <= b;
    layer5_outputs(19) <= b;
    layer5_outputs(20) <= b and not a;
    layer5_outputs(21) <= a and b;
    layer5_outputs(22) <= a or b;
    layer5_outputs(23) <= not a or b;
    layer5_outputs(24) <= not b;
    layer5_outputs(25) <= not a;
    layer5_outputs(26) <= a xor b;
    layer5_outputs(27) <= not a;
    layer5_outputs(28) <= not b;
    layer5_outputs(29) <= not b;
    layer5_outputs(30) <= b and not a;
    layer5_outputs(31) <= not a;
    layer5_outputs(32) <= '0';
    layer5_outputs(33) <= not a or b;
    layer5_outputs(34) <= a or b;
    layer5_outputs(35) <= b;
    layer5_outputs(36) <= a xor b;
    layer5_outputs(37) <= not b;
    layer5_outputs(38) <= not b or a;
    layer5_outputs(39) <= not b;
    layer5_outputs(40) <= b and not a;
    layer5_outputs(41) <= b;
    layer5_outputs(42) <= b and not a;
    layer5_outputs(43) <= a and not b;
    layer5_outputs(44) <= a and b;
    layer5_outputs(45) <= a xor b;
    layer5_outputs(46) <= not (a xor b);
    layer5_outputs(47) <= not a or b;
    layer5_outputs(48) <= not b;
    layer5_outputs(49) <= not b;
    layer5_outputs(50) <= not a or b;
    layer5_outputs(51) <= a or b;
    layer5_outputs(52) <= a;
    layer5_outputs(53) <= b and not a;
    layer5_outputs(54) <= b and not a;
    layer5_outputs(55) <= b;
    layer5_outputs(56) <= not (a and b);
    layer5_outputs(57) <= a and not b;
    layer5_outputs(58) <= not a or b;
    layer5_outputs(59) <= not (a and b);
    layer5_outputs(60) <= not b;
    layer5_outputs(61) <= not a;
    layer5_outputs(62) <= not (a or b);
    layer5_outputs(63) <= not b or a;
    layer5_outputs(64) <= not (a or b);
    layer5_outputs(65) <= a xor b;
    layer5_outputs(66) <= not (a and b);
    layer5_outputs(67) <= '1';
    layer5_outputs(68) <= a xor b;
    layer5_outputs(69) <= not (a or b);
    layer5_outputs(70) <= not b;
    layer5_outputs(71) <= not (a or b);
    layer5_outputs(72) <= not a;
    layer5_outputs(73) <= not (a xor b);
    layer5_outputs(74) <= a;
    layer5_outputs(75) <= a xor b;
    layer5_outputs(76) <= not b;
    layer5_outputs(77) <= a and b;
    layer5_outputs(78) <= a;
    layer5_outputs(79) <= a xor b;
    layer5_outputs(80) <= b and not a;
    layer5_outputs(81) <= not a;
    layer5_outputs(82) <= a or b;
    layer5_outputs(83) <= a;
    layer5_outputs(84) <= not a or b;
    layer5_outputs(85) <= a or b;
    layer5_outputs(86) <= b;
    layer5_outputs(87) <= b and not a;
    layer5_outputs(88) <= not (a or b);
    layer5_outputs(89) <= not b;
    layer5_outputs(90) <= not b;
    layer5_outputs(91) <= not a;
    layer5_outputs(92) <= a or b;
    layer5_outputs(93) <= not a;
    layer5_outputs(94) <= a or b;
    layer5_outputs(95) <= not b;
    layer5_outputs(96) <= a and b;
    layer5_outputs(97) <= a xor b;
    layer5_outputs(98) <= not (a and b);
    layer5_outputs(99) <= a or b;
    layer5_outputs(100) <= not (a and b);
    layer5_outputs(101) <= a or b;
    layer5_outputs(102) <= a and b;
    layer5_outputs(103) <= a and b;
    layer5_outputs(104) <= not a or b;
    layer5_outputs(105) <= not b;
    layer5_outputs(106) <= not b;
    layer5_outputs(107) <= b and not a;
    layer5_outputs(108) <= not (a or b);
    layer5_outputs(109) <= a and not b;
    layer5_outputs(110) <= a;
    layer5_outputs(111) <= not b or a;
    layer5_outputs(112) <= not (a xor b);
    layer5_outputs(113) <= not b;
    layer5_outputs(114) <= b;
    layer5_outputs(115) <= a and not b;
    layer5_outputs(116) <= not b;
    layer5_outputs(117) <= b;
    layer5_outputs(118) <= b;
    layer5_outputs(119) <= not (a xor b);
    layer5_outputs(120) <= not a;
    layer5_outputs(121) <= not a;
    layer5_outputs(122) <= not b;
    layer5_outputs(123) <= a xor b;
    layer5_outputs(124) <= a and b;
    layer5_outputs(125) <= b and not a;
    layer5_outputs(126) <= not (a xor b);
    layer5_outputs(127) <= a and b;
    layer5_outputs(128) <= '1';
    layer5_outputs(129) <= not (a xor b);
    layer5_outputs(130) <= a;
    layer5_outputs(131) <= a;
    layer5_outputs(132) <= a xor b;
    layer5_outputs(133) <= not b;
    layer5_outputs(134) <= not a or b;
    layer5_outputs(135) <= b;
    layer5_outputs(136) <= not a or b;
    layer5_outputs(137) <= not a;
    layer5_outputs(138) <= not (a or b);
    layer5_outputs(139) <= not b;
    layer5_outputs(140) <= '1';
    layer5_outputs(141) <= not (a or b);
    layer5_outputs(142) <= not a;
    layer5_outputs(143) <= not b or a;
    layer5_outputs(144) <= not (a xor b);
    layer5_outputs(145) <= not a;
    layer5_outputs(146) <= not b;
    layer5_outputs(147) <= a;
    layer5_outputs(148) <= a and b;
    layer5_outputs(149) <= a xor b;
    layer5_outputs(150) <= a or b;
    layer5_outputs(151) <= not (a and b);
    layer5_outputs(152) <= not b or a;
    layer5_outputs(153) <= b and not a;
    layer5_outputs(154) <= a;
    layer5_outputs(155) <= not b;
    layer5_outputs(156) <= a and b;
    layer5_outputs(157) <= a and not b;
    layer5_outputs(158) <= a;
    layer5_outputs(159) <= b;
    layer5_outputs(160) <= b;
    layer5_outputs(161) <= not (a or b);
    layer5_outputs(162) <= b and not a;
    layer5_outputs(163) <= not (a and b);
    layer5_outputs(164) <= not a;
    layer5_outputs(165) <= not b or a;
    layer5_outputs(166) <= not a;
    layer5_outputs(167) <= not b or a;
    layer5_outputs(168) <= b;
    layer5_outputs(169) <= not b;
    layer5_outputs(170) <= not (a and b);
    layer5_outputs(171) <= '0';
    layer5_outputs(172) <= not a or b;
    layer5_outputs(173) <= a and not b;
    layer5_outputs(174) <= not a or b;
    layer5_outputs(175) <= b;
    layer5_outputs(176) <= not (a xor b);
    layer5_outputs(177) <= b;
    layer5_outputs(178) <= a and not b;
    layer5_outputs(179) <= a and not b;
    layer5_outputs(180) <= a and b;
    layer5_outputs(181) <= a;
    layer5_outputs(182) <= b;
    layer5_outputs(183) <= a;
    layer5_outputs(184) <= b;
    layer5_outputs(185) <= a or b;
    layer5_outputs(186) <= b;
    layer5_outputs(187) <= a and b;
    layer5_outputs(188) <= a and b;
    layer5_outputs(189) <= a and not b;
    layer5_outputs(190) <= not a;
    layer5_outputs(191) <= a;
    layer5_outputs(192) <= not (a xor b);
    layer5_outputs(193) <= not (a or b);
    layer5_outputs(194) <= a or b;
    layer5_outputs(195) <= a;
    layer5_outputs(196) <= not (a xor b);
    layer5_outputs(197) <= not b or a;
    layer5_outputs(198) <= b;
    layer5_outputs(199) <= not a;
    layer5_outputs(200) <= a;
    layer5_outputs(201) <= not a or b;
    layer5_outputs(202) <= not a;
    layer5_outputs(203) <= not a;
    layer5_outputs(204) <= not b;
    layer5_outputs(205) <= not b;
    layer5_outputs(206) <= not a or b;
    layer5_outputs(207) <= not (a xor b);
    layer5_outputs(208) <= not (a or b);
    layer5_outputs(209) <= a;
    layer5_outputs(210) <= b and not a;
    layer5_outputs(211) <= not a or b;
    layer5_outputs(212) <= a and b;
    layer5_outputs(213) <= not a;
    layer5_outputs(214) <= a;
    layer5_outputs(215) <= b and not a;
    layer5_outputs(216) <= not a;
    layer5_outputs(217) <= a and not b;
    layer5_outputs(218) <= '1';
    layer5_outputs(219) <= a and not b;
    layer5_outputs(220) <= not a;
    layer5_outputs(221) <= a;
    layer5_outputs(222) <= not a or b;
    layer5_outputs(223) <= b;
    layer5_outputs(224) <= not a;
    layer5_outputs(225) <= a xor b;
    layer5_outputs(226) <= not b;
    layer5_outputs(227) <= a and b;
    layer5_outputs(228) <= '0';
    layer5_outputs(229) <= not b;
    layer5_outputs(230) <= not (a or b);
    layer5_outputs(231) <= not b;
    layer5_outputs(232) <= '0';
    layer5_outputs(233) <= not b;
    layer5_outputs(234) <= not b;
    layer5_outputs(235) <= '0';
    layer5_outputs(236) <= a;
    layer5_outputs(237) <= a or b;
    layer5_outputs(238) <= b and not a;
    layer5_outputs(239) <= not a;
    layer5_outputs(240) <= a;
    layer5_outputs(241) <= a and b;
    layer5_outputs(242) <= b;
    layer5_outputs(243) <= b and not a;
    layer5_outputs(244) <= not b;
    layer5_outputs(245) <= not b or a;
    layer5_outputs(246) <= a or b;
    layer5_outputs(247) <= not a or b;
    layer5_outputs(248) <= b;
    layer5_outputs(249) <= not (a and b);
    layer5_outputs(250) <= not b;
    layer5_outputs(251) <= not b;
    layer5_outputs(252) <= not b or a;
    layer5_outputs(253) <= not (a xor b);
    layer5_outputs(254) <= a;
    layer5_outputs(255) <= not a or b;
    layer5_outputs(256) <= not (a xor b);
    layer5_outputs(257) <= not b;
    layer5_outputs(258) <= not (a xor b);
    layer5_outputs(259) <= not (a or b);
    layer5_outputs(260) <= not (a and b);
    layer5_outputs(261) <= a and not b;
    layer5_outputs(262) <= a or b;
    layer5_outputs(263) <= a;
    layer5_outputs(264) <= a;
    layer5_outputs(265) <= a and not b;
    layer5_outputs(266) <= b;
    layer5_outputs(267) <= a xor b;
    layer5_outputs(268) <= not (a xor b);
    layer5_outputs(269) <= b;
    layer5_outputs(270) <= not (a xor b);
    layer5_outputs(271) <= a or b;
    layer5_outputs(272) <= a;
    layer5_outputs(273) <= a xor b;
    layer5_outputs(274) <= a and b;
    layer5_outputs(275) <= a;
    layer5_outputs(276) <= b and not a;
    layer5_outputs(277) <= b and not a;
    layer5_outputs(278) <= a and b;
    layer5_outputs(279) <= b and not a;
    layer5_outputs(280) <= a xor b;
    layer5_outputs(281) <= not a;
    layer5_outputs(282) <= a and b;
    layer5_outputs(283) <= b and not a;
    layer5_outputs(284) <= not (a and b);
    layer5_outputs(285) <= not b or a;
    layer5_outputs(286) <= a or b;
    layer5_outputs(287) <= not b;
    layer5_outputs(288) <= b;
    layer5_outputs(289) <= not a;
    layer5_outputs(290) <= b;
    layer5_outputs(291) <= a;
    layer5_outputs(292) <= '1';
    layer5_outputs(293) <= a;
    layer5_outputs(294) <= not a or b;
    layer5_outputs(295) <= not b;
    layer5_outputs(296) <= a;
    layer5_outputs(297) <= not (a or b);
    layer5_outputs(298) <= b and not a;
    layer5_outputs(299) <= not b or a;
    layer5_outputs(300) <= b;
    layer5_outputs(301) <= not (a xor b);
    layer5_outputs(302) <= not (a xor b);
    layer5_outputs(303) <= a or b;
    layer5_outputs(304) <= a;
    layer5_outputs(305) <= not (a xor b);
    layer5_outputs(306) <= a;
    layer5_outputs(307) <= not a;
    layer5_outputs(308) <= not a or b;
    layer5_outputs(309) <= a;
    layer5_outputs(310) <= a and b;
    layer5_outputs(311) <= a xor b;
    layer5_outputs(312) <= not b or a;
    layer5_outputs(313) <= not (a xor b);
    layer5_outputs(314) <= not b or a;
    layer5_outputs(315) <= not b;
    layer5_outputs(316) <= not a or b;
    layer5_outputs(317) <= not a;
    layer5_outputs(318) <= a and not b;
    layer5_outputs(319) <= '1';
    layer5_outputs(320) <= b and not a;
    layer5_outputs(321) <= b;
    layer5_outputs(322) <= not (a or b);
    layer5_outputs(323) <= a;
    layer5_outputs(324) <= not a;
    layer5_outputs(325) <= not a;
    layer5_outputs(326) <= not b;
    layer5_outputs(327) <= not a;
    layer5_outputs(328) <= not b or a;
    layer5_outputs(329) <= b;
    layer5_outputs(330) <= not a;
    layer5_outputs(331) <= b and not a;
    layer5_outputs(332) <= b;
    layer5_outputs(333) <= a or b;
    layer5_outputs(334) <= b;
    layer5_outputs(335) <= not (a and b);
    layer5_outputs(336) <= not a or b;
    layer5_outputs(337) <= b and not a;
    layer5_outputs(338) <= b;
    layer5_outputs(339) <= not a or b;
    layer5_outputs(340) <= b;
    layer5_outputs(341) <= not (a or b);
    layer5_outputs(342) <= not a;
    layer5_outputs(343) <= not (a xor b);
    layer5_outputs(344) <= a xor b;
    layer5_outputs(345) <= not a or b;
    layer5_outputs(346) <= not (a xor b);
    layer5_outputs(347) <= a;
    layer5_outputs(348) <= b and not a;
    layer5_outputs(349) <= a;
    layer5_outputs(350) <= b;
    layer5_outputs(351) <= a xor b;
    layer5_outputs(352) <= not a or b;
    layer5_outputs(353) <= not a;
    layer5_outputs(354) <= b;
    layer5_outputs(355) <= not a;
    layer5_outputs(356) <= not b;
    layer5_outputs(357) <= not b;
    layer5_outputs(358) <= not (a or b);
    layer5_outputs(359) <= a;
    layer5_outputs(360) <= not b or a;
    layer5_outputs(361) <= not (a xor b);
    layer5_outputs(362) <= a and not b;
    layer5_outputs(363) <= b;
    layer5_outputs(364) <= a;
    layer5_outputs(365) <= a or b;
    layer5_outputs(366) <= not (a or b);
    layer5_outputs(367) <= a xor b;
    layer5_outputs(368) <= not (a or b);
    layer5_outputs(369) <= b and not a;
    layer5_outputs(370) <= b and not a;
    layer5_outputs(371) <= '1';
    layer5_outputs(372) <= a;
    layer5_outputs(373) <= not b;
    layer5_outputs(374) <= a xor b;
    layer5_outputs(375) <= a;
    layer5_outputs(376) <= b;
    layer5_outputs(377) <= a;
    layer5_outputs(378) <= not b;
    layer5_outputs(379) <= not (a xor b);
    layer5_outputs(380) <= a;
    layer5_outputs(381) <= not (a xor b);
    layer5_outputs(382) <= b and not a;
    layer5_outputs(383) <= a and not b;
    layer5_outputs(384) <= not b;
    layer5_outputs(385) <= not a;
    layer5_outputs(386) <= not (a or b);
    layer5_outputs(387) <= not b;
    layer5_outputs(388) <= not a;
    layer5_outputs(389) <= a and b;
    layer5_outputs(390) <= a or b;
    layer5_outputs(391) <= a and b;
    layer5_outputs(392) <= a or b;
    layer5_outputs(393) <= b;
    layer5_outputs(394) <= a and b;
    layer5_outputs(395) <= not a or b;
    layer5_outputs(396) <= not b;
    layer5_outputs(397) <= not a;
    layer5_outputs(398) <= not b;
    layer5_outputs(399) <= a and not b;
    layer5_outputs(400) <= not (a or b);
    layer5_outputs(401) <= a;
    layer5_outputs(402) <= not a;
    layer5_outputs(403) <= not b or a;
    layer5_outputs(404) <= a;
    layer5_outputs(405) <= not a or b;
    layer5_outputs(406) <= not (a and b);
    layer5_outputs(407) <= not b;
    layer5_outputs(408) <= '1';
    layer5_outputs(409) <= a;
    layer5_outputs(410) <= b;
    layer5_outputs(411) <= not (a and b);
    layer5_outputs(412) <= b and not a;
    layer5_outputs(413) <= b;
    layer5_outputs(414) <= b;
    layer5_outputs(415) <= not b;
    layer5_outputs(416) <= not a or b;
    layer5_outputs(417) <= a and not b;
    layer5_outputs(418) <= not (a xor b);
    layer5_outputs(419) <= not b or a;
    layer5_outputs(420) <= b;
    layer5_outputs(421) <= b;
    layer5_outputs(422) <= not b;
    layer5_outputs(423) <= a xor b;
    layer5_outputs(424) <= not a;
    layer5_outputs(425) <= not b or a;
    layer5_outputs(426) <= not a;
    layer5_outputs(427) <= b;
    layer5_outputs(428) <= a or b;
    layer5_outputs(429) <= '1';
    layer5_outputs(430) <= b;
    layer5_outputs(431) <= '0';
    layer5_outputs(432) <= b;
    layer5_outputs(433) <= a and not b;
    layer5_outputs(434) <= a;
    layer5_outputs(435) <= not a;
    layer5_outputs(436) <= a and b;
    layer5_outputs(437) <= a and not b;
    layer5_outputs(438) <= a xor b;
    layer5_outputs(439) <= not (a or b);
    layer5_outputs(440) <= not (a or b);
    layer5_outputs(441) <= not (a xor b);
    layer5_outputs(442) <= not (a or b);
    layer5_outputs(443) <= a or b;
    layer5_outputs(444) <= not b or a;
    layer5_outputs(445) <= not b or a;
    layer5_outputs(446) <= b;
    layer5_outputs(447) <= not a or b;
    layer5_outputs(448) <= not (a or b);
    layer5_outputs(449) <= not (a xor b);
    layer5_outputs(450) <= not (a or b);
    layer5_outputs(451) <= b;
    layer5_outputs(452) <= not a or b;
    layer5_outputs(453) <= b and not a;
    layer5_outputs(454) <= not a or b;
    layer5_outputs(455) <= not b;
    layer5_outputs(456) <= not (a and b);
    layer5_outputs(457) <= not (a and b);
    layer5_outputs(458) <= b;
    layer5_outputs(459) <= a;
    layer5_outputs(460) <= not b;
    layer5_outputs(461) <= b;
    layer5_outputs(462) <= not (a or b);
    layer5_outputs(463) <= b;
    layer5_outputs(464) <= a or b;
    layer5_outputs(465) <= b;
    layer5_outputs(466) <= not a;
    layer5_outputs(467) <= a and not b;
    layer5_outputs(468) <= not a;
    layer5_outputs(469) <= not b;
    layer5_outputs(470) <= b;
    layer5_outputs(471) <= not (a xor b);
    layer5_outputs(472) <= not a or b;
    layer5_outputs(473) <= b and not a;
    layer5_outputs(474) <= not a;
    layer5_outputs(475) <= not b;
    layer5_outputs(476) <= not b;
    layer5_outputs(477) <= a xor b;
    layer5_outputs(478) <= a and not b;
    layer5_outputs(479) <= b;
    layer5_outputs(480) <= b and not a;
    layer5_outputs(481) <= not a;
    layer5_outputs(482) <= b;
    layer5_outputs(483) <= b;
    layer5_outputs(484) <= not (a or b);
    layer5_outputs(485) <= not b or a;
    layer5_outputs(486) <= not a;
    layer5_outputs(487) <= not b;
    layer5_outputs(488) <= a or b;
    layer5_outputs(489) <= not b;
    layer5_outputs(490) <= not (a or b);
    layer5_outputs(491) <= not b;
    layer5_outputs(492) <= a;
    layer5_outputs(493) <= b and not a;
    layer5_outputs(494) <= not a;
    layer5_outputs(495) <= not a or b;
    layer5_outputs(496) <= b;
    layer5_outputs(497) <= not b;
    layer5_outputs(498) <= b and not a;
    layer5_outputs(499) <= not b;
    layer5_outputs(500) <= b and not a;
    layer5_outputs(501) <= not (a and b);
    layer5_outputs(502) <= a and b;
    layer5_outputs(503) <= a and b;
    layer5_outputs(504) <= b;
    layer5_outputs(505) <= b and not a;
    layer5_outputs(506) <= not (a and b);
    layer5_outputs(507) <= a and not b;
    layer5_outputs(508) <= b;
    layer5_outputs(509) <= not b;
    layer5_outputs(510) <= not a;
    layer5_outputs(511) <= not a or b;
    layer5_outputs(512) <= '1';
    layer5_outputs(513) <= b;
    layer5_outputs(514) <= a xor b;
    layer5_outputs(515) <= not (a or b);
    layer5_outputs(516) <= not (a and b);
    layer5_outputs(517) <= not b;
    layer5_outputs(518) <= not a;
    layer5_outputs(519) <= not (a or b);
    layer5_outputs(520) <= b;
    layer5_outputs(521) <= a or b;
    layer5_outputs(522) <= not (a xor b);
    layer5_outputs(523) <= not b;
    layer5_outputs(524) <= not a or b;
    layer5_outputs(525) <= a and b;
    layer5_outputs(526) <= not b;
    layer5_outputs(527) <= not b;
    layer5_outputs(528) <= not a;
    layer5_outputs(529) <= not a;
    layer5_outputs(530) <= a xor b;
    layer5_outputs(531) <= b;
    layer5_outputs(532) <= not a;
    layer5_outputs(533) <= b;
    layer5_outputs(534) <= not (a or b);
    layer5_outputs(535) <= a xor b;
    layer5_outputs(536) <= b and not a;
    layer5_outputs(537) <= a;
    layer5_outputs(538) <= '0';
    layer5_outputs(539) <= a xor b;
    layer5_outputs(540) <= not a or b;
    layer5_outputs(541) <= a xor b;
    layer5_outputs(542) <= not (a or b);
    layer5_outputs(543) <= a and b;
    layer5_outputs(544) <= not a;
    layer5_outputs(545) <= b;
    layer5_outputs(546) <= a or b;
    layer5_outputs(547) <= a and b;
    layer5_outputs(548) <= a or b;
    layer5_outputs(549) <= a and not b;
    layer5_outputs(550) <= not (a or b);
    layer5_outputs(551) <= b;
    layer5_outputs(552) <= a xor b;
    layer5_outputs(553) <= not (a or b);
    layer5_outputs(554) <= not (a and b);
    layer5_outputs(555) <= a and b;
    layer5_outputs(556) <= not (a or b);
    layer5_outputs(557) <= b;
    layer5_outputs(558) <= b and not a;
    layer5_outputs(559) <= a xor b;
    layer5_outputs(560) <= not (a and b);
    layer5_outputs(561) <= a;
    layer5_outputs(562) <= not (a or b);
    layer5_outputs(563) <= not b;
    layer5_outputs(564) <= a xor b;
    layer5_outputs(565) <= not b or a;
    layer5_outputs(566) <= not a;
    layer5_outputs(567) <= not (a xor b);
    layer5_outputs(568) <= a xor b;
    layer5_outputs(569) <= not a;
    layer5_outputs(570) <= b and not a;
    layer5_outputs(571) <= a;
    layer5_outputs(572) <= a;
    layer5_outputs(573) <= a xor b;
    layer5_outputs(574) <= not b or a;
    layer5_outputs(575) <= b;
    layer5_outputs(576) <= not (a xor b);
    layer5_outputs(577) <= a and b;
    layer5_outputs(578) <= not a;
    layer5_outputs(579) <= not a;
    layer5_outputs(580) <= b;
    layer5_outputs(581) <= b and not a;
    layer5_outputs(582) <= b;
    layer5_outputs(583) <= b;
    layer5_outputs(584) <= b;
    layer5_outputs(585) <= a or b;
    layer5_outputs(586) <= not b;
    layer5_outputs(587) <= not (a and b);
    layer5_outputs(588) <= b;
    layer5_outputs(589) <= not b;
    layer5_outputs(590) <= a;
    layer5_outputs(591) <= not a or b;
    layer5_outputs(592) <= not a;
    layer5_outputs(593) <= not (a and b);
    layer5_outputs(594) <= a xor b;
    layer5_outputs(595) <= a;
    layer5_outputs(596) <= b and not a;
    layer5_outputs(597) <= b and not a;
    layer5_outputs(598) <= a or b;
    layer5_outputs(599) <= a;
    layer5_outputs(600) <= a or b;
    layer5_outputs(601) <= a;
    layer5_outputs(602) <= a;
    layer5_outputs(603) <= b;
    layer5_outputs(604) <= b;
    layer5_outputs(605) <= not a;
    layer5_outputs(606) <= not b;
    layer5_outputs(607) <= a xor b;
    layer5_outputs(608) <= a or b;
    layer5_outputs(609) <= a and b;
    layer5_outputs(610) <= a xor b;
    layer5_outputs(611) <= b and not a;
    layer5_outputs(612) <= not a;
    layer5_outputs(613) <= not (a xor b);
    layer5_outputs(614) <= not (a xor b);
    layer5_outputs(615) <= b;
    layer5_outputs(616) <= a;
    layer5_outputs(617) <= b;
    layer5_outputs(618) <= not b;
    layer5_outputs(619) <= b;
    layer5_outputs(620) <= '1';
    layer5_outputs(621) <= not a or b;
    layer5_outputs(622) <= not (a or b);
    layer5_outputs(623) <= a and not b;
    layer5_outputs(624) <= b and not a;
    layer5_outputs(625) <= b;
    layer5_outputs(626) <= not b;
    layer5_outputs(627) <= b;
    layer5_outputs(628) <= a and b;
    layer5_outputs(629) <= a;
    layer5_outputs(630) <= not (a or b);
    layer5_outputs(631) <= not (a or b);
    layer5_outputs(632) <= a and b;
    layer5_outputs(633) <= a and not b;
    layer5_outputs(634) <= b;
    layer5_outputs(635) <= a and b;
    layer5_outputs(636) <= not a;
    layer5_outputs(637) <= not b;
    layer5_outputs(638) <= a and b;
    layer5_outputs(639) <= not (a or b);
    layer5_outputs(640) <= not a or b;
    layer5_outputs(641) <= b;
    layer5_outputs(642) <= b;
    layer5_outputs(643) <= a or b;
    layer5_outputs(644) <= not b;
    layer5_outputs(645) <= b;
    layer5_outputs(646) <= a and b;
    layer5_outputs(647) <= not b;
    layer5_outputs(648) <= not b;
    layer5_outputs(649) <= a and b;
    layer5_outputs(650) <= not a;
    layer5_outputs(651) <= a;
    layer5_outputs(652) <= a xor b;
    layer5_outputs(653) <= b and not a;
    layer5_outputs(654) <= not a;
    layer5_outputs(655) <= '0';
    layer5_outputs(656) <= not a or b;
    layer5_outputs(657) <= a xor b;
    layer5_outputs(658) <= a;
    layer5_outputs(659) <= b;
    layer5_outputs(660) <= not b;
    layer5_outputs(661) <= a and not b;
    layer5_outputs(662) <= a and b;
    layer5_outputs(663) <= b and not a;
    layer5_outputs(664) <= not a;
    layer5_outputs(665) <= a and b;
    layer5_outputs(666) <= not b or a;
    layer5_outputs(667) <= not a;
    layer5_outputs(668) <= not (a or b);
    layer5_outputs(669) <= a;
    layer5_outputs(670) <= not (a or b);
    layer5_outputs(671) <= a and not b;
    layer5_outputs(672) <= a and b;
    layer5_outputs(673) <= a;
    layer5_outputs(674) <= a and not b;
    layer5_outputs(675) <= not a;
    layer5_outputs(676) <= not a;
    layer5_outputs(677) <= a and not b;
    layer5_outputs(678) <= not (a or b);
    layer5_outputs(679) <= not b;
    layer5_outputs(680) <= a and not b;
    layer5_outputs(681) <= a;
    layer5_outputs(682) <= not a;
    layer5_outputs(683) <= not a;
    layer5_outputs(684) <= '0';
    layer5_outputs(685) <= not (a or b);
    layer5_outputs(686) <= not b or a;
    layer5_outputs(687) <= b;
    layer5_outputs(688) <= b;
    layer5_outputs(689) <= not a;
    layer5_outputs(690) <= not a;
    layer5_outputs(691) <= not (a and b);
    layer5_outputs(692) <= b and not a;
    layer5_outputs(693) <= not (a and b);
    layer5_outputs(694) <= a and not b;
    layer5_outputs(695) <= not (a and b);
    layer5_outputs(696) <= a or b;
    layer5_outputs(697) <= b;
    layer5_outputs(698) <= b;
    layer5_outputs(699) <= not a or b;
    layer5_outputs(700) <= not a or b;
    layer5_outputs(701) <= not a;
    layer5_outputs(702) <= a and not b;
    layer5_outputs(703) <= b;
    layer5_outputs(704) <= a;
    layer5_outputs(705) <= b;
    layer5_outputs(706) <= not (a xor b);
    layer5_outputs(707) <= not b;
    layer5_outputs(708) <= a and not b;
    layer5_outputs(709) <= a and b;
    layer5_outputs(710) <= not b;
    layer5_outputs(711) <= not (a and b);
    layer5_outputs(712) <= a xor b;
    layer5_outputs(713) <= not a or b;
    layer5_outputs(714) <= not a or b;
    layer5_outputs(715) <= not b or a;
    layer5_outputs(716) <= a xor b;
    layer5_outputs(717) <= not b or a;
    layer5_outputs(718) <= not a;
    layer5_outputs(719) <= a;
    layer5_outputs(720) <= a;
    layer5_outputs(721) <= a;
    layer5_outputs(722) <= not b;
    layer5_outputs(723) <= not a;
    layer5_outputs(724) <= a xor b;
    layer5_outputs(725) <= not a or b;
    layer5_outputs(726) <= '0';
    layer5_outputs(727) <= not b or a;
    layer5_outputs(728) <= not (a or b);
    layer5_outputs(729) <= a xor b;
    layer5_outputs(730) <= a and not b;
    layer5_outputs(731) <= a and b;
    layer5_outputs(732) <= a xor b;
    layer5_outputs(733) <= a or b;
    layer5_outputs(734) <= a xor b;
    layer5_outputs(735) <= a;
    layer5_outputs(736) <= a and not b;
    layer5_outputs(737) <= not (a xor b);
    layer5_outputs(738) <= not a;
    layer5_outputs(739) <= not (a or b);
    layer5_outputs(740) <= a xor b;
    layer5_outputs(741) <= not (a or b);
    layer5_outputs(742) <= not a;
    layer5_outputs(743) <= not a;
    layer5_outputs(744) <= '1';
    layer5_outputs(745) <= a;
    layer5_outputs(746) <= not (a and b);
    layer5_outputs(747) <= not a;
    layer5_outputs(748) <= b and not a;
    layer5_outputs(749) <= b;
    layer5_outputs(750) <= not b;
    layer5_outputs(751) <= not b or a;
    layer5_outputs(752) <= not a or b;
    layer5_outputs(753) <= a;
    layer5_outputs(754) <= not (a xor b);
    layer5_outputs(755) <= b;
    layer5_outputs(756) <= a;
    layer5_outputs(757) <= a and not b;
    layer5_outputs(758) <= not b;
    layer5_outputs(759) <= not b or a;
    layer5_outputs(760) <= a;
    layer5_outputs(761) <= a and b;
    layer5_outputs(762) <= not a;
    layer5_outputs(763) <= not (a xor b);
    layer5_outputs(764) <= not a;
    layer5_outputs(765) <= a;
    layer5_outputs(766) <= b;
    layer5_outputs(767) <= b;
    layer5_outputs(768) <= b and not a;
    layer5_outputs(769) <= not b or a;
    layer5_outputs(770) <= a;
    layer5_outputs(771) <= a and b;
    layer5_outputs(772) <= b and not a;
    layer5_outputs(773) <= not (a xor b);
    layer5_outputs(774) <= not b;
    layer5_outputs(775) <= not (a or b);
    layer5_outputs(776) <= b and not a;
    layer5_outputs(777) <= a or b;
    layer5_outputs(778) <= a or b;
    layer5_outputs(779) <= not b or a;
    layer5_outputs(780) <= not (a and b);
    layer5_outputs(781) <= not a;
    layer5_outputs(782) <= not (a and b);
    layer5_outputs(783) <= '1';
    layer5_outputs(784) <= not b;
    layer5_outputs(785) <= not b;
    layer5_outputs(786) <= not b or a;
    layer5_outputs(787) <= a or b;
    layer5_outputs(788) <= not b;
    layer5_outputs(789) <= not (a xor b);
    layer5_outputs(790) <= a and not b;
    layer5_outputs(791) <= b;
    layer5_outputs(792) <= not b or a;
    layer5_outputs(793) <= a and not b;
    layer5_outputs(794) <= not (a xor b);
    layer5_outputs(795) <= not a;
    layer5_outputs(796) <= b;
    layer5_outputs(797) <= a;
    layer5_outputs(798) <= not a or b;
    layer5_outputs(799) <= not (a and b);
    layer5_outputs(800) <= not a or b;
    layer5_outputs(801) <= not b;
    layer5_outputs(802) <= a xor b;
    layer5_outputs(803) <= a and not b;
    layer5_outputs(804) <= b;
    layer5_outputs(805) <= b;
    layer5_outputs(806) <= a;
    layer5_outputs(807) <= not b or a;
    layer5_outputs(808) <= a;
    layer5_outputs(809) <= not b;
    layer5_outputs(810) <= a;
    layer5_outputs(811) <= not (a xor b);
    layer5_outputs(812) <= not (a or b);
    layer5_outputs(813) <= not (a xor b);
    layer5_outputs(814) <= a or b;
    layer5_outputs(815) <= a;
    layer5_outputs(816) <= not b;
    layer5_outputs(817) <= not a;
    layer5_outputs(818) <= a;
    layer5_outputs(819) <= a xor b;
    layer5_outputs(820) <= b and not a;
    layer5_outputs(821) <= not a;
    layer5_outputs(822) <= a;
    layer5_outputs(823) <= a xor b;
    layer5_outputs(824) <= b and not a;
    layer5_outputs(825) <= a;
    layer5_outputs(826) <= not (a xor b);
    layer5_outputs(827) <= a;
    layer5_outputs(828) <= b;
    layer5_outputs(829) <= not a;
    layer5_outputs(830) <= a xor b;
    layer5_outputs(831) <= '1';
    layer5_outputs(832) <= b;
    layer5_outputs(833) <= not (a and b);
    layer5_outputs(834) <= not (a xor b);
    layer5_outputs(835) <= not (a and b);
    layer5_outputs(836) <= not (a and b);
    layer5_outputs(837) <= b and not a;
    layer5_outputs(838) <= not b or a;
    layer5_outputs(839) <= not a;
    layer5_outputs(840) <= a or b;
    layer5_outputs(841) <= not a or b;
    layer5_outputs(842) <= a or b;
    layer5_outputs(843) <= a;
    layer5_outputs(844) <= not a;
    layer5_outputs(845) <= b;
    layer5_outputs(846) <= b;
    layer5_outputs(847) <= not a;
    layer5_outputs(848) <= b and not a;
    layer5_outputs(849) <= not b;
    layer5_outputs(850) <= a and b;
    layer5_outputs(851) <= not b;
    layer5_outputs(852) <= not b;
    layer5_outputs(853) <= a and b;
    layer5_outputs(854) <= not (a or b);
    layer5_outputs(855) <= '1';
    layer5_outputs(856) <= a;
    layer5_outputs(857) <= not a;
    layer5_outputs(858) <= a or b;
    layer5_outputs(859) <= a;
    layer5_outputs(860) <= not b;
    layer5_outputs(861) <= not a;
    layer5_outputs(862) <= not b;
    layer5_outputs(863) <= not (a or b);
    layer5_outputs(864) <= not a;
    layer5_outputs(865) <= a xor b;
    layer5_outputs(866) <= not b;
    layer5_outputs(867) <= '0';
    layer5_outputs(868) <= not (a or b);
    layer5_outputs(869) <= b;
    layer5_outputs(870) <= a;
    layer5_outputs(871) <= not b;
    layer5_outputs(872) <= not b;
    layer5_outputs(873) <= not a or b;
    layer5_outputs(874) <= b and not a;
    layer5_outputs(875) <= a or b;
    layer5_outputs(876) <= a or b;
    layer5_outputs(877) <= not (a xor b);
    layer5_outputs(878) <= not a;
    layer5_outputs(879) <= not a;
    layer5_outputs(880) <= not (a xor b);
    layer5_outputs(881) <= not b;
    layer5_outputs(882) <= a or b;
    layer5_outputs(883) <= a xor b;
    layer5_outputs(884) <= not a;
    layer5_outputs(885) <= not (a and b);
    layer5_outputs(886) <= b;
    layer5_outputs(887) <= not (a xor b);
    layer5_outputs(888) <= '1';
    layer5_outputs(889) <= not a;
    layer5_outputs(890) <= a and b;
    layer5_outputs(891) <= not (a and b);
    layer5_outputs(892) <= not (a or b);
    layer5_outputs(893) <= not a;
    layer5_outputs(894) <= not b;
    layer5_outputs(895) <= not (a and b);
    layer5_outputs(896) <= b;
    layer5_outputs(897) <= not b;
    layer5_outputs(898) <= not a;
    layer5_outputs(899) <= not a;
    layer5_outputs(900) <= not b or a;
    layer5_outputs(901) <= not a;
    layer5_outputs(902) <= a xor b;
    layer5_outputs(903) <= not (a and b);
    layer5_outputs(904) <= not b;
    layer5_outputs(905) <= a;
    layer5_outputs(906) <= b;
    layer5_outputs(907) <= not b or a;
    layer5_outputs(908) <= not a;
    layer5_outputs(909) <= not a;
    layer5_outputs(910) <= '0';
    layer5_outputs(911) <= not b;
    layer5_outputs(912) <= not a;
    layer5_outputs(913) <= a and b;
    layer5_outputs(914) <= not b;
    layer5_outputs(915) <= not a;
    layer5_outputs(916) <= not a or b;
    layer5_outputs(917) <= not b;
    layer5_outputs(918) <= not b;
    layer5_outputs(919) <= not b;
    layer5_outputs(920) <= a and not b;
    layer5_outputs(921) <= not a;
    layer5_outputs(922) <= not a;
    layer5_outputs(923) <= b;
    layer5_outputs(924) <= not a;
    layer5_outputs(925) <= a and not b;
    layer5_outputs(926) <= a;
    layer5_outputs(927) <= b and not a;
    layer5_outputs(928) <= a or b;
    layer5_outputs(929) <= a;
    layer5_outputs(930) <= a xor b;
    layer5_outputs(931) <= not b;
    layer5_outputs(932) <= a or b;
    layer5_outputs(933) <= not a;
    layer5_outputs(934) <= b;
    layer5_outputs(935) <= not b or a;
    layer5_outputs(936) <= b;
    layer5_outputs(937) <= not (a and b);
    layer5_outputs(938) <= a or b;
    layer5_outputs(939) <= b;
    layer5_outputs(940) <= not b or a;
    layer5_outputs(941) <= a and b;
    layer5_outputs(942) <= a or b;
    layer5_outputs(943) <= a;
    layer5_outputs(944) <= b;
    layer5_outputs(945) <= b and not a;
    layer5_outputs(946) <= a;
    layer5_outputs(947) <= a;
    layer5_outputs(948) <= not a;
    layer5_outputs(949) <= a;
    layer5_outputs(950) <= not a;
    layer5_outputs(951) <= b;
    layer5_outputs(952) <= not b;
    layer5_outputs(953) <= not a;
    layer5_outputs(954) <= a xor b;
    layer5_outputs(955) <= not b;
    layer5_outputs(956) <= b;
    layer5_outputs(957) <= b and not a;
    layer5_outputs(958) <= b and not a;
    layer5_outputs(959) <= not (a xor b);
    layer5_outputs(960) <= a xor b;
    layer5_outputs(961) <= b;
    layer5_outputs(962) <= a and not b;
    layer5_outputs(963) <= not (a xor b);
    layer5_outputs(964) <= a;
    layer5_outputs(965) <= not (a or b);
    layer5_outputs(966) <= not a;
    layer5_outputs(967) <= not a;
    layer5_outputs(968) <= not (a and b);
    layer5_outputs(969) <= not a;
    layer5_outputs(970) <= a and not b;
    layer5_outputs(971) <= b;
    layer5_outputs(972) <= b;
    layer5_outputs(973) <= not (a or b);
    layer5_outputs(974) <= not (a or b);
    layer5_outputs(975) <= not (a and b);
    layer5_outputs(976) <= not b;
    layer5_outputs(977) <= a;
    layer5_outputs(978) <= b;
    layer5_outputs(979) <= not b;
    layer5_outputs(980) <= a or b;
    layer5_outputs(981) <= b;
    layer5_outputs(982) <= a and not b;
    layer5_outputs(983) <= a;
    layer5_outputs(984) <= b;
    layer5_outputs(985) <= not b;
    layer5_outputs(986) <= not a;
    layer5_outputs(987) <= not a;
    layer5_outputs(988) <= b;
    layer5_outputs(989) <= a;
    layer5_outputs(990) <= not (a and b);
    layer5_outputs(991) <= a and not b;
    layer5_outputs(992) <= not a;
    layer5_outputs(993) <= not a;
    layer5_outputs(994) <= not b;
    layer5_outputs(995) <= not b;
    layer5_outputs(996) <= a;
    layer5_outputs(997) <= a;
    layer5_outputs(998) <= not a or b;
    layer5_outputs(999) <= b;
    layer5_outputs(1000) <= a;
    layer5_outputs(1001) <= b;
    layer5_outputs(1002) <= a and b;
    layer5_outputs(1003) <= b and not a;
    layer5_outputs(1004) <= not b;
    layer5_outputs(1005) <= not b;
    layer5_outputs(1006) <= a;
    layer5_outputs(1007) <= a or b;
    layer5_outputs(1008) <= a;
    layer5_outputs(1009) <= not (a xor b);
    layer5_outputs(1010) <= not a or b;
    layer5_outputs(1011) <= a or b;
    layer5_outputs(1012) <= a xor b;
    layer5_outputs(1013) <= not a;
    layer5_outputs(1014) <= a or b;
    layer5_outputs(1015) <= b;
    layer5_outputs(1016) <= a xor b;
    layer5_outputs(1017) <= not a;
    layer5_outputs(1018) <= not (a and b);
    layer5_outputs(1019) <= not b or a;
    layer5_outputs(1020) <= a;
    layer5_outputs(1021) <= b and not a;
    layer5_outputs(1022) <= not b;
    layer5_outputs(1023) <= a and not b;
    layer5_outputs(1024) <= b;
    layer5_outputs(1025) <= not b or a;
    layer5_outputs(1026) <= not (a or b);
    layer5_outputs(1027) <= not b or a;
    layer5_outputs(1028) <= b;
    layer5_outputs(1029) <= not a;
    layer5_outputs(1030) <= not b;
    layer5_outputs(1031) <= a and b;
    layer5_outputs(1032) <= a;
    layer5_outputs(1033) <= a and b;
    layer5_outputs(1034) <= a and b;
    layer5_outputs(1035) <= b;
    layer5_outputs(1036) <= b;
    layer5_outputs(1037) <= not (a and b);
    layer5_outputs(1038) <= not b;
    layer5_outputs(1039) <= b;
    layer5_outputs(1040) <= not (a xor b);
    layer5_outputs(1041) <= a;
    layer5_outputs(1042) <= not (a xor b);
    layer5_outputs(1043) <= not b;
    layer5_outputs(1044) <= a and not b;
    layer5_outputs(1045) <= not b;
    layer5_outputs(1046) <= b;
    layer5_outputs(1047) <= not b;
    layer5_outputs(1048) <= a and not b;
    layer5_outputs(1049) <= not (a xor b);
    layer5_outputs(1050) <= not (a xor b);
    layer5_outputs(1051) <= not (a or b);
    layer5_outputs(1052) <= '1';
    layer5_outputs(1053) <= not (a xor b);
    layer5_outputs(1054) <= a xor b;
    layer5_outputs(1055) <= not a;
    layer5_outputs(1056) <= not a;
    layer5_outputs(1057) <= not (a and b);
    layer5_outputs(1058) <= a;
    layer5_outputs(1059) <= a and not b;
    layer5_outputs(1060) <= a and b;
    layer5_outputs(1061) <= not a;
    layer5_outputs(1062) <= not (a xor b);
    layer5_outputs(1063) <= not b;
    layer5_outputs(1064) <= a;
    layer5_outputs(1065) <= a or b;
    layer5_outputs(1066) <= b and not a;
    layer5_outputs(1067) <= not (a xor b);
    layer5_outputs(1068) <= a and not b;
    layer5_outputs(1069) <= a;
    layer5_outputs(1070) <= not a or b;
    layer5_outputs(1071) <= a;
    layer5_outputs(1072) <= not (a or b);
    layer5_outputs(1073) <= not (a or b);
    layer5_outputs(1074) <= a and b;
    layer5_outputs(1075) <= a and b;
    layer5_outputs(1076) <= not (a xor b);
    layer5_outputs(1077) <= a;
    layer5_outputs(1078) <= not a or b;
    layer5_outputs(1079) <= '1';
    layer5_outputs(1080) <= b;
    layer5_outputs(1081) <= not b;
    layer5_outputs(1082) <= a xor b;
    layer5_outputs(1083) <= a or b;
    layer5_outputs(1084) <= a;
    layer5_outputs(1085) <= b and not a;
    layer5_outputs(1086) <= a xor b;
    layer5_outputs(1087) <= not a;
    layer5_outputs(1088) <= not a;
    layer5_outputs(1089) <= b;
    layer5_outputs(1090) <= not a;
    layer5_outputs(1091) <= a and not b;
    layer5_outputs(1092) <= not (a or b);
    layer5_outputs(1093) <= not (a xor b);
    layer5_outputs(1094) <= not a;
    layer5_outputs(1095) <= not (a and b);
    layer5_outputs(1096) <= not a;
    layer5_outputs(1097) <= not (a xor b);
    layer5_outputs(1098) <= not b or a;
    layer5_outputs(1099) <= b and not a;
    layer5_outputs(1100) <= not (a and b);
    layer5_outputs(1101) <= a or b;
    layer5_outputs(1102) <= a;
    layer5_outputs(1103) <= not (a xor b);
    layer5_outputs(1104) <= b;
    layer5_outputs(1105) <= a and b;
    layer5_outputs(1106) <= not a or b;
    layer5_outputs(1107) <= b;
    layer5_outputs(1108) <= a;
    layer5_outputs(1109) <= not b;
    layer5_outputs(1110) <= a and b;
    layer5_outputs(1111) <= b;
    layer5_outputs(1112) <= b and not a;
    layer5_outputs(1113) <= a and b;
    layer5_outputs(1114) <= not a;
    layer5_outputs(1115) <= a and not b;
    layer5_outputs(1116) <= a;
    layer5_outputs(1117) <= not a;
    layer5_outputs(1118) <= a and not b;
    layer5_outputs(1119) <= b;
    layer5_outputs(1120) <= not a;
    layer5_outputs(1121) <= a and b;
    layer5_outputs(1122) <= a and b;
    layer5_outputs(1123) <= a and b;
    layer5_outputs(1124) <= b;
    layer5_outputs(1125) <= a and b;
    layer5_outputs(1126) <= a and b;
    layer5_outputs(1127) <= a and not b;
    layer5_outputs(1128) <= a;
    layer5_outputs(1129) <= a xor b;
    layer5_outputs(1130) <= a or b;
    layer5_outputs(1131) <= not (a or b);
    layer5_outputs(1132) <= b;
    layer5_outputs(1133) <= a or b;
    layer5_outputs(1134) <= not (a or b);
    layer5_outputs(1135) <= not a;
    layer5_outputs(1136) <= not a;
    layer5_outputs(1137) <= a or b;
    layer5_outputs(1138) <= not a;
    layer5_outputs(1139) <= not (a xor b);
    layer5_outputs(1140) <= not (a and b);
    layer5_outputs(1141) <= a;
    layer5_outputs(1142) <= a;
    layer5_outputs(1143) <= not b or a;
    layer5_outputs(1144) <= not b;
    layer5_outputs(1145) <= not a or b;
    layer5_outputs(1146) <= not (a xor b);
    layer5_outputs(1147) <= a and b;
    layer5_outputs(1148) <= not (a and b);
    layer5_outputs(1149) <= a and b;
    layer5_outputs(1150) <= not a or b;
    layer5_outputs(1151) <= a;
    layer5_outputs(1152) <= b;
    layer5_outputs(1153) <= '1';
    layer5_outputs(1154) <= a and b;
    layer5_outputs(1155) <= a;
    layer5_outputs(1156) <= not a or b;
    layer5_outputs(1157) <= b and not a;
    layer5_outputs(1158) <= not a;
    layer5_outputs(1159) <= not a or b;
    layer5_outputs(1160) <= a and not b;
    layer5_outputs(1161) <= a and not b;
    layer5_outputs(1162) <= not b;
    layer5_outputs(1163) <= a or b;
    layer5_outputs(1164) <= a;
    layer5_outputs(1165) <= a;
    layer5_outputs(1166) <= b;
    layer5_outputs(1167) <= a and not b;
    layer5_outputs(1168) <= a;
    layer5_outputs(1169) <= a;
    layer5_outputs(1170) <= not (a xor b);
    layer5_outputs(1171) <= not b;
    layer5_outputs(1172) <= b;
    layer5_outputs(1173) <= not a;
    layer5_outputs(1174) <= not b;
    layer5_outputs(1175) <= a;
    layer5_outputs(1176) <= a;
    layer5_outputs(1177) <= a xor b;
    layer5_outputs(1178) <= not a or b;
    layer5_outputs(1179) <= a xor b;
    layer5_outputs(1180) <= a and b;
    layer5_outputs(1181) <= not (a and b);
    layer5_outputs(1182) <= a xor b;
    layer5_outputs(1183) <= a and b;
    layer5_outputs(1184) <= not (a or b);
    layer5_outputs(1185) <= a and not b;
    layer5_outputs(1186) <= a and not b;
    layer5_outputs(1187) <= not (a and b);
    layer5_outputs(1188) <= b and not a;
    layer5_outputs(1189) <= not a;
    layer5_outputs(1190) <= a xor b;
    layer5_outputs(1191) <= not b;
    layer5_outputs(1192) <= b;
    layer5_outputs(1193) <= a;
    layer5_outputs(1194) <= a;
    layer5_outputs(1195) <= b;
    layer5_outputs(1196) <= not a or b;
    layer5_outputs(1197) <= a or b;
    layer5_outputs(1198) <= not a or b;
    layer5_outputs(1199) <= not (a xor b);
    layer5_outputs(1200) <= a;
    layer5_outputs(1201) <= a and b;
    layer5_outputs(1202) <= a xor b;
    layer5_outputs(1203) <= b and not a;
    layer5_outputs(1204) <= not a;
    layer5_outputs(1205) <= b;
    layer5_outputs(1206) <= not b;
    layer5_outputs(1207) <= a and not b;
    layer5_outputs(1208) <= not b;
    layer5_outputs(1209) <= a;
    layer5_outputs(1210) <= not (a xor b);
    layer5_outputs(1211) <= a;
    layer5_outputs(1212) <= b;
    layer5_outputs(1213) <= not (a and b);
    layer5_outputs(1214) <= not a;
    layer5_outputs(1215) <= not a or b;
    layer5_outputs(1216) <= b;
    layer5_outputs(1217) <= b;
    layer5_outputs(1218) <= not b;
    layer5_outputs(1219) <= not b or a;
    layer5_outputs(1220) <= a;
    layer5_outputs(1221) <= not a;
    layer5_outputs(1222) <= a;
    layer5_outputs(1223) <= not (a and b);
    layer5_outputs(1224) <= not a;
    layer5_outputs(1225) <= a;
    layer5_outputs(1226) <= a;
    layer5_outputs(1227) <= not a or b;
    layer5_outputs(1228) <= a xor b;
    layer5_outputs(1229) <= not (a or b);
    layer5_outputs(1230) <= b;
    layer5_outputs(1231) <= a;
    layer5_outputs(1232) <= not b or a;
    layer5_outputs(1233) <= a xor b;
    layer5_outputs(1234) <= not b;
    layer5_outputs(1235) <= a;
    layer5_outputs(1236) <= a or b;
    layer5_outputs(1237) <= not (a xor b);
    layer5_outputs(1238) <= a;
    layer5_outputs(1239) <= not (a xor b);
    layer5_outputs(1240) <= not (a xor b);
    layer5_outputs(1241) <= a;
    layer5_outputs(1242) <= a and not b;
    layer5_outputs(1243) <= a;
    layer5_outputs(1244) <= not a or b;
    layer5_outputs(1245) <= b;
    layer5_outputs(1246) <= not a;
    layer5_outputs(1247) <= not a;
    layer5_outputs(1248) <= not (a and b);
    layer5_outputs(1249) <= not a;
    layer5_outputs(1250) <= a and b;
    layer5_outputs(1251) <= '0';
    layer5_outputs(1252) <= not b;
    layer5_outputs(1253) <= not (a or b);
    layer5_outputs(1254) <= a xor b;
    layer5_outputs(1255) <= a;
    layer5_outputs(1256) <= a xor b;
    layer5_outputs(1257) <= b and not a;
    layer5_outputs(1258) <= not a;
    layer5_outputs(1259) <= a xor b;
    layer5_outputs(1260) <= not a or b;
    layer5_outputs(1261) <= '1';
    layer5_outputs(1262) <= b and not a;
    layer5_outputs(1263) <= not a;
    layer5_outputs(1264) <= not b or a;
    layer5_outputs(1265) <= not b or a;
    layer5_outputs(1266) <= not (a xor b);
    layer5_outputs(1267) <= not b;
    layer5_outputs(1268) <= not a;
    layer5_outputs(1269) <= not a or b;
    layer5_outputs(1270) <= a and not b;
    layer5_outputs(1271) <= not a;
    layer5_outputs(1272) <= not b or a;
    layer5_outputs(1273) <= b;
    layer5_outputs(1274) <= not a or b;
    layer5_outputs(1275) <= not (a xor b);
    layer5_outputs(1276) <= a and b;
    layer5_outputs(1277) <= not b;
    layer5_outputs(1278) <= a or b;
    layer5_outputs(1279) <= not a;
    layer5_outputs(1280) <= not a;
    layer5_outputs(1281) <= '0';
    layer5_outputs(1282) <= not b;
    layer5_outputs(1283) <= a xor b;
    layer5_outputs(1284) <= not a;
    layer5_outputs(1285) <= not b;
    layer5_outputs(1286) <= a xor b;
    layer5_outputs(1287) <= a or b;
    layer5_outputs(1288) <= b and not a;
    layer5_outputs(1289) <= b;
    layer5_outputs(1290) <= not a or b;
    layer5_outputs(1291) <= a;
    layer5_outputs(1292) <= b;
    layer5_outputs(1293) <= not a or b;
    layer5_outputs(1294) <= a and b;
    layer5_outputs(1295) <= not b;
    layer5_outputs(1296) <= not b or a;
    layer5_outputs(1297) <= not a;
    layer5_outputs(1298) <= b and not a;
    layer5_outputs(1299) <= a xor b;
    layer5_outputs(1300) <= not a;
    layer5_outputs(1301) <= a;
    layer5_outputs(1302) <= b;
    layer5_outputs(1303) <= b;
    layer5_outputs(1304) <= not a;
    layer5_outputs(1305) <= not b or a;
    layer5_outputs(1306) <= not a;
    layer5_outputs(1307) <= b and not a;
    layer5_outputs(1308) <= not a;
    layer5_outputs(1309) <= not (a and b);
    layer5_outputs(1310) <= b;
    layer5_outputs(1311) <= not (a xor b);
    layer5_outputs(1312) <= not b;
    layer5_outputs(1313) <= not b;
    layer5_outputs(1314) <= a;
    layer5_outputs(1315) <= not (a or b);
    layer5_outputs(1316) <= a xor b;
    layer5_outputs(1317) <= a;
    layer5_outputs(1318) <= a and not b;
    layer5_outputs(1319) <= not b;
    layer5_outputs(1320) <= not b;
    layer5_outputs(1321) <= not (a and b);
    layer5_outputs(1322) <= a;
    layer5_outputs(1323) <= a;
    layer5_outputs(1324) <= a;
    layer5_outputs(1325) <= not (a xor b);
    layer5_outputs(1326) <= not (a and b);
    layer5_outputs(1327) <= not a;
    layer5_outputs(1328) <= not (a or b);
    layer5_outputs(1329) <= not b or a;
    layer5_outputs(1330) <= b and not a;
    layer5_outputs(1331) <= not a;
    layer5_outputs(1332) <= not (a or b);
    layer5_outputs(1333) <= not a or b;
    layer5_outputs(1334) <= not (a or b);
    layer5_outputs(1335) <= b and not a;
    layer5_outputs(1336) <= a xor b;
    layer5_outputs(1337) <= a;
    layer5_outputs(1338) <= a or b;
    layer5_outputs(1339) <= not a;
    layer5_outputs(1340) <= not b;
    layer5_outputs(1341) <= not a;
    layer5_outputs(1342) <= b;
    layer5_outputs(1343) <= a or b;
    layer5_outputs(1344) <= a and not b;
    layer5_outputs(1345) <= a and not b;
    layer5_outputs(1346) <= a;
    layer5_outputs(1347) <= not (a and b);
    layer5_outputs(1348) <= not b;
    layer5_outputs(1349) <= not (a or b);
    layer5_outputs(1350) <= a;
    layer5_outputs(1351) <= not b or a;
    layer5_outputs(1352) <= a and not b;
    layer5_outputs(1353) <= not (a xor b);
    layer5_outputs(1354) <= not b;
    layer5_outputs(1355) <= b and not a;
    layer5_outputs(1356) <= not (a and b);
    layer5_outputs(1357) <= not a;
    layer5_outputs(1358) <= not a;
    layer5_outputs(1359) <= '1';
    layer5_outputs(1360) <= not a or b;
    layer5_outputs(1361) <= a;
    layer5_outputs(1362) <= not a or b;
    layer5_outputs(1363) <= not a or b;
    layer5_outputs(1364) <= not a;
    layer5_outputs(1365) <= b and not a;
    layer5_outputs(1366) <= not (a xor b);
    layer5_outputs(1367) <= a;
    layer5_outputs(1368) <= a;
    layer5_outputs(1369) <= b;
    layer5_outputs(1370) <= not (a and b);
    layer5_outputs(1371) <= b and not a;
    layer5_outputs(1372) <= a;
    layer5_outputs(1373) <= not (a and b);
    layer5_outputs(1374) <= not (a xor b);
    layer5_outputs(1375) <= a;
    layer5_outputs(1376) <= not b;
    layer5_outputs(1377) <= b and not a;
    layer5_outputs(1378) <= not (a xor b);
    layer5_outputs(1379) <= not a;
    layer5_outputs(1380) <= a;
    layer5_outputs(1381) <= not b;
    layer5_outputs(1382) <= not (a or b);
    layer5_outputs(1383) <= not b;
    layer5_outputs(1384) <= b;
    layer5_outputs(1385) <= a and not b;
    layer5_outputs(1386) <= b;
    layer5_outputs(1387) <= not (a xor b);
    layer5_outputs(1388) <= not b;
    layer5_outputs(1389) <= a xor b;
    layer5_outputs(1390) <= not b;
    layer5_outputs(1391) <= not b;
    layer5_outputs(1392) <= b;
    layer5_outputs(1393) <= a;
    layer5_outputs(1394) <= '0';
    layer5_outputs(1395) <= a and b;
    layer5_outputs(1396) <= '0';
    layer5_outputs(1397) <= a;
    layer5_outputs(1398) <= not (a and b);
    layer5_outputs(1399) <= b;
    layer5_outputs(1400) <= a xor b;
    layer5_outputs(1401) <= a;
    layer5_outputs(1402) <= not a;
    layer5_outputs(1403) <= b;
    layer5_outputs(1404) <= not a;
    layer5_outputs(1405) <= a;
    layer5_outputs(1406) <= '0';
    layer5_outputs(1407) <= a or b;
    layer5_outputs(1408) <= not (a or b);
    layer5_outputs(1409) <= a and not b;
    layer5_outputs(1410) <= b;
    layer5_outputs(1411) <= a or b;
    layer5_outputs(1412) <= a;
    layer5_outputs(1413) <= not (a or b);
    layer5_outputs(1414) <= not a or b;
    layer5_outputs(1415) <= not a;
    layer5_outputs(1416) <= a xor b;
    layer5_outputs(1417) <= not (a and b);
    layer5_outputs(1418) <= not a;
    layer5_outputs(1419) <= not a;
    layer5_outputs(1420) <= not a;
    layer5_outputs(1421) <= not (a and b);
    layer5_outputs(1422) <= not b;
    layer5_outputs(1423) <= a;
    layer5_outputs(1424) <= b and not a;
    layer5_outputs(1425) <= a xor b;
    layer5_outputs(1426) <= a and not b;
    layer5_outputs(1427) <= a xor b;
    layer5_outputs(1428) <= '1';
    layer5_outputs(1429) <= not b;
    layer5_outputs(1430) <= b and not a;
    layer5_outputs(1431) <= not a;
    layer5_outputs(1432) <= not a;
    layer5_outputs(1433) <= not (a xor b);
    layer5_outputs(1434) <= not a or b;
    layer5_outputs(1435) <= b;
    layer5_outputs(1436) <= a xor b;
    layer5_outputs(1437) <= not b;
    layer5_outputs(1438) <= a;
    layer5_outputs(1439) <= not b;
    layer5_outputs(1440) <= b and not a;
    layer5_outputs(1441) <= not a;
    layer5_outputs(1442) <= a or b;
    layer5_outputs(1443) <= a;
    layer5_outputs(1444) <= not a;
    layer5_outputs(1445) <= not (a xor b);
    layer5_outputs(1446) <= a;
    layer5_outputs(1447) <= a and not b;
    layer5_outputs(1448) <= b and not a;
    layer5_outputs(1449) <= a;
    layer5_outputs(1450) <= not b;
    layer5_outputs(1451) <= not b or a;
    layer5_outputs(1452) <= a and not b;
    layer5_outputs(1453) <= not b;
    layer5_outputs(1454) <= not b;
    layer5_outputs(1455) <= not a;
    layer5_outputs(1456) <= not a;
    layer5_outputs(1457) <= a or b;
    layer5_outputs(1458) <= a and b;
    layer5_outputs(1459) <= not (a or b);
    layer5_outputs(1460) <= a;
    layer5_outputs(1461) <= '0';
    layer5_outputs(1462) <= b;
    layer5_outputs(1463) <= not (a xor b);
    layer5_outputs(1464) <= not (a or b);
    layer5_outputs(1465) <= not a;
    layer5_outputs(1466) <= not (a or b);
    layer5_outputs(1467) <= a and not b;
    layer5_outputs(1468) <= b and not a;
    layer5_outputs(1469) <= not (a and b);
    layer5_outputs(1470) <= not (a xor b);
    layer5_outputs(1471) <= b;
    layer5_outputs(1472) <= not (a xor b);
    layer5_outputs(1473) <= b;
    layer5_outputs(1474) <= b;
    layer5_outputs(1475) <= a or b;
    layer5_outputs(1476) <= a;
    layer5_outputs(1477) <= not a;
    layer5_outputs(1478) <= not (a and b);
    layer5_outputs(1479) <= not b or a;
    layer5_outputs(1480) <= b;
    layer5_outputs(1481) <= not (a xor b);
    layer5_outputs(1482) <= b;
    layer5_outputs(1483) <= a xor b;
    layer5_outputs(1484) <= a xor b;
    layer5_outputs(1485) <= a;
    layer5_outputs(1486) <= not a;
    layer5_outputs(1487) <= a;
    layer5_outputs(1488) <= a xor b;
    layer5_outputs(1489) <= not (a and b);
    layer5_outputs(1490) <= not (a xor b);
    layer5_outputs(1491) <= a xor b;
    layer5_outputs(1492) <= not (a xor b);
    layer5_outputs(1493) <= not a;
    layer5_outputs(1494) <= not b;
    layer5_outputs(1495) <= a or b;
    layer5_outputs(1496) <= not a;
    layer5_outputs(1497) <= a or b;
    layer5_outputs(1498) <= b;
    layer5_outputs(1499) <= a xor b;
    layer5_outputs(1500) <= not (a xor b);
    layer5_outputs(1501) <= '1';
    layer5_outputs(1502) <= '0';
    layer5_outputs(1503) <= not a;
    layer5_outputs(1504) <= not (a xor b);
    layer5_outputs(1505) <= not a or b;
    layer5_outputs(1506) <= not a or b;
    layer5_outputs(1507) <= not (a and b);
    layer5_outputs(1508) <= '0';
    layer5_outputs(1509) <= a xor b;
    layer5_outputs(1510) <= not b;
    layer5_outputs(1511) <= a;
    layer5_outputs(1512) <= not b;
    layer5_outputs(1513) <= not (a xor b);
    layer5_outputs(1514) <= not b;
    layer5_outputs(1515) <= a;
    layer5_outputs(1516) <= not b;
    layer5_outputs(1517) <= not (a or b);
    layer5_outputs(1518) <= not b;
    layer5_outputs(1519) <= not (a xor b);
    layer5_outputs(1520) <= not (a and b);
    layer5_outputs(1521) <= b;
    layer5_outputs(1522) <= b;
    layer5_outputs(1523) <= b;
    layer5_outputs(1524) <= not b;
    layer5_outputs(1525) <= not a;
    layer5_outputs(1526) <= not b;
    layer5_outputs(1527) <= not (a xor b);
    layer5_outputs(1528) <= not b;
    layer5_outputs(1529) <= a;
    layer5_outputs(1530) <= a;
    layer5_outputs(1531) <= not (a or b);
    layer5_outputs(1532) <= a and not b;
    layer5_outputs(1533) <= a xor b;
    layer5_outputs(1534) <= not a;
    layer5_outputs(1535) <= a or b;
    layer5_outputs(1536) <= not (a and b);
    layer5_outputs(1537) <= not a or b;
    layer5_outputs(1538) <= a;
    layer5_outputs(1539) <= a xor b;
    layer5_outputs(1540) <= not a;
    layer5_outputs(1541) <= a or b;
    layer5_outputs(1542) <= not (a or b);
    layer5_outputs(1543) <= not a or b;
    layer5_outputs(1544) <= a xor b;
    layer5_outputs(1545) <= a xor b;
    layer5_outputs(1546) <= a or b;
    layer5_outputs(1547) <= b and not a;
    layer5_outputs(1548) <= not a;
    layer5_outputs(1549) <= a and not b;
    layer5_outputs(1550) <= a and not b;
    layer5_outputs(1551) <= not (a xor b);
    layer5_outputs(1552) <= not b;
    layer5_outputs(1553) <= not a or b;
    layer5_outputs(1554) <= a;
    layer5_outputs(1555) <= b;
    layer5_outputs(1556) <= a and b;
    layer5_outputs(1557) <= b;
    layer5_outputs(1558) <= not (a xor b);
    layer5_outputs(1559) <= not b;
    layer5_outputs(1560) <= not b;
    layer5_outputs(1561) <= not a;
    layer5_outputs(1562) <= a xor b;
    layer5_outputs(1563) <= not b or a;
    layer5_outputs(1564) <= a xor b;
    layer5_outputs(1565) <= a;
    layer5_outputs(1566) <= not (a xor b);
    layer5_outputs(1567) <= not (a xor b);
    layer5_outputs(1568) <= a and not b;
    layer5_outputs(1569) <= not b or a;
    layer5_outputs(1570) <= b and not a;
    layer5_outputs(1571) <= not a;
    layer5_outputs(1572) <= not b;
    layer5_outputs(1573) <= a and b;
    layer5_outputs(1574) <= a and not b;
    layer5_outputs(1575) <= b and not a;
    layer5_outputs(1576) <= not a;
    layer5_outputs(1577) <= b;
    layer5_outputs(1578) <= a and b;
    layer5_outputs(1579) <= not b;
    layer5_outputs(1580) <= not b;
    layer5_outputs(1581) <= not a;
    layer5_outputs(1582) <= not (a or b);
    layer5_outputs(1583) <= not b;
    layer5_outputs(1584) <= a;
    layer5_outputs(1585) <= not a or b;
    layer5_outputs(1586) <= not b;
    layer5_outputs(1587) <= a;
    layer5_outputs(1588) <= b;
    layer5_outputs(1589) <= not (a or b);
    layer5_outputs(1590) <= a xor b;
    layer5_outputs(1591) <= a;
    layer5_outputs(1592) <= b and not a;
    layer5_outputs(1593) <= not (a or b);
    layer5_outputs(1594) <= '0';
    layer5_outputs(1595) <= not a;
    layer5_outputs(1596) <= not a or b;
    layer5_outputs(1597) <= a;
    layer5_outputs(1598) <= not b;
    layer5_outputs(1599) <= a and not b;
    layer5_outputs(1600) <= not b;
    layer5_outputs(1601) <= a;
    layer5_outputs(1602) <= b and not a;
    layer5_outputs(1603) <= b;
    layer5_outputs(1604) <= a and not b;
    layer5_outputs(1605) <= b;
    layer5_outputs(1606) <= not (a and b);
    layer5_outputs(1607) <= not (a or b);
    layer5_outputs(1608) <= not a or b;
    layer5_outputs(1609) <= not a;
    layer5_outputs(1610) <= a xor b;
    layer5_outputs(1611) <= b and not a;
    layer5_outputs(1612) <= a and b;
    layer5_outputs(1613) <= b;
    layer5_outputs(1614) <= a and not b;
    layer5_outputs(1615) <= a or b;
    layer5_outputs(1616) <= a xor b;
    layer5_outputs(1617) <= a;
    layer5_outputs(1618) <= a;
    layer5_outputs(1619) <= not (a or b);
    layer5_outputs(1620) <= b;
    layer5_outputs(1621) <= a xor b;
    layer5_outputs(1622) <= not b;
    layer5_outputs(1623) <= a and not b;
    layer5_outputs(1624) <= not (a and b);
    layer5_outputs(1625) <= not b;
    layer5_outputs(1626) <= b;
    layer5_outputs(1627) <= '1';
    layer5_outputs(1628) <= b;
    layer5_outputs(1629) <= a;
    layer5_outputs(1630) <= a;
    layer5_outputs(1631) <= a;
    layer5_outputs(1632) <= not a or b;
    layer5_outputs(1633) <= not a or b;
    layer5_outputs(1634) <= a xor b;
    layer5_outputs(1635) <= a or b;
    layer5_outputs(1636) <= b and not a;
    layer5_outputs(1637) <= a;
    layer5_outputs(1638) <= not a;
    layer5_outputs(1639) <= a xor b;
    layer5_outputs(1640) <= a;
    layer5_outputs(1641) <= b;
    layer5_outputs(1642) <= not b;
    layer5_outputs(1643) <= not b;
    layer5_outputs(1644) <= b;
    layer5_outputs(1645) <= a and not b;
    layer5_outputs(1646) <= b;
    layer5_outputs(1647) <= not (a xor b);
    layer5_outputs(1648) <= b;
    layer5_outputs(1649) <= a;
    layer5_outputs(1650) <= not (a or b);
    layer5_outputs(1651) <= '0';
    layer5_outputs(1652) <= a xor b;
    layer5_outputs(1653) <= a and not b;
    layer5_outputs(1654) <= a;
    layer5_outputs(1655) <= not a;
    layer5_outputs(1656) <= a and b;
    layer5_outputs(1657) <= not (a or b);
    layer5_outputs(1658) <= not b;
    layer5_outputs(1659) <= b;
    layer5_outputs(1660) <= a xor b;
    layer5_outputs(1661) <= not (a xor b);
    layer5_outputs(1662) <= a xor b;
    layer5_outputs(1663) <= a or b;
    layer5_outputs(1664) <= a;
    layer5_outputs(1665) <= b and not a;
    layer5_outputs(1666) <= a xor b;
    layer5_outputs(1667) <= not (a xor b);
    layer5_outputs(1668) <= a;
    layer5_outputs(1669) <= b;
    layer5_outputs(1670) <= not (a xor b);
    layer5_outputs(1671) <= not b;
    layer5_outputs(1672) <= a;
    layer5_outputs(1673) <= not a;
    layer5_outputs(1674) <= a and b;
    layer5_outputs(1675) <= not (a or b);
    layer5_outputs(1676) <= a or b;
    layer5_outputs(1677) <= a and b;
    layer5_outputs(1678) <= not b or a;
    layer5_outputs(1679) <= a;
    layer5_outputs(1680) <= not b;
    layer5_outputs(1681) <= a and b;
    layer5_outputs(1682) <= a;
    layer5_outputs(1683) <= a and b;
    layer5_outputs(1684) <= b;
    layer5_outputs(1685) <= not b;
    layer5_outputs(1686) <= not (a xor b);
    layer5_outputs(1687) <= a xor b;
    layer5_outputs(1688) <= not b;
    layer5_outputs(1689) <= not (a and b);
    layer5_outputs(1690) <= b and not a;
    layer5_outputs(1691) <= not a;
    layer5_outputs(1692) <= not b or a;
    layer5_outputs(1693) <= a xor b;
    layer5_outputs(1694) <= not b;
    layer5_outputs(1695) <= not b or a;
    layer5_outputs(1696) <= not b;
    layer5_outputs(1697) <= a and not b;
    layer5_outputs(1698) <= a xor b;
    layer5_outputs(1699) <= a and not b;
    layer5_outputs(1700) <= not b;
    layer5_outputs(1701) <= a;
    layer5_outputs(1702) <= b;
    layer5_outputs(1703) <= a or b;
    layer5_outputs(1704) <= b;
    layer5_outputs(1705) <= not (a xor b);
    layer5_outputs(1706) <= a or b;
    layer5_outputs(1707) <= not (a or b);
    layer5_outputs(1708) <= not (a and b);
    layer5_outputs(1709) <= not a;
    layer5_outputs(1710) <= '0';
    layer5_outputs(1711) <= not b or a;
    layer5_outputs(1712) <= not b;
    layer5_outputs(1713) <= not (a xor b);
    layer5_outputs(1714) <= not b;
    layer5_outputs(1715) <= not a;
    layer5_outputs(1716) <= not (a xor b);
    layer5_outputs(1717) <= not a;
    layer5_outputs(1718) <= not (a xor b);
    layer5_outputs(1719) <= not b;
    layer5_outputs(1720) <= not (a xor b);
    layer5_outputs(1721) <= b;
    layer5_outputs(1722) <= b and not a;
    layer5_outputs(1723) <= not b or a;
    layer5_outputs(1724) <= not b;
    layer5_outputs(1725) <= not (a and b);
    layer5_outputs(1726) <= not a;
    layer5_outputs(1727) <= not a;
    layer5_outputs(1728) <= not a or b;
    layer5_outputs(1729) <= a or b;
    layer5_outputs(1730) <= a;
    layer5_outputs(1731) <= a and not b;
    layer5_outputs(1732) <= not b or a;
    layer5_outputs(1733) <= a;
    layer5_outputs(1734) <= b and not a;
    layer5_outputs(1735) <= not (a xor b);
    layer5_outputs(1736) <= a xor b;
    layer5_outputs(1737) <= not a;
    layer5_outputs(1738) <= b;
    layer5_outputs(1739) <= a and b;
    layer5_outputs(1740) <= a xor b;
    layer5_outputs(1741) <= not b or a;
    layer5_outputs(1742) <= not (a or b);
    layer5_outputs(1743) <= a and b;
    layer5_outputs(1744) <= a xor b;
    layer5_outputs(1745) <= a and not b;
    layer5_outputs(1746) <= not (a or b);
    layer5_outputs(1747) <= b;
    layer5_outputs(1748) <= a or b;
    layer5_outputs(1749) <= a and b;
    layer5_outputs(1750) <= not a;
    layer5_outputs(1751) <= a or b;
    layer5_outputs(1752) <= not (a or b);
    layer5_outputs(1753) <= not a;
    layer5_outputs(1754) <= not a;
    layer5_outputs(1755) <= not b or a;
    layer5_outputs(1756) <= not (a and b);
    layer5_outputs(1757) <= a;
    layer5_outputs(1758) <= a or b;
    layer5_outputs(1759) <= b;
    layer5_outputs(1760) <= not (a and b);
    layer5_outputs(1761) <= b;
    layer5_outputs(1762) <= not (a or b);
    layer5_outputs(1763) <= b and not a;
    layer5_outputs(1764) <= '0';
    layer5_outputs(1765) <= not b;
    layer5_outputs(1766) <= b;
    layer5_outputs(1767) <= not (a or b);
    layer5_outputs(1768) <= a xor b;
    layer5_outputs(1769) <= not b;
    layer5_outputs(1770) <= not (a xor b);
    layer5_outputs(1771) <= b;
    layer5_outputs(1772) <= a;
    layer5_outputs(1773) <= a and b;
    layer5_outputs(1774) <= not b;
    layer5_outputs(1775) <= a;
    layer5_outputs(1776) <= not (a xor b);
    layer5_outputs(1777) <= a or b;
    layer5_outputs(1778) <= '0';
    layer5_outputs(1779) <= a xor b;
    layer5_outputs(1780) <= a and not b;
    layer5_outputs(1781) <= not b;
    layer5_outputs(1782) <= not a or b;
    layer5_outputs(1783) <= not a;
    layer5_outputs(1784) <= not (a xor b);
    layer5_outputs(1785) <= b;
    layer5_outputs(1786) <= not (a and b);
    layer5_outputs(1787) <= not b or a;
    layer5_outputs(1788) <= not a;
    layer5_outputs(1789) <= not a;
    layer5_outputs(1790) <= b and not a;
    layer5_outputs(1791) <= not b;
    layer5_outputs(1792) <= a and not b;
    layer5_outputs(1793) <= not a;
    layer5_outputs(1794) <= not b;
    layer5_outputs(1795) <= b and not a;
    layer5_outputs(1796) <= not b;
    layer5_outputs(1797) <= not (a and b);
    layer5_outputs(1798) <= a and b;
    layer5_outputs(1799) <= not b;
    layer5_outputs(1800) <= a;
    layer5_outputs(1801) <= not a;
    layer5_outputs(1802) <= not a;
    layer5_outputs(1803) <= a;
    layer5_outputs(1804) <= not (a xor b);
    layer5_outputs(1805) <= not b;
    layer5_outputs(1806) <= not a;
    layer5_outputs(1807) <= not b;
    layer5_outputs(1808) <= not (a xor b);
    layer5_outputs(1809) <= a and not b;
    layer5_outputs(1810) <= not a or b;
    layer5_outputs(1811) <= not a;
    layer5_outputs(1812) <= not b;
    layer5_outputs(1813) <= a or b;
    layer5_outputs(1814) <= '0';
    layer5_outputs(1815) <= '1';
    layer5_outputs(1816) <= a;
    layer5_outputs(1817) <= a;
    layer5_outputs(1818) <= a or b;
    layer5_outputs(1819) <= not (a and b);
    layer5_outputs(1820) <= not a;
    layer5_outputs(1821) <= b;
    layer5_outputs(1822) <= a and b;
    layer5_outputs(1823) <= not a or b;
    layer5_outputs(1824) <= a xor b;
    layer5_outputs(1825) <= b;
    layer5_outputs(1826) <= not b;
    layer5_outputs(1827) <= a;
    layer5_outputs(1828) <= not b or a;
    layer5_outputs(1829) <= b and not a;
    layer5_outputs(1830) <= b;
    layer5_outputs(1831) <= not b;
    layer5_outputs(1832) <= not (a xor b);
    layer5_outputs(1833) <= b;
    layer5_outputs(1834) <= not (a xor b);
    layer5_outputs(1835) <= a;
    layer5_outputs(1836) <= a and b;
    layer5_outputs(1837) <= a or b;
    layer5_outputs(1838) <= b;
    layer5_outputs(1839) <= a and not b;
    layer5_outputs(1840) <= a xor b;
    layer5_outputs(1841) <= b;
    layer5_outputs(1842) <= a;
    layer5_outputs(1843) <= not a or b;
    layer5_outputs(1844) <= not b;
    layer5_outputs(1845) <= a and b;
    layer5_outputs(1846) <= not b or a;
    layer5_outputs(1847) <= a xor b;
    layer5_outputs(1848) <= not b or a;
    layer5_outputs(1849) <= not a;
    layer5_outputs(1850) <= not a;
    layer5_outputs(1851) <= not (a and b);
    layer5_outputs(1852) <= not (a or b);
    layer5_outputs(1853) <= a or b;
    layer5_outputs(1854) <= b and not a;
    layer5_outputs(1855) <= not (a or b);
    layer5_outputs(1856) <= not b;
    layer5_outputs(1857) <= a;
    layer5_outputs(1858) <= a;
    layer5_outputs(1859) <= '0';
    layer5_outputs(1860) <= b;
    layer5_outputs(1861) <= a;
    layer5_outputs(1862) <= a xor b;
    layer5_outputs(1863) <= b;
    layer5_outputs(1864) <= not b;
    layer5_outputs(1865) <= a;
    layer5_outputs(1866) <= a xor b;
    layer5_outputs(1867) <= a xor b;
    layer5_outputs(1868) <= a and not b;
    layer5_outputs(1869) <= not b or a;
    layer5_outputs(1870) <= b;
    layer5_outputs(1871) <= b;
    layer5_outputs(1872) <= '0';
    layer5_outputs(1873) <= not (a or b);
    layer5_outputs(1874) <= not (a or b);
    layer5_outputs(1875) <= '0';
    layer5_outputs(1876) <= b;
    layer5_outputs(1877) <= a;
    layer5_outputs(1878) <= b;
    layer5_outputs(1879) <= b;
    layer5_outputs(1880) <= b and not a;
    layer5_outputs(1881) <= not a;
    layer5_outputs(1882) <= not (a xor b);
    layer5_outputs(1883) <= not b;
    layer5_outputs(1884) <= not a;
    layer5_outputs(1885) <= a and not b;
    layer5_outputs(1886) <= a or b;
    layer5_outputs(1887) <= not (a or b);
    layer5_outputs(1888) <= not (a and b);
    layer5_outputs(1889) <= not (a and b);
    layer5_outputs(1890) <= not b or a;
    layer5_outputs(1891) <= not a or b;
    layer5_outputs(1892) <= not (a xor b);
    layer5_outputs(1893) <= not b;
    layer5_outputs(1894) <= a;
    layer5_outputs(1895) <= not (a xor b);
    layer5_outputs(1896) <= a;
    layer5_outputs(1897) <= not (a and b);
    layer5_outputs(1898) <= not (a or b);
    layer5_outputs(1899) <= a and not b;
    layer5_outputs(1900) <= a or b;
    layer5_outputs(1901) <= not a or b;
    layer5_outputs(1902) <= a or b;
    layer5_outputs(1903) <= a and b;
    layer5_outputs(1904) <= not a;
    layer5_outputs(1905) <= b;
    layer5_outputs(1906) <= a;
    layer5_outputs(1907) <= b and not a;
    layer5_outputs(1908) <= not b or a;
    layer5_outputs(1909) <= a;
    layer5_outputs(1910) <= not (a and b);
    layer5_outputs(1911) <= b;
    layer5_outputs(1912) <= a and b;
    layer5_outputs(1913) <= not b or a;
    layer5_outputs(1914) <= a and b;
    layer5_outputs(1915) <= not b or a;
    layer5_outputs(1916) <= not a or b;
    layer5_outputs(1917) <= not a;
    layer5_outputs(1918) <= a or b;
    layer5_outputs(1919) <= b;
    layer5_outputs(1920) <= a;
    layer5_outputs(1921) <= b and not a;
    layer5_outputs(1922) <= b;
    layer5_outputs(1923) <= b;
    layer5_outputs(1924) <= not b;
    layer5_outputs(1925) <= b and not a;
    layer5_outputs(1926) <= a or b;
    layer5_outputs(1927) <= not (a and b);
    layer5_outputs(1928) <= not a;
    layer5_outputs(1929) <= a xor b;
    layer5_outputs(1930) <= a;
    layer5_outputs(1931) <= not b;
    layer5_outputs(1932) <= not (a and b);
    layer5_outputs(1933) <= not a or b;
    layer5_outputs(1934) <= a and not b;
    layer5_outputs(1935) <= not (a xor b);
    layer5_outputs(1936) <= not (a or b);
    layer5_outputs(1937) <= a or b;
    layer5_outputs(1938) <= a or b;
    layer5_outputs(1939) <= not a or b;
    layer5_outputs(1940) <= b and not a;
    layer5_outputs(1941) <= a;
    layer5_outputs(1942) <= a or b;
    layer5_outputs(1943) <= not a or b;
    layer5_outputs(1944) <= not b or a;
    layer5_outputs(1945) <= not b;
    layer5_outputs(1946) <= not b or a;
    layer5_outputs(1947) <= not a;
    layer5_outputs(1948) <= a or b;
    layer5_outputs(1949) <= b;
    layer5_outputs(1950) <= not (a xor b);
    layer5_outputs(1951) <= not (a or b);
    layer5_outputs(1952) <= a or b;
    layer5_outputs(1953) <= b;
    layer5_outputs(1954) <= a xor b;
    layer5_outputs(1955) <= not a;
    layer5_outputs(1956) <= a xor b;
    layer5_outputs(1957) <= not b;
    layer5_outputs(1958) <= b;
    layer5_outputs(1959) <= b;
    layer5_outputs(1960) <= b;
    layer5_outputs(1961) <= not b or a;
    layer5_outputs(1962) <= not b or a;
    layer5_outputs(1963) <= not b;
    layer5_outputs(1964) <= a and not b;
    layer5_outputs(1965) <= not a;
    layer5_outputs(1966) <= a;
    layer5_outputs(1967) <= not a;
    layer5_outputs(1968) <= not (a or b);
    layer5_outputs(1969) <= a;
    layer5_outputs(1970) <= not (a or b);
    layer5_outputs(1971) <= a;
    layer5_outputs(1972) <= not b;
    layer5_outputs(1973) <= '0';
    layer5_outputs(1974) <= a and not b;
    layer5_outputs(1975) <= not (a xor b);
    layer5_outputs(1976) <= not a;
    layer5_outputs(1977) <= b and not a;
    layer5_outputs(1978) <= a;
    layer5_outputs(1979) <= a;
    layer5_outputs(1980) <= not (a and b);
    layer5_outputs(1981) <= not (a and b);
    layer5_outputs(1982) <= '0';
    layer5_outputs(1983) <= not (a xor b);
    layer5_outputs(1984) <= not a;
    layer5_outputs(1985) <= not a;
    layer5_outputs(1986) <= not b or a;
    layer5_outputs(1987) <= not (a and b);
    layer5_outputs(1988) <= b;
    layer5_outputs(1989) <= a;
    layer5_outputs(1990) <= not (a xor b);
    layer5_outputs(1991) <= a;
    layer5_outputs(1992) <= b;
    layer5_outputs(1993) <= not b or a;
    layer5_outputs(1994) <= not (a and b);
    layer5_outputs(1995) <= b and not a;
    layer5_outputs(1996) <= not (a xor b);
    layer5_outputs(1997) <= a or b;
    layer5_outputs(1998) <= a;
    layer5_outputs(1999) <= a;
    layer5_outputs(2000) <= a xor b;
    layer5_outputs(2001) <= not b;
    layer5_outputs(2002) <= a xor b;
    layer5_outputs(2003) <= not b;
    layer5_outputs(2004) <= a;
    layer5_outputs(2005) <= not a;
    layer5_outputs(2006) <= not b;
    layer5_outputs(2007) <= a;
    layer5_outputs(2008) <= not b;
    layer5_outputs(2009) <= not (a or b);
    layer5_outputs(2010) <= a and not b;
    layer5_outputs(2011) <= not a;
    layer5_outputs(2012) <= not (a or b);
    layer5_outputs(2013) <= not (a or b);
    layer5_outputs(2014) <= not a or b;
    layer5_outputs(2015) <= not b;
    layer5_outputs(2016) <= a and not b;
    layer5_outputs(2017) <= not b;
    layer5_outputs(2018) <= not b;
    layer5_outputs(2019) <= b and not a;
    layer5_outputs(2020) <= not b or a;
    layer5_outputs(2021) <= a and not b;
    layer5_outputs(2022) <= a xor b;
    layer5_outputs(2023) <= a or b;
    layer5_outputs(2024) <= not b;
    layer5_outputs(2025) <= b;
    layer5_outputs(2026) <= '0';
    layer5_outputs(2027) <= not (a and b);
    layer5_outputs(2028) <= a;
    layer5_outputs(2029) <= not a;
    layer5_outputs(2030) <= a xor b;
    layer5_outputs(2031) <= not a;
    layer5_outputs(2032) <= not b;
    layer5_outputs(2033) <= a;
    layer5_outputs(2034) <= a;
    layer5_outputs(2035) <= a;
    layer5_outputs(2036) <= not (a xor b);
    layer5_outputs(2037) <= not b;
    layer5_outputs(2038) <= not b;
    layer5_outputs(2039) <= b;
    layer5_outputs(2040) <= not a;
    layer5_outputs(2041) <= not a;
    layer5_outputs(2042) <= not (a or b);
    layer5_outputs(2043) <= not b;
    layer5_outputs(2044) <= not a;
    layer5_outputs(2045) <= b;
    layer5_outputs(2046) <= not b;
    layer5_outputs(2047) <= b;
    layer5_outputs(2048) <= a;
    layer5_outputs(2049) <= not (a xor b);
    layer5_outputs(2050) <= a;
    layer5_outputs(2051) <= not a or b;
    layer5_outputs(2052) <= b and not a;
    layer5_outputs(2053) <= not a;
    layer5_outputs(2054) <= b;
    layer5_outputs(2055) <= a or b;
    layer5_outputs(2056) <= a or b;
    layer5_outputs(2057) <= b and not a;
    layer5_outputs(2058) <= a xor b;
    layer5_outputs(2059) <= not a;
    layer5_outputs(2060) <= not a;
    layer5_outputs(2061) <= not a;
    layer5_outputs(2062) <= not (a xor b);
    layer5_outputs(2063) <= a;
    layer5_outputs(2064) <= a;
    layer5_outputs(2065) <= a;
    layer5_outputs(2066) <= a;
    layer5_outputs(2067) <= b;
    layer5_outputs(2068) <= a;
    layer5_outputs(2069) <= not b;
    layer5_outputs(2070) <= a;
    layer5_outputs(2071) <= b;
    layer5_outputs(2072) <= a and b;
    layer5_outputs(2073) <= not b or a;
    layer5_outputs(2074) <= not b;
    layer5_outputs(2075) <= not a;
    layer5_outputs(2076) <= b;
    layer5_outputs(2077) <= not a;
    layer5_outputs(2078) <= b and not a;
    layer5_outputs(2079) <= b;
    layer5_outputs(2080) <= b;
    layer5_outputs(2081) <= a or b;
    layer5_outputs(2082) <= not b;
    layer5_outputs(2083) <= b;
    layer5_outputs(2084) <= not (a and b);
    layer5_outputs(2085) <= a xor b;
    layer5_outputs(2086) <= a or b;
    layer5_outputs(2087) <= not a or b;
    layer5_outputs(2088) <= a xor b;
    layer5_outputs(2089) <= not b;
    layer5_outputs(2090) <= not a or b;
    layer5_outputs(2091) <= not a;
    layer5_outputs(2092) <= a or b;
    layer5_outputs(2093) <= not b;
    layer5_outputs(2094) <= a;
    layer5_outputs(2095) <= not (a xor b);
    layer5_outputs(2096) <= b;
    layer5_outputs(2097) <= a and b;
    layer5_outputs(2098) <= a;
    layer5_outputs(2099) <= a xor b;
    layer5_outputs(2100) <= not (a or b);
    layer5_outputs(2101) <= not (a xor b);
    layer5_outputs(2102) <= b;
    layer5_outputs(2103) <= a and b;
    layer5_outputs(2104) <= not b or a;
    layer5_outputs(2105) <= not b;
    layer5_outputs(2106) <= a;
    layer5_outputs(2107) <= a xor b;
    layer5_outputs(2108) <= b;
    layer5_outputs(2109) <= not b;
    layer5_outputs(2110) <= not (a xor b);
    layer5_outputs(2111) <= b;
    layer5_outputs(2112) <= b;
    layer5_outputs(2113) <= a and b;
    layer5_outputs(2114) <= a;
    layer5_outputs(2115) <= a or b;
    layer5_outputs(2116) <= a or b;
    layer5_outputs(2117) <= a;
    layer5_outputs(2118) <= not b;
    layer5_outputs(2119) <= b and not a;
    layer5_outputs(2120) <= a;
    layer5_outputs(2121) <= a and not b;
    layer5_outputs(2122) <= a;
    layer5_outputs(2123) <= not b or a;
    layer5_outputs(2124) <= not b;
    layer5_outputs(2125) <= b;
    layer5_outputs(2126) <= a xor b;
    layer5_outputs(2127) <= a and not b;
    layer5_outputs(2128) <= a and b;
    layer5_outputs(2129) <= b;
    layer5_outputs(2130) <= a and not b;
    layer5_outputs(2131) <= not a;
    layer5_outputs(2132) <= a;
    layer5_outputs(2133) <= a and b;
    layer5_outputs(2134) <= not (a and b);
    layer5_outputs(2135) <= not a or b;
    layer5_outputs(2136) <= not b;
    layer5_outputs(2137) <= not a or b;
    layer5_outputs(2138) <= not b;
    layer5_outputs(2139) <= a or b;
    layer5_outputs(2140) <= not b;
    layer5_outputs(2141) <= not (a or b);
    layer5_outputs(2142) <= not a;
    layer5_outputs(2143) <= not a;
    layer5_outputs(2144) <= not a or b;
    layer5_outputs(2145) <= b;
    layer5_outputs(2146) <= not (a or b);
    layer5_outputs(2147) <= not a or b;
    layer5_outputs(2148) <= a;
    layer5_outputs(2149) <= not b;
    layer5_outputs(2150) <= a or b;
    layer5_outputs(2151) <= not a or b;
    layer5_outputs(2152) <= not a;
    layer5_outputs(2153) <= not (a or b);
    layer5_outputs(2154) <= b;
    layer5_outputs(2155) <= a or b;
    layer5_outputs(2156) <= not b;
    layer5_outputs(2157) <= not a;
    layer5_outputs(2158) <= not a;
    layer5_outputs(2159) <= a;
    layer5_outputs(2160) <= not b;
    layer5_outputs(2161) <= b;
    layer5_outputs(2162) <= b;
    layer5_outputs(2163) <= not (a and b);
    layer5_outputs(2164) <= a and b;
    layer5_outputs(2165) <= a or b;
    layer5_outputs(2166) <= not (a and b);
    layer5_outputs(2167) <= a and not b;
    layer5_outputs(2168) <= a and not b;
    layer5_outputs(2169) <= a and not b;
    layer5_outputs(2170) <= not b;
    layer5_outputs(2171) <= a xor b;
    layer5_outputs(2172) <= '0';
    layer5_outputs(2173) <= not b or a;
    layer5_outputs(2174) <= a xor b;
    layer5_outputs(2175) <= not a;
    layer5_outputs(2176) <= not b;
    layer5_outputs(2177) <= not b or a;
    layer5_outputs(2178) <= not b;
    layer5_outputs(2179) <= b;
    layer5_outputs(2180) <= a;
    layer5_outputs(2181) <= not a or b;
    layer5_outputs(2182) <= a or b;
    layer5_outputs(2183) <= not b;
    layer5_outputs(2184) <= a;
    layer5_outputs(2185) <= b;
    layer5_outputs(2186) <= a or b;
    layer5_outputs(2187) <= a and b;
    layer5_outputs(2188) <= a;
    layer5_outputs(2189) <= a or b;
    layer5_outputs(2190) <= a xor b;
    layer5_outputs(2191) <= b;
    layer5_outputs(2192) <= not a;
    layer5_outputs(2193) <= a;
    layer5_outputs(2194) <= a xor b;
    layer5_outputs(2195) <= not (a xor b);
    layer5_outputs(2196) <= not (a and b);
    layer5_outputs(2197) <= not (a and b);
    layer5_outputs(2198) <= not b;
    layer5_outputs(2199) <= not b;
    layer5_outputs(2200) <= a;
    layer5_outputs(2201) <= a xor b;
    layer5_outputs(2202) <= '1';
    layer5_outputs(2203) <= not b;
    layer5_outputs(2204) <= b;
    layer5_outputs(2205) <= b and not a;
    layer5_outputs(2206) <= not b;
    layer5_outputs(2207) <= not (a or b);
    layer5_outputs(2208) <= '0';
    layer5_outputs(2209) <= not b or a;
    layer5_outputs(2210) <= a and b;
    layer5_outputs(2211) <= not (a xor b);
    layer5_outputs(2212) <= not a or b;
    layer5_outputs(2213) <= a xor b;
    layer5_outputs(2214) <= not (a and b);
    layer5_outputs(2215) <= not a or b;
    layer5_outputs(2216) <= a or b;
    layer5_outputs(2217) <= not a;
    layer5_outputs(2218) <= a xor b;
    layer5_outputs(2219) <= not a;
    layer5_outputs(2220) <= not b or a;
    layer5_outputs(2221) <= not a or b;
    layer5_outputs(2222) <= b;
    layer5_outputs(2223) <= b;
    layer5_outputs(2224) <= b;
    layer5_outputs(2225) <= b and not a;
    layer5_outputs(2226) <= a or b;
    layer5_outputs(2227) <= a xor b;
    layer5_outputs(2228) <= b and not a;
    layer5_outputs(2229) <= b;
    layer5_outputs(2230) <= a;
    layer5_outputs(2231) <= a or b;
    layer5_outputs(2232) <= not (a or b);
    layer5_outputs(2233) <= a and not b;
    layer5_outputs(2234) <= not (a xor b);
    layer5_outputs(2235) <= b and not a;
    layer5_outputs(2236) <= a and not b;
    layer5_outputs(2237) <= not b;
    layer5_outputs(2238) <= not b;
    layer5_outputs(2239) <= a xor b;
    layer5_outputs(2240) <= not a;
    layer5_outputs(2241) <= b;
    layer5_outputs(2242) <= b and not a;
    layer5_outputs(2243) <= not (a xor b);
    layer5_outputs(2244) <= not (a and b);
    layer5_outputs(2245) <= a;
    layer5_outputs(2246) <= not b or a;
    layer5_outputs(2247) <= not a;
    layer5_outputs(2248) <= a;
    layer5_outputs(2249) <= b and not a;
    layer5_outputs(2250) <= a and b;
    layer5_outputs(2251) <= not (a and b);
    layer5_outputs(2252) <= not a;
    layer5_outputs(2253) <= not (a or b);
    layer5_outputs(2254) <= not b;
    layer5_outputs(2255) <= a;
    layer5_outputs(2256) <= not (a xor b);
    layer5_outputs(2257) <= not b;
    layer5_outputs(2258) <= a;
    layer5_outputs(2259) <= not (a and b);
    layer5_outputs(2260) <= b and not a;
    layer5_outputs(2261) <= b;
    layer5_outputs(2262) <= b;
    layer5_outputs(2263) <= a and b;
    layer5_outputs(2264) <= not b;
    layer5_outputs(2265) <= a and not b;
    layer5_outputs(2266) <= not b;
    layer5_outputs(2267) <= a and b;
    layer5_outputs(2268) <= a;
    layer5_outputs(2269) <= a;
    layer5_outputs(2270) <= '1';
    layer5_outputs(2271) <= not b;
    layer5_outputs(2272) <= a;
    layer5_outputs(2273) <= not (a and b);
    layer5_outputs(2274) <= not (a or b);
    layer5_outputs(2275) <= '1';
    layer5_outputs(2276) <= not a or b;
    layer5_outputs(2277) <= not b or a;
    layer5_outputs(2278) <= not (a and b);
    layer5_outputs(2279) <= not a;
    layer5_outputs(2280) <= not (a and b);
    layer5_outputs(2281) <= a and b;
    layer5_outputs(2282) <= not b;
    layer5_outputs(2283) <= b;
    layer5_outputs(2284) <= not b;
    layer5_outputs(2285) <= a;
    layer5_outputs(2286) <= '1';
    layer5_outputs(2287) <= '0';
    layer5_outputs(2288) <= a;
    layer5_outputs(2289) <= b and not a;
    layer5_outputs(2290) <= not b;
    layer5_outputs(2291) <= b;
    layer5_outputs(2292) <= not a;
    layer5_outputs(2293) <= not (a xor b);
    layer5_outputs(2294) <= not b or a;
    layer5_outputs(2295) <= not b;
    layer5_outputs(2296) <= b;
    layer5_outputs(2297) <= a;
    layer5_outputs(2298) <= b;
    layer5_outputs(2299) <= not a or b;
    layer5_outputs(2300) <= not b or a;
    layer5_outputs(2301) <= not b or a;
    layer5_outputs(2302) <= not b;
    layer5_outputs(2303) <= b;
    layer5_outputs(2304) <= a;
    layer5_outputs(2305) <= not a;
    layer5_outputs(2306) <= b and not a;
    layer5_outputs(2307) <= not (a and b);
    layer5_outputs(2308) <= a;
    layer5_outputs(2309) <= not (a or b);
    layer5_outputs(2310) <= b;
    layer5_outputs(2311) <= a;
    layer5_outputs(2312) <= not (a or b);
    layer5_outputs(2313) <= not b or a;
    layer5_outputs(2314) <= a xor b;
    layer5_outputs(2315) <= b and not a;
    layer5_outputs(2316) <= a and b;
    layer5_outputs(2317) <= a and b;
    layer5_outputs(2318) <= not a;
    layer5_outputs(2319) <= a and not b;
    layer5_outputs(2320) <= not (a xor b);
    layer5_outputs(2321) <= not a;
    layer5_outputs(2322) <= a and not b;
    layer5_outputs(2323) <= not b or a;
    layer5_outputs(2324) <= b and not a;
    layer5_outputs(2325) <= not (a or b);
    layer5_outputs(2326) <= not a;
    layer5_outputs(2327) <= a xor b;
    layer5_outputs(2328) <= a and not b;
    layer5_outputs(2329) <= not b;
    layer5_outputs(2330) <= b and not a;
    layer5_outputs(2331) <= a and b;
    layer5_outputs(2332) <= not (a and b);
    layer5_outputs(2333) <= a or b;
    layer5_outputs(2334) <= not a or b;
    layer5_outputs(2335) <= not b or a;
    layer5_outputs(2336) <= '0';
    layer5_outputs(2337) <= a xor b;
    layer5_outputs(2338) <= not (a xor b);
    layer5_outputs(2339) <= not a or b;
    layer5_outputs(2340) <= not b;
    layer5_outputs(2341) <= b;
    layer5_outputs(2342) <= not b or a;
    layer5_outputs(2343) <= a;
    layer5_outputs(2344) <= a;
    layer5_outputs(2345) <= not a;
    layer5_outputs(2346) <= b and not a;
    layer5_outputs(2347) <= not a;
    layer5_outputs(2348) <= not a;
    layer5_outputs(2349) <= a;
    layer5_outputs(2350) <= not (a and b);
    layer5_outputs(2351) <= a and b;
    layer5_outputs(2352) <= b;
    layer5_outputs(2353) <= not b;
    layer5_outputs(2354) <= b;
    layer5_outputs(2355) <= b;
    layer5_outputs(2356) <= not a;
    layer5_outputs(2357) <= a;
    layer5_outputs(2358) <= a;
    layer5_outputs(2359) <= b;
    layer5_outputs(2360) <= b and not a;
    layer5_outputs(2361) <= b and not a;
    layer5_outputs(2362) <= b and not a;
    layer5_outputs(2363) <= not b;
    layer5_outputs(2364) <= not (a and b);
    layer5_outputs(2365) <= '0';
    layer5_outputs(2366) <= a xor b;
    layer5_outputs(2367) <= not a;
    layer5_outputs(2368) <= a xor b;
    layer5_outputs(2369) <= a;
    layer5_outputs(2370) <= a and not b;
    layer5_outputs(2371) <= '1';
    layer5_outputs(2372) <= not a;
    layer5_outputs(2373) <= not a;
    layer5_outputs(2374) <= not b;
    layer5_outputs(2375) <= not b;
    layer5_outputs(2376) <= not a;
    layer5_outputs(2377) <= b;
    layer5_outputs(2378) <= not b;
    layer5_outputs(2379) <= not a;
    layer5_outputs(2380) <= not b;
    layer5_outputs(2381) <= b and not a;
    layer5_outputs(2382) <= not b;
    layer5_outputs(2383) <= not (a or b);
    layer5_outputs(2384) <= b;
    layer5_outputs(2385) <= b;
    layer5_outputs(2386) <= a xor b;
    layer5_outputs(2387) <= not a or b;
    layer5_outputs(2388) <= not (a or b);
    layer5_outputs(2389) <= a;
    layer5_outputs(2390) <= b;
    layer5_outputs(2391) <= a or b;
    layer5_outputs(2392) <= not b;
    layer5_outputs(2393) <= not (a or b);
    layer5_outputs(2394) <= not (a xor b);
    layer5_outputs(2395) <= not b;
    layer5_outputs(2396) <= '0';
    layer5_outputs(2397) <= not (a and b);
    layer5_outputs(2398) <= not b;
    layer5_outputs(2399) <= a or b;
    layer5_outputs(2400) <= b;
    layer5_outputs(2401) <= a;
    layer5_outputs(2402) <= b;
    layer5_outputs(2403) <= a and b;
    layer5_outputs(2404) <= a;
    layer5_outputs(2405) <= a and not b;
    layer5_outputs(2406) <= not b;
    layer5_outputs(2407) <= not (a xor b);
    layer5_outputs(2408) <= b;
    layer5_outputs(2409) <= not a or b;
    layer5_outputs(2410) <= not b;
    layer5_outputs(2411) <= not b or a;
    layer5_outputs(2412) <= not (a and b);
    layer5_outputs(2413) <= b;
    layer5_outputs(2414) <= b;
    layer5_outputs(2415) <= a;
    layer5_outputs(2416) <= not a or b;
    layer5_outputs(2417) <= not b or a;
    layer5_outputs(2418) <= b and not a;
    layer5_outputs(2419) <= a xor b;
    layer5_outputs(2420) <= not b or a;
    layer5_outputs(2421) <= not b;
    layer5_outputs(2422) <= not (a and b);
    layer5_outputs(2423) <= not b;
    layer5_outputs(2424) <= b and not a;
    layer5_outputs(2425) <= a or b;
    layer5_outputs(2426) <= b;
    layer5_outputs(2427) <= not (a or b);
    layer5_outputs(2428) <= not b or a;
    layer5_outputs(2429) <= a;
    layer5_outputs(2430) <= a and b;
    layer5_outputs(2431) <= not b;
    layer5_outputs(2432) <= a and not b;
    layer5_outputs(2433) <= not a;
    layer5_outputs(2434) <= a and not b;
    layer5_outputs(2435) <= not (a or b);
    layer5_outputs(2436) <= a xor b;
    layer5_outputs(2437) <= a and not b;
    layer5_outputs(2438) <= a;
    layer5_outputs(2439) <= not a or b;
    layer5_outputs(2440) <= a and b;
    layer5_outputs(2441) <= b;
    layer5_outputs(2442) <= a or b;
    layer5_outputs(2443) <= b;
    layer5_outputs(2444) <= a;
    layer5_outputs(2445) <= b;
    layer5_outputs(2446) <= not a;
    layer5_outputs(2447) <= a and not b;
    layer5_outputs(2448) <= not a;
    layer5_outputs(2449) <= not b;
    layer5_outputs(2450) <= not a or b;
    layer5_outputs(2451) <= not a or b;
    layer5_outputs(2452) <= a and not b;
    layer5_outputs(2453) <= not (a and b);
    layer5_outputs(2454) <= not a;
    layer5_outputs(2455) <= b and not a;
    layer5_outputs(2456) <= b and not a;
    layer5_outputs(2457) <= a or b;
    layer5_outputs(2458) <= b;
    layer5_outputs(2459) <= not b;
    layer5_outputs(2460) <= b;
    layer5_outputs(2461) <= a;
    layer5_outputs(2462) <= b and not a;
    layer5_outputs(2463) <= not (a xor b);
    layer5_outputs(2464) <= a;
    layer5_outputs(2465) <= not (a xor b);
    layer5_outputs(2466) <= a xor b;
    layer5_outputs(2467) <= not (a or b);
    layer5_outputs(2468) <= not a;
    layer5_outputs(2469) <= not b or a;
    layer5_outputs(2470) <= not b or a;
    layer5_outputs(2471) <= not a;
    layer5_outputs(2472) <= not b;
    layer5_outputs(2473) <= not b;
    layer5_outputs(2474) <= not b;
    layer5_outputs(2475) <= not (a or b);
    layer5_outputs(2476) <= not (a xor b);
    layer5_outputs(2477) <= not a;
    layer5_outputs(2478) <= not (a and b);
    layer5_outputs(2479) <= a or b;
    layer5_outputs(2480) <= a;
    layer5_outputs(2481) <= not (a or b);
    layer5_outputs(2482) <= not b;
    layer5_outputs(2483) <= a;
    layer5_outputs(2484) <= b;
    layer5_outputs(2485) <= not b;
    layer5_outputs(2486) <= not (a or b);
    layer5_outputs(2487) <= not a;
    layer5_outputs(2488) <= a and b;
    layer5_outputs(2489) <= a and b;
    layer5_outputs(2490) <= a;
    layer5_outputs(2491) <= not a;
    layer5_outputs(2492) <= not b;
    layer5_outputs(2493) <= not a;
    layer5_outputs(2494) <= not b;
    layer5_outputs(2495) <= a or b;
    layer5_outputs(2496) <= not a or b;
    layer5_outputs(2497) <= a xor b;
    layer5_outputs(2498) <= not b;
    layer5_outputs(2499) <= not b;
    layer5_outputs(2500) <= not (a or b);
    layer5_outputs(2501) <= not a;
    layer5_outputs(2502) <= a or b;
    layer5_outputs(2503) <= not (a xor b);
    layer5_outputs(2504) <= '0';
    layer5_outputs(2505) <= '1';
    layer5_outputs(2506) <= not a;
    layer5_outputs(2507) <= not a or b;
    layer5_outputs(2508) <= not b;
    layer5_outputs(2509) <= not b;
    layer5_outputs(2510) <= not a;
    layer5_outputs(2511) <= a or b;
    layer5_outputs(2512) <= not (a or b);
    layer5_outputs(2513) <= b;
    layer5_outputs(2514) <= not a;
    layer5_outputs(2515) <= a or b;
    layer5_outputs(2516) <= not a or b;
    layer5_outputs(2517) <= a xor b;
    layer5_outputs(2518) <= not b;
    layer5_outputs(2519) <= a;
    layer5_outputs(2520) <= not b;
    layer5_outputs(2521) <= not a;
    layer5_outputs(2522) <= not b or a;
    layer5_outputs(2523) <= not (a or b);
    layer5_outputs(2524) <= a xor b;
    layer5_outputs(2525) <= a or b;
    layer5_outputs(2526) <= not a or b;
    layer5_outputs(2527) <= not b;
    layer5_outputs(2528) <= not (a xor b);
    layer5_outputs(2529) <= a;
    layer5_outputs(2530) <= not (a or b);
    layer5_outputs(2531) <= b;
    layer5_outputs(2532) <= a and b;
    layer5_outputs(2533) <= b and not a;
    layer5_outputs(2534) <= not (a xor b);
    layer5_outputs(2535) <= not (a xor b);
    layer5_outputs(2536) <= not (a xor b);
    layer5_outputs(2537) <= a;
    layer5_outputs(2538) <= b;
    layer5_outputs(2539) <= a xor b;
    layer5_outputs(2540) <= not (a or b);
    layer5_outputs(2541) <= not (a xor b);
    layer5_outputs(2542) <= not a;
    layer5_outputs(2543) <= not b;
    layer5_outputs(2544) <= not (a or b);
    layer5_outputs(2545) <= a and not b;
    layer5_outputs(2546) <= not (a or b);
    layer5_outputs(2547) <= a xor b;
    layer5_outputs(2548) <= a and not b;
    layer5_outputs(2549) <= a and b;
    layer5_outputs(2550) <= b and not a;
    layer5_outputs(2551) <= not (a or b);
    layer5_outputs(2552) <= a or b;
    layer5_outputs(2553) <= '0';
    layer5_outputs(2554) <= not a or b;
    layer5_outputs(2555) <= '1';
    layer5_outputs(2556) <= not b;
    layer5_outputs(2557) <= not a;
    layer5_outputs(2558) <= not b or a;
    layer5_outputs(2559) <= a;
    layer5_outputs(2560) <= not a;
    layer5_outputs(2561) <= b;
    layer5_outputs(2562) <= a xor b;
    layer5_outputs(2563) <= b and not a;
    layer5_outputs(2564) <= a;
    layer5_outputs(2565) <= b;
    layer5_outputs(2566) <= not (a xor b);
    layer5_outputs(2567) <= not b or a;
    layer5_outputs(2568) <= b;
    layer5_outputs(2569) <= a or b;
    layer5_outputs(2570) <= not b or a;
    layer5_outputs(2571) <= a and b;
    layer5_outputs(2572) <= not a;
    layer5_outputs(2573) <= b;
    layer5_outputs(2574) <= b;
    layer5_outputs(2575) <= b and not a;
    layer5_outputs(2576) <= not (a or b);
    layer5_outputs(2577) <= not a;
    layer5_outputs(2578) <= b and not a;
    layer5_outputs(2579) <= not b;
    layer5_outputs(2580) <= not a or b;
    layer5_outputs(2581) <= '0';
    layer5_outputs(2582) <= a xor b;
    layer5_outputs(2583) <= not a;
    layer5_outputs(2584) <= not a or b;
    layer5_outputs(2585) <= not b;
    layer5_outputs(2586) <= a and b;
    layer5_outputs(2587) <= b;
    layer5_outputs(2588) <= '0';
    layer5_outputs(2589) <= b;
    layer5_outputs(2590) <= b;
    layer5_outputs(2591) <= a and b;
    layer5_outputs(2592) <= a;
    layer5_outputs(2593) <= not b;
    layer5_outputs(2594) <= not b;
    layer5_outputs(2595) <= b;
    layer5_outputs(2596) <= a;
    layer5_outputs(2597) <= a;
    layer5_outputs(2598) <= a;
    layer5_outputs(2599) <= a or b;
    layer5_outputs(2600) <= not (a and b);
    layer5_outputs(2601) <= a;
    layer5_outputs(2602) <= not b;
    layer5_outputs(2603) <= a and not b;
    layer5_outputs(2604) <= a and not b;
    layer5_outputs(2605) <= not b;
    layer5_outputs(2606) <= not (a xor b);
    layer5_outputs(2607) <= not b;
    layer5_outputs(2608) <= not a or b;
    layer5_outputs(2609) <= a;
    layer5_outputs(2610) <= a and not b;
    layer5_outputs(2611) <= b;
    layer5_outputs(2612) <= not b or a;
    layer5_outputs(2613) <= not b;
    layer5_outputs(2614) <= not (a and b);
    layer5_outputs(2615) <= not b;
    layer5_outputs(2616) <= not a or b;
    layer5_outputs(2617) <= not (a or b);
    layer5_outputs(2618) <= not b;
    layer5_outputs(2619) <= not a;
    layer5_outputs(2620) <= not a or b;
    layer5_outputs(2621) <= b;
    layer5_outputs(2622) <= not a;
    layer5_outputs(2623) <= b;
    layer5_outputs(2624) <= b;
    layer5_outputs(2625) <= a and not b;
    layer5_outputs(2626) <= not a or b;
    layer5_outputs(2627) <= not b or a;
    layer5_outputs(2628) <= not a;
    layer5_outputs(2629) <= a or b;
    layer5_outputs(2630) <= b;
    layer5_outputs(2631) <= not b;
    layer5_outputs(2632) <= not b or a;
    layer5_outputs(2633) <= b and not a;
    layer5_outputs(2634) <= '1';
    layer5_outputs(2635) <= a and b;
    layer5_outputs(2636) <= a or b;
    layer5_outputs(2637) <= a;
    layer5_outputs(2638) <= not a;
    layer5_outputs(2639) <= b;
    layer5_outputs(2640) <= a or b;
    layer5_outputs(2641) <= a;
    layer5_outputs(2642) <= a;
    layer5_outputs(2643) <= a xor b;
    layer5_outputs(2644) <= b;
    layer5_outputs(2645) <= not a;
    layer5_outputs(2646) <= a xor b;
    layer5_outputs(2647) <= a;
    layer5_outputs(2648) <= not a or b;
    layer5_outputs(2649) <= not a;
    layer5_outputs(2650) <= a xor b;
    layer5_outputs(2651) <= a;
    layer5_outputs(2652) <= not a;
    layer5_outputs(2653) <= not (a and b);
    layer5_outputs(2654) <= a or b;
    layer5_outputs(2655) <= b;
    layer5_outputs(2656) <= not (a xor b);
    layer5_outputs(2657) <= a xor b;
    layer5_outputs(2658) <= not b;
    layer5_outputs(2659) <= not (a and b);
    layer5_outputs(2660) <= a or b;
    layer5_outputs(2661) <= b;
    layer5_outputs(2662) <= a or b;
    layer5_outputs(2663) <= not (a or b);
    layer5_outputs(2664) <= not (a or b);
    layer5_outputs(2665) <= a;
    layer5_outputs(2666) <= not (a and b);
    layer5_outputs(2667) <= a or b;
    layer5_outputs(2668) <= b;
    layer5_outputs(2669) <= b and not a;
    layer5_outputs(2670) <= b;
    layer5_outputs(2671) <= not b;
    layer5_outputs(2672) <= b and not a;
    layer5_outputs(2673) <= a;
    layer5_outputs(2674) <= not (a xor b);
    layer5_outputs(2675) <= b;
    layer5_outputs(2676) <= a and b;
    layer5_outputs(2677) <= not (a and b);
    layer5_outputs(2678) <= not a;
    layer5_outputs(2679) <= b;
    layer5_outputs(2680) <= not (a or b);
    layer5_outputs(2681) <= a or b;
    layer5_outputs(2682) <= not b or a;
    layer5_outputs(2683) <= not (a and b);
    layer5_outputs(2684) <= not (a and b);
    layer5_outputs(2685) <= a and not b;
    layer5_outputs(2686) <= a;
    layer5_outputs(2687) <= not a;
    layer5_outputs(2688) <= not a or b;
    layer5_outputs(2689) <= not (a or b);
    layer5_outputs(2690) <= a;
    layer5_outputs(2691) <= b;
    layer5_outputs(2692) <= not (a and b);
    layer5_outputs(2693) <= a;
    layer5_outputs(2694) <= not (a and b);
    layer5_outputs(2695) <= not (a or b);
    layer5_outputs(2696) <= a and not b;
    layer5_outputs(2697) <= a xor b;
    layer5_outputs(2698) <= a xor b;
    layer5_outputs(2699) <= not a;
    layer5_outputs(2700) <= b;
    layer5_outputs(2701) <= a or b;
    layer5_outputs(2702) <= not b or a;
    layer5_outputs(2703) <= a;
    layer5_outputs(2704) <= not (a and b);
    layer5_outputs(2705) <= a xor b;
    layer5_outputs(2706) <= not b;
    layer5_outputs(2707) <= a and b;
    layer5_outputs(2708) <= b;
    layer5_outputs(2709) <= not (a or b);
    layer5_outputs(2710) <= b;
    layer5_outputs(2711) <= not b or a;
    layer5_outputs(2712) <= not a;
    layer5_outputs(2713) <= b;
    layer5_outputs(2714) <= not b or a;
    layer5_outputs(2715) <= a and b;
    layer5_outputs(2716) <= a xor b;
    layer5_outputs(2717) <= a or b;
    layer5_outputs(2718) <= a;
    layer5_outputs(2719) <= a and b;
    layer5_outputs(2720) <= a xor b;
    layer5_outputs(2721) <= '0';
    layer5_outputs(2722) <= not b;
    layer5_outputs(2723) <= b;
    layer5_outputs(2724) <= a;
    layer5_outputs(2725) <= a or b;
    layer5_outputs(2726) <= a and b;
    layer5_outputs(2727) <= a or b;
    layer5_outputs(2728) <= a xor b;
    layer5_outputs(2729) <= not b;
    layer5_outputs(2730) <= a and b;
    layer5_outputs(2731) <= a and not b;
    layer5_outputs(2732) <= not b;
    layer5_outputs(2733) <= not (a or b);
    layer5_outputs(2734) <= b;
    layer5_outputs(2735) <= not b or a;
    layer5_outputs(2736) <= not (a and b);
    layer5_outputs(2737) <= a;
    layer5_outputs(2738) <= a or b;
    layer5_outputs(2739) <= a xor b;
    layer5_outputs(2740) <= not b or a;
    layer5_outputs(2741) <= not a;
    layer5_outputs(2742) <= not (a and b);
    layer5_outputs(2743) <= a;
    layer5_outputs(2744) <= not a;
    layer5_outputs(2745) <= a or b;
    layer5_outputs(2746) <= b;
    layer5_outputs(2747) <= not b;
    layer5_outputs(2748) <= b;
    layer5_outputs(2749) <= a;
    layer5_outputs(2750) <= not (a and b);
    layer5_outputs(2751) <= not (a xor b);
    layer5_outputs(2752) <= a;
    layer5_outputs(2753) <= not (a xor b);
    layer5_outputs(2754) <= a xor b;
    layer5_outputs(2755) <= b;
    layer5_outputs(2756) <= a and not b;
    layer5_outputs(2757) <= b;
    layer5_outputs(2758) <= b;
    layer5_outputs(2759) <= not b;
    layer5_outputs(2760) <= b;
    layer5_outputs(2761) <= not a;
    layer5_outputs(2762) <= not (a xor b);
    layer5_outputs(2763) <= b;
    layer5_outputs(2764) <= a and not b;
    layer5_outputs(2765) <= not (a and b);
    layer5_outputs(2766) <= not (a and b);
    layer5_outputs(2767) <= a and b;
    layer5_outputs(2768) <= a and not b;
    layer5_outputs(2769) <= not a or b;
    layer5_outputs(2770) <= b and not a;
    layer5_outputs(2771) <= not a;
    layer5_outputs(2772) <= not a or b;
    layer5_outputs(2773) <= not b or a;
    layer5_outputs(2774) <= not a;
    layer5_outputs(2775) <= a and not b;
    layer5_outputs(2776) <= b;
    layer5_outputs(2777) <= b;
    layer5_outputs(2778) <= not (a xor b);
    layer5_outputs(2779) <= a;
    layer5_outputs(2780) <= not a or b;
    layer5_outputs(2781) <= not b;
    layer5_outputs(2782) <= not b;
    layer5_outputs(2783) <= not (a or b);
    layer5_outputs(2784) <= not b;
    layer5_outputs(2785) <= not b;
    layer5_outputs(2786) <= a xor b;
    layer5_outputs(2787) <= a and not b;
    layer5_outputs(2788) <= not a;
    layer5_outputs(2789) <= not b or a;
    layer5_outputs(2790) <= not a or b;
    layer5_outputs(2791) <= '0';
    layer5_outputs(2792) <= not (a xor b);
    layer5_outputs(2793) <= not b;
    layer5_outputs(2794) <= a;
    layer5_outputs(2795) <= not a or b;
    layer5_outputs(2796) <= not a;
    layer5_outputs(2797) <= b;
    layer5_outputs(2798) <= b;
    layer5_outputs(2799) <= not a or b;
    layer5_outputs(2800) <= b;
    layer5_outputs(2801) <= not b or a;
    layer5_outputs(2802) <= b;
    layer5_outputs(2803) <= not b;
    layer5_outputs(2804) <= not b;
    layer5_outputs(2805) <= not (a or b);
    layer5_outputs(2806) <= not b;
    layer5_outputs(2807) <= not b or a;
    layer5_outputs(2808) <= not a;
    layer5_outputs(2809) <= b;
    layer5_outputs(2810) <= a and b;
    layer5_outputs(2811) <= not a or b;
    layer5_outputs(2812) <= not a or b;
    layer5_outputs(2813) <= b;
    layer5_outputs(2814) <= a and not b;
    layer5_outputs(2815) <= a xor b;
    layer5_outputs(2816) <= a xor b;
    layer5_outputs(2817) <= not b;
    layer5_outputs(2818) <= a and b;
    layer5_outputs(2819) <= not (a or b);
    layer5_outputs(2820) <= a;
    layer5_outputs(2821) <= a and b;
    layer5_outputs(2822) <= a and not b;
    layer5_outputs(2823) <= a and b;
    layer5_outputs(2824) <= a;
    layer5_outputs(2825) <= not (a xor b);
    layer5_outputs(2826) <= a xor b;
    layer5_outputs(2827) <= not a;
    layer5_outputs(2828) <= a;
    layer5_outputs(2829) <= not (a or b);
    layer5_outputs(2830) <= a xor b;
    layer5_outputs(2831) <= not b;
    layer5_outputs(2832) <= a and b;
    layer5_outputs(2833) <= a;
    layer5_outputs(2834) <= b and not a;
    layer5_outputs(2835) <= not (a and b);
    layer5_outputs(2836) <= a and b;
    layer5_outputs(2837) <= b;
    layer5_outputs(2838) <= not (a and b);
    layer5_outputs(2839) <= a or b;
    layer5_outputs(2840) <= b;
    layer5_outputs(2841) <= '1';
    layer5_outputs(2842) <= not a or b;
    layer5_outputs(2843) <= a or b;
    layer5_outputs(2844) <= a and not b;
    layer5_outputs(2845) <= a or b;
    layer5_outputs(2846) <= b;
    layer5_outputs(2847) <= a xor b;
    layer5_outputs(2848) <= a and b;
    layer5_outputs(2849) <= not (a and b);
    layer5_outputs(2850) <= not b;
    layer5_outputs(2851) <= b and not a;
    layer5_outputs(2852) <= not a or b;
    layer5_outputs(2853) <= not (a or b);
    layer5_outputs(2854) <= not b;
    layer5_outputs(2855) <= a or b;
    layer5_outputs(2856) <= not b;
    layer5_outputs(2857) <= not a;
    layer5_outputs(2858) <= a and not b;
    layer5_outputs(2859) <= not a;
    layer5_outputs(2860) <= a and b;
    layer5_outputs(2861) <= b;
    layer5_outputs(2862) <= not a;
    layer5_outputs(2863) <= a and not b;
    layer5_outputs(2864) <= a and b;
    layer5_outputs(2865) <= not (a xor b);
    layer5_outputs(2866) <= a xor b;
    layer5_outputs(2867) <= not (a or b);
    layer5_outputs(2868) <= not a;
    layer5_outputs(2869) <= not b;
    layer5_outputs(2870) <= a and not b;
    layer5_outputs(2871) <= a xor b;
    layer5_outputs(2872) <= not a;
    layer5_outputs(2873) <= a xor b;
    layer5_outputs(2874) <= not (a and b);
    layer5_outputs(2875) <= a and b;
    layer5_outputs(2876) <= not b;
    layer5_outputs(2877) <= b;
    layer5_outputs(2878) <= b;
    layer5_outputs(2879) <= b;
    layer5_outputs(2880) <= not (a xor b);
    layer5_outputs(2881) <= not b;
    layer5_outputs(2882) <= not a or b;
    layer5_outputs(2883) <= not b;
    layer5_outputs(2884) <= not (a and b);
    layer5_outputs(2885) <= a;
    layer5_outputs(2886) <= b;
    layer5_outputs(2887) <= b and not a;
    layer5_outputs(2888) <= not a;
    layer5_outputs(2889) <= a xor b;
    layer5_outputs(2890) <= a xor b;
    layer5_outputs(2891) <= not b;
    layer5_outputs(2892) <= not (a or b);
    layer5_outputs(2893) <= not b;
    layer5_outputs(2894) <= '1';
    layer5_outputs(2895) <= not (a xor b);
    layer5_outputs(2896) <= not (a and b);
    layer5_outputs(2897) <= not b;
    layer5_outputs(2898) <= not (a and b);
    layer5_outputs(2899) <= b;
    layer5_outputs(2900) <= not a;
    layer5_outputs(2901) <= a;
    layer5_outputs(2902) <= '1';
    layer5_outputs(2903) <= a;
    layer5_outputs(2904) <= not a;
    layer5_outputs(2905) <= not a;
    layer5_outputs(2906) <= a xor b;
    layer5_outputs(2907) <= not b;
    layer5_outputs(2908) <= not b;
    layer5_outputs(2909) <= a and b;
    layer5_outputs(2910) <= not b;
    layer5_outputs(2911) <= a;
    layer5_outputs(2912) <= not a;
    layer5_outputs(2913) <= a xor b;
    layer5_outputs(2914) <= not a or b;
    layer5_outputs(2915) <= not (a or b);
    layer5_outputs(2916) <= not b;
    layer5_outputs(2917) <= not a;
    layer5_outputs(2918) <= a or b;
    layer5_outputs(2919) <= a and b;
    layer5_outputs(2920) <= a and not b;
    layer5_outputs(2921) <= a;
    layer5_outputs(2922) <= a;
    layer5_outputs(2923) <= not b;
    layer5_outputs(2924) <= a or b;
    layer5_outputs(2925) <= '1';
    layer5_outputs(2926) <= a and b;
    layer5_outputs(2927) <= a and b;
    layer5_outputs(2928) <= not a;
    layer5_outputs(2929) <= not (a or b);
    layer5_outputs(2930) <= not (a or b);
    layer5_outputs(2931) <= not (a xor b);
    layer5_outputs(2932) <= a and not b;
    layer5_outputs(2933) <= not (a xor b);
    layer5_outputs(2934) <= not b or a;
    layer5_outputs(2935) <= not a;
    layer5_outputs(2936) <= b and not a;
    layer5_outputs(2937) <= not b;
    layer5_outputs(2938) <= a;
    layer5_outputs(2939) <= not b;
    layer5_outputs(2940) <= not (a and b);
    layer5_outputs(2941) <= not b;
    layer5_outputs(2942) <= not (a or b);
    layer5_outputs(2943) <= a;
    layer5_outputs(2944) <= b;
    layer5_outputs(2945) <= a;
    layer5_outputs(2946) <= b and not a;
    layer5_outputs(2947) <= '0';
    layer5_outputs(2948) <= a or b;
    layer5_outputs(2949) <= not b;
    layer5_outputs(2950) <= not (a xor b);
    layer5_outputs(2951) <= not b;
    layer5_outputs(2952) <= a or b;
    layer5_outputs(2953) <= not (a and b);
    layer5_outputs(2954) <= not (a xor b);
    layer5_outputs(2955) <= b;
    layer5_outputs(2956) <= not b;
    layer5_outputs(2957) <= not b;
    layer5_outputs(2958) <= not (a and b);
    layer5_outputs(2959) <= a and b;
    layer5_outputs(2960) <= not (a xor b);
    layer5_outputs(2961) <= not (a xor b);
    layer5_outputs(2962) <= not b;
    layer5_outputs(2963) <= a;
    layer5_outputs(2964) <= b;
    layer5_outputs(2965) <= b;
    layer5_outputs(2966) <= b;
    layer5_outputs(2967) <= not b or a;
    layer5_outputs(2968) <= a xor b;
    layer5_outputs(2969) <= a and b;
    layer5_outputs(2970) <= not a;
    layer5_outputs(2971) <= not a;
    layer5_outputs(2972) <= not a;
    layer5_outputs(2973) <= a and not b;
    layer5_outputs(2974) <= not b or a;
    layer5_outputs(2975) <= not (a xor b);
    layer5_outputs(2976) <= a and b;
    layer5_outputs(2977) <= not a;
    layer5_outputs(2978) <= a and b;
    layer5_outputs(2979) <= not a;
    layer5_outputs(2980) <= b;
    layer5_outputs(2981) <= b and not a;
    layer5_outputs(2982) <= b;
    layer5_outputs(2983) <= a;
    layer5_outputs(2984) <= a and b;
    layer5_outputs(2985) <= not a or b;
    layer5_outputs(2986) <= not b;
    layer5_outputs(2987) <= a and not b;
    layer5_outputs(2988) <= b;
    layer5_outputs(2989) <= b and not a;
    layer5_outputs(2990) <= b;
    layer5_outputs(2991) <= b;
    layer5_outputs(2992) <= a and b;
    layer5_outputs(2993) <= a xor b;
    layer5_outputs(2994) <= not (a xor b);
    layer5_outputs(2995) <= a or b;
    layer5_outputs(2996) <= not b;
    layer5_outputs(2997) <= not a;
    layer5_outputs(2998) <= a;
    layer5_outputs(2999) <= not a;
    layer5_outputs(3000) <= not b;
    layer5_outputs(3001) <= a;
    layer5_outputs(3002) <= not (a or b);
    layer5_outputs(3003) <= a;
    layer5_outputs(3004) <= not (a xor b);
    layer5_outputs(3005) <= a or b;
    layer5_outputs(3006) <= not (a or b);
    layer5_outputs(3007) <= b;
    layer5_outputs(3008) <= a xor b;
    layer5_outputs(3009) <= a;
    layer5_outputs(3010) <= a or b;
    layer5_outputs(3011) <= b and not a;
    layer5_outputs(3012) <= not b;
    layer5_outputs(3013) <= b;
    layer5_outputs(3014) <= not a;
    layer5_outputs(3015) <= a and not b;
    layer5_outputs(3016) <= a;
    layer5_outputs(3017) <= a;
    layer5_outputs(3018) <= a and not b;
    layer5_outputs(3019) <= not b or a;
    layer5_outputs(3020) <= not (a and b);
    layer5_outputs(3021) <= not b;
    layer5_outputs(3022) <= not a or b;
    layer5_outputs(3023) <= not b;
    layer5_outputs(3024) <= a or b;
    layer5_outputs(3025) <= a xor b;
    layer5_outputs(3026) <= not a;
    layer5_outputs(3027) <= b;
    layer5_outputs(3028) <= a and not b;
    layer5_outputs(3029) <= not (a and b);
    layer5_outputs(3030) <= not b or a;
    layer5_outputs(3031) <= a;
    layer5_outputs(3032) <= '1';
    layer5_outputs(3033) <= b;
    layer5_outputs(3034) <= not (a and b);
    layer5_outputs(3035) <= a xor b;
    layer5_outputs(3036) <= a;
    layer5_outputs(3037) <= a;
    layer5_outputs(3038) <= not (a and b);
    layer5_outputs(3039) <= not a;
    layer5_outputs(3040) <= not b;
    layer5_outputs(3041) <= a;
    layer5_outputs(3042) <= a xor b;
    layer5_outputs(3043) <= not a;
    layer5_outputs(3044) <= not (a or b);
    layer5_outputs(3045) <= b and not a;
    layer5_outputs(3046) <= b;
    layer5_outputs(3047) <= a and b;
    layer5_outputs(3048) <= a or b;
    layer5_outputs(3049) <= not (a xor b);
    layer5_outputs(3050) <= not b;
    layer5_outputs(3051) <= b;
    layer5_outputs(3052) <= b;
    layer5_outputs(3053) <= not (a xor b);
    layer5_outputs(3054) <= b;
    layer5_outputs(3055) <= a or b;
    layer5_outputs(3056) <= not a;
    layer5_outputs(3057) <= not a;
    layer5_outputs(3058) <= not a or b;
    layer5_outputs(3059) <= not b;
    layer5_outputs(3060) <= not b;
    layer5_outputs(3061) <= not a;
    layer5_outputs(3062) <= not (a xor b);
    layer5_outputs(3063) <= not a;
    layer5_outputs(3064) <= not a;
    layer5_outputs(3065) <= not (a xor b);
    layer5_outputs(3066) <= b;
    layer5_outputs(3067) <= not (a or b);
    layer5_outputs(3068) <= b and not a;
    layer5_outputs(3069) <= not a or b;
    layer5_outputs(3070) <= '1';
    layer5_outputs(3071) <= not (a xor b);
    layer5_outputs(3072) <= a;
    layer5_outputs(3073) <= not a;
    layer5_outputs(3074) <= b and not a;
    layer5_outputs(3075) <= not (a or b);
    layer5_outputs(3076) <= a and not b;
    layer5_outputs(3077) <= not a;
    layer5_outputs(3078) <= not (a xor b);
    layer5_outputs(3079) <= not a;
    layer5_outputs(3080) <= not a;
    layer5_outputs(3081) <= b;
    layer5_outputs(3082) <= b;
    layer5_outputs(3083) <= not (a and b);
    layer5_outputs(3084) <= b;
    layer5_outputs(3085) <= not (a and b);
    layer5_outputs(3086) <= b;
    layer5_outputs(3087) <= not (a xor b);
    layer5_outputs(3088) <= not (a xor b);
    layer5_outputs(3089) <= a;
    layer5_outputs(3090) <= a;
    layer5_outputs(3091) <= not (a or b);
    layer5_outputs(3092) <= a xor b;
    layer5_outputs(3093) <= a;
    layer5_outputs(3094) <= not (a xor b);
    layer5_outputs(3095) <= '1';
    layer5_outputs(3096) <= not (a xor b);
    layer5_outputs(3097) <= not (a xor b);
    layer5_outputs(3098) <= b and not a;
    layer5_outputs(3099) <= not (a xor b);
    layer5_outputs(3100) <= a xor b;
    layer5_outputs(3101) <= not (a or b);
    layer5_outputs(3102) <= b and not a;
    layer5_outputs(3103) <= not b;
    layer5_outputs(3104) <= a and not b;
    layer5_outputs(3105) <= not b;
    layer5_outputs(3106) <= a;
    layer5_outputs(3107) <= a;
    layer5_outputs(3108) <= a or b;
    layer5_outputs(3109) <= a or b;
    layer5_outputs(3110) <= b and not a;
    layer5_outputs(3111) <= b;
    layer5_outputs(3112) <= a xor b;
    layer5_outputs(3113) <= a or b;
    layer5_outputs(3114) <= not b or a;
    layer5_outputs(3115) <= not b or a;
    layer5_outputs(3116) <= not a;
    layer5_outputs(3117) <= not a;
    layer5_outputs(3118) <= not (a or b);
    layer5_outputs(3119) <= not (a xor b);
    layer5_outputs(3120) <= not (a or b);
    layer5_outputs(3121) <= not (a xor b);
    layer5_outputs(3122) <= b and not a;
    layer5_outputs(3123) <= not (a and b);
    layer5_outputs(3124) <= not (a xor b);
    layer5_outputs(3125) <= a xor b;
    layer5_outputs(3126) <= a and not b;
    layer5_outputs(3127) <= not b;
    layer5_outputs(3128) <= not a;
    layer5_outputs(3129) <= not a;
    layer5_outputs(3130) <= a;
    layer5_outputs(3131) <= not (a xor b);
    layer5_outputs(3132) <= a;
    layer5_outputs(3133) <= not (a and b);
    layer5_outputs(3134) <= not a;
    layer5_outputs(3135) <= a;
    layer5_outputs(3136) <= a and not b;
    layer5_outputs(3137) <= b;
    layer5_outputs(3138) <= not (a or b);
    layer5_outputs(3139) <= not b;
    layer5_outputs(3140) <= not (a or b);
    layer5_outputs(3141) <= a;
    layer5_outputs(3142) <= not b;
    layer5_outputs(3143) <= not (a or b);
    layer5_outputs(3144) <= not a;
    layer5_outputs(3145) <= not a;
    layer5_outputs(3146) <= a or b;
    layer5_outputs(3147) <= not a;
    layer5_outputs(3148) <= a or b;
    layer5_outputs(3149) <= a and b;
    layer5_outputs(3150) <= a or b;
    layer5_outputs(3151) <= a and b;
    layer5_outputs(3152) <= a;
    layer5_outputs(3153) <= b and not a;
    layer5_outputs(3154) <= a;
    layer5_outputs(3155) <= not b;
    layer5_outputs(3156) <= not b;
    layer5_outputs(3157) <= '1';
    layer5_outputs(3158) <= not (a and b);
    layer5_outputs(3159) <= a;
    layer5_outputs(3160) <= a;
    layer5_outputs(3161) <= not a;
    layer5_outputs(3162) <= not b;
    layer5_outputs(3163) <= not a;
    layer5_outputs(3164) <= b;
    layer5_outputs(3165) <= a and b;
    layer5_outputs(3166) <= b;
    layer5_outputs(3167) <= not a;
    layer5_outputs(3168) <= not b;
    layer5_outputs(3169) <= not a;
    layer5_outputs(3170) <= a or b;
    layer5_outputs(3171) <= not b or a;
    layer5_outputs(3172) <= a xor b;
    layer5_outputs(3173) <= a xor b;
    layer5_outputs(3174) <= a;
    layer5_outputs(3175) <= not b or a;
    layer5_outputs(3176) <= not (a or b);
    layer5_outputs(3177) <= not a or b;
    layer5_outputs(3178) <= not a;
    layer5_outputs(3179) <= not a;
    layer5_outputs(3180) <= b;
    layer5_outputs(3181) <= not (a and b);
    layer5_outputs(3182) <= not (a xor b);
    layer5_outputs(3183) <= b;
    layer5_outputs(3184) <= not b;
    layer5_outputs(3185) <= a;
    layer5_outputs(3186) <= a and not b;
    layer5_outputs(3187) <= not b;
    layer5_outputs(3188) <= a;
    layer5_outputs(3189) <= not (a xor b);
    layer5_outputs(3190) <= not a or b;
    layer5_outputs(3191) <= b;
    layer5_outputs(3192) <= not b;
    layer5_outputs(3193) <= a and not b;
    layer5_outputs(3194) <= a and b;
    layer5_outputs(3195) <= not a;
    layer5_outputs(3196) <= b;
    layer5_outputs(3197) <= not b;
    layer5_outputs(3198) <= not b;
    layer5_outputs(3199) <= not b;
    layer5_outputs(3200) <= not b or a;
    layer5_outputs(3201) <= a and b;
    layer5_outputs(3202) <= not b;
    layer5_outputs(3203) <= not (a or b);
    layer5_outputs(3204) <= b;
    layer5_outputs(3205) <= not a;
    layer5_outputs(3206) <= not (a or b);
    layer5_outputs(3207) <= not (a xor b);
    layer5_outputs(3208) <= a and b;
    layer5_outputs(3209) <= not b;
    layer5_outputs(3210) <= not b;
    layer5_outputs(3211) <= not (a xor b);
    layer5_outputs(3212) <= not (a or b);
    layer5_outputs(3213) <= not (a and b);
    layer5_outputs(3214) <= not b or a;
    layer5_outputs(3215) <= not b;
    layer5_outputs(3216) <= a or b;
    layer5_outputs(3217) <= a and b;
    layer5_outputs(3218) <= b;
    layer5_outputs(3219) <= a xor b;
    layer5_outputs(3220) <= a;
    layer5_outputs(3221) <= a and b;
    layer5_outputs(3222) <= not b or a;
    layer5_outputs(3223) <= '1';
    layer5_outputs(3224) <= b;
    layer5_outputs(3225) <= not (a xor b);
    layer5_outputs(3226) <= not (a and b);
    layer5_outputs(3227) <= b and not a;
    layer5_outputs(3228) <= b and not a;
    layer5_outputs(3229) <= a;
    layer5_outputs(3230) <= not (a xor b);
    layer5_outputs(3231) <= not (a and b);
    layer5_outputs(3232) <= a;
    layer5_outputs(3233) <= not a;
    layer5_outputs(3234) <= '0';
    layer5_outputs(3235) <= a;
    layer5_outputs(3236) <= a;
    layer5_outputs(3237) <= a;
    layer5_outputs(3238) <= a and b;
    layer5_outputs(3239) <= b;
    layer5_outputs(3240) <= not (a xor b);
    layer5_outputs(3241) <= not b or a;
    layer5_outputs(3242) <= a and b;
    layer5_outputs(3243) <= not a or b;
    layer5_outputs(3244) <= not (a or b);
    layer5_outputs(3245) <= not a;
    layer5_outputs(3246) <= a or b;
    layer5_outputs(3247) <= a xor b;
    layer5_outputs(3248) <= not (a xor b);
    layer5_outputs(3249) <= a;
    layer5_outputs(3250) <= a and not b;
    layer5_outputs(3251) <= not b;
    layer5_outputs(3252) <= b and not a;
    layer5_outputs(3253) <= a or b;
    layer5_outputs(3254) <= not (a or b);
    layer5_outputs(3255) <= a;
    layer5_outputs(3256) <= not (a and b);
    layer5_outputs(3257) <= not b;
    layer5_outputs(3258) <= a xor b;
    layer5_outputs(3259) <= not a;
    layer5_outputs(3260) <= b and not a;
    layer5_outputs(3261) <= b and not a;
    layer5_outputs(3262) <= a;
    layer5_outputs(3263) <= a;
    layer5_outputs(3264) <= a or b;
    layer5_outputs(3265) <= b;
    layer5_outputs(3266) <= a and b;
    layer5_outputs(3267) <= b;
    layer5_outputs(3268) <= b;
    layer5_outputs(3269) <= not b or a;
    layer5_outputs(3270) <= a and not b;
    layer5_outputs(3271) <= b and not a;
    layer5_outputs(3272) <= not (a and b);
    layer5_outputs(3273) <= not (a xor b);
    layer5_outputs(3274) <= b and not a;
    layer5_outputs(3275) <= not a;
    layer5_outputs(3276) <= not (a or b);
    layer5_outputs(3277) <= not a or b;
    layer5_outputs(3278) <= not (a xor b);
    layer5_outputs(3279) <= not b;
    layer5_outputs(3280) <= a;
    layer5_outputs(3281) <= a;
    layer5_outputs(3282) <= not (a xor b);
    layer5_outputs(3283) <= a;
    layer5_outputs(3284) <= a xor b;
    layer5_outputs(3285) <= not (a or b);
    layer5_outputs(3286) <= a and b;
    layer5_outputs(3287) <= not b;
    layer5_outputs(3288) <= not (a xor b);
    layer5_outputs(3289) <= not b;
    layer5_outputs(3290) <= not (a xor b);
    layer5_outputs(3291) <= b;
    layer5_outputs(3292) <= b and not a;
    layer5_outputs(3293) <= a and not b;
    layer5_outputs(3294) <= a xor b;
    layer5_outputs(3295) <= '0';
    layer5_outputs(3296) <= not b;
    layer5_outputs(3297) <= a;
    layer5_outputs(3298) <= a and b;
    layer5_outputs(3299) <= '0';
    layer5_outputs(3300) <= not b;
    layer5_outputs(3301) <= a and not b;
    layer5_outputs(3302) <= a or b;
    layer5_outputs(3303) <= a;
    layer5_outputs(3304) <= not (a xor b);
    layer5_outputs(3305) <= not a;
    layer5_outputs(3306) <= '1';
    layer5_outputs(3307) <= a and not b;
    layer5_outputs(3308) <= b;
    layer5_outputs(3309) <= a;
    layer5_outputs(3310) <= a and not b;
    layer5_outputs(3311) <= not (a and b);
    layer5_outputs(3312) <= not (a and b);
    layer5_outputs(3313) <= not b;
    layer5_outputs(3314) <= not (a or b);
    layer5_outputs(3315) <= not (a xor b);
    layer5_outputs(3316) <= b;
    layer5_outputs(3317) <= not b;
    layer5_outputs(3318) <= not a or b;
    layer5_outputs(3319) <= a and not b;
    layer5_outputs(3320) <= not (a and b);
    layer5_outputs(3321) <= b and not a;
    layer5_outputs(3322) <= a xor b;
    layer5_outputs(3323) <= a;
    layer5_outputs(3324) <= a or b;
    layer5_outputs(3325) <= b;
    layer5_outputs(3326) <= not b or a;
    layer5_outputs(3327) <= b and not a;
    layer5_outputs(3328) <= not b or a;
    layer5_outputs(3329) <= b and not a;
    layer5_outputs(3330) <= a;
    layer5_outputs(3331) <= not (a or b);
    layer5_outputs(3332) <= a xor b;
    layer5_outputs(3333) <= b and not a;
    layer5_outputs(3334) <= not (a xor b);
    layer5_outputs(3335) <= not b;
    layer5_outputs(3336) <= b;
    layer5_outputs(3337) <= not (a xor b);
    layer5_outputs(3338) <= a xor b;
    layer5_outputs(3339) <= not a or b;
    layer5_outputs(3340) <= b;
    layer5_outputs(3341) <= not a or b;
    layer5_outputs(3342) <= a and b;
    layer5_outputs(3343) <= not b;
    layer5_outputs(3344) <= b;
    layer5_outputs(3345) <= not (a xor b);
    layer5_outputs(3346) <= not b;
    layer5_outputs(3347) <= b;
    layer5_outputs(3348) <= not b or a;
    layer5_outputs(3349) <= a;
    layer5_outputs(3350) <= a xor b;
    layer5_outputs(3351) <= not b;
    layer5_outputs(3352) <= not (a xor b);
    layer5_outputs(3353) <= not (a or b);
    layer5_outputs(3354) <= a or b;
    layer5_outputs(3355) <= a or b;
    layer5_outputs(3356) <= not (a and b);
    layer5_outputs(3357) <= not a;
    layer5_outputs(3358) <= b and not a;
    layer5_outputs(3359) <= not (a and b);
    layer5_outputs(3360) <= not (a and b);
    layer5_outputs(3361) <= a;
    layer5_outputs(3362) <= not (a xor b);
    layer5_outputs(3363) <= a;
    layer5_outputs(3364) <= not a;
    layer5_outputs(3365) <= not a;
    layer5_outputs(3366) <= b and not a;
    layer5_outputs(3367) <= not b or a;
    layer5_outputs(3368) <= not (a or b);
    layer5_outputs(3369) <= a;
    layer5_outputs(3370) <= not a or b;
    layer5_outputs(3371) <= a xor b;
    layer5_outputs(3372) <= not a or b;
    layer5_outputs(3373) <= not a;
    layer5_outputs(3374) <= not (a xor b);
    layer5_outputs(3375) <= a xor b;
    layer5_outputs(3376) <= not (a xor b);
    layer5_outputs(3377) <= b;
    layer5_outputs(3378) <= not b;
    layer5_outputs(3379) <= not a;
    layer5_outputs(3380) <= a and not b;
    layer5_outputs(3381) <= a and not b;
    layer5_outputs(3382) <= not b;
    layer5_outputs(3383) <= a;
    layer5_outputs(3384) <= b;
    layer5_outputs(3385) <= not b;
    layer5_outputs(3386) <= b;
    layer5_outputs(3387) <= a or b;
    layer5_outputs(3388) <= not (a xor b);
    layer5_outputs(3389) <= b;
    layer5_outputs(3390) <= not a;
    layer5_outputs(3391) <= a;
    layer5_outputs(3392) <= a and b;
    layer5_outputs(3393) <= not b;
    layer5_outputs(3394) <= a and not b;
    layer5_outputs(3395) <= b;
    layer5_outputs(3396) <= not (a or b);
    layer5_outputs(3397) <= b;
    layer5_outputs(3398) <= not (a and b);
    layer5_outputs(3399) <= a or b;
    layer5_outputs(3400) <= b;
    layer5_outputs(3401) <= '1';
    layer5_outputs(3402) <= '0';
    layer5_outputs(3403) <= not b;
    layer5_outputs(3404) <= a or b;
    layer5_outputs(3405) <= a;
    layer5_outputs(3406) <= not a;
    layer5_outputs(3407) <= a;
    layer5_outputs(3408) <= not b or a;
    layer5_outputs(3409) <= not b;
    layer5_outputs(3410) <= a and not b;
    layer5_outputs(3411) <= not b or a;
    layer5_outputs(3412) <= b;
    layer5_outputs(3413) <= not b;
    layer5_outputs(3414) <= a or b;
    layer5_outputs(3415) <= a and b;
    layer5_outputs(3416) <= a or b;
    layer5_outputs(3417) <= not a;
    layer5_outputs(3418) <= not (a and b);
    layer5_outputs(3419) <= b;
    layer5_outputs(3420) <= not b;
    layer5_outputs(3421) <= not (a and b);
    layer5_outputs(3422) <= a and not b;
    layer5_outputs(3423) <= a or b;
    layer5_outputs(3424) <= not b or a;
    layer5_outputs(3425) <= not (a xor b);
    layer5_outputs(3426) <= b and not a;
    layer5_outputs(3427) <= a;
    layer5_outputs(3428) <= not (a xor b);
    layer5_outputs(3429) <= a;
    layer5_outputs(3430) <= not b or a;
    layer5_outputs(3431) <= a;
    layer5_outputs(3432) <= a xor b;
    layer5_outputs(3433) <= b;
    layer5_outputs(3434) <= not (a or b);
    layer5_outputs(3435) <= '0';
    layer5_outputs(3436) <= not b or a;
    layer5_outputs(3437) <= a and b;
    layer5_outputs(3438) <= not (a and b);
    layer5_outputs(3439) <= a;
    layer5_outputs(3440) <= not (a or b);
    layer5_outputs(3441) <= not b;
    layer5_outputs(3442) <= '1';
    layer5_outputs(3443) <= not (a and b);
    layer5_outputs(3444) <= a or b;
    layer5_outputs(3445) <= b;
    layer5_outputs(3446) <= not b;
    layer5_outputs(3447) <= not (a or b);
    layer5_outputs(3448) <= b;
    layer5_outputs(3449) <= '1';
    layer5_outputs(3450) <= a;
    layer5_outputs(3451) <= not (a and b);
    layer5_outputs(3452) <= b and not a;
    layer5_outputs(3453) <= not a or b;
    layer5_outputs(3454) <= a xor b;
    layer5_outputs(3455) <= not (a and b);
    layer5_outputs(3456) <= a;
    layer5_outputs(3457) <= a or b;
    layer5_outputs(3458) <= a and b;
    layer5_outputs(3459) <= not a;
    layer5_outputs(3460) <= b;
    layer5_outputs(3461) <= b;
    layer5_outputs(3462) <= not (a xor b);
    layer5_outputs(3463) <= a and not b;
    layer5_outputs(3464) <= a;
    layer5_outputs(3465) <= not b;
    layer5_outputs(3466) <= a and b;
    layer5_outputs(3467) <= a;
    layer5_outputs(3468) <= not b;
    layer5_outputs(3469) <= a;
    layer5_outputs(3470) <= a;
    layer5_outputs(3471) <= not (a and b);
    layer5_outputs(3472) <= a and not b;
    layer5_outputs(3473) <= not (a xor b);
    layer5_outputs(3474) <= a or b;
    layer5_outputs(3475) <= a and b;
    layer5_outputs(3476) <= not a or b;
    layer5_outputs(3477) <= b;
    layer5_outputs(3478) <= a xor b;
    layer5_outputs(3479) <= a or b;
    layer5_outputs(3480) <= not b or a;
    layer5_outputs(3481) <= b;
    layer5_outputs(3482) <= not (a and b);
    layer5_outputs(3483) <= not (a or b);
    layer5_outputs(3484) <= not a or b;
    layer5_outputs(3485) <= a and b;
    layer5_outputs(3486) <= a;
    layer5_outputs(3487) <= not a or b;
    layer5_outputs(3488) <= a xor b;
    layer5_outputs(3489) <= b;
    layer5_outputs(3490) <= not a or b;
    layer5_outputs(3491) <= '0';
    layer5_outputs(3492) <= not a;
    layer5_outputs(3493) <= a;
    layer5_outputs(3494) <= not b;
    layer5_outputs(3495) <= not b or a;
    layer5_outputs(3496) <= not a;
    layer5_outputs(3497) <= a and b;
    layer5_outputs(3498) <= not b;
    layer5_outputs(3499) <= not a;
    layer5_outputs(3500) <= not (a and b);
    layer5_outputs(3501) <= not b;
    layer5_outputs(3502) <= not (a xor b);
    layer5_outputs(3503) <= a;
    layer5_outputs(3504) <= a and not b;
    layer5_outputs(3505) <= not b;
    layer5_outputs(3506) <= not (a or b);
    layer5_outputs(3507) <= not a or b;
    layer5_outputs(3508) <= not (a xor b);
    layer5_outputs(3509) <= b and not a;
    layer5_outputs(3510) <= a and not b;
    layer5_outputs(3511) <= '0';
    layer5_outputs(3512) <= not b or a;
    layer5_outputs(3513) <= not (a or b);
    layer5_outputs(3514) <= not a;
    layer5_outputs(3515) <= not a or b;
    layer5_outputs(3516) <= a;
    layer5_outputs(3517) <= a and not b;
    layer5_outputs(3518) <= not (a xor b);
    layer5_outputs(3519) <= not b;
    layer5_outputs(3520) <= not a or b;
    layer5_outputs(3521) <= not (a and b);
    layer5_outputs(3522) <= a and b;
    layer5_outputs(3523) <= not a;
    layer5_outputs(3524) <= a and not b;
    layer5_outputs(3525) <= a or b;
    layer5_outputs(3526) <= not b;
    layer5_outputs(3527) <= not b;
    layer5_outputs(3528) <= b;
    layer5_outputs(3529) <= a;
    layer5_outputs(3530) <= not a or b;
    layer5_outputs(3531) <= a and not b;
    layer5_outputs(3532) <= a and b;
    layer5_outputs(3533) <= not (a and b);
    layer5_outputs(3534) <= a and not b;
    layer5_outputs(3535) <= not a or b;
    layer5_outputs(3536) <= a xor b;
    layer5_outputs(3537) <= a and not b;
    layer5_outputs(3538) <= not a or b;
    layer5_outputs(3539) <= a;
    layer5_outputs(3540) <= not b or a;
    layer5_outputs(3541) <= not b;
    layer5_outputs(3542) <= not a;
    layer5_outputs(3543) <= not (a and b);
    layer5_outputs(3544) <= not (a and b);
    layer5_outputs(3545) <= not b;
    layer5_outputs(3546) <= a;
    layer5_outputs(3547) <= a;
    layer5_outputs(3548) <= a;
    layer5_outputs(3549) <= a;
    layer5_outputs(3550) <= a or b;
    layer5_outputs(3551) <= a or b;
    layer5_outputs(3552) <= not (a xor b);
    layer5_outputs(3553) <= not a;
    layer5_outputs(3554) <= not b or a;
    layer5_outputs(3555) <= b and not a;
    layer5_outputs(3556) <= not a or b;
    layer5_outputs(3557) <= a and b;
    layer5_outputs(3558) <= b;
    layer5_outputs(3559) <= not b;
    layer5_outputs(3560) <= a;
    layer5_outputs(3561) <= not b;
    layer5_outputs(3562) <= a and not b;
    layer5_outputs(3563) <= a or b;
    layer5_outputs(3564) <= b;
    layer5_outputs(3565) <= b;
    layer5_outputs(3566) <= not b;
    layer5_outputs(3567) <= a and not b;
    layer5_outputs(3568) <= a and not b;
    layer5_outputs(3569) <= b;
    layer5_outputs(3570) <= a;
    layer5_outputs(3571) <= a and not b;
    layer5_outputs(3572) <= not (a or b);
    layer5_outputs(3573) <= b;
    layer5_outputs(3574) <= a;
    layer5_outputs(3575) <= not b or a;
    layer5_outputs(3576) <= a and b;
    layer5_outputs(3577) <= not b;
    layer5_outputs(3578) <= a;
    layer5_outputs(3579) <= not a;
    layer5_outputs(3580) <= not a or b;
    layer5_outputs(3581) <= not b;
    layer5_outputs(3582) <= a;
    layer5_outputs(3583) <= a and not b;
    layer5_outputs(3584) <= a and b;
    layer5_outputs(3585) <= b;
    layer5_outputs(3586) <= not b;
    layer5_outputs(3587) <= not b or a;
    layer5_outputs(3588) <= not (a or b);
    layer5_outputs(3589) <= a;
    layer5_outputs(3590) <= '0';
    layer5_outputs(3591) <= b;
    layer5_outputs(3592) <= not a or b;
    layer5_outputs(3593) <= not b;
    layer5_outputs(3594) <= not b or a;
    layer5_outputs(3595) <= a;
    layer5_outputs(3596) <= not (a or b);
    layer5_outputs(3597) <= a and not b;
    layer5_outputs(3598) <= not (a xor b);
    layer5_outputs(3599) <= a and not b;
    layer5_outputs(3600) <= a;
    layer5_outputs(3601) <= not (a and b);
    layer5_outputs(3602) <= not b;
    layer5_outputs(3603) <= not b;
    layer5_outputs(3604) <= not a or b;
    layer5_outputs(3605) <= a xor b;
    layer5_outputs(3606) <= not (a xor b);
    layer5_outputs(3607) <= not b or a;
    layer5_outputs(3608) <= a;
    layer5_outputs(3609) <= a;
    layer5_outputs(3610) <= not b or a;
    layer5_outputs(3611) <= a;
    layer5_outputs(3612) <= not a or b;
    layer5_outputs(3613) <= not (a and b);
    layer5_outputs(3614) <= not (a xor b);
    layer5_outputs(3615) <= '0';
    layer5_outputs(3616) <= b;
    layer5_outputs(3617) <= b;
    layer5_outputs(3618) <= a;
    layer5_outputs(3619) <= not a or b;
    layer5_outputs(3620) <= a and b;
    layer5_outputs(3621) <= not b or a;
    layer5_outputs(3622) <= not (a and b);
    layer5_outputs(3623) <= a or b;
    layer5_outputs(3624) <= a;
    layer5_outputs(3625) <= not (a or b);
    layer5_outputs(3626) <= b;
    layer5_outputs(3627) <= b;
    layer5_outputs(3628) <= b;
    layer5_outputs(3629) <= not a or b;
    layer5_outputs(3630) <= not a or b;
    layer5_outputs(3631) <= not a or b;
    layer5_outputs(3632) <= not (a xor b);
    layer5_outputs(3633) <= not (a and b);
    layer5_outputs(3634) <= not b;
    layer5_outputs(3635) <= a xor b;
    layer5_outputs(3636) <= not b or a;
    layer5_outputs(3637) <= a or b;
    layer5_outputs(3638) <= not (a and b);
    layer5_outputs(3639) <= '1';
    layer5_outputs(3640) <= not a;
    layer5_outputs(3641) <= a and b;
    layer5_outputs(3642) <= b;
    layer5_outputs(3643) <= not b or a;
    layer5_outputs(3644) <= not (a or b);
    layer5_outputs(3645) <= a;
    layer5_outputs(3646) <= not (a xor b);
    layer5_outputs(3647) <= not a;
    layer5_outputs(3648) <= not (a and b);
    layer5_outputs(3649) <= b;
    layer5_outputs(3650) <= a or b;
    layer5_outputs(3651) <= not b;
    layer5_outputs(3652) <= '1';
    layer5_outputs(3653) <= not b;
    layer5_outputs(3654) <= b;
    layer5_outputs(3655) <= not (a and b);
    layer5_outputs(3656) <= a xor b;
    layer5_outputs(3657) <= not a;
    layer5_outputs(3658) <= a and b;
    layer5_outputs(3659) <= a xor b;
    layer5_outputs(3660) <= not (a or b);
    layer5_outputs(3661) <= not a;
    layer5_outputs(3662) <= a xor b;
    layer5_outputs(3663) <= a;
    layer5_outputs(3664) <= a and b;
    layer5_outputs(3665) <= not b;
    layer5_outputs(3666) <= a and not b;
    layer5_outputs(3667) <= not a;
    layer5_outputs(3668) <= not b;
    layer5_outputs(3669) <= not a;
    layer5_outputs(3670) <= b;
    layer5_outputs(3671) <= not (a or b);
    layer5_outputs(3672) <= not (a or b);
    layer5_outputs(3673) <= a and b;
    layer5_outputs(3674) <= not (a xor b);
    layer5_outputs(3675) <= a;
    layer5_outputs(3676) <= b;
    layer5_outputs(3677) <= b;
    layer5_outputs(3678) <= not b;
    layer5_outputs(3679) <= not (a or b);
    layer5_outputs(3680) <= not (a xor b);
    layer5_outputs(3681) <= not a;
    layer5_outputs(3682) <= b;
    layer5_outputs(3683) <= not a;
    layer5_outputs(3684) <= not a or b;
    layer5_outputs(3685) <= '0';
    layer5_outputs(3686) <= not (a xor b);
    layer5_outputs(3687) <= a xor b;
    layer5_outputs(3688) <= not (a and b);
    layer5_outputs(3689) <= not a or b;
    layer5_outputs(3690) <= b;
    layer5_outputs(3691) <= not b;
    layer5_outputs(3692) <= not (a or b);
    layer5_outputs(3693) <= b;
    layer5_outputs(3694) <= not (a xor b);
    layer5_outputs(3695) <= not a;
    layer5_outputs(3696) <= a;
    layer5_outputs(3697) <= not b;
    layer5_outputs(3698) <= not b;
    layer5_outputs(3699) <= a;
    layer5_outputs(3700) <= b;
    layer5_outputs(3701) <= a and not b;
    layer5_outputs(3702) <= not a;
    layer5_outputs(3703) <= not a or b;
    layer5_outputs(3704) <= a or b;
    layer5_outputs(3705) <= not (a or b);
    layer5_outputs(3706) <= not a;
    layer5_outputs(3707) <= not b;
    layer5_outputs(3708) <= not a or b;
    layer5_outputs(3709) <= not (a xor b);
    layer5_outputs(3710) <= not b;
    layer5_outputs(3711) <= not b or a;
    layer5_outputs(3712) <= '0';
    layer5_outputs(3713) <= not (a or b);
    layer5_outputs(3714) <= a xor b;
    layer5_outputs(3715) <= not b or a;
    layer5_outputs(3716) <= a and b;
    layer5_outputs(3717) <= not a;
    layer5_outputs(3718) <= a;
    layer5_outputs(3719) <= b;
    layer5_outputs(3720) <= not a;
    layer5_outputs(3721) <= not a;
    layer5_outputs(3722) <= not b;
    layer5_outputs(3723) <= a xor b;
    layer5_outputs(3724) <= not (a xor b);
    layer5_outputs(3725) <= not b;
    layer5_outputs(3726) <= a or b;
    layer5_outputs(3727) <= not (a xor b);
    layer5_outputs(3728) <= b;
    layer5_outputs(3729) <= a or b;
    layer5_outputs(3730) <= a xor b;
    layer5_outputs(3731) <= a xor b;
    layer5_outputs(3732) <= not (a or b);
    layer5_outputs(3733) <= not a;
    layer5_outputs(3734) <= not b;
    layer5_outputs(3735) <= not b;
    layer5_outputs(3736) <= not b;
    layer5_outputs(3737) <= not a;
    layer5_outputs(3738) <= a and not b;
    layer5_outputs(3739) <= not a;
    layer5_outputs(3740) <= a and b;
    layer5_outputs(3741) <= b and not a;
    layer5_outputs(3742) <= b;
    layer5_outputs(3743) <= b and not a;
    layer5_outputs(3744) <= a xor b;
    layer5_outputs(3745) <= a or b;
    layer5_outputs(3746) <= not a;
    layer5_outputs(3747) <= a xor b;
    layer5_outputs(3748) <= b;
    layer5_outputs(3749) <= not a or b;
    layer5_outputs(3750) <= b;
    layer5_outputs(3751) <= not (a and b);
    layer5_outputs(3752) <= not b;
    layer5_outputs(3753) <= not (a xor b);
    layer5_outputs(3754) <= not (a xor b);
    layer5_outputs(3755) <= b and not a;
    layer5_outputs(3756) <= not b or a;
    layer5_outputs(3757) <= not (a and b);
    layer5_outputs(3758) <= not b;
    layer5_outputs(3759) <= a;
    layer5_outputs(3760) <= not b or a;
    layer5_outputs(3761) <= a or b;
    layer5_outputs(3762) <= not a or b;
    layer5_outputs(3763) <= a and not b;
    layer5_outputs(3764) <= not a;
    layer5_outputs(3765) <= not (a or b);
    layer5_outputs(3766) <= not a;
    layer5_outputs(3767) <= a and not b;
    layer5_outputs(3768) <= not a;
    layer5_outputs(3769) <= not (a xor b);
    layer5_outputs(3770) <= a;
    layer5_outputs(3771) <= not a;
    layer5_outputs(3772) <= a or b;
    layer5_outputs(3773) <= not a;
    layer5_outputs(3774) <= b;
    layer5_outputs(3775) <= not a or b;
    layer5_outputs(3776) <= not (a and b);
    layer5_outputs(3777) <= b;
    layer5_outputs(3778) <= a xor b;
    layer5_outputs(3779) <= a or b;
    layer5_outputs(3780) <= not b;
    layer5_outputs(3781) <= a or b;
    layer5_outputs(3782) <= a;
    layer5_outputs(3783) <= not (a xor b);
    layer5_outputs(3784) <= b and not a;
    layer5_outputs(3785) <= a and b;
    layer5_outputs(3786) <= not b;
    layer5_outputs(3787) <= not (a xor b);
    layer5_outputs(3788) <= not a;
    layer5_outputs(3789) <= not (a xor b);
    layer5_outputs(3790) <= a;
    layer5_outputs(3791) <= not (a or b);
    layer5_outputs(3792) <= not b;
    layer5_outputs(3793) <= not (a and b);
    layer5_outputs(3794) <= a and not b;
    layer5_outputs(3795) <= a;
    layer5_outputs(3796) <= a;
    layer5_outputs(3797) <= not (a and b);
    layer5_outputs(3798) <= b;
    layer5_outputs(3799) <= not b or a;
    layer5_outputs(3800) <= not (a xor b);
    layer5_outputs(3801) <= not b or a;
    layer5_outputs(3802) <= b and not a;
    layer5_outputs(3803) <= a and b;
    layer5_outputs(3804) <= not (a xor b);
    layer5_outputs(3805) <= not a;
    layer5_outputs(3806) <= not b or a;
    layer5_outputs(3807) <= b and not a;
    layer5_outputs(3808) <= a;
    layer5_outputs(3809) <= not b;
    layer5_outputs(3810) <= not a or b;
    layer5_outputs(3811) <= not a;
    layer5_outputs(3812) <= b;
    layer5_outputs(3813) <= not b or a;
    layer5_outputs(3814) <= not (a xor b);
    layer5_outputs(3815) <= a and not b;
    layer5_outputs(3816) <= not b;
    layer5_outputs(3817) <= not (a or b);
    layer5_outputs(3818) <= a;
    layer5_outputs(3819) <= a;
    layer5_outputs(3820) <= not (a or b);
    layer5_outputs(3821) <= not (a or b);
    layer5_outputs(3822) <= a xor b;
    layer5_outputs(3823) <= b;
    layer5_outputs(3824) <= not a or b;
    layer5_outputs(3825) <= not a;
    layer5_outputs(3826) <= not b;
    layer5_outputs(3827) <= b and not a;
    layer5_outputs(3828) <= b and not a;
    layer5_outputs(3829) <= not (a and b);
    layer5_outputs(3830) <= a;
    layer5_outputs(3831) <= not a;
    layer5_outputs(3832) <= not (a xor b);
    layer5_outputs(3833) <= not b or a;
    layer5_outputs(3834) <= a xor b;
    layer5_outputs(3835) <= not a;
    layer5_outputs(3836) <= not b;
    layer5_outputs(3837) <= not (a xor b);
    layer5_outputs(3838) <= not a;
    layer5_outputs(3839) <= a and b;
    layer5_outputs(3840) <= a and not b;
    layer5_outputs(3841) <= b;
    layer5_outputs(3842) <= a xor b;
    layer5_outputs(3843) <= not a;
    layer5_outputs(3844) <= '1';
    layer5_outputs(3845) <= not b or a;
    layer5_outputs(3846) <= b;
    layer5_outputs(3847) <= a and b;
    layer5_outputs(3848) <= a and b;
    layer5_outputs(3849) <= not b;
    layer5_outputs(3850) <= not b;
    layer5_outputs(3851) <= b;
    layer5_outputs(3852) <= a and b;
    layer5_outputs(3853) <= a;
    layer5_outputs(3854) <= b;
    layer5_outputs(3855) <= not b;
    layer5_outputs(3856) <= not b;
    layer5_outputs(3857) <= not (a or b);
    layer5_outputs(3858) <= not b;
    layer5_outputs(3859) <= b;
    layer5_outputs(3860) <= not a;
    layer5_outputs(3861) <= a;
    layer5_outputs(3862) <= not a;
    layer5_outputs(3863) <= not b or a;
    layer5_outputs(3864) <= '1';
    layer5_outputs(3865) <= a and b;
    layer5_outputs(3866) <= not a or b;
    layer5_outputs(3867) <= b and not a;
    layer5_outputs(3868) <= not b or a;
    layer5_outputs(3869) <= not a;
    layer5_outputs(3870) <= b and not a;
    layer5_outputs(3871) <= b;
    layer5_outputs(3872) <= not a;
    layer5_outputs(3873) <= not b or a;
    layer5_outputs(3874) <= not b;
    layer5_outputs(3875) <= a xor b;
    layer5_outputs(3876) <= not (a and b);
    layer5_outputs(3877) <= not (a or b);
    layer5_outputs(3878) <= a or b;
    layer5_outputs(3879) <= not (a and b);
    layer5_outputs(3880) <= not (a and b);
    layer5_outputs(3881) <= not a;
    layer5_outputs(3882) <= not (a and b);
    layer5_outputs(3883) <= not a;
    layer5_outputs(3884) <= not b;
    layer5_outputs(3885) <= a xor b;
    layer5_outputs(3886) <= a xor b;
    layer5_outputs(3887) <= not a;
    layer5_outputs(3888) <= not b;
    layer5_outputs(3889) <= not a or b;
    layer5_outputs(3890) <= a xor b;
    layer5_outputs(3891) <= a or b;
    layer5_outputs(3892) <= a or b;
    layer5_outputs(3893) <= a and not b;
    layer5_outputs(3894) <= b;
    layer5_outputs(3895) <= a xor b;
    layer5_outputs(3896) <= not b;
    layer5_outputs(3897) <= '0';
    layer5_outputs(3898) <= a or b;
    layer5_outputs(3899) <= not (a or b);
    layer5_outputs(3900) <= a xor b;
    layer5_outputs(3901) <= b;
    layer5_outputs(3902) <= not (a or b);
    layer5_outputs(3903) <= a or b;
    layer5_outputs(3904) <= a;
    layer5_outputs(3905) <= not b;
    layer5_outputs(3906) <= b and not a;
    layer5_outputs(3907) <= b and not a;
    layer5_outputs(3908) <= not b;
    layer5_outputs(3909) <= a;
    layer5_outputs(3910) <= a or b;
    layer5_outputs(3911) <= not a;
    layer5_outputs(3912) <= b;
    layer5_outputs(3913) <= a xor b;
    layer5_outputs(3914) <= a or b;
    layer5_outputs(3915) <= not (a or b);
    layer5_outputs(3916) <= a and b;
    layer5_outputs(3917) <= not b;
    layer5_outputs(3918) <= not a;
    layer5_outputs(3919) <= not a or b;
    layer5_outputs(3920) <= a xor b;
    layer5_outputs(3921) <= b;
    layer5_outputs(3922) <= not (a and b);
    layer5_outputs(3923) <= not (a and b);
    layer5_outputs(3924) <= a;
    layer5_outputs(3925) <= a and b;
    layer5_outputs(3926) <= a and not b;
    layer5_outputs(3927) <= a and b;
    layer5_outputs(3928) <= not a;
    layer5_outputs(3929) <= not b or a;
    layer5_outputs(3930) <= not a;
    layer5_outputs(3931) <= not a;
    layer5_outputs(3932) <= not b;
    layer5_outputs(3933) <= not a;
    layer5_outputs(3934) <= a and b;
    layer5_outputs(3935) <= a or b;
    layer5_outputs(3936) <= a xor b;
    layer5_outputs(3937) <= b;
    layer5_outputs(3938) <= not a;
    layer5_outputs(3939) <= b and not a;
    layer5_outputs(3940) <= not b;
    layer5_outputs(3941) <= not b or a;
    layer5_outputs(3942) <= a;
    layer5_outputs(3943) <= not b;
    layer5_outputs(3944) <= not (a and b);
    layer5_outputs(3945) <= b;
    layer5_outputs(3946) <= a xor b;
    layer5_outputs(3947) <= b;
    layer5_outputs(3948) <= not (a or b);
    layer5_outputs(3949) <= not (a and b);
    layer5_outputs(3950) <= a and not b;
    layer5_outputs(3951) <= not a or b;
    layer5_outputs(3952) <= not (a and b);
    layer5_outputs(3953) <= not b;
    layer5_outputs(3954) <= a;
    layer5_outputs(3955) <= a and not b;
    layer5_outputs(3956) <= not (a or b);
    layer5_outputs(3957) <= not (a xor b);
    layer5_outputs(3958) <= not a;
    layer5_outputs(3959) <= a or b;
    layer5_outputs(3960) <= not (a or b);
    layer5_outputs(3961) <= a and b;
    layer5_outputs(3962) <= b;
    layer5_outputs(3963) <= not b;
    layer5_outputs(3964) <= not b or a;
    layer5_outputs(3965) <= not a or b;
    layer5_outputs(3966) <= a xor b;
    layer5_outputs(3967) <= not b or a;
    layer5_outputs(3968) <= not a;
    layer5_outputs(3969) <= not b;
    layer5_outputs(3970) <= b and not a;
    layer5_outputs(3971) <= not a;
    layer5_outputs(3972) <= not a;
    layer5_outputs(3973) <= not b or a;
    layer5_outputs(3974) <= not b;
    layer5_outputs(3975) <= not a or b;
    layer5_outputs(3976) <= not b;
    layer5_outputs(3977) <= a and not b;
    layer5_outputs(3978) <= not (a and b);
    layer5_outputs(3979) <= a or b;
    layer5_outputs(3980) <= not a or b;
    layer5_outputs(3981) <= a and b;
    layer5_outputs(3982) <= a xor b;
    layer5_outputs(3983) <= not a;
    layer5_outputs(3984) <= not a;
    layer5_outputs(3985) <= b;
    layer5_outputs(3986) <= b;
    layer5_outputs(3987) <= not (a or b);
    layer5_outputs(3988) <= a;
    layer5_outputs(3989) <= not a or b;
    layer5_outputs(3990) <= not (a and b);
    layer5_outputs(3991) <= not (a xor b);
    layer5_outputs(3992) <= not a;
    layer5_outputs(3993) <= a;
    layer5_outputs(3994) <= a or b;
    layer5_outputs(3995) <= b;
    layer5_outputs(3996) <= b and not a;
    layer5_outputs(3997) <= not b;
    layer5_outputs(3998) <= not b;
    layer5_outputs(3999) <= not b;
    layer5_outputs(4000) <= b;
    layer5_outputs(4001) <= b;
    layer5_outputs(4002) <= not b;
    layer5_outputs(4003) <= a;
    layer5_outputs(4004) <= not b;
    layer5_outputs(4005) <= not (a xor b);
    layer5_outputs(4006) <= a;
    layer5_outputs(4007) <= a and not b;
    layer5_outputs(4008) <= not b;
    layer5_outputs(4009) <= not (a xor b);
    layer5_outputs(4010) <= not b;
    layer5_outputs(4011) <= not (a xor b);
    layer5_outputs(4012) <= b and not a;
    layer5_outputs(4013) <= b;
    layer5_outputs(4014) <= not a;
    layer5_outputs(4015) <= not (a xor b);
    layer5_outputs(4016) <= b;
    layer5_outputs(4017) <= '0';
    layer5_outputs(4018) <= a xor b;
    layer5_outputs(4019) <= b and not a;
    layer5_outputs(4020) <= b and not a;
    layer5_outputs(4021) <= not b;
    layer5_outputs(4022) <= a and not b;
    layer5_outputs(4023) <= not b;
    layer5_outputs(4024) <= not b;
    layer5_outputs(4025) <= not b;
    layer5_outputs(4026) <= a;
    layer5_outputs(4027) <= not (a and b);
    layer5_outputs(4028) <= not b;
    layer5_outputs(4029) <= b;
    layer5_outputs(4030) <= b;
    layer5_outputs(4031) <= not (a or b);
    layer5_outputs(4032) <= a or b;
    layer5_outputs(4033) <= not b;
    layer5_outputs(4034) <= not (a xor b);
    layer5_outputs(4035) <= not b;
    layer5_outputs(4036) <= not (a and b);
    layer5_outputs(4037) <= '0';
    layer5_outputs(4038) <= a;
    layer5_outputs(4039) <= b and not a;
    layer5_outputs(4040) <= a or b;
    layer5_outputs(4041) <= not a;
    layer5_outputs(4042) <= not b or a;
    layer5_outputs(4043) <= a xor b;
    layer5_outputs(4044) <= a and not b;
    layer5_outputs(4045) <= b;
    layer5_outputs(4046) <= not (a xor b);
    layer5_outputs(4047) <= a xor b;
    layer5_outputs(4048) <= b;
    layer5_outputs(4049) <= a xor b;
    layer5_outputs(4050) <= a;
    layer5_outputs(4051) <= not (a xor b);
    layer5_outputs(4052) <= a and not b;
    layer5_outputs(4053) <= not b or a;
    layer5_outputs(4054) <= not a or b;
    layer5_outputs(4055) <= a;
    layer5_outputs(4056) <= a and b;
    layer5_outputs(4057) <= not (a xor b);
    layer5_outputs(4058) <= not b;
    layer5_outputs(4059) <= not b or a;
    layer5_outputs(4060) <= b and not a;
    layer5_outputs(4061) <= not (a and b);
    layer5_outputs(4062) <= not b;
    layer5_outputs(4063) <= not a or b;
    layer5_outputs(4064) <= not (a and b);
    layer5_outputs(4065) <= not b or a;
    layer5_outputs(4066) <= not b;
    layer5_outputs(4067) <= not a;
    layer5_outputs(4068) <= not b;
    layer5_outputs(4069) <= a and b;
    layer5_outputs(4070) <= a;
    layer5_outputs(4071) <= not b or a;
    layer5_outputs(4072) <= a;
    layer5_outputs(4073) <= a xor b;
    layer5_outputs(4074) <= not a;
    layer5_outputs(4075) <= not (a and b);
    layer5_outputs(4076) <= not a;
    layer5_outputs(4077) <= a;
    layer5_outputs(4078) <= b;
    layer5_outputs(4079) <= not a;
    layer5_outputs(4080) <= not (a or b);
    layer5_outputs(4081) <= '0';
    layer5_outputs(4082) <= not a;
    layer5_outputs(4083) <= a and b;
    layer5_outputs(4084) <= a xor b;
    layer5_outputs(4085) <= not (a and b);
    layer5_outputs(4086) <= not a;
    layer5_outputs(4087) <= not a;
    layer5_outputs(4088) <= not b;
    layer5_outputs(4089) <= b;
    layer5_outputs(4090) <= not a;
    layer5_outputs(4091) <= a and not b;
    layer5_outputs(4092) <= not b;
    layer5_outputs(4093) <= b and not a;
    layer5_outputs(4094) <= not a or b;
    layer5_outputs(4095) <= a;
    layer5_outputs(4096) <= a and not b;
    layer5_outputs(4097) <= a or b;
    layer5_outputs(4098) <= b;
    layer5_outputs(4099) <= not b or a;
    layer5_outputs(4100) <= not b;
    layer5_outputs(4101) <= a;
    layer5_outputs(4102) <= not (a or b);
    layer5_outputs(4103) <= not a;
    layer5_outputs(4104) <= b;
    layer5_outputs(4105) <= not a;
    layer5_outputs(4106) <= a xor b;
    layer5_outputs(4107) <= a;
    layer5_outputs(4108) <= b;
    layer5_outputs(4109) <= a xor b;
    layer5_outputs(4110) <= not (a or b);
    layer5_outputs(4111) <= not b;
    layer5_outputs(4112) <= b and not a;
    layer5_outputs(4113) <= not (a xor b);
    layer5_outputs(4114) <= a and b;
    layer5_outputs(4115) <= not b;
    layer5_outputs(4116) <= not (a or b);
    layer5_outputs(4117) <= a;
    layer5_outputs(4118) <= a and not b;
    layer5_outputs(4119) <= not a;
    layer5_outputs(4120) <= a or b;
    layer5_outputs(4121) <= b;
    layer5_outputs(4122) <= not b;
    layer5_outputs(4123) <= not a;
    layer5_outputs(4124) <= not b or a;
    layer5_outputs(4125) <= not b;
    layer5_outputs(4126) <= a and b;
    layer5_outputs(4127) <= not b or a;
    layer5_outputs(4128) <= a xor b;
    layer5_outputs(4129) <= not b;
    layer5_outputs(4130) <= a or b;
    layer5_outputs(4131) <= not a;
    layer5_outputs(4132) <= a and b;
    layer5_outputs(4133) <= not (a xor b);
    layer5_outputs(4134) <= not b;
    layer5_outputs(4135) <= not (a xor b);
    layer5_outputs(4136) <= a;
    layer5_outputs(4137) <= not a;
    layer5_outputs(4138) <= not (a xor b);
    layer5_outputs(4139) <= not b;
    layer5_outputs(4140) <= not a;
    layer5_outputs(4141) <= a and b;
    layer5_outputs(4142) <= a or b;
    layer5_outputs(4143) <= not a or b;
    layer5_outputs(4144) <= a and b;
    layer5_outputs(4145) <= not a;
    layer5_outputs(4146) <= not a;
    layer5_outputs(4147) <= not b;
    layer5_outputs(4148) <= b;
    layer5_outputs(4149) <= not (a xor b);
    layer5_outputs(4150) <= b;
    layer5_outputs(4151) <= a;
    layer5_outputs(4152) <= a or b;
    layer5_outputs(4153) <= not a;
    layer5_outputs(4154) <= a;
    layer5_outputs(4155) <= a;
    layer5_outputs(4156) <= b;
    layer5_outputs(4157) <= a;
    layer5_outputs(4158) <= not b;
    layer5_outputs(4159) <= b;
    layer5_outputs(4160) <= not a;
    layer5_outputs(4161) <= not a or b;
    layer5_outputs(4162) <= not b or a;
    layer5_outputs(4163) <= b;
    layer5_outputs(4164) <= not a or b;
    layer5_outputs(4165) <= not a or b;
    layer5_outputs(4166) <= not b;
    layer5_outputs(4167) <= not (a and b);
    layer5_outputs(4168) <= b;
    layer5_outputs(4169) <= not a or b;
    layer5_outputs(4170) <= not (a or b);
    layer5_outputs(4171) <= not (a xor b);
    layer5_outputs(4172) <= not (a and b);
    layer5_outputs(4173) <= not a or b;
    layer5_outputs(4174) <= a;
    layer5_outputs(4175) <= not b;
    layer5_outputs(4176) <= b;
    layer5_outputs(4177) <= not a;
    layer5_outputs(4178) <= a;
    layer5_outputs(4179) <= not b or a;
    layer5_outputs(4180) <= not b;
    layer5_outputs(4181) <= not (a or b);
    layer5_outputs(4182) <= not a;
    layer5_outputs(4183) <= not a;
    layer5_outputs(4184) <= not (a and b);
    layer5_outputs(4185) <= a and b;
    layer5_outputs(4186) <= a;
    layer5_outputs(4187) <= not (a xor b);
    layer5_outputs(4188) <= a;
    layer5_outputs(4189) <= a xor b;
    layer5_outputs(4190) <= not (a and b);
    layer5_outputs(4191) <= not b or a;
    layer5_outputs(4192) <= b;
    layer5_outputs(4193) <= b;
    layer5_outputs(4194) <= a and not b;
    layer5_outputs(4195) <= a and b;
    layer5_outputs(4196) <= not (a xor b);
    layer5_outputs(4197) <= not a or b;
    layer5_outputs(4198) <= '1';
    layer5_outputs(4199) <= not (a and b);
    layer5_outputs(4200) <= a;
    layer5_outputs(4201) <= not a;
    layer5_outputs(4202) <= not a;
    layer5_outputs(4203) <= not b;
    layer5_outputs(4204) <= a xor b;
    layer5_outputs(4205) <= a and not b;
    layer5_outputs(4206) <= a xor b;
    layer5_outputs(4207) <= a or b;
    layer5_outputs(4208) <= not (a and b);
    layer5_outputs(4209) <= a;
    layer5_outputs(4210) <= a and b;
    layer5_outputs(4211) <= a;
    layer5_outputs(4212) <= not a;
    layer5_outputs(4213) <= not a;
    layer5_outputs(4214) <= a;
    layer5_outputs(4215) <= a and b;
    layer5_outputs(4216) <= b and not a;
    layer5_outputs(4217) <= not b or a;
    layer5_outputs(4218) <= a xor b;
    layer5_outputs(4219) <= not (a or b);
    layer5_outputs(4220) <= b and not a;
    layer5_outputs(4221) <= not a;
    layer5_outputs(4222) <= b;
    layer5_outputs(4223) <= b;
    layer5_outputs(4224) <= not (a xor b);
    layer5_outputs(4225) <= a xor b;
    layer5_outputs(4226) <= not a;
    layer5_outputs(4227) <= not a;
    layer5_outputs(4228) <= not b or a;
    layer5_outputs(4229) <= not (a xor b);
    layer5_outputs(4230) <= not b;
    layer5_outputs(4231) <= not (a or b);
    layer5_outputs(4232) <= not (a or b);
    layer5_outputs(4233) <= b and not a;
    layer5_outputs(4234) <= a or b;
    layer5_outputs(4235) <= not b or a;
    layer5_outputs(4236) <= not b or a;
    layer5_outputs(4237) <= a;
    layer5_outputs(4238) <= not a;
    layer5_outputs(4239) <= not a;
    layer5_outputs(4240) <= b and not a;
    layer5_outputs(4241) <= a xor b;
    layer5_outputs(4242) <= a;
    layer5_outputs(4243) <= b;
    layer5_outputs(4244) <= b;
    layer5_outputs(4245) <= b;
    layer5_outputs(4246) <= not b;
    layer5_outputs(4247) <= a;
    layer5_outputs(4248) <= b and not a;
    layer5_outputs(4249) <= b;
    layer5_outputs(4250) <= not a;
    layer5_outputs(4251) <= a xor b;
    layer5_outputs(4252) <= b and not a;
    layer5_outputs(4253) <= not b or a;
    layer5_outputs(4254) <= a;
    layer5_outputs(4255) <= a;
    layer5_outputs(4256) <= not a or b;
    layer5_outputs(4257) <= not a;
    layer5_outputs(4258) <= not b;
    layer5_outputs(4259) <= a xor b;
    layer5_outputs(4260) <= a and not b;
    layer5_outputs(4261) <= a xor b;
    layer5_outputs(4262) <= a or b;
    layer5_outputs(4263) <= b and not a;
    layer5_outputs(4264) <= a and b;
    layer5_outputs(4265) <= a or b;
    layer5_outputs(4266) <= b and not a;
    layer5_outputs(4267) <= b;
    layer5_outputs(4268) <= '1';
    layer5_outputs(4269) <= not b;
    layer5_outputs(4270) <= not a or b;
    layer5_outputs(4271) <= not (a and b);
    layer5_outputs(4272) <= not a;
    layer5_outputs(4273) <= a;
    layer5_outputs(4274) <= not b;
    layer5_outputs(4275) <= not a or b;
    layer5_outputs(4276) <= a;
    layer5_outputs(4277) <= not a;
    layer5_outputs(4278) <= a and b;
    layer5_outputs(4279) <= b;
    layer5_outputs(4280) <= a and not b;
    layer5_outputs(4281) <= not a;
    layer5_outputs(4282) <= b;
    layer5_outputs(4283) <= b and not a;
    layer5_outputs(4284) <= b and not a;
    layer5_outputs(4285) <= a;
    layer5_outputs(4286) <= a;
    layer5_outputs(4287) <= a xor b;
    layer5_outputs(4288) <= not a;
    layer5_outputs(4289) <= not b or a;
    layer5_outputs(4290) <= b and not a;
    layer5_outputs(4291) <= b;
    layer5_outputs(4292) <= a or b;
    layer5_outputs(4293) <= b;
    layer5_outputs(4294) <= b and not a;
    layer5_outputs(4295) <= not (a or b);
    layer5_outputs(4296) <= a and b;
    layer5_outputs(4297) <= not (a or b);
    layer5_outputs(4298) <= not a or b;
    layer5_outputs(4299) <= a xor b;
    layer5_outputs(4300) <= a xor b;
    layer5_outputs(4301) <= a xor b;
    layer5_outputs(4302) <= a and not b;
    layer5_outputs(4303) <= not a;
    layer5_outputs(4304) <= not a;
    layer5_outputs(4305) <= not b;
    layer5_outputs(4306) <= not b;
    layer5_outputs(4307) <= not (a xor b);
    layer5_outputs(4308) <= not b;
    layer5_outputs(4309) <= not b;
    layer5_outputs(4310) <= not a;
    layer5_outputs(4311) <= not b;
    layer5_outputs(4312) <= a xor b;
    layer5_outputs(4313) <= a and not b;
    layer5_outputs(4314) <= b;
    layer5_outputs(4315) <= a;
    layer5_outputs(4316) <= not b or a;
    layer5_outputs(4317) <= not b;
    layer5_outputs(4318) <= not a or b;
    layer5_outputs(4319) <= b;
    layer5_outputs(4320) <= not a;
    layer5_outputs(4321) <= b;
    layer5_outputs(4322) <= not a;
    layer5_outputs(4323) <= not (a and b);
    layer5_outputs(4324) <= not a;
    layer5_outputs(4325) <= a xor b;
    layer5_outputs(4326) <= not a;
    layer5_outputs(4327) <= a or b;
    layer5_outputs(4328) <= a or b;
    layer5_outputs(4329) <= not b;
    layer5_outputs(4330) <= a;
    layer5_outputs(4331) <= b and not a;
    layer5_outputs(4332) <= not a;
    layer5_outputs(4333) <= not b or a;
    layer5_outputs(4334) <= a xor b;
    layer5_outputs(4335) <= b and not a;
    layer5_outputs(4336) <= '0';
    layer5_outputs(4337) <= '0';
    layer5_outputs(4338) <= not (a and b);
    layer5_outputs(4339) <= a xor b;
    layer5_outputs(4340) <= b and not a;
    layer5_outputs(4341) <= b and not a;
    layer5_outputs(4342) <= not (a and b);
    layer5_outputs(4343) <= not a;
    layer5_outputs(4344) <= a;
    layer5_outputs(4345) <= a;
    layer5_outputs(4346) <= not (a or b);
    layer5_outputs(4347) <= not a;
    layer5_outputs(4348) <= not a;
    layer5_outputs(4349) <= not b;
    layer5_outputs(4350) <= b;
    layer5_outputs(4351) <= not b or a;
    layer5_outputs(4352) <= b;
    layer5_outputs(4353) <= a xor b;
    layer5_outputs(4354) <= a;
    layer5_outputs(4355) <= not b;
    layer5_outputs(4356) <= a or b;
    layer5_outputs(4357) <= b;
    layer5_outputs(4358) <= a and b;
    layer5_outputs(4359) <= not b or a;
    layer5_outputs(4360) <= not (a xor b);
    layer5_outputs(4361) <= not a;
    layer5_outputs(4362) <= not (a and b);
    layer5_outputs(4363) <= a xor b;
    layer5_outputs(4364) <= b and not a;
    layer5_outputs(4365) <= not b;
    layer5_outputs(4366) <= a;
    layer5_outputs(4367) <= b;
    layer5_outputs(4368) <= not b;
    layer5_outputs(4369) <= not (a and b);
    layer5_outputs(4370) <= a or b;
    layer5_outputs(4371) <= b;
    layer5_outputs(4372) <= not a;
    layer5_outputs(4373) <= a or b;
    layer5_outputs(4374) <= a;
    layer5_outputs(4375) <= b;
    layer5_outputs(4376) <= not b;
    layer5_outputs(4377) <= not a;
    layer5_outputs(4378) <= not (a and b);
    layer5_outputs(4379) <= a or b;
    layer5_outputs(4380) <= not b or a;
    layer5_outputs(4381) <= b and not a;
    layer5_outputs(4382) <= not (a or b);
    layer5_outputs(4383) <= not b;
    layer5_outputs(4384) <= b and not a;
    layer5_outputs(4385) <= a xor b;
    layer5_outputs(4386) <= not a;
    layer5_outputs(4387) <= a;
    layer5_outputs(4388) <= a and not b;
    layer5_outputs(4389) <= a and not b;
    layer5_outputs(4390) <= b and not a;
    layer5_outputs(4391) <= b and not a;
    layer5_outputs(4392) <= b;
    layer5_outputs(4393) <= not a or b;
    layer5_outputs(4394) <= not a;
    layer5_outputs(4395) <= a;
    layer5_outputs(4396) <= not b;
    layer5_outputs(4397) <= b;
    layer5_outputs(4398) <= not a or b;
    layer5_outputs(4399) <= not a;
    layer5_outputs(4400) <= not a;
    layer5_outputs(4401) <= not (a xor b);
    layer5_outputs(4402) <= not a or b;
    layer5_outputs(4403) <= not (a or b);
    layer5_outputs(4404) <= not (a xor b);
    layer5_outputs(4405) <= b;
    layer5_outputs(4406) <= not a or b;
    layer5_outputs(4407) <= not a;
    layer5_outputs(4408) <= not a;
    layer5_outputs(4409) <= a;
    layer5_outputs(4410) <= a;
    layer5_outputs(4411) <= a or b;
    layer5_outputs(4412) <= not (a and b);
    layer5_outputs(4413) <= a xor b;
    layer5_outputs(4414) <= not (a or b);
    layer5_outputs(4415) <= a and not b;
    layer5_outputs(4416) <= a and not b;
    layer5_outputs(4417) <= a;
    layer5_outputs(4418) <= not b;
    layer5_outputs(4419) <= not (a xor b);
    layer5_outputs(4420) <= a;
    layer5_outputs(4421) <= a and b;
    layer5_outputs(4422) <= not (a xor b);
    layer5_outputs(4423) <= a;
    layer5_outputs(4424) <= a or b;
    layer5_outputs(4425) <= a;
    layer5_outputs(4426) <= a;
    layer5_outputs(4427) <= not b;
    layer5_outputs(4428) <= not a or b;
    layer5_outputs(4429) <= a xor b;
    layer5_outputs(4430) <= a or b;
    layer5_outputs(4431) <= not a;
    layer5_outputs(4432) <= not (a and b);
    layer5_outputs(4433) <= a;
    layer5_outputs(4434) <= b and not a;
    layer5_outputs(4435) <= a and not b;
    layer5_outputs(4436) <= '1';
    layer5_outputs(4437) <= not a;
    layer5_outputs(4438) <= a xor b;
    layer5_outputs(4439) <= a xor b;
    layer5_outputs(4440) <= b and not a;
    layer5_outputs(4441) <= not b;
    layer5_outputs(4442) <= b and not a;
    layer5_outputs(4443) <= a and not b;
    layer5_outputs(4444) <= a xor b;
    layer5_outputs(4445) <= b;
    layer5_outputs(4446) <= a and not b;
    layer5_outputs(4447) <= a;
    layer5_outputs(4448) <= b;
    layer5_outputs(4449) <= not a;
    layer5_outputs(4450) <= a;
    layer5_outputs(4451) <= not b;
    layer5_outputs(4452) <= not (a or b);
    layer5_outputs(4453) <= not a;
    layer5_outputs(4454) <= '0';
    layer5_outputs(4455) <= '0';
    layer5_outputs(4456) <= b;
    layer5_outputs(4457) <= not (a xor b);
    layer5_outputs(4458) <= a xor b;
    layer5_outputs(4459) <= b;
    layer5_outputs(4460) <= not b;
    layer5_outputs(4461) <= not a;
    layer5_outputs(4462) <= b;
    layer5_outputs(4463) <= not a;
    layer5_outputs(4464) <= a and not b;
    layer5_outputs(4465) <= b and not a;
    layer5_outputs(4466) <= not b;
    layer5_outputs(4467) <= not b;
    layer5_outputs(4468) <= a;
    layer5_outputs(4469) <= not b;
    layer5_outputs(4470) <= a xor b;
    layer5_outputs(4471) <= b;
    layer5_outputs(4472) <= not a;
    layer5_outputs(4473) <= b;
    layer5_outputs(4474) <= not a;
    layer5_outputs(4475) <= b;
    layer5_outputs(4476) <= a or b;
    layer5_outputs(4477) <= not b;
    layer5_outputs(4478) <= not a or b;
    layer5_outputs(4479) <= not (a and b);
    layer5_outputs(4480) <= b;
    layer5_outputs(4481) <= not (a xor b);
    layer5_outputs(4482) <= b;
    layer5_outputs(4483) <= not (a xor b);
    layer5_outputs(4484) <= a and b;
    layer5_outputs(4485) <= a or b;
    layer5_outputs(4486) <= not (a or b);
    layer5_outputs(4487) <= a xor b;
    layer5_outputs(4488) <= a and b;
    layer5_outputs(4489) <= a;
    layer5_outputs(4490) <= not (a and b);
    layer5_outputs(4491) <= b;
    layer5_outputs(4492) <= not (a or b);
    layer5_outputs(4493) <= b and not a;
    layer5_outputs(4494) <= not a or b;
    layer5_outputs(4495) <= b;
    layer5_outputs(4496) <= not (a and b);
    layer5_outputs(4497) <= a xor b;
    layer5_outputs(4498) <= not (a and b);
    layer5_outputs(4499) <= a;
    layer5_outputs(4500) <= b and not a;
    layer5_outputs(4501) <= '0';
    layer5_outputs(4502) <= b;
    layer5_outputs(4503) <= not a or b;
    layer5_outputs(4504) <= not a;
    layer5_outputs(4505) <= not (a xor b);
    layer5_outputs(4506) <= b;
    layer5_outputs(4507) <= not a;
    layer5_outputs(4508) <= a;
    layer5_outputs(4509) <= b;
    layer5_outputs(4510) <= not a;
    layer5_outputs(4511) <= a;
    layer5_outputs(4512) <= b;
    layer5_outputs(4513) <= a;
    layer5_outputs(4514) <= not b or a;
    layer5_outputs(4515) <= not (a or b);
    layer5_outputs(4516) <= b;
    layer5_outputs(4517) <= not a;
    layer5_outputs(4518) <= not b;
    layer5_outputs(4519) <= not b or a;
    layer5_outputs(4520) <= b and not a;
    layer5_outputs(4521) <= not a or b;
    layer5_outputs(4522) <= b;
    layer5_outputs(4523) <= a and not b;
    layer5_outputs(4524) <= not a;
    layer5_outputs(4525) <= not b or a;
    layer5_outputs(4526) <= b;
    layer5_outputs(4527) <= b;
    layer5_outputs(4528) <= a;
    layer5_outputs(4529) <= b;
    layer5_outputs(4530) <= not a;
    layer5_outputs(4531) <= not b or a;
    layer5_outputs(4532) <= not b;
    layer5_outputs(4533) <= '1';
    layer5_outputs(4534) <= not b;
    layer5_outputs(4535) <= a xor b;
    layer5_outputs(4536) <= not (a and b);
    layer5_outputs(4537) <= a xor b;
    layer5_outputs(4538) <= a xor b;
    layer5_outputs(4539) <= not b;
    layer5_outputs(4540) <= not b;
    layer5_outputs(4541) <= b and not a;
    layer5_outputs(4542) <= a xor b;
    layer5_outputs(4543) <= b and not a;
    layer5_outputs(4544) <= a xor b;
    layer5_outputs(4545) <= not (a and b);
    layer5_outputs(4546) <= not a or b;
    layer5_outputs(4547) <= not (a and b);
    layer5_outputs(4548) <= not b;
    layer5_outputs(4549) <= a and not b;
    layer5_outputs(4550) <= not b;
    layer5_outputs(4551) <= a;
    layer5_outputs(4552) <= not (a or b);
    layer5_outputs(4553) <= a;
    layer5_outputs(4554) <= not a;
    layer5_outputs(4555) <= a and b;
    layer5_outputs(4556) <= not a;
    layer5_outputs(4557) <= a xor b;
    layer5_outputs(4558) <= '0';
    layer5_outputs(4559) <= not (a and b);
    layer5_outputs(4560) <= not b or a;
    layer5_outputs(4561) <= '0';
    layer5_outputs(4562) <= not b;
    layer5_outputs(4563) <= a and not b;
    layer5_outputs(4564) <= b;
    layer5_outputs(4565) <= not (a xor b);
    layer5_outputs(4566) <= not a;
    layer5_outputs(4567) <= not a;
    layer5_outputs(4568) <= '1';
    layer5_outputs(4569) <= b;
    layer5_outputs(4570) <= a and not b;
    layer5_outputs(4571) <= not b or a;
    layer5_outputs(4572) <= not a or b;
    layer5_outputs(4573) <= not b;
    layer5_outputs(4574) <= not (a xor b);
    layer5_outputs(4575) <= a and not b;
    layer5_outputs(4576) <= not (a or b);
    layer5_outputs(4577) <= b and not a;
    layer5_outputs(4578) <= a;
    layer5_outputs(4579) <= a and not b;
    layer5_outputs(4580) <= not a or b;
    layer5_outputs(4581) <= not a or b;
    layer5_outputs(4582) <= a or b;
    layer5_outputs(4583) <= not a;
    layer5_outputs(4584) <= a or b;
    layer5_outputs(4585) <= '1';
    layer5_outputs(4586) <= not a;
    layer5_outputs(4587) <= a and not b;
    layer5_outputs(4588) <= a;
    layer5_outputs(4589) <= b;
    layer5_outputs(4590) <= a;
    layer5_outputs(4591) <= '0';
    layer5_outputs(4592) <= not (a or b);
    layer5_outputs(4593) <= not (a xor b);
    layer5_outputs(4594) <= not a;
    layer5_outputs(4595) <= a and not b;
    layer5_outputs(4596) <= a or b;
    layer5_outputs(4597) <= b and not a;
    layer5_outputs(4598) <= a;
    layer5_outputs(4599) <= a xor b;
    layer5_outputs(4600) <= a and not b;
    layer5_outputs(4601) <= not a;
    layer5_outputs(4602) <= not b;
    layer5_outputs(4603) <= a and not b;
    layer5_outputs(4604) <= a;
    layer5_outputs(4605) <= a;
    layer5_outputs(4606) <= a;
    layer5_outputs(4607) <= not (a or b);
    layer5_outputs(4608) <= not (a and b);
    layer5_outputs(4609) <= not a;
    layer5_outputs(4610) <= b;
    layer5_outputs(4611) <= a;
    layer5_outputs(4612) <= a;
    layer5_outputs(4613) <= not a;
    layer5_outputs(4614) <= a and not b;
    layer5_outputs(4615) <= b;
    layer5_outputs(4616) <= b and not a;
    layer5_outputs(4617) <= a;
    layer5_outputs(4618) <= not b;
    layer5_outputs(4619) <= not a;
    layer5_outputs(4620) <= not (a or b);
    layer5_outputs(4621) <= a;
    layer5_outputs(4622) <= not (a or b);
    layer5_outputs(4623) <= b;
    layer5_outputs(4624) <= a and b;
    layer5_outputs(4625) <= not b or a;
    layer5_outputs(4626) <= b;
    layer5_outputs(4627) <= not b;
    layer5_outputs(4628) <= b;
    layer5_outputs(4629) <= a and b;
    layer5_outputs(4630) <= b;
    layer5_outputs(4631) <= not a or b;
    layer5_outputs(4632) <= '1';
    layer5_outputs(4633) <= not b or a;
    layer5_outputs(4634) <= b and not a;
    layer5_outputs(4635) <= '1';
    layer5_outputs(4636) <= a;
    layer5_outputs(4637) <= a xor b;
    layer5_outputs(4638) <= not b;
    layer5_outputs(4639) <= not b or a;
    layer5_outputs(4640) <= a;
    layer5_outputs(4641) <= not (a and b);
    layer5_outputs(4642) <= not b;
    layer5_outputs(4643) <= not b or a;
    layer5_outputs(4644) <= b and not a;
    layer5_outputs(4645) <= a xor b;
    layer5_outputs(4646) <= not (a or b);
    layer5_outputs(4647) <= b and not a;
    layer5_outputs(4648) <= a and not b;
    layer5_outputs(4649) <= b;
    layer5_outputs(4650) <= not b;
    layer5_outputs(4651) <= b;
    layer5_outputs(4652) <= not b or a;
    layer5_outputs(4653) <= not (a or b);
    layer5_outputs(4654) <= not a;
    layer5_outputs(4655) <= not (a and b);
    layer5_outputs(4656) <= not a;
    layer5_outputs(4657) <= not b;
    layer5_outputs(4658) <= a and b;
    layer5_outputs(4659) <= not a;
    layer5_outputs(4660) <= b and not a;
    layer5_outputs(4661) <= b;
    layer5_outputs(4662) <= a xor b;
    layer5_outputs(4663) <= not a or b;
    layer5_outputs(4664) <= a or b;
    layer5_outputs(4665) <= not a;
    layer5_outputs(4666) <= a or b;
    layer5_outputs(4667) <= b;
    layer5_outputs(4668) <= a and b;
    layer5_outputs(4669) <= not (a xor b);
    layer5_outputs(4670) <= a;
    layer5_outputs(4671) <= a or b;
    layer5_outputs(4672) <= a or b;
    layer5_outputs(4673) <= not a;
    layer5_outputs(4674) <= b and not a;
    layer5_outputs(4675) <= not (a and b);
    layer5_outputs(4676) <= not (a or b);
    layer5_outputs(4677) <= a and not b;
    layer5_outputs(4678) <= a;
    layer5_outputs(4679) <= not b or a;
    layer5_outputs(4680) <= b;
    layer5_outputs(4681) <= not (a or b);
    layer5_outputs(4682) <= b and not a;
    layer5_outputs(4683) <= a;
    layer5_outputs(4684) <= b;
    layer5_outputs(4685) <= a and not b;
    layer5_outputs(4686) <= not b;
    layer5_outputs(4687) <= not (a xor b);
    layer5_outputs(4688) <= b;
    layer5_outputs(4689) <= not a;
    layer5_outputs(4690) <= not (a or b);
    layer5_outputs(4691) <= not b;
    layer5_outputs(4692) <= not (a xor b);
    layer5_outputs(4693) <= not a;
    layer5_outputs(4694) <= '0';
    layer5_outputs(4695) <= b;
    layer5_outputs(4696) <= a;
    layer5_outputs(4697) <= not a or b;
    layer5_outputs(4698) <= not (a and b);
    layer5_outputs(4699) <= not b;
    layer5_outputs(4700) <= not a;
    layer5_outputs(4701) <= not a or b;
    layer5_outputs(4702) <= a and b;
    layer5_outputs(4703) <= not (a and b);
    layer5_outputs(4704) <= a;
    layer5_outputs(4705) <= not b;
    layer5_outputs(4706) <= a xor b;
    layer5_outputs(4707) <= a and b;
    layer5_outputs(4708) <= a and not b;
    layer5_outputs(4709) <= not a;
    layer5_outputs(4710) <= not b;
    layer5_outputs(4711) <= a xor b;
    layer5_outputs(4712) <= b;
    layer5_outputs(4713) <= not (a xor b);
    layer5_outputs(4714) <= not a;
    layer5_outputs(4715) <= a and b;
    layer5_outputs(4716) <= a;
    layer5_outputs(4717) <= not a or b;
    layer5_outputs(4718) <= a and b;
    layer5_outputs(4719) <= not b;
    layer5_outputs(4720) <= a;
    layer5_outputs(4721) <= not a;
    layer5_outputs(4722) <= not b or a;
    layer5_outputs(4723) <= not (a xor b);
    layer5_outputs(4724) <= b;
    layer5_outputs(4725) <= not (a xor b);
    layer5_outputs(4726) <= not b;
    layer5_outputs(4727) <= a and b;
    layer5_outputs(4728) <= not (a and b);
    layer5_outputs(4729) <= not (a or b);
    layer5_outputs(4730) <= not (a or b);
    layer5_outputs(4731) <= b;
    layer5_outputs(4732) <= not a or b;
    layer5_outputs(4733) <= not (a xor b);
    layer5_outputs(4734) <= not a;
    layer5_outputs(4735) <= not a;
    layer5_outputs(4736) <= not (a xor b);
    layer5_outputs(4737) <= a;
    layer5_outputs(4738) <= a xor b;
    layer5_outputs(4739) <= not (a or b);
    layer5_outputs(4740) <= a;
    layer5_outputs(4741) <= b;
    layer5_outputs(4742) <= b;
    layer5_outputs(4743) <= b;
    layer5_outputs(4744) <= a;
    layer5_outputs(4745) <= not a;
    layer5_outputs(4746) <= b;
    layer5_outputs(4747) <= not b;
    layer5_outputs(4748) <= a xor b;
    layer5_outputs(4749) <= a and b;
    layer5_outputs(4750) <= a and b;
    layer5_outputs(4751) <= not a;
    layer5_outputs(4752) <= not b;
    layer5_outputs(4753) <= b and not a;
    layer5_outputs(4754) <= a and b;
    layer5_outputs(4755) <= not b or a;
    layer5_outputs(4756) <= a xor b;
    layer5_outputs(4757) <= b;
    layer5_outputs(4758) <= not (a or b);
    layer5_outputs(4759) <= a;
    layer5_outputs(4760) <= not a or b;
    layer5_outputs(4761) <= not (a or b);
    layer5_outputs(4762) <= not a;
    layer5_outputs(4763) <= not b or a;
    layer5_outputs(4764) <= not a or b;
    layer5_outputs(4765) <= a and b;
    layer5_outputs(4766) <= not (a xor b);
    layer5_outputs(4767) <= not (a or b);
    layer5_outputs(4768) <= b;
    layer5_outputs(4769) <= not b;
    layer5_outputs(4770) <= a and not b;
    layer5_outputs(4771) <= a;
    layer5_outputs(4772) <= b;
    layer5_outputs(4773) <= not a;
    layer5_outputs(4774) <= not a;
    layer5_outputs(4775) <= not a or b;
    layer5_outputs(4776) <= b and not a;
    layer5_outputs(4777) <= b;
    layer5_outputs(4778) <= not (a or b);
    layer5_outputs(4779) <= not b or a;
    layer5_outputs(4780) <= not (a xor b);
    layer5_outputs(4781) <= a and not b;
    layer5_outputs(4782) <= not (a or b);
    layer5_outputs(4783) <= not b or a;
    layer5_outputs(4784) <= not b;
    layer5_outputs(4785) <= not b;
    layer5_outputs(4786) <= b and not a;
    layer5_outputs(4787) <= not a;
    layer5_outputs(4788) <= a;
    layer5_outputs(4789) <= a and not b;
    layer5_outputs(4790) <= not a;
    layer5_outputs(4791) <= a;
    layer5_outputs(4792) <= not (a xor b);
    layer5_outputs(4793) <= b and not a;
    layer5_outputs(4794) <= a xor b;
    layer5_outputs(4795) <= not a;
    layer5_outputs(4796) <= not a;
    layer5_outputs(4797) <= '0';
    layer5_outputs(4798) <= not b;
    layer5_outputs(4799) <= not (a and b);
    layer5_outputs(4800) <= not (a and b);
    layer5_outputs(4801) <= '1';
    layer5_outputs(4802) <= a or b;
    layer5_outputs(4803) <= a and not b;
    layer5_outputs(4804) <= b and not a;
    layer5_outputs(4805) <= not (a and b);
    layer5_outputs(4806) <= a and not b;
    layer5_outputs(4807) <= a;
    layer5_outputs(4808) <= '1';
    layer5_outputs(4809) <= not b;
    layer5_outputs(4810) <= a xor b;
    layer5_outputs(4811) <= a and not b;
    layer5_outputs(4812) <= a;
    layer5_outputs(4813) <= not b;
    layer5_outputs(4814) <= b and not a;
    layer5_outputs(4815) <= a and not b;
    layer5_outputs(4816) <= not (a or b);
    layer5_outputs(4817) <= b and not a;
    layer5_outputs(4818) <= a xor b;
    layer5_outputs(4819) <= b;
    layer5_outputs(4820) <= a or b;
    layer5_outputs(4821) <= b and not a;
    layer5_outputs(4822) <= not b;
    layer5_outputs(4823) <= b;
    layer5_outputs(4824) <= a and not b;
    layer5_outputs(4825) <= '1';
    layer5_outputs(4826) <= a;
    layer5_outputs(4827) <= not b;
    layer5_outputs(4828) <= a;
    layer5_outputs(4829) <= a;
    layer5_outputs(4830) <= not (a and b);
    layer5_outputs(4831) <= '0';
    layer5_outputs(4832) <= not a;
    layer5_outputs(4833) <= not b;
    layer5_outputs(4834) <= a;
    layer5_outputs(4835) <= not a;
    layer5_outputs(4836) <= not b;
    layer5_outputs(4837) <= not a;
    layer5_outputs(4838) <= a and b;
    layer5_outputs(4839) <= b and not a;
    layer5_outputs(4840) <= a or b;
    layer5_outputs(4841) <= b;
    layer5_outputs(4842) <= '1';
    layer5_outputs(4843) <= not (a xor b);
    layer5_outputs(4844) <= b;
    layer5_outputs(4845) <= b;
    layer5_outputs(4846) <= not (a and b);
    layer5_outputs(4847) <= not b or a;
    layer5_outputs(4848) <= not (a xor b);
    layer5_outputs(4849) <= a and b;
    layer5_outputs(4850) <= not a;
    layer5_outputs(4851) <= a;
    layer5_outputs(4852) <= '1';
    layer5_outputs(4853) <= a and b;
    layer5_outputs(4854) <= a or b;
    layer5_outputs(4855) <= not a or b;
    layer5_outputs(4856) <= b;
    layer5_outputs(4857) <= not b or a;
    layer5_outputs(4858) <= not b;
    layer5_outputs(4859) <= a;
    layer5_outputs(4860) <= b;
    layer5_outputs(4861) <= not (a and b);
    layer5_outputs(4862) <= b;
    layer5_outputs(4863) <= b;
    layer5_outputs(4864) <= a xor b;
    layer5_outputs(4865) <= not b;
    layer5_outputs(4866) <= b;
    layer5_outputs(4867) <= a;
    layer5_outputs(4868) <= not (a xor b);
    layer5_outputs(4869) <= not b;
    layer5_outputs(4870) <= not b or a;
    layer5_outputs(4871) <= b;
    layer5_outputs(4872) <= not b;
    layer5_outputs(4873) <= not b;
    layer5_outputs(4874) <= b and not a;
    layer5_outputs(4875) <= b and not a;
    layer5_outputs(4876) <= not b;
    layer5_outputs(4877) <= not (a xor b);
    layer5_outputs(4878) <= a or b;
    layer5_outputs(4879) <= a or b;
    layer5_outputs(4880) <= a and not b;
    layer5_outputs(4881) <= not b;
    layer5_outputs(4882) <= not b;
    layer5_outputs(4883) <= b and not a;
    layer5_outputs(4884) <= not (a and b);
    layer5_outputs(4885) <= not b or a;
    layer5_outputs(4886) <= a xor b;
    layer5_outputs(4887) <= b and not a;
    layer5_outputs(4888) <= b;
    layer5_outputs(4889) <= a or b;
    layer5_outputs(4890) <= not a;
    layer5_outputs(4891) <= a xor b;
    layer5_outputs(4892) <= a and b;
    layer5_outputs(4893) <= a;
    layer5_outputs(4894) <= not b;
    layer5_outputs(4895) <= not (a or b);
    layer5_outputs(4896) <= b;
    layer5_outputs(4897) <= not b or a;
    layer5_outputs(4898) <= a xor b;
    layer5_outputs(4899) <= not (a xor b);
    layer5_outputs(4900) <= not b or a;
    layer5_outputs(4901) <= a;
    layer5_outputs(4902) <= a;
    layer5_outputs(4903) <= not (a xor b);
    layer5_outputs(4904) <= a;
    layer5_outputs(4905) <= a xor b;
    layer5_outputs(4906) <= a;
    layer5_outputs(4907) <= not a;
    layer5_outputs(4908) <= a xor b;
    layer5_outputs(4909) <= a and not b;
    layer5_outputs(4910) <= not b;
    layer5_outputs(4911) <= not b;
    layer5_outputs(4912) <= not a;
    layer5_outputs(4913) <= not a or b;
    layer5_outputs(4914) <= not b;
    layer5_outputs(4915) <= not b or a;
    layer5_outputs(4916) <= '0';
    layer5_outputs(4917) <= a and not b;
    layer5_outputs(4918) <= b;
    layer5_outputs(4919) <= b;
    layer5_outputs(4920) <= a;
    layer5_outputs(4921) <= not b or a;
    layer5_outputs(4922) <= b;
    layer5_outputs(4923) <= not b;
    layer5_outputs(4924) <= '1';
    layer5_outputs(4925) <= a and b;
    layer5_outputs(4926) <= not b;
    layer5_outputs(4927) <= b and not a;
    layer5_outputs(4928) <= b and not a;
    layer5_outputs(4929) <= a;
    layer5_outputs(4930) <= a;
    layer5_outputs(4931) <= a and b;
    layer5_outputs(4932) <= a and b;
    layer5_outputs(4933) <= b;
    layer5_outputs(4934) <= a;
    layer5_outputs(4935) <= not (a or b);
    layer5_outputs(4936) <= b;
    layer5_outputs(4937) <= not b or a;
    layer5_outputs(4938) <= b;
    layer5_outputs(4939) <= not a;
    layer5_outputs(4940) <= a;
    layer5_outputs(4941) <= not b;
    layer5_outputs(4942) <= b and not a;
    layer5_outputs(4943) <= b;
    layer5_outputs(4944) <= not (a xor b);
    layer5_outputs(4945) <= b and not a;
    layer5_outputs(4946) <= not b;
    layer5_outputs(4947) <= not b;
    layer5_outputs(4948) <= not b or a;
    layer5_outputs(4949) <= a and not b;
    layer5_outputs(4950) <= not b or a;
    layer5_outputs(4951) <= not (a xor b);
    layer5_outputs(4952) <= '0';
    layer5_outputs(4953) <= a or b;
    layer5_outputs(4954) <= not a or b;
    layer5_outputs(4955) <= '0';
    layer5_outputs(4956) <= a and not b;
    layer5_outputs(4957) <= a and not b;
    layer5_outputs(4958) <= a and b;
    layer5_outputs(4959) <= not (a xor b);
    layer5_outputs(4960) <= not a;
    layer5_outputs(4961) <= '1';
    layer5_outputs(4962) <= b and not a;
    layer5_outputs(4963) <= not b or a;
    layer5_outputs(4964) <= not (a xor b);
    layer5_outputs(4965) <= '1';
    layer5_outputs(4966) <= b and not a;
    layer5_outputs(4967) <= a and not b;
    layer5_outputs(4968) <= a xor b;
    layer5_outputs(4969) <= not (a and b);
    layer5_outputs(4970) <= a;
    layer5_outputs(4971) <= not b or a;
    layer5_outputs(4972) <= b and not a;
    layer5_outputs(4973) <= a and b;
    layer5_outputs(4974) <= not a;
    layer5_outputs(4975) <= a xor b;
    layer5_outputs(4976) <= not (a xor b);
    layer5_outputs(4977) <= not a;
    layer5_outputs(4978) <= not b;
    layer5_outputs(4979) <= not (a xor b);
    layer5_outputs(4980) <= not (a and b);
    layer5_outputs(4981) <= '1';
    layer5_outputs(4982) <= a xor b;
    layer5_outputs(4983) <= not (a xor b);
    layer5_outputs(4984) <= a;
    layer5_outputs(4985) <= not a;
    layer5_outputs(4986) <= a xor b;
    layer5_outputs(4987) <= not b;
    layer5_outputs(4988) <= not b or a;
    layer5_outputs(4989) <= a or b;
    layer5_outputs(4990) <= not (a and b);
    layer5_outputs(4991) <= not a;
    layer5_outputs(4992) <= not b;
    layer5_outputs(4993) <= not b;
    layer5_outputs(4994) <= a xor b;
    layer5_outputs(4995) <= not a;
    layer5_outputs(4996) <= not (a xor b);
    layer5_outputs(4997) <= a and not b;
    layer5_outputs(4998) <= not b;
    layer5_outputs(4999) <= not b or a;
    layer5_outputs(5000) <= '1';
    layer5_outputs(5001) <= not b;
    layer5_outputs(5002) <= b and not a;
    layer5_outputs(5003) <= not (a xor b);
    layer5_outputs(5004) <= not (a xor b);
    layer5_outputs(5005) <= b and not a;
    layer5_outputs(5006) <= a or b;
    layer5_outputs(5007) <= a and b;
    layer5_outputs(5008) <= not a;
    layer5_outputs(5009) <= not b;
    layer5_outputs(5010) <= b;
    layer5_outputs(5011) <= '1';
    layer5_outputs(5012) <= b and not a;
    layer5_outputs(5013) <= '0';
    layer5_outputs(5014) <= not (a xor b);
    layer5_outputs(5015) <= not b or a;
    layer5_outputs(5016) <= a xor b;
    layer5_outputs(5017) <= not b;
    layer5_outputs(5018) <= a xor b;
    layer5_outputs(5019) <= a;
    layer5_outputs(5020) <= a;
    layer5_outputs(5021) <= not a;
    layer5_outputs(5022) <= a and b;
    layer5_outputs(5023) <= not a or b;
    layer5_outputs(5024) <= a;
    layer5_outputs(5025) <= a;
    layer5_outputs(5026) <= not (a xor b);
    layer5_outputs(5027) <= b;
    layer5_outputs(5028) <= a and b;
    layer5_outputs(5029) <= a xor b;
    layer5_outputs(5030) <= b;
    layer5_outputs(5031) <= not (a xor b);
    layer5_outputs(5032) <= b;
    layer5_outputs(5033) <= a;
    layer5_outputs(5034) <= b;
    layer5_outputs(5035) <= not (a or b);
    layer5_outputs(5036) <= '1';
    layer5_outputs(5037) <= not a;
    layer5_outputs(5038) <= not (a or b);
    layer5_outputs(5039) <= a and b;
    layer5_outputs(5040) <= not (a or b);
    layer5_outputs(5041) <= not (a and b);
    layer5_outputs(5042) <= a xor b;
    layer5_outputs(5043) <= not (a or b);
    layer5_outputs(5044) <= not a or b;
    layer5_outputs(5045) <= not b;
    layer5_outputs(5046) <= b;
    layer5_outputs(5047) <= b and not a;
    layer5_outputs(5048) <= b;
    layer5_outputs(5049) <= not a;
    layer5_outputs(5050) <= not (a or b);
    layer5_outputs(5051) <= not (a or b);
    layer5_outputs(5052) <= a;
    layer5_outputs(5053) <= a xor b;
    layer5_outputs(5054) <= a and b;
    layer5_outputs(5055) <= a xor b;
    layer5_outputs(5056) <= a xor b;
    layer5_outputs(5057) <= a;
    layer5_outputs(5058) <= not a;
    layer5_outputs(5059) <= not (a xor b);
    layer5_outputs(5060) <= a;
    layer5_outputs(5061) <= '0';
    layer5_outputs(5062) <= b;
    layer5_outputs(5063) <= not b;
    layer5_outputs(5064) <= not a or b;
    layer5_outputs(5065) <= a xor b;
    layer5_outputs(5066) <= b;
    layer5_outputs(5067) <= a xor b;
    layer5_outputs(5068) <= not a or b;
    layer5_outputs(5069) <= not a;
    layer5_outputs(5070) <= not b;
    layer5_outputs(5071) <= not a or b;
    layer5_outputs(5072) <= b;
    layer5_outputs(5073) <= not a;
    layer5_outputs(5074) <= not a;
    layer5_outputs(5075) <= a or b;
    layer5_outputs(5076) <= a and b;
    layer5_outputs(5077) <= not (a xor b);
    layer5_outputs(5078) <= not (a or b);
    layer5_outputs(5079) <= a and not b;
    layer5_outputs(5080) <= not (a or b);
    layer5_outputs(5081) <= not a;
    layer5_outputs(5082) <= not b;
    layer5_outputs(5083) <= not b or a;
    layer5_outputs(5084) <= b and not a;
    layer5_outputs(5085) <= a xor b;
    layer5_outputs(5086) <= not b;
    layer5_outputs(5087) <= not b or a;
    layer5_outputs(5088) <= not a or b;
    layer5_outputs(5089) <= a;
    layer5_outputs(5090) <= a and not b;
    layer5_outputs(5091) <= not a;
    layer5_outputs(5092) <= a xor b;
    layer5_outputs(5093) <= not b or a;
    layer5_outputs(5094) <= a and not b;
    layer5_outputs(5095) <= not a;
    layer5_outputs(5096) <= not b;
    layer5_outputs(5097) <= not a;
    layer5_outputs(5098) <= b;
    layer5_outputs(5099) <= not (a and b);
    layer5_outputs(5100) <= not (a or b);
    layer5_outputs(5101) <= '0';
    layer5_outputs(5102) <= '0';
    layer5_outputs(5103) <= not b;
    layer5_outputs(5104) <= b;
    layer5_outputs(5105) <= not (a and b);
    layer5_outputs(5106) <= a xor b;
    layer5_outputs(5107) <= b and not a;
    layer5_outputs(5108) <= b and not a;
    layer5_outputs(5109) <= not b or a;
    layer5_outputs(5110) <= a or b;
    layer5_outputs(5111) <= a xor b;
    layer5_outputs(5112) <= a or b;
    layer5_outputs(5113) <= a;
    layer5_outputs(5114) <= b and not a;
    layer5_outputs(5115) <= not b;
    layer5_outputs(5116) <= not a;
    layer5_outputs(5117) <= a;
    layer5_outputs(5118) <= not (a xor b);
    layer5_outputs(5119) <= a and b;
    layer5_outputs(5120) <= b;
    layer5_outputs(5121) <= b and not a;
    layer5_outputs(5122) <= not (a or b);
    layer5_outputs(5123) <= not (a or b);
    layer5_outputs(5124) <= b;
    layer5_outputs(5125) <= not b;
    layer5_outputs(5126) <= b and not a;
    layer5_outputs(5127) <= a and b;
    layer5_outputs(5128) <= b;
    layer5_outputs(5129) <= a xor b;
    layer5_outputs(5130) <= a and not b;
    layer5_outputs(5131) <= not b;
    layer5_outputs(5132) <= not a;
    layer5_outputs(5133) <= b and not a;
    layer5_outputs(5134) <= '0';
    layer5_outputs(5135) <= b;
    layer5_outputs(5136) <= b;
    layer5_outputs(5137) <= not (a and b);
    layer5_outputs(5138) <= not b;
    layer5_outputs(5139) <= b and not a;
    layer5_outputs(5140) <= a and not b;
    layer5_outputs(5141) <= a or b;
    layer5_outputs(5142) <= not a or b;
    layer5_outputs(5143) <= not b or a;
    layer5_outputs(5144) <= b;
    layer5_outputs(5145) <= not b;
    layer5_outputs(5146) <= not a;
    layer5_outputs(5147) <= b;
    layer5_outputs(5148) <= not b or a;
    layer5_outputs(5149) <= not a;
    layer5_outputs(5150) <= a and not b;
    layer5_outputs(5151) <= b;
    layer5_outputs(5152) <= '0';
    layer5_outputs(5153) <= not (a xor b);
    layer5_outputs(5154) <= a and b;
    layer5_outputs(5155) <= not a;
    layer5_outputs(5156) <= not (a xor b);
    layer5_outputs(5157) <= b and not a;
    layer5_outputs(5158) <= a or b;
    layer5_outputs(5159) <= a;
    layer5_outputs(5160) <= b;
    layer5_outputs(5161) <= not b;
    layer5_outputs(5162) <= b;
    layer5_outputs(5163) <= '0';
    layer5_outputs(5164) <= not b;
    layer5_outputs(5165) <= a;
    layer5_outputs(5166) <= '1';
    layer5_outputs(5167) <= a;
    layer5_outputs(5168) <= not (a or b);
    layer5_outputs(5169) <= not b;
    layer5_outputs(5170) <= a;
    layer5_outputs(5171) <= not b;
    layer5_outputs(5172) <= not b;
    layer5_outputs(5173) <= b;
    layer5_outputs(5174) <= a and b;
    layer5_outputs(5175) <= not a;
    layer5_outputs(5176) <= not b;
    layer5_outputs(5177) <= not b or a;
    layer5_outputs(5178) <= a xor b;
    layer5_outputs(5179) <= a;
    layer5_outputs(5180) <= a and not b;
    layer5_outputs(5181) <= a and b;
    layer5_outputs(5182) <= b;
    layer5_outputs(5183) <= not b;
    layer5_outputs(5184) <= b and not a;
    layer5_outputs(5185) <= not (a and b);
    layer5_outputs(5186) <= a xor b;
    layer5_outputs(5187) <= not b;
    layer5_outputs(5188) <= not (a xor b);
    layer5_outputs(5189) <= not b or a;
    layer5_outputs(5190) <= '1';
    layer5_outputs(5191) <= b;
    layer5_outputs(5192) <= not b or a;
    layer5_outputs(5193) <= a and not b;
    layer5_outputs(5194) <= a;
    layer5_outputs(5195) <= not b or a;
    layer5_outputs(5196) <= a xor b;
    layer5_outputs(5197) <= a xor b;
    layer5_outputs(5198) <= not a or b;
    layer5_outputs(5199) <= '0';
    layer5_outputs(5200) <= a;
    layer5_outputs(5201) <= b;
    layer5_outputs(5202) <= not (a or b);
    layer5_outputs(5203) <= not b;
    layer5_outputs(5204) <= a or b;
    layer5_outputs(5205) <= b;
    layer5_outputs(5206) <= a;
    layer5_outputs(5207) <= a xor b;
    layer5_outputs(5208) <= not b;
    layer5_outputs(5209) <= not a;
    layer5_outputs(5210) <= not b;
    layer5_outputs(5211) <= not (a xor b);
    layer5_outputs(5212) <= b and not a;
    layer5_outputs(5213) <= not a;
    layer5_outputs(5214) <= not b;
    layer5_outputs(5215) <= not b;
    layer5_outputs(5216) <= not b;
    layer5_outputs(5217) <= a;
    layer5_outputs(5218) <= a;
    layer5_outputs(5219) <= not (a or b);
    layer5_outputs(5220) <= not b or a;
    layer5_outputs(5221) <= b;
    layer5_outputs(5222) <= not (a or b);
    layer5_outputs(5223) <= a and not b;
    layer5_outputs(5224) <= not (a or b);
    layer5_outputs(5225) <= not b;
    layer5_outputs(5226) <= not a;
    layer5_outputs(5227) <= a and not b;
    layer5_outputs(5228) <= a and b;
    layer5_outputs(5229) <= not (a xor b);
    layer5_outputs(5230) <= not a;
    layer5_outputs(5231) <= not a or b;
    layer5_outputs(5232) <= not b;
    layer5_outputs(5233) <= not (a or b);
    layer5_outputs(5234) <= a or b;
    layer5_outputs(5235) <= a or b;
    layer5_outputs(5236) <= not b;
    layer5_outputs(5237) <= b and not a;
    layer5_outputs(5238) <= not (a or b);
    layer5_outputs(5239) <= not a or b;
    layer5_outputs(5240) <= '1';
    layer5_outputs(5241) <= not (a xor b);
    layer5_outputs(5242) <= b;
    layer5_outputs(5243) <= not a or b;
    layer5_outputs(5244) <= a and b;
    layer5_outputs(5245) <= not (a and b);
    layer5_outputs(5246) <= a;
    layer5_outputs(5247) <= a xor b;
    layer5_outputs(5248) <= not (a xor b);
    layer5_outputs(5249) <= a;
    layer5_outputs(5250) <= not b;
    layer5_outputs(5251) <= b and not a;
    layer5_outputs(5252) <= b;
    layer5_outputs(5253) <= a xor b;
    layer5_outputs(5254) <= b and not a;
    layer5_outputs(5255) <= not (a xor b);
    layer5_outputs(5256) <= a;
    layer5_outputs(5257) <= a xor b;
    layer5_outputs(5258) <= not (a or b);
    layer5_outputs(5259) <= not b;
    layer5_outputs(5260) <= b;
    layer5_outputs(5261) <= b;
    layer5_outputs(5262) <= b;
    layer5_outputs(5263) <= not a;
    layer5_outputs(5264) <= a;
    layer5_outputs(5265) <= not a;
    layer5_outputs(5266) <= a xor b;
    layer5_outputs(5267) <= not (a xor b);
    layer5_outputs(5268) <= not b;
    layer5_outputs(5269) <= not b;
    layer5_outputs(5270) <= not (a or b);
    layer5_outputs(5271) <= b;
    layer5_outputs(5272) <= not b;
    layer5_outputs(5273) <= a or b;
    layer5_outputs(5274) <= a or b;
    layer5_outputs(5275) <= a or b;
    layer5_outputs(5276) <= not a;
    layer5_outputs(5277) <= a and not b;
    layer5_outputs(5278) <= not b;
    layer5_outputs(5279) <= a;
    layer5_outputs(5280) <= a xor b;
    layer5_outputs(5281) <= a or b;
    layer5_outputs(5282) <= not (a or b);
    layer5_outputs(5283) <= not b or a;
    layer5_outputs(5284) <= b and not a;
    layer5_outputs(5285) <= a;
    layer5_outputs(5286) <= not b;
    layer5_outputs(5287) <= a;
    layer5_outputs(5288) <= b;
    layer5_outputs(5289) <= a;
    layer5_outputs(5290) <= a and b;
    layer5_outputs(5291) <= a;
    layer5_outputs(5292) <= b and not a;
    layer5_outputs(5293) <= b;
    layer5_outputs(5294) <= a;
    layer5_outputs(5295) <= a;
    layer5_outputs(5296) <= not a;
    layer5_outputs(5297) <= a;
    layer5_outputs(5298) <= a and b;
    layer5_outputs(5299) <= '0';
    layer5_outputs(5300) <= not a;
    layer5_outputs(5301) <= not a or b;
    layer5_outputs(5302) <= not a;
    layer5_outputs(5303) <= not b or a;
    layer5_outputs(5304) <= '0';
    layer5_outputs(5305) <= not a;
    layer5_outputs(5306) <= not b or a;
    layer5_outputs(5307) <= not (a xor b);
    layer5_outputs(5308) <= b and not a;
    layer5_outputs(5309) <= not (a xor b);
    layer5_outputs(5310) <= a and not b;
    layer5_outputs(5311) <= a and not b;
    layer5_outputs(5312) <= b;
    layer5_outputs(5313) <= not (a xor b);
    layer5_outputs(5314) <= not a;
    layer5_outputs(5315) <= a and b;
    layer5_outputs(5316) <= not (a or b);
    layer5_outputs(5317) <= a and b;
    layer5_outputs(5318) <= a;
    layer5_outputs(5319) <= a xor b;
    layer5_outputs(5320) <= not b;
    layer5_outputs(5321) <= not a;
    layer5_outputs(5322) <= not (a or b);
    layer5_outputs(5323) <= not b;
    layer5_outputs(5324) <= a;
    layer5_outputs(5325) <= not a;
    layer5_outputs(5326) <= not a;
    layer5_outputs(5327) <= a and b;
    layer5_outputs(5328) <= a or b;
    layer5_outputs(5329) <= b;
    layer5_outputs(5330) <= not (a xor b);
    layer5_outputs(5331) <= a or b;
    layer5_outputs(5332) <= b and not a;
    layer5_outputs(5333) <= not a;
    layer5_outputs(5334) <= not a or b;
    layer5_outputs(5335) <= not (a and b);
    layer5_outputs(5336) <= not a;
    layer5_outputs(5337) <= a;
    layer5_outputs(5338) <= not b;
    layer5_outputs(5339) <= not (a and b);
    layer5_outputs(5340) <= b;
    layer5_outputs(5341) <= not b or a;
    layer5_outputs(5342) <= a and not b;
    layer5_outputs(5343) <= a;
    layer5_outputs(5344) <= not a;
    layer5_outputs(5345) <= b;
    layer5_outputs(5346) <= not (a xor b);
    layer5_outputs(5347) <= b and not a;
    layer5_outputs(5348) <= not a;
    layer5_outputs(5349) <= a and b;
    layer5_outputs(5350) <= '1';
    layer5_outputs(5351) <= not a;
    layer5_outputs(5352) <= not (a or b);
    layer5_outputs(5353) <= a;
    layer5_outputs(5354) <= a and not b;
    layer5_outputs(5355) <= not a or b;
    layer5_outputs(5356) <= b and not a;
    layer5_outputs(5357) <= not a;
    layer5_outputs(5358) <= b;
    layer5_outputs(5359) <= b and not a;
    layer5_outputs(5360) <= not (a or b);
    layer5_outputs(5361) <= '0';
    layer5_outputs(5362) <= a;
    layer5_outputs(5363) <= a or b;
    layer5_outputs(5364) <= not (a xor b);
    layer5_outputs(5365) <= not a;
    layer5_outputs(5366) <= '1';
    layer5_outputs(5367) <= b;
    layer5_outputs(5368) <= a and b;
    layer5_outputs(5369) <= a and not b;
    layer5_outputs(5370) <= b and not a;
    layer5_outputs(5371) <= b;
    layer5_outputs(5372) <= not (a xor b);
    layer5_outputs(5373) <= b;
    layer5_outputs(5374) <= not a;
    layer5_outputs(5375) <= not a or b;
    layer5_outputs(5376) <= not b;
    layer5_outputs(5377) <= not b or a;
    layer5_outputs(5378) <= '1';
    layer5_outputs(5379) <= not (a xor b);
    layer5_outputs(5380) <= a and b;
    layer5_outputs(5381) <= not a or b;
    layer5_outputs(5382) <= not b;
    layer5_outputs(5383) <= not a;
    layer5_outputs(5384) <= a or b;
    layer5_outputs(5385) <= a;
    layer5_outputs(5386) <= '1';
    layer5_outputs(5387) <= '0';
    layer5_outputs(5388) <= not a;
    layer5_outputs(5389) <= b and not a;
    layer5_outputs(5390) <= a or b;
    layer5_outputs(5391) <= not b;
    layer5_outputs(5392) <= a or b;
    layer5_outputs(5393) <= not (a and b);
    layer5_outputs(5394) <= a xor b;
    layer5_outputs(5395) <= not b or a;
    layer5_outputs(5396) <= '1';
    layer5_outputs(5397) <= not (a and b);
    layer5_outputs(5398) <= a xor b;
    layer5_outputs(5399) <= not (a xor b);
    layer5_outputs(5400) <= a and b;
    layer5_outputs(5401) <= not b;
    layer5_outputs(5402) <= not b;
    layer5_outputs(5403) <= a;
    layer5_outputs(5404) <= b and not a;
    layer5_outputs(5405) <= not a;
    layer5_outputs(5406) <= not (a or b);
    layer5_outputs(5407) <= '1';
    layer5_outputs(5408) <= a and not b;
    layer5_outputs(5409) <= not (a or b);
    layer5_outputs(5410) <= a or b;
    layer5_outputs(5411) <= b;
    layer5_outputs(5412) <= a and not b;
    layer5_outputs(5413) <= a xor b;
    layer5_outputs(5414) <= a;
    layer5_outputs(5415) <= not a;
    layer5_outputs(5416) <= b and not a;
    layer5_outputs(5417) <= a and not b;
    layer5_outputs(5418) <= b;
    layer5_outputs(5419) <= b;
    layer5_outputs(5420) <= b;
    layer5_outputs(5421) <= not a;
    layer5_outputs(5422) <= a;
    layer5_outputs(5423) <= a or b;
    layer5_outputs(5424) <= not (a or b);
    layer5_outputs(5425) <= b and not a;
    layer5_outputs(5426) <= not (a or b);
    layer5_outputs(5427) <= a and b;
    layer5_outputs(5428) <= a and b;
    layer5_outputs(5429) <= not (a xor b);
    layer5_outputs(5430) <= a xor b;
    layer5_outputs(5431) <= not a;
    layer5_outputs(5432) <= not a or b;
    layer5_outputs(5433) <= not a;
    layer5_outputs(5434) <= not a;
    layer5_outputs(5435) <= a;
    layer5_outputs(5436) <= a;
    layer5_outputs(5437) <= a or b;
    layer5_outputs(5438) <= b and not a;
    layer5_outputs(5439) <= not b;
    layer5_outputs(5440) <= not b;
    layer5_outputs(5441) <= '1';
    layer5_outputs(5442) <= not a or b;
    layer5_outputs(5443) <= a and b;
    layer5_outputs(5444) <= b and not a;
    layer5_outputs(5445) <= b;
    layer5_outputs(5446) <= not (a and b);
    layer5_outputs(5447) <= b;
    layer5_outputs(5448) <= a or b;
    layer5_outputs(5449) <= not b;
    layer5_outputs(5450) <= not a or b;
    layer5_outputs(5451) <= not (a xor b);
    layer5_outputs(5452) <= not (a xor b);
    layer5_outputs(5453) <= not (a xor b);
    layer5_outputs(5454) <= a xor b;
    layer5_outputs(5455) <= not (a and b);
    layer5_outputs(5456) <= a;
    layer5_outputs(5457) <= a xor b;
    layer5_outputs(5458) <= a and b;
    layer5_outputs(5459) <= not a;
    layer5_outputs(5460) <= not a;
    layer5_outputs(5461) <= b;
    layer5_outputs(5462) <= a or b;
    layer5_outputs(5463) <= not b;
    layer5_outputs(5464) <= b and not a;
    layer5_outputs(5465) <= not a or b;
    layer5_outputs(5466) <= a xor b;
    layer5_outputs(5467) <= a;
    layer5_outputs(5468) <= a xor b;
    layer5_outputs(5469) <= b;
    layer5_outputs(5470) <= not b;
    layer5_outputs(5471) <= not a;
    layer5_outputs(5472) <= not b or a;
    layer5_outputs(5473) <= b;
    layer5_outputs(5474) <= not a or b;
    layer5_outputs(5475) <= a and not b;
    layer5_outputs(5476) <= not a or b;
    layer5_outputs(5477) <= not b;
    layer5_outputs(5478) <= not b;
    layer5_outputs(5479) <= not a;
    layer5_outputs(5480) <= a or b;
    layer5_outputs(5481) <= not (a xor b);
    layer5_outputs(5482) <= not (a xor b);
    layer5_outputs(5483) <= not (a xor b);
    layer5_outputs(5484) <= not a;
    layer5_outputs(5485) <= b;
    layer5_outputs(5486) <= not (a or b);
    layer5_outputs(5487) <= not a;
    layer5_outputs(5488) <= a and b;
    layer5_outputs(5489) <= a;
    layer5_outputs(5490) <= not (a and b);
    layer5_outputs(5491) <= not (a xor b);
    layer5_outputs(5492) <= a and b;
    layer5_outputs(5493) <= not a;
    layer5_outputs(5494) <= not b;
    layer5_outputs(5495) <= a;
    layer5_outputs(5496) <= a and not b;
    layer5_outputs(5497) <= a xor b;
    layer5_outputs(5498) <= b;
    layer5_outputs(5499) <= not (a or b);
    layer5_outputs(5500) <= a;
    layer5_outputs(5501) <= not a;
    layer5_outputs(5502) <= a or b;
    layer5_outputs(5503) <= not b or a;
    layer5_outputs(5504) <= a and not b;
    layer5_outputs(5505) <= not b;
    layer5_outputs(5506) <= not a;
    layer5_outputs(5507) <= not b;
    layer5_outputs(5508) <= a and not b;
    layer5_outputs(5509) <= a and b;
    layer5_outputs(5510) <= not b;
    layer5_outputs(5511) <= not (a xor b);
    layer5_outputs(5512) <= a and not b;
    layer5_outputs(5513) <= b;
    layer5_outputs(5514) <= b;
    layer5_outputs(5515) <= not a or b;
    layer5_outputs(5516) <= a or b;
    layer5_outputs(5517) <= not (a and b);
    layer5_outputs(5518) <= a or b;
    layer5_outputs(5519) <= b;
    layer5_outputs(5520) <= '0';
    layer5_outputs(5521) <= a xor b;
    layer5_outputs(5522) <= not (a and b);
    layer5_outputs(5523) <= a and b;
    layer5_outputs(5524) <= b and not a;
    layer5_outputs(5525) <= a and not b;
    layer5_outputs(5526) <= b and not a;
    layer5_outputs(5527) <= not (a and b);
    layer5_outputs(5528) <= not b or a;
    layer5_outputs(5529) <= not (a or b);
    layer5_outputs(5530) <= a and b;
    layer5_outputs(5531) <= not b;
    layer5_outputs(5532) <= not (a or b);
    layer5_outputs(5533) <= a and not b;
    layer5_outputs(5534) <= b;
    layer5_outputs(5535) <= not (a xor b);
    layer5_outputs(5536) <= a and b;
    layer5_outputs(5537) <= a xor b;
    layer5_outputs(5538) <= b;
    layer5_outputs(5539) <= b;
    layer5_outputs(5540) <= not b or a;
    layer5_outputs(5541) <= b;
    layer5_outputs(5542) <= b;
    layer5_outputs(5543) <= a;
    layer5_outputs(5544) <= b;
    layer5_outputs(5545) <= not (a or b);
    layer5_outputs(5546) <= b;
    layer5_outputs(5547) <= b;
    layer5_outputs(5548) <= not (a xor b);
    layer5_outputs(5549) <= not a or b;
    layer5_outputs(5550) <= not (a or b);
    layer5_outputs(5551) <= not a or b;
    layer5_outputs(5552) <= not a;
    layer5_outputs(5553) <= a and not b;
    layer5_outputs(5554) <= a or b;
    layer5_outputs(5555) <= not (a xor b);
    layer5_outputs(5556) <= not (a and b);
    layer5_outputs(5557) <= a and not b;
    layer5_outputs(5558) <= not a;
    layer5_outputs(5559) <= a and b;
    layer5_outputs(5560) <= a;
    layer5_outputs(5561) <= not b;
    layer5_outputs(5562) <= a;
    layer5_outputs(5563) <= a;
    layer5_outputs(5564) <= a or b;
    layer5_outputs(5565) <= b and not a;
    layer5_outputs(5566) <= not b;
    layer5_outputs(5567) <= a;
    layer5_outputs(5568) <= not a or b;
    layer5_outputs(5569) <= a;
    layer5_outputs(5570) <= a and not b;
    layer5_outputs(5571) <= b;
    layer5_outputs(5572) <= a;
    layer5_outputs(5573) <= a xor b;
    layer5_outputs(5574) <= a and not b;
    layer5_outputs(5575) <= a and not b;
    layer5_outputs(5576) <= not (a and b);
    layer5_outputs(5577) <= a or b;
    layer5_outputs(5578) <= not b;
    layer5_outputs(5579) <= a and b;
    layer5_outputs(5580) <= b;
    layer5_outputs(5581) <= not (a xor b);
    layer5_outputs(5582) <= a or b;
    layer5_outputs(5583) <= a and not b;
    layer5_outputs(5584) <= '0';
    layer5_outputs(5585) <= a and not b;
    layer5_outputs(5586) <= b;
    layer5_outputs(5587) <= '0';
    layer5_outputs(5588) <= not a or b;
    layer5_outputs(5589) <= not a or b;
    layer5_outputs(5590) <= a xor b;
    layer5_outputs(5591) <= not a or b;
    layer5_outputs(5592) <= a xor b;
    layer5_outputs(5593) <= not b;
    layer5_outputs(5594) <= a and b;
    layer5_outputs(5595) <= a;
    layer5_outputs(5596) <= b;
    layer5_outputs(5597) <= not (a and b);
    layer5_outputs(5598) <= a;
    layer5_outputs(5599) <= not a;
    layer5_outputs(5600) <= not (a xor b);
    layer5_outputs(5601) <= not (a and b);
    layer5_outputs(5602) <= b;
    layer5_outputs(5603) <= not a;
    layer5_outputs(5604) <= a or b;
    layer5_outputs(5605) <= not b;
    layer5_outputs(5606) <= not b;
    layer5_outputs(5607) <= b;
    layer5_outputs(5608) <= b;
    layer5_outputs(5609) <= not b;
    layer5_outputs(5610) <= a;
    layer5_outputs(5611) <= b;
    layer5_outputs(5612) <= a xor b;
    layer5_outputs(5613) <= a and not b;
    layer5_outputs(5614) <= b;
    layer5_outputs(5615) <= a;
    layer5_outputs(5616) <= not (a xor b);
    layer5_outputs(5617) <= a;
    layer5_outputs(5618) <= not a or b;
    layer5_outputs(5619) <= not a;
    layer5_outputs(5620) <= not (a and b);
    layer5_outputs(5621) <= not (a or b);
    layer5_outputs(5622) <= not a;
    layer5_outputs(5623) <= a xor b;
    layer5_outputs(5624) <= a xor b;
    layer5_outputs(5625) <= a and not b;
    layer5_outputs(5626) <= not (a xor b);
    layer5_outputs(5627) <= '0';
    layer5_outputs(5628) <= not b or a;
    layer5_outputs(5629) <= a;
    layer5_outputs(5630) <= a or b;
    layer5_outputs(5631) <= not (a xor b);
    layer5_outputs(5632) <= a xor b;
    layer5_outputs(5633) <= not (a and b);
    layer5_outputs(5634) <= not a or b;
    layer5_outputs(5635) <= not a or b;
    layer5_outputs(5636) <= not a;
    layer5_outputs(5637) <= not a;
    layer5_outputs(5638) <= not (a and b);
    layer5_outputs(5639) <= not (a or b);
    layer5_outputs(5640) <= not a;
    layer5_outputs(5641) <= not b;
    layer5_outputs(5642) <= not b or a;
    layer5_outputs(5643) <= a;
    layer5_outputs(5644) <= '0';
    layer5_outputs(5645) <= not a;
    layer5_outputs(5646) <= b;
    layer5_outputs(5647) <= a and not b;
    layer5_outputs(5648) <= not a;
    layer5_outputs(5649) <= not (a and b);
    layer5_outputs(5650) <= not a;
    layer5_outputs(5651) <= not b;
    layer5_outputs(5652) <= '1';
    layer5_outputs(5653) <= not a;
    layer5_outputs(5654) <= b;
    layer5_outputs(5655) <= not a or b;
    layer5_outputs(5656) <= a xor b;
    layer5_outputs(5657) <= b;
    layer5_outputs(5658) <= a xor b;
    layer5_outputs(5659) <= not (a and b);
    layer5_outputs(5660) <= not b or a;
    layer5_outputs(5661) <= b and not a;
    layer5_outputs(5662) <= b;
    layer5_outputs(5663) <= not (a xor b);
    layer5_outputs(5664) <= not b;
    layer5_outputs(5665) <= not a;
    layer5_outputs(5666) <= a;
    layer5_outputs(5667) <= not (a xor b);
    layer5_outputs(5668) <= not a;
    layer5_outputs(5669) <= b;
    layer5_outputs(5670) <= b;
    layer5_outputs(5671) <= not b or a;
    layer5_outputs(5672) <= b and not a;
    layer5_outputs(5673) <= not a;
    layer5_outputs(5674) <= a or b;
    layer5_outputs(5675) <= a;
    layer5_outputs(5676) <= not a;
    layer5_outputs(5677) <= not (a and b);
    layer5_outputs(5678) <= not b or a;
    layer5_outputs(5679) <= a or b;
    layer5_outputs(5680) <= a and not b;
    layer5_outputs(5681) <= a xor b;
    layer5_outputs(5682) <= not b;
    layer5_outputs(5683) <= not a or b;
    layer5_outputs(5684) <= not (a or b);
    layer5_outputs(5685) <= a;
    layer5_outputs(5686) <= not a or b;
    layer5_outputs(5687) <= not a;
    layer5_outputs(5688) <= a xor b;
    layer5_outputs(5689) <= not a;
    layer5_outputs(5690) <= not (a or b);
    layer5_outputs(5691) <= a;
    layer5_outputs(5692) <= a and not b;
    layer5_outputs(5693) <= a and b;
    layer5_outputs(5694) <= a and not b;
    layer5_outputs(5695) <= b and not a;
    layer5_outputs(5696) <= not b;
    layer5_outputs(5697) <= not b;
    layer5_outputs(5698) <= not a;
    layer5_outputs(5699) <= a;
    layer5_outputs(5700) <= a and not b;
    layer5_outputs(5701) <= not a;
    layer5_outputs(5702) <= not a or b;
    layer5_outputs(5703) <= not b;
    layer5_outputs(5704) <= not a or b;
    layer5_outputs(5705) <= not (a xor b);
    layer5_outputs(5706) <= not (a and b);
    layer5_outputs(5707) <= not (a and b);
    layer5_outputs(5708) <= not b;
    layer5_outputs(5709) <= a or b;
    layer5_outputs(5710) <= not (a and b);
    layer5_outputs(5711) <= b and not a;
    layer5_outputs(5712) <= a and not b;
    layer5_outputs(5713) <= a or b;
    layer5_outputs(5714) <= a and not b;
    layer5_outputs(5715) <= not a;
    layer5_outputs(5716) <= a and not b;
    layer5_outputs(5717) <= not a or b;
    layer5_outputs(5718) <= not b;
    layer5_outputs(5719) <= not b;
    layer5_outputs(5720) <= a;
    layer5_outputs(5721) <= not b or a;
    layer5_outputs(5722) <= not a;
    layer5_outputs(5723) <= not b;
    layer5_outputs(5724) <= not a;
    layer5_outputs(5725) <= a;
    layer5_outputs(5726) <= a;
    layer5_outputs(5727) <= not b or a;
    layer5_outputs(5728) <= not (a xor b);
    layer5_outputs(5729) <= a;
    layer5_outputs(5730) <= b and not a;
    layer5_outputs(5731) <= a and not b;
    layer5_outputs(5732) <= not a;
    layer5_outputs(5733) <= not (a and b);
    layer5_outputs(5734) <= a or b;
    layer5_outputs(5735) <= a or b;
    layer5_outputs(5736) <= a;
    layer5_outputs(5737) <= not b or a;
    layer5_outputs(5738) <= not b;
    layer5_outputs(5739) <= not b or a;
    layer5_outputs(5740) <= not b;
    layer5_outputs(5741) <= not a;
    layer5_outputs(5742) <= a;
    layer5_outputs(5743) <= not (a xor b);
    layer5_outputs(5744) <= not (a xor b);
    layer5_outputs(5745) <= not (a or b);
    layer5_outputs(5746) <= not b or a;
    layer5_outputs(5747) <= not b;
    layer5_outputs(5748) <= a;
    layer5_outputs(5749) <= b;
    layer5_outputs(5750) <= a xor b;
    layer5_outputs(5751) <= a;
    layer5_outputs(5752) <= a and b;
    layer5_outputs(5753) <= not a;
    layer5_outputs(5754) <= a or b;
    layer5_outputs(5755) <= not b;
    layer5_outputs(5756) <= not (a xor b);
    layer5_outputs(5757) <= not (a and b);
    layer5_outputs(5758) <= not a;
    layer5_outputs(5759) <= a;
    layer5_outputs(5760) <= not (a and b);
    layer5_outputs(5761) <= not (a or b);
    layer5_outputs(5762) <= not (a xor b);
    layer5_outputs(5763) <= not b;
    layer5_outputs(5764) <= a or b;
    layer5_outputs(5765) <= not a;
    layer5_outputs(5766) <= not a;
    layer5_outputs(5767) <= not (a or b);
    layer5_outputs(5768) <= a and not b;
    layer5_outputs(5769) <= b;
    layer5_outputs(5770) <= a and b;
    layer5_outputs(5771) <= a and not b;
    layer5_outputs(5772) <= not a;
    layer5_outputs(5773) <= not a;
    layer5_outputs(5774) <= b;
    layer5_outputs(5775) <= not a or b;
    layer5_outputs(5776) <= not (a xor b);
    layer5_outputs(5777) <= not b;
    layer5_outputs(5778) <= not (a and b);
    layer5_outputs(5779) <= b and not a;
    layer5_outputs(5780) <= not b;
    layer5_outputs(5781) <= a or b;
    layer5_outputs(5782) <= a and not b;
    layer5_outputs(5783) <= a;
    layer5_outputs(5784) <= a xor b;
    layer5_outputs(5785) <= '1';
    layer5_outputs(5786) <= not a;
    layer5_outputs(5787) <= a;
    layer5_outputs(5788) <= not a;
    layer5_outputs(5789) <= not (a or b);
    layer5_outputs(5790) <= not (a xor b);
    layer5_outputs(5791) <= a;
    layer5_outputs(5792) <= not a or b;
    layer5_outputs(5793) <= not (a and b);
    layer5_outputs(5794) <= a xor b;
    layer5_outputs(5795) <= b;
    layer5_outputs(5796) <= '1';
    layer5_outputs(5797) <= b and not a;
    layer5_outputs(5798) <= a;
    layer5_outputs(5799) <= a;
    layer5_outputs(5800) <= a xor b;
    layer5_outputs(5801) <= not (a or b);
    layer5_outputs(5802) <= not a or b;
    layer5_outputs(5803) <= not b or a;
    layer5_outputs(5804) <= not (a or b);
    layer5_outputs(5805) <= b;
    layer5_outputs(5806) <= a;
    layer5_outputs(5807) <= not (a and b);
    layer5_outputs(5808) <= not b;
    layer5_outputs(5809) <= b;
    layer5_outputs(5810) <= not b;
    layer5_outputs(5811) <= a;
    layer5_outputs(5812) <= a and not b;
    layer5_outputs(5813) <= b;
    layer5_outputs(5814) <= b;
    layer5_outputs(5815) <= not (a and b);
    layer5_outputs(5816) <= a;
    layer5_outputs(5817) <= a;
    layer5_outputs(5818) <= not b or a;
    layer5_outputs(5819) <= not (a or b);
    layer5_outputs(5820) <= not b or a;
    layer5_outputs(5821) <= not b;
    layer5_outputs(5822) <= not b or a;
    layer5_outputs(5823) <= a or b;
    layer5_outputs(5824) <= b and not a;
    layer5_outputs(5825) <= not a;
    layer5_outputs(5826) <= not (a and b);
    layer5_outputs(5827) <= not b or a;
    layer5_outputs(5828) <= a xor b;
    layer5_outputs(5829) <= b and not a;
    layer5_outputs(5830) <= not b;
    layer5_outputs(5831) <= not (a or b);
    layer5_outputs(5832) <= not (a xor b);
    layer5_outputs(5833) <= b;
    layer5_outputs(5834) <= '0';
    layer5_outputs(5835) <= not a;
    layer5_outputs(5836) <= a and b;
    layer5_outputs(5837) <= a;
    layer5_outputs(5838) <= not (a and b);
    layer5_outputs(5839) <= not (a xor b);
    layer5_outputs(5840) <= not b;
    layer5_outputs(5841) <= b and not a;
    layer5_outputs(5842) <= not a;
    layer5_outputs(5843) <= b and not a;
    layer5_outputs(5844) <= a and not b;
    layer5_outputs(5845) <= b;
    layer5_outputs(5846) <= not a or b;
    layer5_outputs(5847) <= b;
    layer5_outputs(5848) <= b;
    layer5_outputs(5849) <= not a or b;
    layer5_outputs(5850) <= a xor b;
    layer5_outputs(5851) <= a xor b;
    layer5_outputs(5852) <= not (a and b);
    layer5_outputs(5853) <= a;
    layer5_outputs(5854) <= b;
    layer5_outputs(5855) <= not (a xor b);
    layer5_outputs(5856) <= not (a xor b);
    layer5_outputs(5857) <= not a;
    layer5_outputs(5858) <= not b;
    layer5_outputs(5859) <= b;
    layer5_outputs(5860) <= a and b;
    layer5_outputs(5861) <= not a or b;
    layer5_outputs(5862) <= b and not a;
    layer5_outputs(5863) <= not b;
    layer5_outputs(5864) <= not a or b;
    layer5_outputs(5865) <= not a;
    layer5_outputs(5866) <= a xor b;
    layer5_outputs(5867) <= not (a and b);
    layer5_outputs(5868) <= not b or a;
    layer5_outputs(5869) <= not b or a;
    layer5_outputs(5870) <= a and not b;
    layer5_outputs(5871) <= a xor b;
    layer5_outputs(5872) <= not (a xor b);
    layer5_outputs(5873) <= a;
    layer5_outputs(5874) <= not a;
    layer5_outputs(5875) <= not (a xor b);
    layer5_outputs(5876) <= not b;
    layer5_outputs(5877) <= a and b;
    layer5_outputs(5878) <= not a;
    layer5_outputs(5879) <= not (a or b);
    layer5_outputs(5880) <= not a;
    layer5_outputs(5881) <= a and b;
    layer5_outputs(5882) <= b and not a;
    layer5_outputs(5883) <= a;
    layer5_outputs(5884) <= not a or b;
    layer5_outputs(5885) <= a;
    layer5_outputs(5886) <= not a;
    layer5_outputs(5887) <= not (a xor b);
    layer5_outputs(5888) <= not a;
    layer5_outputs(5889) <= b and not a;
    layer5_outputs(5890) <= not b;
    layer5_outputs(5891) <= not a;
    layer5_outputs(5892) <= not (a or b);
    layer5_outputs(5893) <= not b or a;
    layer5_outputs(5894) <= not a;
    layer5_outputs(5895) <= not b or a;
    layer5_outputs(5896) <= b and not a;
    layer5_outputs(5897) <= not (a xor b);
    layer5_outputs(5898) <= a xor b;
    layer5_outputs(5899) <= b;
    layer5_outputs(5900) <= b;
    layer5_outputs(5901) <= not a;
    layer5_outputs(5902) <= a or b;
    layer5_outputs(5903) <= '1';
    layer5_outputs(5904) <= a xor b;
    layer5_outputs(5905) <= not a;
    layer5_outputs(5906) <= not a;
    layer5_outputs(5907) <= not (a and b);
    layer5_outputs(5908) <= not a or b;
    layer5_outputs(5909) <= b;
    layer5_outputs(5910) <= not b;
    layer5_outputs(5911) <= a and not b;
    layer5_outputs(5912) <= not (a xor b);
    layer5_outputs(5913) <= not a;
    layer5_outputs(5914) <= not (a xor b);
    layer5_outputs(5915) <= not (a xor b);
    layer5_outputs(5916) <= not (a and b);
    layer5_outputs(5917) <= b and not a;
    layer5_outputs(5918) <= not (a xor b);
    layer5_outputs(5919) <= not a;
    layer5_outputs(5920) <= not (a and b);
    layer5_outputs(5921) <= a and not b;
    layer5_outputs(5922) <= not a or b;
    layer5_outputs(5923) <= not a or b;
    layer5_outputs(5924) <= not (a xor b);
    layer5_outputs(5925) <= not (a and b);
    layer5_outputs(5926) <= '0';
    layer5_outputs(5927) <= a and not b;
    layer5_outputs(5928) <= not b;
    layer5_outputs(5929) <= not a;
    layer5_outputs(5930) <= not a or b;
    layer5_outputs(5931) <= b;
    layer5_outputs(5932) <= '0';
    layer5_outputs(5933) <= a xor b;
    layer5_outputs(5934) <= not b;
    layer5_outputs(5935) <= b;
    layer5_outputs(5936) <= a xor b;
    layer5_outputs(5937) <= not b;
    layer5_outputs(5938) <= a;
    layer5_outputs(5939) <= b;
    layer5_outputs(5940) <= a and b;
    layer5_outputs(5941) <= not a;
    layer5_outputs(5942) <= not a;
    layer5_outputs(5943) <= a and b;
    layer5_outputs(5944) <= not a;
    layer5_outputs(5945) <= not b or a;
    layer5_outputs(5946) <= b;
    layer5_outputs(5947) <= not (a or b);
    layer5_outputs(5948) <= not a or b;
    layer5_outputs(5949) <= not (a and b);
    layer5_outputs(5950) <= not b;
    layer5_outputs(5951) <= b and not a;
    layer5_outputs(5952) <= a and b;
    layer5_outputs(5953) <= not b;
    layer5_outputs(5954) <= b and not a;
    layer5_outputs(5955) <= b and not a;
    layer5_outputs(5956) <= b;
    layer5_outputs(5957) <= a xor b;
    layer5_outputs(5958) <= not a or b;
    layer5_outputs(5959) <= b and not a;
    layer5_outputs(5960) <= not b;
    layer5_outputs(5961) <= b;
    layer5_outputs(5962) <= not a;
    layer5_outputs(5963) <= not b;
    layer5_outputs(5964) <= not (a and b);
    layer5_outputs(5965) <= b and not a;
    layer5_outputs(5966) <= b;
    layer5_outputs(5967) <= not a;
    layer5_outputs(5968) <= b;
    layer5_outputs(5969) <= b;
    layer5_outputs(5970) <= not b;
    layer5_outputs(5971) <= not (a or b);
    layer5_outputs(5972) <= not a;
    layer5_outputs(5973) <= not (a xor b);
    layer5_outputs(5974) <= not (a and b);
    layer5_outputs(5975) <= a;
    layer5_outputs(5976) <= b;
    layer5_outputs(5977) <= b;
    layer5_outputs(5978) <= not a;
    layer5_outputs(5979) <= a or b;
    layer5_outputs(5980) <= not a;
    layer5_outputs(5981) <= not a;
    layer5_outputs(5982) <= not b;
    layer5_outputs(5983) <= a;
    layer5_outputs(5984) <= a and not b;
    layer5_outputs(5985) <= not b;
    layer5_outputs(5986) <= a or b;
    layer5_outputs(5987) <= a and b;
    layer5_outputs(5988) <= not (a and b);
    layer5_outputs(5989) <= a;
    layer5_outputs(5990) <= not (a and b);
    layer5_outputs(5991) <= a;
    layer5_outputs(5992) <= not (a xor b);
    layer5_outputs(5993) <= a and not b;
    layer5_outputs(5994) <= a or b;
    layer5_outputs(5995) <= a and not b;
    layer5_outputs(5996) <= not b;
    layer5_outputs(5997) <= not (a xor b);
    layer5_outputs(5998) <= b;
    layer5_outputs(5999) <= a and not b;
    layer5_outputs(6000) <= b;
    layer5_outputs(6001) <= b;
    layer5_outputs(6002) <= a xor b;
    layer5_outputs(6003) <= not b;
    layer5_outputs(6004) <= a xor b;
    layer5_outputs(6005) <= a and b;
    layer5_outputs(6006) <= a xor b;
    layer5_outputs(6007) <= not (a xor b);
    layer5_outputs(6008) <= b;
    layer5_outputs(6009) <= b and not a;
    layer5_outputs(6010) <= a;
    layer5_outputs(6011) <= not (a or b);
    layer5_outputs(6012) <= b;
    layer5_outputs(6013) <= not (a xor b);
    layer5_outputs(6014) <= not a;
    layer5_outputs(6015) <= b;
    layer5_outputs(6016) <= not a or b;
    layer5_outputs(6017) <= not b or a;
    layer5_outputs(6018) <= not a;
    layer5_outputs(6019) <= not (a xor b);
    layer5_outputs(6020) <= a or b;
    layer5_outputs(6021) <= not (a xor b);
    layer5_outputs(6022) <= not a;
    layer5_outputs(6023) <= not b or a;
    layer5_outputs(6024) <= a;
    layer5_outputs(6025) <= a xor b;
    layer5_outputs(6026) <= a xor b;
    layer5_outputs(6027) <= a xor b;
    layer5_outputs(6028) <= not a;
    layer5_outputs(6029) <= not b;
    layer5_outputs(6030) <= a;
    layer5_outputs(6031) <= b;
    layer5_outputs(6032) <= a and not b;
    layer5_outputs(6033) <= b;
    layer5_outputs(6034) <= not (a and b);
    layer5_outputs(6035) <= a or b;
    layer5_outputs(6036) <= a xor b;
    layer5_outputs(6037) <= not (a xor b);
    layer5_outputs(6038) <= not a;
    layer5_outputs(6039) <= a xor b;
    layer5_outputs(6040) <= not b or a;
    layer5_outputs(6041) <= not b;
    layer5_outputs(6042) <= not b;
    layer5_outputs(6043) <= a or b;
    layer5_outputs(6044) <= a;
    layer5_outputs(6045) <= a;
    layer5_outputs(6046) <= b and not a;
    layer5_outputs(6047) <= a;
    layer5_outputs(6048) <= a;
    layer5_outputs(6049) <= b and not a;
    layer5_outputs(6050) <= b;
    layer5_outputs(6051) <= not a;
    layer5_outputs(6052) <= not (a and b);
    layer5_outputs(6053) <= b and not a;
    layer5_outputs(6054) <= not (a or b);
    layer5_outputs(6055) <= not b or a;
    layer5_outputs(6056) <= a and not b;
    layer5_outputs(6057) <= b and not a;
    layer5_outputs(6058) <= not a;
    layer5_outputs(6059) <= not a or b;
    layer5_outputs(6060) <= not a or b;
    layer5_outputs(6061) <= not a;
    layer5_outputs(6062) <= not b;
    layer5_outputs(6063) <= a and not b;
    layer5_outputs(6064) <= not (a or b);
    layer5_outputs(6065) <= not a or b;
    layer5_outputs(6066) <= a xor b;
    layer5_outputs(6067) <= not a;
    layer5_outputs(6068) <= not a or b;
    layer5_outputs(6069) <= a;
    layer5_outputs(6070) <= a and not b;
    layer5_outputs(6071) <= a;
    layer5_outputs(6072) <= not b;
    layer5_outputs(6073) <= a;
    layer5_outputs(6074) <= not (a or b);
    layer5_outputs(6075) <= not (a or b);
    layer5_outputs(6076) <= not a or b;
    layer5_outputs(6077) <= b;
    layer5_outputs(6078) <= b and not a;
    layer5_outputs(6079) <= not a;
    layer5_outputs(6080) <= not a or b;
    layer5_outputs(6081) <= not (a and b);
    layer5_outputs(6082) <= not (a xor b);
    layer5_outputs(6083) <= b and not a;
    layer5_outputs(6084) <= not a;
    layer5_outputs(6085) <= not (a xor b);
    layer5_outputs(6086) <= b;
    layer5_outputs(6087) <= a and not b;
    layer5_outputs(6088) <= not a;
    layer5_outputs(6089) <= a;
    layer5_outputs(6090) <= not b;
    layer5_outputs(6091) <= not (a xor b);
    layer5_outputs(6092) <= a and not b;
    layer5_outputs(6093) <= not a;
    layer5_outputs(6094) <= not (a and b);
    layer5_outputs(6095) <= '0';
    layer5_outputs(6096) <= not a;
    layer5_outputs(6097) <= b;
    layer5_outputs(6098) <= not (a xor b);
    layer5_outputs(6099) <= a and b;
    layer5_outputs(6100) <= not (a or b);
    layer5_outputs(6101) <= not (a xor b);
    layer5_outputs(6102) <= b;
    layer5_outputs(6103) <= a;
    layer5_outputs(6104) <= '0';
    layer5_outputs(6105) <= not a or b;
    layer5_outputs(6106) <= not (a or b);
    layer5_outputs(6107) <= a or b;
    layer5_outputs(6108) <= not a;
    layer5_outputs(6109) <= not a;
    layer5_outputs(6110) <= b and not a;
    layer5_outputs(6111) <= not a;
    layer5_outputs(6112) <= '0';
    layer5_outputs(6113) <= not (a and b);
    layer5_outputs(6114) <= not a;
    layer5_outputs(6115) <= not (a or b);
    layer5_outputs(6116) <= a xor b;
    layer5_outputs(6117) <= a;
    layer5_outputs(6118) <= b;
    layer5_outputs(6119) <= not (a xor b);
    layer5_outputs(6120) <= b and not a;
    layer5_outputs(6121) <= not (a xor b);
    layer5_outputs(6122) <= not a;
    layer5_outputs(6123) <= b and not a;
    layer5_outputs(6124) <= b and not a;
    layer5_outputs(6125) <= a and b;
    layer5_outputs(6126) <= not (a xor b);
    layer5_outputs(6127) <= not (a and b);
    layer5_outputs(6128) <= a;
    layer5_outputs(6129) <= a;
    layer5_outputs(6130) <= a and b;
    layer5_outputs(6131) <= not b;
    layer5_outputs(6132) <= not b or a;
    layer5_outputs(6133) <= not (a and b);
    layer5_outputs(6134) <= b;
    layer5_outputs(6135) <= not b;
    layer5_outputs(6136) <= a and not b;
    layer5_outputs(6137) <= b;
    layer5_outputs(6138) <= not b;
    layer5_outputs(6139) <= not (a xor b);
    layer5_outputs(6140) <= not a or b;
    layer5_outputs(6141) <= not (a and b);
    layer5_outputs(6142) <= not b;
    layer5_outputs(6143) <= not (a xor b);
    layer5_outputs(6144) <= not b;
    layer5_outputs(6145) <= b;
    layer5_outputs(6146) <= b;
    layer5_outputs(6147) <= not (a or b);
    layer5_outputs(6148) <= b and not a;
    layer5_outputs(6149) <= a;
    layer5_outputs(6150) <= not a;
    layer5_outputs(6151) <= a and b;
    layer5_outputs(6152) <= a and b;
    layer5_outputs(6153) <= not b;
    layer5_outputs(6154) <= not (a and b);
    layer5_outputs(6155) <= not a;
    layer5_outputs(6156) <= '1';
    layer5_outputs(6157) <= not b or a;
    layer5_outputs(6158) <= not (a xor b);
    layer5_outputs(6159) <= b;
    layer5_outputs(6160) <= a and b;
    layer5_outputs(6161) <= not a;
    layer5_outputs(6162) <= not a;
    layer5_outputs(6163) <= not b or a;
    layer5_outputs(6164) <= not b;
    layer5_outputs(6165) <= a;
    layer5_outputs(6166) <= not a;
    layer5_outputs(6167) <= a;
    layer5_outputs(6168) <= not b or a;
    layer5_outputs(6169) <= not b;
    layer5_outputs(6170) <= a xor b;
    layer5_outputs(6171) <= not b;
    layer5_outputs(6172) <= a and not b;
    layer5_outputs(6173) <= not a;
    layer5_outputs(6174) <= a;
    layer5_outputs(6175) <= not (a and b);
    layer5_outputs(6176) <= not a;
    layer5_outputs(6177) <= not a;
    layer5_outputs(6178) <= a;
    layer5_outputs(6179) <= b and not a;
    layer5_outputs(6180) <= not (a or b);
    layer5_outputs(6181) <= not a;
    layer5_outputs(6182) <= a xor b;
    layer5_outputs(6183) <= a and not b;
    layer5_outputs(6184) <= not a;
    layer5_outputs(6185) <= '0';
    layer5_outputs(6186) <= a and b;
    layer5_outputs(6187) <= a;
    layer5_outputs(6188) <= not (a xor b);
    layer5_outputs(6189) <= a or b;
    layer5_outputs(6190) <= not (a xor b);
    layer5_outputs(6191) <= a;
    layer5_outputs(6192) <= a;
    layer5_outputs(6193) <= not b;
    layer5_outputs(6194) <= not (a xor b);
    layer5_outputs(6195) <= b;
    layer5_outputs(6196) <= a;
    layer5_outputs(6197) <= not (a and b);
    layer5_outputs(6198) <= not b;
    layer5_outputs(6199) <= '1';
    layer5_outputs(6200) <= b;
    layer5_outputs(6201) <= b;
    layer5_outputs(6202) <= a;
    layer5_outputs(6203) <= b and not a;
    layer5_outputs(6204) <= not a;
    layer5_outputs(6205) <= not (a and b);
    layer5_outputs(6206) <= not (a or b);
    layer5_outputs(6207) <= a;
    layer5_outputs(6208) <= not (a xor b);
    layer5_outputs(6209) <= b;
    layer5_outputs(6210) <= a and not b;
    layer5_outputs(6211) <= not a;
    layer5_outputs(6212) <= not a;
    layer5_outputs(6213) <= not (a or b);
    layer5_outputs(6214) <= a and not b;
    layer5_outputs(6215) <= not a or b;
    layer5_outputs(6216) <= '0';
    layer5_outputs(6217) <= not (a or b);
    layer5_outputs(6218) <= not (a and b);
    layer5_outputs(6219) <= a xor b;
    layer5_outputs(6220) <= b;
    layer5_outputs(6221) <= not b;
    layer5_outputs(6222) <= a xor b;
    layer5_outputs(6223) <= a;
    layer5_outputs(6224) <= not (a or b);
    layer5_outputs(6225) <= not b;
    layer5_outputs(6226) <= b;
    layer5_outputs(6227) <= a;
    layer5_outputs(6228) <= a;
    layer5_outputs(6229) <= b;
    layer5_outputs(6230) <= a;
    layer5_outputs(6231) <= not (a xor b);
    layer5_outputs(6232) <= not (a xor b);
    layer5_outputs(6233) <= b;
    layer5_outputs(6234) <= a;
    layer5_outputs(6235) <= not (a or b);
    layer5_outputs(6236) <= a or b;
    layer5_outputs(6237) <= not a;
    layer5_outputs(6238) <= a xor b;
    layer5_outputs(6239) <= not (a xor b);
    layer5_outputs(6240) <= not a;
    layer5_outputs(6241) <= not (a xor b);
    layer5_outputs(6242) <= a and b;
    layer5_outputs(6243) <= a and b;
    layer5_outputs(6244) <= a;
    layer5_outputs(6245) <= not (a and b);
    layer5_outputs(6246) <= not a;
    layer5_outputs(6247) <= not a;
    layer5_outputs(6248) <= a and not b;
    layer5_outputs(6249) <= not (a xor b);
    layer5_outputs(6250) <= b;
    layer5_outputs(6251) <= not b or a;
    layer5_outputs(6252) <= a and not b;
    layer5_outputs(6253) <= not a;
    layer5_outputs(6254) <= not b;
    layer5_outputs(6255) <= a and b;
    layer5_outputs(6256) <= not a;
    layer5_outputs(6257) <= a and not b;
    layer5_outputs(6258) <= b;
    layer5_outputs(6259) <= a or b;
    layer5_outputs(6260) <= not b or a;
    layer5_outputs(6261) <= not (a xor b);
    layer5_outputs(6262) <= not (a or b);
    layer5_outputs(6263) <= not (a and b);
    layer5_outputs(6264) <= not a or b;
    layer5_outputs(6265) <= b and not a;
    layer5_outputs(6266) <= a;
    layer5_outputs(6267) <= b;
    layer5_outputs(6268) <= a;
    layer5_outputs(6269) <= a;
    layer5_outputs(6270) <= not (a and b);
    layer5_outputs(6271) <= '1';
    layer5_outputs(6272) <= not (a xor b);
    layer5_outputs(6273) <= not a;
    layer5_outputs(6274) <= a;
    layer5_outputs(6275) <= not a;
    layer5_outputs(6276) <= a;
    layer5_outputs(6277) <= not (a or b);
    layer5_outputs(6278) <= a;
    layer5_outputs(6279) <= not a;
    layer5_outputs(6280) <= a or b;
    layer5_outputs(6281) <= a and b;
    layer5_outputs(6282) <= not b;
    layer5_outputs(6283) <= b;
    layer5_outputs(6284) <= a;
    layer5_outputs(6285) <= not b;
    layer5_outputs(6286) <= a and b;
    layer5_outputs(6287) <= not (a xor b);
    layer5_outputs(6288) <= a xor b;
    layer5_outputs(6289) <= not (a xor b);
    layer5_outputs(6290) <= not a;
    layer5_outputs(6291) <= not a;
    layer5_outputs(6292) <= not (a and b);
    layer5_outputs(6293) <= not b;
    layer5_outputs(6294) <= a and not b;
    layer5_outputs(6295) <= a;
    layer5_outputs(6296) <= '0';
    layer5_outputs(6297) <= not b or a;
    layer5_outputs(6298) <= not a;
    layer5_outputs(6299) <= not b or a;
    layer5_outputs(6300) <= a or b;
    layer5_outputs(6301) <= b;
    layer5_outputs(6302) <= not (a and b);
    layer5_outputs(6303) <= '1';
    layer5_outputs(6304) <= not a;
    layer5_outputs(6305) <= a and b;
    layer5_outputs(6306) <= not b;
    layer5_outputs(6307) <= b;
    layer5_outputs(6308) <= a;
    layer5_outputs(6309) <= b;
    layer5_outputs(6310) <= not (a or b);
    layer5_outputs(6311) <= b and not a;
    layer5_outputs(6312) <= a xor b;
    layer5_outputs(6313) <= b;
    layer5_outputs(6314) <= not (a xor b);
    layer5_outputs(6315) <= a;
    layer5_outputs(6316) <= not (a xor b);
    layer5_outputs(6317) <= not b or a;
    layer5_outputs(6318) <= b;
    layer5_outputs(6319) <= b;
    layer5_outputs(6320) <= a and not b;
    layer5_outputs(6321) <= a;
    layer5_outputs(6322) <= a;
    layer5_outputs(6323) <= a or b;
    layer5_outputs(6324) <= not a;
    layer5_outputs(6325) <= not a;
    layer5_outputs(6326) <= not b;
    layer5_outputs(6327) <= a;
    layer5_outputs(6328) <= not b;
    layer5_outputs(6329) <= not (a and b);
    layer5_outputs(6330) <= a xor b;
    layer5_outputs(6331) <= not (a or b);
    layer5_outputs(6332) <= not b or a;
    layer5_outputs(6333) <= a and not b;
    layer5_outputs(6334) <= a xor b;
    layer5_outputs(6335) <= b and not a;
    layer5_outputs(6336) <= a;
    layer5_outputs(6337) <= a;
    layer5_outputs(6338) <= not (a or b);
    layer5_outputs(6339) <= not b;
    layer5_outputs(6340) <= b and not a;
    layer5_outputs(6341) <= not b or a;
    layer5_outputs(6342) <= a;
    layer5_outputs(6343) <= b;
    layer5_outputs(6344) <= not a or b;
    layer5_outputs(6345) <= a;
    layer5_outputs(6346) <= not b or a;
    layer5_outputs(6347) <= a or b;
    layer5_outputs(6348) <= not b;
    layer5_outputs(6349) <= not b;
    layer5_outputs(6350) <= not b;
    layer5_outputs(6351) <= b and not a;
    layer5_outputs(6352) <= not a;
    layer5_outputs(6353) <= a xor b;
    layer5_outputs(6354) <= b;
    layer5_outputs(6355) <= '1';
    layer5_outputs(6356) <= a;
    layer5_outputs(6357) <= a and b;
    layer5_outputs(6358) <= not b;
    layer5_outputs(6359) <= not a;
    layer5_outputs(6360) <= not b;
    layer5_outputs(6361) <= not a;
    layer5_outputs(6362) <= not a or b;
    layer5_outputs(6363) <= not (a and b);
    layer5_outputs(6364) <= not b;
    layer5_outputs(6365) <= not (a or b);
    layer5_outputs(6366) <= not b;
    layer5_outputs(6367) <= b and not a;
    layer5_outputs(6368) <= not a or b;
    layer5_outputs(6369) <= a or b;
    layer5_outputs(6370) <= a or b;
    layer5_outputs(6371) <= a or b;
    layer5_outputs(6372) <= a and b;
    layer5_outputs(6373) <= a or b;
    layer5_outputs(6374) <= b;
    layer5_outputs(6375) <= b;
    layer5_outputs(6376) <= not a;
    layer5_outputs(6377) <= not (a or b);
    layer5_outputs(6378) <= a and b;
    layer5_outputs(6379) <= not b;
    layer5_outputs(6380) <= a;
    layer5_outputs(6381) <= b and not a;
    layer5_outputs(6382) <= not b or a;
    layer5_outputs(6383) <= b;
    layer5_outputs(6384) <= not b or a;
    layer5_outputs(6385) <= a;
    layer5_outputs(6386) <= a;
    layer5_outputs(6387) <= not b;
    layer5_outputs(6388) <= a and not b;
    layer5_outputs(6389) <= not (a xor b);
    layer5_outputs(6390) <= a or b;
    layer5_outputs(6391) <= b;
    layer5_outputs(6392) <= not b;
    layer5_outputs(6393) <= not a or b;
    layer5_outputs(6394) <= not (a and b);
    layer5_outputs(6395) <= not a or b;
    layer5_outputs(6396) <= a or b;
    layer5_outputs(6397) <= not a;
    layer5_outputs(6398) <= a;
    layer5_outputs(6399) <= not a;
    layer5_outputs(6400) <= a and b;
    layer5_outputs(6401) <= a;
    layer5_outputs(6402) <= not (a xor b);
    layer5_outputs(6403) <= not a;
    layer5_outputs(6404) <= a;
    layer5_outputs(6405) <= '1';
    layer5_outputs(6406) <= a and not b;
    layer5_outputs(6407) <= not b or a;
    layer5_outputs(6408) <= a;
    layer5_outputs(6409) <= a or b;
    layer5_outputs(6410) <= not b or a;
    layer5_outputs(6411) <= not (a xor b);
    layer5_outputs(6412) <= b;
    layer5_outputs(6413) <= b and not a;
    layer5_outputs(6414) <= not (a or b);
    layer5_outputs(6415) <= a and not b;
    layer5_outputs(6416) <= b;
    layer5_outputs(6417) <= not (a xor b);
    layer5_outputs(6418) <= b;
    layer5_outputs(6419) <= not (a xor b);
    layer5_outputs(6420) <= not b;
    layer5_outputs(6421) <= not (a or b);
    layer5_outputs(6422) <= a or b;
    layer5_outputs(6423) <= b;
    layer5_outputs(6424) <= not b or a;
    layer5_outputs(6425) <= b;
    layer5_outputs(6426) <= not a;
    layer5_outputs(6427) <= a;
    layer5_outputs(6428) <= not (a and b);
    layer5_outputs(6429) <= not b;
    layer5_outputs(6430) <= a and b;
    layer5_outputs(6431) <= not b;
    layer5_outputs(6432) <= not a;
    layer5_outputs(6433) <= not a;
    layer5_outputs(6434) <= not b;
    layer5_outputs(6435) <= a;
    layer5_outputs(6436) <= not (a and b);
    layer5_outputs(6437) <= not (a and b);
    layer5_outputs(6438) <= not a;
    layer5_outputs(6439) <= a xor b;
    layer5_outputs(6440) <= not (a xor b);
    layer5_outputs(6441) <= not (a xor b);
    layer5_outputs(6442) <= a;
    layer5_outputs(6443) <= not b;
    layer5_outputs(6444) <= a;
    layer5_outputs(6445) <= not b;
    layer5_outputs(6446) <= a or b;
    layer5_outputs(6447) <= b;
    layer5_outputs(6448) <= not b or a;
    layer5_outputs(6449) <= b and not a;
    layer5_outputs(6450) <= not b;
    layer5_outputs(6451) <= a;
    layer5_outputs(6452) <= not (a and b);
    layer5_outputs(6453) <= a xor b;
    layer5_outputs(6454) <= b and not a;
    layer5_outputs(6455) <= a;
    layer5_outputs(6456) <= a or b;
    layer5_outputs(6457) <= a xor b;
    layer5_outputs(6458) <= '0';
    layer5_outputs(6459) <= a and b;
    layer5_outputs(6460) <= a;
    layer5_outputs(6461) <= not a;
    layer5_outputs(6462) <= not (a and b);
    layer5_outputs(6463) <= b;
    layer5_outputs(6464) <= a;
    layer5_outputs(6465) <= not (a or b);
    layer5_outputs(6466) <= not (a and b);
    layer5_outputs(6467) <= a and not b;
    layer5_outputs(6468) <= a and not b;
    layer5_outputs(6469) <= not a;
    layer5_outputs(6470) <= a xor b;
    layer5_outputs(6471) <= not (a xor b);
    layer5_outputs(6472) <= a or b;
    layer5_outputs(6473) <= b and not a;
    layer5_outputs(6474) <= not a;
    layer5_outputs(6475) <= a xor b;
    layer5_outputs(6476) <= b and not a;
    layer5_outputs(6477) <= b;
    layer5_outputs(6478) <= a and b;
    layer5_outputs(6479) <= not a;
    layer5_outputs(6480) <= b and not a;
    layer5_outputs(6481) <= a;
    layer5_outputs(6482) <= b and not a;
    layer5_outputs(6483) <= not (a xor b);
    layer5_outputs(6484) <= a xor b;
    layer5_outputs(6485) <= b;
    layer5_outputs(6486) <= not b or a;
    layer5_outputs(6487) <= not b;
    layer5_outputs(6488) <= '0';
    layer5_outputs(6489) <= a or b;
    layer5_outputs(6490) <= b;
    layer5_outputs(6491) <= a and not b;
    layer5_outputs(6492) <= not b or a;
    layer5_outputs(6493) <= not (a xor b);
    layer5_outputs(6494) <= b;
    layer5_outputs(6495) <= not (a xor b);
    layer5_outputs(6496) <= a and not b;
    layer5_outputs(6497) <= a and b;
    layer5_outputs(6498) <= not (a and b);
    layer5_outputs(6499) <= a;
    layer5_outputs(6500) <= b;
    layer5_outputs(6501) <= not (a or b);
    layer5_outputs(6502) <= a or b;
    layer5_outputs(6503) <= '1';
    layer5_outputs(6504) <= b;
    layer5_outputs(6505) <= not (a and b);
    layer5_outputs(6506) <= not (a xor b);
    layer5_outputs(6507) <= not b;
    layer5_outputs(6508) <= a;
    layer5_outputs(6509) <= b;
    layer5_outputs(6510) <= a and b;
    layer5_outputs(6511) <= not a;
    layer5_outputs(6512) <= a xor b;
    layer5_outputs(6513) <= a or b;
    layer5_outputs(6514) <= not (a and b);
    layer5_outputs(6515) <= not (a xor b);
    layer5_outputs(6516) <= a xor b;
    layer5_outputs(6517) <= b;
    layer5_outputs(6518) <= b;
    layer5_outputs(6519) <= not a or b;
    layer5_outputs(6520) <= b;
    layer5_outputs(6521) <= a or b;
    layer5_outputs(6522) <= a xor b;
    layer5_outputs(6523) <= b;
    layer5_outputs(6524) <= not (a and b);
    layer5_outputs(6525) <= a xor b;
    layer5_outputs(6526) <= not (a xor b);
    layer5_outputs(6527) <= not a;
    layer5_outputs(6528) <= not a;
    layer5_outputs(6529) <= a;
    layer5_outputs(6530) <= b;
    layer5_outputs(6531) <= not (a and b);
    layer5_outputs(6532) <= not (a or b);
    layer5_outputs(6533) <= not (a xor b);
    layer5_outputs(6534) <= a;
    layer5_outputs(6535) <= a and not b;
    layer5_outputs(6536) <= a;
    layer5_outputs(6537) <= not b or a;
    layer5_outputs(6538) <= a;
    layer5_outputs(6539) <= not (a xor b);
    layer5_outputs(6540) <= not a;
    layer5_outputs(6541) <= b and not a;
    layer5_outputs(6542) <= not (a xor b);
    layer5_outputs(6543) <= b;
    layer5_outputs(6544) <= not a;
    layer5_outputs(6545) <= a xor b;
    layer5_outputs(6546) <= not b;
    layer5_outputs(6547) <= not (a and b);
    layer5_outputs(6548) <= b;
    layer5_outputs(6549) <= not a or b;
    layer5_outputs(6550) <= '0';
    layer5_outputs(6551) <= b and not a;
    layer5_outputs(6552) <= a;
    layer5_outputs(6553) <= a;
    layer5_outputs(6554) <= not (a xor b);
    layer5_outputs(6555) <= b;
    layer5_outputs(6556) <= a or b;
    layer5_outputs(6557) <= b;
    layer5_outputs(6558) <= not a;
    layer5_outputs(6559) <= a or b;
    layer5_outputs(6560) <= not a;
    layer5_outputs(6561) <= a and not b;
    layer5_outputs(6562) <= '1';
    layer5_outputs(6563) <= a or b;
    layer5_outputs(6564) <= '1';
    layer5_outputs(6565) <= not a;
    layer5_outputs(6566) <= not b or a;
    layer5_outputs(6567) <= b;
    layer5_outputs(6568) <= b;
    layer5_outputs(6569) <= a;
    layer5_outputs(6570) <= a or b;
    layer5_outputs(6571) <= a;
    layer5_outputs(6572) <= not a;
    layer5_outputs(6573) <= a or b;
    layer5_outputs(6574) <= not a;
    layer5_outputs(6575) <= a or b;
    layer5_outputs(6576) <= b and not a;
    layer5_outputs(6577) <= a and not b;
    layer5_outputs(6578) <= b;
    layer5_outputs(6579) <= not b;
    layer5_outputs(6580) <= a;
    layer5_outputs(6581) <= not b or a;
    layer5_outputs(6582) <= a and b;
    layer5_outputs(6583) <= a;
    layer5_outputs(6584) <= not (a xor b);
    layer5_outputs(6585) <= not a or b;
    layer5_outputs(6586) <= not b;
    layer5_outputs(6587) <= a;
    layer5_outputs(6588) <= not (a or b);
    layer5_outputs(6589) <= not b or a;
    layer5_outputs(6590) <= a;
    layer5_outputs(6591) <= not a or b;
    layer5_outputs(6592) <= not b;
    layer5_outputs(6593) <= not b;
    layer5_outputs(6594) <= a xor b;
    layer5_outputs(6595) <= a and not b;
    layer5_outputs(6596) <= '1';
    layer5_outputs(6597) <= not b or a;
    layer5_outputs(6598) <= '1';
    layer5_outputs(6599) <= b;
    layer5_outputs(6600) <= b;
    layer5_outputs(6601) <= b;
    layer5_outputs(6602) <= a or b;
    layer5_outputs(6603) <= not b;
    layer5_outputs(6604) <= a;
    layer5_outputs(6605) <= not b;
    layer5_outputs(6606) <= b;
    layer5_outputs(6607) <= a and not b;
    layer5_outputs(6608) <= a;
    layer5_outputs(6609) <= a or b;
    layer5_outputs(6610) <= a or b;
    layer5_outputs(6611) <= not b or a;
    layer5_outputs(6612) <= not b;
    layer5_outputs(6613) <= a;
    layer5_outputs(6614) <= not (a or b);
    layer5_outputs(6615) <= not b;
    layer5_outputs(6616) <= a xor b;
    layer5_outputs(6617) <= a and b;
    layer5_outputs(6618) <= not a or b;
    layer5_outputs(6619) <= not a;
    layer5_outputs(6620) <= not a or b;
    layer5_outputs(6621) <= b;
    layer5_outputs(6622) <= a or b;
    layer5_outputs(6623) <= '1';
    layer5_outputs(6624) <= a;
    layer5_outputs(6625) <= not a;
    layer5_outputs(6626) <= b;
    layer5_outputs(6627) <= not (a xor b);
    layer5_outputs(6628) <= not b;
    layer5_outputs(6629) <= not b or a;
    layer5_outputs(6630) <= a xor b;
    layer5_outputs(6631) <= not (a xor b);
    layer5_outputs(6632) <= a and b;
    layer5_outputs(6633) <= a or b;
    layer5_outputs(6634) <= not (a xor b);
    layer5_outputs(6635) <= a and b;
    layer5_outputs(6636) <= b;
    layer5_outputs(6637) <= a;
    layer5_outputs(6638) <= not (a or b);
    layer5_outputs(6639) <= b;
    layer5_outputs(6640) <= a or b;
    layer5_outputs(6641) <= a or b;
    layer5_outputs(6642) <= a;
    layer5_outputs(6643) <= a and not b;
    layer5_outputs(6644) <= not a;
    layer5_outputs(6645) <= '1';
    layer5_outputs(6646) <= a and b;
    layer5_outputs(6647) <= a;
    layer5_outputs(6648) <= a and not b;
    layer5_outputs(6649) <= '1';
    layer5_outputs(6650) <= a;
    layer5_outputs(6651) <= not b or a;
    layer5_outputs(6652) <= a;
    layer5_outputs(6653) <= b;
    layer5_outputs(6654) <= not a or b;
    layer5_outputs(6655) <= not (a xor b);
    layer5_outputs(6656) <= not b;
    layer5_outputs(6657) <= b;
    layer5_outputs(6658) <= a and not b;
    layer5_outputs(6659) <= not (a or b);
    layer5_outputs(6660) <= '1';
    layer5_outputs(6661) <= a or b;
    layer5_outputs(6662) <= '1';
    layer5_outputs(6663) <= not (a and b);
    layer5_outputs(6664) <= not b;
    layer5_outputs(6665) <= a;
    layer5_outputs(6666) <= not b;
    layer5_outputs(6667) <= b and not a;
    layer5_outputs(6668) <= not b;
    layer5_outputs(6669) <= not a or b;
    layer5_outputs(6670) <= a and b;
    layer5_outputs(6671) <= not (a or b);
    layer5_outputs(6672) <= not b or a;
    layer5_outputs(6673) <= not (a or b);
    layer5_outputs(6674) <= b;
    layer5_outputs(6675) <= not (a xor b);
    layer5_outputs(6676) <= a;
    layer5_outputs(6677) <= a;
    layer5_outputs(6678) <= not (a xor b);
    layer5_outputs(6679) <= a and not b;
    layer5_outputs(6680) <= not b;
    layer5_outputs(6681) <= b;
    layer5_outputs(6682) <= a xor b;
    layer5_outputs(6683) <= not (a xor b);
    layer5_outputs(6684) <= not a;
    layer5_outputs(6685) <= not a;
    layer5_outputs(6686) <= '1';
    layer5_outputs(6687) <= not a;
    layer5_outputs(6688) <= a and not b;
    layer5_outputs(6689) <= a and not b;
    layer5_outputs(6690) <= not a;
    layer5_outputs(6691) <= '1';
    layer5_outputs(6692) <= b;
    layer5_outputs(6693) <= not (a and b);
    layer5_outputs(6694) <= a;
    layer5_outputs(6695) <= not (a and b);
    layer5_outputs(6696) <= not (a xor b);
    layer5_outputs(6697) <= a xor b;
    layer5_outputs(6698) <= b;
    layer5_outputs(6699) <= '0';
    layer5_outputs(6700) <= a and b;
    layer5_outputs(6701) <= not (a or b);
    layer5_outputs(6702) <= a;
    layer5_outputs(6703) <= not (a xor b);
    layer5_outputs(6704) <= not b or a;
    layer5_outputs(6705) <= not (a xor b);
    layer5_outputs(6706) <= a and not b;
    layer5_outputs(6707) <= '0';
    layer5_outputs(6708) <= b;
    layer5_outputs(6709) <= a xor b;
    layer5_outputs(6710) <= not b;
    layer5_outputs(6711) <= a and b;
    layer5_outputs(6712) <= not (a and b);
    layer5_outputs(6713) <= '1';
    layer5_outputs(6714) <= b;
    layer5_outputs(6715) <= not a;
    layer5_outputs(6716) <= a;
    layer5_outputs(6717) <= b;
    layer5_outputs(6718) <= not a;
    layer5_outputs(6719) <= b and not a;
    layer5_outputs(6720) <= not a;
    layer5_outputs(6721) <= not (a or b);
    layer5_outputs(6722) <= not (a and b);
    layer5_outputs(6723) <= not b or a;
    layer5_outputs(6724) <= b and not a;
    layer5_outputs(6725) <= not (a and b);
    layer5_outputs(6726) <= a xor b;
    layer5_outputs(6727) <= a and not b;
    layer5_outputs(6728) <= not (a and b);
    layer5_outputs(6729) <= b and not a;
    layer5_outputs(6730) <= not a;
    layer5_outputs(6731) <= b and not a;
    layer5_outputs(6732) <= a and not b;
    layer5_outputs(6733) <= b;
    layer5_outputs(6734) <= b;
    layer5_outputs(6735) <= not a;
    layer5_outputs(6736) <= a and not b;
    layer5_outputs(6737) <= a;
    layer5_outputs(6738) <= a or b;
    layer5_outputs(6739) <= not (a or b);
    layer5_outputs(6740) <= not b;
    layer5_outputs(6741) <= a;
    layer5_outputs(6742) <= not (a or b);
    layer5_outputs(6743) <= not a;
    layer5_outputs(6744) <= b;
    layer5_outputs(6745) <= b;
    layer5_outputs(6746) <= not b;
    layer5_outputs(6747) <= not b;
    layer5_outputs(6748) <= not a;
    layer5_outputs(6749) <= b;
    layer5_outputs(6750) <= not b;
    layer5_outputs(6751) <= not a;
    layer5_outputs(6752) <= '1';
    layer5_outputs(6753) <= a xor b;
    layer5_outputs(6754) <= not a;
    layer5_outputs(6755) <= b;
    layer5_outputs(6756) <= a xor b;
    layer5_outputs(6757) <= '0';
    layer5_outputs(6758) <= a;
    layer5_outputs(6759) <= a;
    layer5_outputs(6760) <= a and b;
    layer5_outputs(6761) <= a xor b;
    layer5_outputs(6762) <= a;
    layer5_outputs(6763) <= not (a or b);
    layer5_outputs(6764) <= not (a xor b);
    layer5_outputs(6765) <= not (a or b);
    layer5_outputs(6766) <= not a;
    layer5_outputs(6767) <= b;
    layer5_outputs(6768) <= not a;
    layer5_outputs(6769) <= a and b;
    layer5_outputs(6770) <= not b;
    layer5_outputs(6771) <= not (a xor b);
    layer5_outputs(6772) <= not (a or b);
    layer5_outputs(6773) <= b;
    layer5_outputs(6774) <= not a or b;
    layer5_outputs(6775) <= not (a xor b);
    layer5_outputs(6776) <= not b or a;
    layer5_outputs(6777) <= not a;
    layer5_outputs(6778) <= not b;
    layer5_outputs(6779) <= not b;
    layer5_outputs(6780) <= not (a and b);
    layer5_outputs(6781) <= a xor b;
    layer5_outputs(6782) <= not (a and b);
    layer5_outputs(6783) <= b and not a;
    layer5_outputs(6784) <= not a;
    layer5_outputs(6785) <= b;
    layer5_outputs(6786) <= not (a xor b);
    layer5_outputs(6787) <= not b;
    layer5_outputs(6788) <= not b;
    layer5_outputs(6789) <= a or b;
    layer5_outputs(6790) <= not (a xor b);
    layer5_outputs(6791) <= not b;
    layer5_outputs(6792) <= a;
    layer5_outputs(6793) <= not b;
    layer5_outputs(6794) <= a and b;
    layer5_outputs(6795) <= not a;
    layer5_outputs(6796) <= a xor b;
    layer5_outputs(6797) <= not (a xor b);
    layer5_outputs(6798) <= not b or a;
    layer5_outputs(6799) <= a or b;
    layer5_outputs(6800) <= '0';
    layer5_outputs(6801) <= not (a xor b);
    layer5_outputs(6802) <= not a;
    layer5_outputs(6803) <= not b or a;
    layer5_outputs(6804) <= not b;
    layer5_outputs(6805) <= a;
    layer5_outputs(6806) <= not (a or b);
    layer5_outputs(6807) <= not (a and b);
    layer5_outputs(6808) <= not a or b;
    layer5_outputs(6809) <= not b;
    layer5_outputs(6810) <= a and b;
    layer5_outputs(6811) <= b;
    layer5_outputs(6812) <= b;
    layer5_outputs(6813) <= not (a and b);
    layer5_outputs(6814) <= '1';
    layer5_outputs(6815) <= not b or a;
    layer5_outputs(6816) <= not (a and b);
    layer5_outputs(6817) <= a and b;
    layer5_outputs(6818) <= a or b;
    layer5_outputs(6819) <= a;
    layer5_outputs(6820) <= not a or b;
    layer5_outputs(6821) <= '1';
    layer5_outputs(6822) <= not b or a;
    layer5_outputs(6823) <= not a;
    layer5_outputs(6824) <= not a or b;
    layer5_outputs(6825) <= b;
    layer5_outputs(6826) <= a or b;
    layer5_outputs(6827) <= a xor b;
    layer5_outputs(6828) <= not b;
    layer5_outputs(6829) <= not b;
    layer5_outputs(6830) <= not a;
    layer5_outputs(6831) <= not (a or b);
    layer5_outputs(6832) <= not a or b;
    layer5_outputs(6833) <= a and b;
    layer5_outputs(6834) <= not a;
    layer5_outputs(6835) <= a and b;
    layer5_outputs(6836) <= not (a xor b);
    layer5_outputs(6837) <= not (a or b);
    layer5_outputs(6838) <= b;
    layer5_outputs(6839) <= not (a or b);
    layer5_outputs(6840) <= not b or a;
    layer5_outputs(6841) <= not b;
    layer5_outputs(6842) <= not (a and b);
    layer5_outputs(6843) <= not b;
    layer5_outputs(6844) <= b;
    layer5_outputs(6845) <= not a;
    layer5_outputs(6846) <= a xor b;
    layer5_outputs(6847) <= not a;
    layer5_outputs(6848) <= b;
    layer5_outputs(6849) <= not a;
    layer5_outputs(6850) <= not b or a;
    layer5_outputs(6851) <= a;
    layer5_outputs(6852) <= not a or b;
    layer5_outputs(6853) <= a or b;
    layer5_outputs(6854) <= not a or b;
    layer5_outputs(6855) <= not (a xor b);
    layer5_outputs(6856) <= b;
    layer5_outputs(6857) <= not (a and b);
    layer5_outputs(6858) <= not a or b;
    layer5_outputs(6859) <= a xor b;
    layer5_outputs(6860) <= a and not b;
    layer5_outputs(6861) <= not a;
    layer5_outputs(6862) <= not a;
    layer5_outputs(6863) <= b;
    layer5_outputs(6864) <= b;
    layer5_outputs(6865) <= not b;
    layer5_outputs(6866) <= not (a xor b);
    layer5_outputs(6867) <= not b;
    layer5_outputs(6868) <= not a;
    layer5_outputs(6869) <= not (a or b);
    layer5_outputs(6870) <= not a or b;
    layer5_outputs(6871) <= a and not b;
    layer5_outputs(6872) <= b;
    layer5_outputs(6873) <= a;
    layer5_outputs(6874) <= a;
    layer5_outputs(6875) <= not (a and b);
    layer5_outputs(6876) <= a xor b;
    layer5_outputs(6877) <= a xor b;
    layer5_outputs(6878) <= not b;
    layer5_outputs(6879) <= a and not b;
    layer5_outputs(6880) <= a;
    layer5_outputs(6881) <= a xor b;
    layer5_outputs(6882) <= not a;
    layer5_outputs(6883) <= b;
    layer5_outputs(6884) <= a and b;
    layer5_outputs(6885) <= not b;
    layer5_outputs(6886) <= a;
    layer5_outputs(6887) <= b;
    layer5_outputs(6888) <= not a;
    layer5_outputs(6889) <= a;
    layer5_outputs(6890) <= not b or a;
    layer5_outputs(6891) <= not (a and b);
    layer5_outputs(6892) <= not a or b;
    layer5_outputs(6893) <= not a or b;
    layer5_outputs(6894) <= not (a or b);
    layer5_outputs(6895) <= not b;
    layer5_outputs(6896) <= not (a xor b);
    layer5_outputs(6897) <= a xor b;
    layer5_outputs(6898) <= not a;
    layer5_outputs(6899) <= b and not a;
    layer5_outputs(6900) <= not (a and b);
    layer5_outputs(6901) <= b;
    layer5_outputs(6902) <= b;
    layer5_outputs(6903) <= a xor b;
    layer5_outputs(6904) <= not (a xor b);
    layer5_outputs(6905) <= a and not b;
    layer5_outputs(6906) <= b;
    layer5_outputs(6907) <= not a;
    layer5_outputs(6908) <= not a;
    layer5_outputs(6909) <= a;
    layer5_outputs(6910) <= a and b;
    layer5_outputs(6911) <= a and not b;
    layer5_outputs(6912) <= a or b;
    layer5_outputs(6913) <= not (a xor b);
    layer5_outputs(6914) <= b;
    layer5_outputs(6915) <= not a;
    layer5_outputs(6916) <= b and not a;
    layer5_outputs(6917) <= not (a xor b);
    layer5_outputs(6918) <= b and not a;
    layer5_outputs(6919) <= b;
    layer5_outputs(6920) <= b and not a;
    layer5_outputs(6921) <= '1';
    layer5_outputs(6922) <= b;
    layer5_outputs(6923) <= not (a xor b);
    layer5_outputs(6924) <= not (a and b);
    layer5_outputs(6925) <= not b;
    layer5_outputs(6926) <= not a;
    layer5_outputs(6927) <= not (a and b);
    layer5_outputs(6928) <= not (a or b);
    layer5_outputs(6929) <= not a or b;
    layer5_outputs(6930) <= a and not b;
    layer5_outputs(6931) <= not a;
    layer5_outputs(6932) <= not (a and b);
    layer5_outputs(6933) <= b and not a;
    layer5_outputs(6934) <= b and not a;
    layer5_outputs(6935) <= not a;
    layer5_outputs(6936) <= b;
    layer5_outputs(6937) <= not a;
    layer5_outputs(6938) <= a xor b;
    layer5_outputs(6939) <= not a or b;
    layer5_outputs(6940) <= not b or a;
    layer5_outputs(6941) <= not a;
    layer5_outputs(6942) <= not b;
    layer5_outputs(6943) <= b;
    layer5_outputs(6944) <= a and not b;
    layer5_outputs(6945) <= a or b;
    layer5_outputs(6946) <= not a;
    layer5_outputs(6947) <= not a or b;
    layer5_outputs(6948) <= not (a xor b);
    layer5_outputs(6949) <= a xor b;
    layer5_outputs(6950) <= a or b;
    layer5_outputs(6951) <= not (a and b);
    layer5_outputs(6952) <= not b;
    layer5_outputs(6953) <= a xor b;
    layer5_outputs(6954) <= not b;
    layer5_outputs(6955) <= not a;
    layer5_outputs(6956) <= not b or a;
    layer5_outputs(6957) <= a xor b;
    layer5_outputs(6958) <= a and not b;
    layer5_outputs(6959) <= not b or a;
    layer5_outputs(6960) <= a and not b;
    layer5_outputs(6961) <= a;
    layer5_outputs(6962) <= b;
    layer5_outputs(6963) <= b;
    layer5_outputs(6964) <= a xor b;
    layer5_outputs(6965) <= a or b;
    layer5_outputs(6966) <= '0';
    layer5_outputs(6967) <= a or b;
    layer5_outputs(6968) <= a and b;
    layer5_outputs(6969) <= not b;
    layer5_outputs(6970) <= not (a xor b);
    layer5_outputs(6971) <= not (a and b);
    layer5_outputs(6972) <= b;
    layer5_outputs(6973) <= not a;
    layer5_outputs(6974) <= b;
    layer5_outputs(6975) <= b;
    layer5_outputs(6976) <= a;
    layer5_outputs(6977) <= not (a xor b);
    layer5_outputs(6978) <= not b;
    layer5_outputs(6979) <= not (a or b);
    layer5_outputs(6980) <= a or b;
    layer5_outputs(6981) <= b and not a;
    layer5_outputs(6982) <= a or b;
    layer5_outputs(6983) <= b;
    layer5_outputs(6984) <= a xor b;
    layer5_outputs(6985) <= not a;
    layer5_outputs(6986) <= not a;
    layer5_outputs(6987) <= not (a or b);
    layer5_outputs(6988) <= a and not b;
    layer5_outputs(6989) <= not a or b;
    layer5_outputs(6990) <= not (a xor b);
    layer5_outputs(6991) <= b;
    layer5_outputs(6992) <= not (a and b);
    layer5_outputs(6993) <= not (a xor b);
    layer5_outputs(6994) <= a;
    layer5_outputs(6995) <= not b or a;
    layer5_outputs(6996) <= b;
    layer5_outputs(6997) <= not (a xor b);
    layer5_outputs(6998) <= not b;
    layer5_outputs(6999) <= a and b;
    layer5_outputs(7000) <= a;
    layer5_outputs(7001) <= not (a or b);
    layer5_outputs(7002) <= not b;
    layer5_outputs(7003) <= a;
    layer5_outputs(7004) <= b;
    layer5_outputs(7005) <= not a;
    layer5_outputs(7006) <= not a;
    layer5_outputs(7007) <= b;
    layer5_outputs(7008) <= a;
    layer5_outputs(7009) <= b;
    layer5_outputs(7010) <= a and b;
    layer5_outputs(7011) <= not (a and b);
    layer5_outputs(7012) <= not (a xor b);
    layer5_outputs(7013) <= a and b;
    layer5_outputs(7014) <= a and b;
    layer5_outputs(7015) <= not b;
    layer5_outputs(7016) <= '1';
    layer5_outputs(7017) <= not a;
    layer5_outputs(7018) <= not (a xor b);
    layer5_outputs(7019) <= not b;
    layer5_outputs(7020) <= a;
    layer5_outputs(7021) <= not (a or b);
    layer5_outputs(7022) <= not b;
    layer5_outputs(7023) <= not b;
    layer5_outputs(7024) <= not b;
    layer5_outputs(7025) <= not (a and b);
    layer5_outputs(7026) <= a;
    layer5_outputs(7027) <= not b;
    layer5_outputs(7028) <= b and not a;
    layer5_outputs(7029) <= not b;
    layer5_outputs(7030) <= not b or a;
    layer5_outputs(7031) <= a xor b;
    layer5_outputs(7032) <= a and b;
    layer5_outputs(7033) <= a and b;
    layer5_outputs(7034) <= b;
    layer5_outputs(7035) <= a;
    layer5_outputs(7036) <= a and b;
    layer5_outputs(7037) <= not b or a;
    layer5_outputs(7038) <= not b;
    layer5_outputs(7039) <= not (a and b);
    layer5_outputs(7040) <= not b;
    layer5_outputs(7041) <= a and not b;
    layer5_outputs(7042) <= not (a xor b);
    layer5_outputs(7043) <= not b or a;
    layer5_outputs(7044) <= b;
    layer5_outputs(7045) <= a and not b;
    layer5_outputs(7046) <= not b;
    layer5_outputs(7047) <= not b or a;
    layer5_outputs(7048) <= not (a or b);
    layer5_outputs(7049) <= not b;
    layer5_outputs(7050) <= a xor b;
    layer5_outputs(7051) <= not a or b;
    layer5_outputs(7052) <= not a or b;
    layer5_outputs(7053) <= not b;
    layer5_outputs(7054) <= not b or a;
    layer5_outputs(7055) <= a;
    layer5_outputs(7056) <= a;
    layer5_outputs(7057) <= b;
    layer5_outputs(7058) <= not (a and b);
    layer5_outputs(7059) <= not a;
    layer5_outputs(7060) <= a;
    layer5_outputs(7061) <= a and b;
    layer5_outputs(7062) <= not b or a;
    layer5_outputs(7063) <= a;
    layer5_outputs(7064) <= not b;
    layer5_outputs(7065) <= a and not b;
    layer5_outputs(7066) <= a or b;
    layer5_outputs(7067) <= not (a xor b);
    layer5_outputs(7068) <= a or b;
    layer5_outputs(7069) <= b and not a;
    layer5_outputs(7070) <= '0';
    layer5_outputs(7071) <= a;
    layer5_outputs(7072) <= '0';
    layer5_outputs(7073) <= not (a xor b);
    layer5_outputs(7074) <= a;
    layer5_outputs(7075) <= not (a xor b);
    layer5_outputs(7076) <= not b;
    layer5_outputs(7077) <= not a or b;
    layer5_outputs(7078) <= not b or a;
    layer5_outputs(7079) <= b;
    layer5_outputs(7080) <= a and b;
    layer5_outputs(7081) <= not b;
    layer5_outputs(7082) <= b and not a;
    layer5_outputs(7083) <= not (a xor b);
    layer5_outputs(7084) <= not (a and b);
    layer5_outputs(7085) <= b;
    layer5_outputs(7086) <= not (a and b);
    layer5_outputs(7087) <= not (a xor b);
    layer5_outputs(7088) <= not a;
    layer5_outputs(7089) <= a;
    layer5_outputs(7090) <= a and b;
    layer5_outputs(7091) <= a or b;
    layer5_outputs(7092) <= not a;
    layer5_outputs(7093) <= b and not a;
    layer5_outputs(7094) <= not (a or b);
    layer5_outputs(7095) <= not (a and b);
    layer5_outputs(7096) <= not b;
    layer5_outputs(7097) <= not (a or b);
    layer5_outputs(7098) <= not (a and b);
    layer5_outputs(7099) <= a and b;
    layer5_outputs(7100) <= a xor b;
    layer5_outputs(7101) <= not b;
    layer5_outputs(7102) <= b and not a;
    layer5_outputs(7103) <= not b;
    layer5_outputs(7104) <= not b or a;
    layer5_outputs(7105) <= b;
    layer5_outputs(7106) <= not (a and b);
    layer5_outputs(7107) <= not b;
    layer5_outputs(7108) <= '0';
    layer5_outputs(7109) <= not b;
    layer5_outputs(7110) <= a and not b;
    layer5_outputs(7111) <= b;
    layer5_outputs(7112) <= b and not a;
    layer5_outputs(7113) <= b;
    layer5_outputs(7114) <= b and not a;
    layer5_outputs(7115) <= not b;
    layer5_outputs(7116) <= a;
    layer5_outputs(7117) <= a or b;
    layer5_outputs(7118) <= not a;
    layer5_outputs(7119) <= b;
    layer5_outputs(7120) <= a;
    layer5_outputs(7121) <= not b;
    layer5_outputs(7122) <= not (a and b);
    layer5_outputs(7123) <= not (a or b);
    layer5_outputs(7124) <= b;
    layer5_outputs(7125) <= a or b;
    layer5_outputs(7126) <= b;
    layer5_outputs(7127) <= a xor b;
    layer5_outputs(7128) <= a xor b;
    layer5_outputs(7129) <= a;
    layer5_outputs(7130) <= a;
    layer5_outputs(7131) <= b;
    layer5_outputs(7132) <= not a;
    layer5_outputs(7133) <= a;
    layer5_outputs(7134) <= not (a xor b);
    layer5_outputs(7135) <= not (a xor b);
    layer5_outputs(7136) <= not a or b;
    layer5_outputs(7137) <= not a or b;
    layer5_outputs(7138) <= not a;
    layer5_outputs(7139) <= not (a or b);
    layer5_outputs(7140) <= a or b;
    layer5_outputs(7141) <= not (a xor b);
    layer5_outputs(7142) <= not b or a;
    layer5_outputs(7143) <= a xor b;
    layer5_outputs(7144) <= not b;
    layer5_outputs(7145) <= b;
    layer5_outputs(7146) <= not a;
    layer5_outputs(7147) <= not (a and b);
    layer5_outputs(7148) <= b and not a;
    layer5_outputs(7149) <= not a;
    layer5_outputs(7150) <= b;
    layer5_outputs(7151) <= not (a or b);
    layer5_outputs(7152) <= not a or b;
    layer5_outputs(7153) <= not b;
    layer5_outputs(7154) <= not a or b;
    layer5_outputs(7155) <= not b;
    layer5_outputs(7156) <= a;
    layer5_outputs(7157) <= a;
    layer5_outputs(7158) <= not (a xor b);
    layer5_outputs(7159) <= a;
    layer5_outputs(7160) <= not b;
    layer5_outputs(7161) <= a or b;
    layer5_outputs(7162) <= a;
    layer5_outputs(7163) <= b;
    layer5_outputs(7164) <= b;
    layer5_outputs(7165) <= a;
    layer5_outputs(7166) <= not (a xor b);
    layer5_outputs(7167) <= b;
    layer5_outputs(7168) <= not b;
    layer5_outputs(7169) <= a and b;
    layer5_outputs(7170) <= not (a or b);
    layer5_outputs(7171) <= not b or a;
    layer5_outputs(7172) <= not (a and b);
    layer5_outputs(7173) <= a;
    layer5_outputs(7174) <= a;
    layer5_outputs(7175) <= not b;
    layer5_outputs(7176) <= a or b;
    layer5_outputs(7177) <= not a or b;
    layer5_outputs(7178) <= a and not b;
    layer5_outputs(7179) <= not (a xor b);
    layer5_outputs(7180) <= not a or b;
    layer5_outputs(7181) <= a;
    layer5_outputs(7182) <= not (a and b);
    layer5_outputs(7183) <= not a or b;
    layer5_outputs(7184) <= a;
    layer5_outputs(7185) <= b;
    layer5_outputs(7186) <= not b;
    layer5_outputs(7187) <= not (a or b);
    layer5_outputs(7188) <= a;
    layer5_outputs(7189) <= not a or b;
    layer5_outputs(7190) <= not (a or b);
    layer5_outputs(7191) <= a and not b;
    layer5_outputs(7192) <= a;
    layer5_outputs(7193) <= a and not b;
    layer5_outputs(7194) <= not (a or b);
    layer5_outputs(7195) <= b and not a;
    layer5_outputs(7196) <= b;
    layer5_outputs(7197) <= not (a and b);
    layer5_outputs(7198) <= a and b;
    layer5_outputs(7199) <= b;
    layer5_outputs(7200) <= a and not b;
    layer5_outputs(7201) <= not (a xor b);
    layer5_outputs(7202) <= a and b;
    layer5_outputs(7203) <= a;
    layer5_outputs(7204) <= not a;
    layer5_outputs(7205) <= not b;
    layer5_outputs(7206) <= a xor b;
    layer5_outputs(7207) <= not b;
    layer5_outputs(7208) <= not a;
    layer5_outputs(7209) <= a;
    layer5_outputs(7210) <= b;
    layer5_outputs(7211) <= b;
    layer5_outputs(7212) <= not (a xor b);
    layer5_outputs(7213) <= b;
    layer5_outputs(7214) <= not a or b;
    layer5_outputs(7215) <= not b;
    layer5_outputs(7216) <= not a or b;
    layer5_outputs(7217) <= b;
    layer5_outputs(7218) <= not b;
    layer5_outputs(7219) <= not (a and b);
    layer5_outputs(7220) <= a xor b;
    layer5_outputs(7221) <= a and b;
    layer5_outputs(7222) <= b and not a;
    layer5_outputs(7223) <= a or b;
    layer5_outputs(7224) <= not b or a;
    layer5_outputs(7225) <= not a or b;
    layer5_outputs(7226) <= not a or b;
    layer5_outputs(7227) <= not a;
    layer5_outputs(7228) <= a or b;
    layer5_outputs(7229) <= not b or a;
    layer5_outputs(7230) <= not a;
    layer5_outputs(7231) <= not a or b;
    layer5_outputs(7232) <= a and b;
    layer5_outputs(7233) <= b;
    layer5_outputs(7234) <= not a;
    layer5_outputs(7235) <= not (a xor b);
    layer5_outputs(7236) <= not b or a;
    layer5_outputs(7237) <= a;
    layer5_outputs(7238) <= not a;
    layer5_outputs(7239) <= b and not a;
    layer5_outputs(7240) <= a and not b;
    layer5_outputs(7241) <= not (a xor b);
    layer5_outputs(7242) <= not a;
    layer5_outputs(7243) <= '0';
    layer5_outputs(7244) <= a and b;
    layer5_outputs(7245) <= b;
    layer5_outputs(7246) <= not b;
    layer5_outputs(7247) <= not (a xor b);
    layer5_outputs(7248) <= b;
    layer5_outputs(7249) <= not a;
    layer5_outputs(7250) <= b;
    layer5_outputs(7251) <= not a;
    layer5_outputs(7252) <= not b;
    layer5_outputs(7253) <= not (a and b);
    layer5_outputs(7254) <= a;
    layer5_outputs(7255) <= b;
    layer5_outputs(7256) <= a;
    layer5_outputs(7257) <= not b;
    layer5_outputs(7258) <= not (a and b);
    layer5_outputs(7259) <= b and not a;
    layer5_outputs(7260) <= a xor b;
    layer5_outputs(7261) <= b;
    layer5_outputs(7262) <= a xor b;
    layer5_outputs(7263) <= not b;
    layer5_outputs(7264) <= a xor b;
    layer5_outputs(7265) <= b;
    layer5_outputs(7266) <= b and not a;
    layer5_outputs(7267) <= not (a xor b);
    layer5_outputs(7268) <= not b;
    layer5_outputs(7269) <= not (a and b);
    layer5_outputs(7270) <= not (a or b);
    layer5_outputs(7271) <= not a or b;
    layer5_outputs(7272) <= a;
    layer5_outputs(7273) <= not b;
    layer5_outputs(7274) <= not a or b;
    layer5_outputs(7275) <= not a;
    layer5_outputs(7276) <= b and not a;
    layer5_outputs(7277) <= a xor b;
    layer5_outputs(7278) <= not b;
    layer5_outputs(7279) <= not b;
    layer5_outputs(7280) <= b and not a;
    layer5_outputs(7281) <= b and not a;
    layer5_outputs(7282) <= not a;
    layer5_outputs(7283) <= b and not a;
    layer5_outputs(7284) <= a;
    layer5_outputs(7285) <= b;
    layer5_outputs(7286) <= b;
    layer5_outputs(7287) <= not (a xor b);
    layer5_outputs(7288) <= a and not b;
    layer5_outputs(7289) <= not b or a;
    layer5_outputs(7290) <= not b;
    layer5_outputs(7291) <= not a or b;
    layer5_outputs(7292) <= not a;
    layer5_outputs(7293) <= not a or b;
    layer5_outputs(7294) <= a and b;
    layer5_outputs(7295) <= a xor b;
    layer5_outputs(7296) <= b;
    layer5_outputs(7297) <= a or b;
    layer5_outputs(7298) <= not (a xor b);
    layer5_outputs(7299) <= a xor b;
    layer5_outputs(7300) <= not a;
    layer5_outputs(7301) <= a or b;
    layer5_outputs(7302) <= a and not b;
    layer5_outputs(7303) <= not a;
    layer5_outputs(7304) <= not b;
    layer5_outputs(7305) <= b;
    layer5_outputs(7306) <= b;
    layer5_outputs(7307) <= b and not a;
    layer5_outputs(7308) <= a and not b;
    layer5_outputs(7309) <= not b or a;
    layer5_outputs(7310) <= '0';
    layer5_outputs(7311) <= not (a or b);
    layer5_outputs(7312) <= not (a or b);
    layer5_outputs(7313) <= not a;
    layer5_outputs(7314) <= a;
    layer5_outputs(7315) <= a xor b;
    layer5_outputs(7316) <= not b;
    layer5_outputs(7317) <= a or b;
    layer5_outputs(7318) <= a;
    layer5_outputs(7319) <= not b;
    layer5_outputs(7320) <= a xor b;
    layer5_outputs(7321) <= not (a xor b);
    layer5_outputs(7322) <= a xor b;
    layer5_outputs(7323) <= a and b;
    layer5_outputs(7324) <= a and b;
    layer5_outputs(7325) <= not b or a;
    layer5_outputs(7326) <= not b;
    layer5_outputs(7327) <= not b;
    layer5_outputs(7328) <= not a or b;
    layer5_outputs(7329) <= a;
    layer5_outputs(7330) <= not b;
    layer5_outputs(7331) <= a and b;
    layer5_outputs(7332) <= b and not a;
    layer5_outputs(7333) <= not a;
    layer5_outputs(7334) <= not a;
    layer5_outputs(7335) <= not (a xor b);
    layer5_outputs(7336) <= a and b;
    layer5_outputs(7337) <= a or b;
    layer5_outputs(7338) <= not a;
    layer5_outputs(7339) <= not (a xor b);
    layer5_outputs(7340) <= b;
    layer5_outputs(7341) <= not a;
    layer5_outputs(7342) <= not b or a;
    layer5_outputs(7343) <= b and not a;
    layer5_outputs(7344) <= a;
    layer5_outputs(7345) <= a;
    layer5_outputs(7346) <= not (a or b);
    layer5_outputs(7347) <= a and b;
    layer5_outputs(7348) <= a xor b;
    layer5_outputs(7349) <= a xor b;
    layer5_outputs(7350) <= not (a or b);
    layer5_outputs(7351) <= not b;
    layer5_outputs(7352) <= not a or b;
    layer5_outputs(7353) <= a and b;
    layer5_outputs(7354) <= a or b;
    layer5_outputs(7355) <= not b;
    layer5_outputs(7356) <= not (a or b);
    layer5_outputs(7357) <= b;
    layer5_outputs(7358) <= a;
    layer5_outputs(7359) <= not (a xor b);
    layer5_outputs(7360) <= a and not b;
    layer5_outputs(7361) <= a or b;
    layer5_outputs(7362) <= not a;
    layer5_outputs(7363) <= not b or a;
    layer5_outputs(7364) <= not (a or b);
    layer5_outputs(7365) <= a and not b;
    layer5_outputs(7366) <= not (a xor b);
    layer5_outputs(7367) <= not b or a;
    layer5_outputs(7368) <= not (a or b);
    layer5_outputs(7369) <= not a;
    layer5_outputs(7370) <= not a;
    layer5_outputs(7371) <= not b;
    layer5_outputs(7372) <= not a;
    layer5_outputs(7373) <= b and not a;
    layer5_outputs(7374) <= b;
    layer5_outputs(7375) <= b and not a;
    layer5_outputs(7376) <= a xor b;
    layer5_outputs(7377) <= a;
    layer5_outputs(7378) <= not b;
    layer5_outputs(7379) <= not (a or b);
    layer5_outputs(7380) <= not a;
    layer5_outputs(7381) <= a and b;
    layer5_outputs(7382) <= b;
    layer5_outputs(7383) <= not a;
    layer5_outputs(7384) <= not (a and b);
    layer5_outputs(7385) <= not (a or b);
    layer5_outputs(7386) <= not a;
    layer5_outputs(7387) <= a xor b;
    layer5_outputs(7388) <= a;
    layer5_outputs(7389) <= a;
    layer5_outputs(7390) <= not b;
    layer5_outputs(7391) <= b;
    layer5_outputs(7392) <= not (a and b);
    layer5_outputs(7393) <= not a;
    layer5_outputs(7394) <= a;
    layer5_outputs(7395) <= a;
    layer5_outputs(7396) <= not (a or b);
    layer5_outputs(7397) <= a or b;
    layer5_outputs(7398) <= not (a xor b);
    layer5_outputs(7399) <= not a or b;
    layer5_outputs(7400) <= a;
    layer5_outputs(7401) <= a and not b;
    layer5_outputs(7402) <= a xor b;
    layer5_outputs(7403) <= a or b;
    layer5_outputs(7404) <= b;
    layer5_outputs(7405) <= a and not b;
    layer5_outputs(7406) <= '0';
    layer5_outputs(7407) <= not (a or b);
    layer5_outputs(7408) <= not (a or b);
    layer5_outputs(7409) <= not b;
    layer5_outputs(7410) <= '0';
    layer5_outputs(7411) <= not (a xor b);
    layer5_outputs(7412) <= a;
    layer5_outputs(7413) <= not a or b;
    layer5_outputs(7414) <= not a;
    layer5_outputs(7415) <= b and not a;
    layer5_outputs(7416) <= not b or a;
    layer5_outputs(7417) <= a and b;
    layer5_outputs(7418) <= not b or a;
    layer5_outputs(7419) <= not a;
    layer5_outputs(7420) <= not a;
    layer5_outputs(7421) <= not b;
    layer5_outputs(7422) <= not b or a;
    layer5_outputs(7423) <= not b;
    layer5_outputs(7424) <= not a;
    layer5_outputs(7425) <= not (a and b);
    layer5_outputs(7426) <= not a;
    layer5_outputs(7427) <= b;
    layer5_outputs(7428) <= a xor b;
    layer5_outputs(7429) <= a;
    layer5_outputs(7430) <= a and not b;
    layer5_outputs(7431) <= a;
    layer5_outputs(7432) <= not a;
    layer5_outputs(7433) <= b and not a;
    layer5_outputs(7434) <= a;
    layer5_outputs(7435) <= a and b;
    layer5_outputs(7436) <= not (a or b);
    layer5_outputs(7437) <= not b;
    layer5_outputs(7438) <= not b;
    layer5_outputs(7439) <= not b or a;
    layer5_outputs(7440) <= b;
    layer5_outputs(7441) <= a or b;
    layer5_outputs(7442) <= not a;
    layer5_outputs(7443) <= a and b;
    layer5_outputs(7444) <= a or b;
    layer5_outputs(7445) <= b;
    layer5_outputs(7446) <= a;
    layer5_outputs(7447) <= b and not a;
    layer5_outputs(7448) <= b;
    layer5_outputs(7449) <= a xor b;
    layer5_outputs(7450) <= not a;
    layer5_outputs(7451) <= not a;
    layer5_outputs(7452) <= not b;
    layer5_outputs(7453) <= not a;
    layer5_outputs(7454) <= not (a or b);
    layer5_outputs(7455) <= a;
    layer5_outputs(7456) <= a xor b;
    layer5_outputs(7457) <= a;
    layer5_outputs(7458) <= a and b;
    layer5_outputs(7459) <= b;
    layer5_outputs(7460) <= a;
    layer5_outputs(7461) <= not (a and b);
    layer5_outputs(7462) <= not a;
    layer5_outputs(7463) <= not (a and b);
    layer5_outputs(7464) <= not (a and b);
    layer5_outputs(7465) <= a and b;
    layer5_outputs(7466) <= not b;
    layer5_outputs(7467) <= not (a xor b);
    layer5_outputs(7468) <= b;
    layer5_outputs(7469) <= not b or a;
    layer5_outputs(7470) <= a;
    layer5_outputs(7471) <= not a or b;
    layer5_outputs(7472) <= a or b;
    layer5_outputs(7473) <= b;
    layer5_outputs(7474) <= not a;
    layer5_outputs(7475) <= not b or a;
    layer5_outputs(7476) <= a or b;
    layer5_outputs(7477) <= not (a or b);
    layer5_outputs(7478) <= not b;
    layer5_outputs(7479) <= a;
    layer5_outputs(7480) <= a;
    layer5_outputs(7481) <= not (a xor b);
    layer5_outputs(7482) <= not (a or b);
    layer5_outputs(7483) <= not a;
    layer5_outputs(7484) <= not b;
    layer5_outputs(7485) <= a;
    layer5_outputs(7486) <= not a;
    layer5_outputs(7487) <= not b;
    layer5_outputs(7488) <= a;
    layer5_outputs(7489) <= b;
    layer5_outputs(7490) <= a;
    layer5_outputs(7491) <= not b;
    layer5_outputs(7492) <= not (a or b);
    layer5_outputs(7493) <= not (a and b);
    layer5_outputs(7494) <= not a;
    layer5_outputs(7495) <= b and not a;
    layer5_outputs(7496) <= not b;
    layer5_outputs(7497) <= b;
    layer5_outputs(7498) <= a and not b;
    layer5_outputs(7499) <= b;
    layer5_outputs(7500) <= not a;
    layer5_outputs(7501) <= a;
    layer5_outputs(7502) <= a xor b;
    layer5_outputs(7503) <= a;
    layer5_outputs(7504) <= a or b;
    layer5_outputs(7505) <= not b;
    layer5_outputs(7506) <= not a or b;
    layer5_outputs(7507) <= not a or b;
    layer5_outputs(7508) <= not (a or b);
    layer5_outputs(7509) <= not (a or b);
    layer5_outputs(7510) <= b and not a;
    layer5_outputs(7511) <= not a;
    layer5_outputs(7512) <= not (a xor b);
    layer5_outputs(7513) <= not a;
    layer5_outputs(7514) <= a or b;
    layer5_outputs(7515) <= b and not a;
    layer5_outputs(7516) <= a and not b;
    layer5_outputs(7517) <= a or b;
    layer5_outputs(7518) <= b;
    layer5_outputs(7519) <= not b or a;
    layer5_outputs(7520) <= a and not b;
    layer5_outputs(7521) <= not (a xor b);
    layer5_outputs(7522) <= not b or a;
    layer5_outputs(7523) <= a;
    layer5_outputs(7524) <= a xor b;
    layer5_outputs(7525) <= not b;
    layer5_outputs(7526) <= not a or b;
    layer5_outputs(7527) <= not b;
    layer5_outputs(7528) <= a and b;
    layer5_outputs(7529) <= a or b;
    layer5_outputs(7530) <= not (a and b);
    layer5_outputs(7531) <= a and b;
    layer5_outputs(7532) <= b;
    layer5_outputs(7533) <= not a;
    layer5_outputs(7534) <= a xor b;
    layer5_outputs(7535) <= not (a and b);
    layer5_outputs(7536) <= not b;
    layer5_outputs(7537) <= b and not a;
    layer5_outputs(7538) <= b;
    layer5_outputs(7539) <= not b or a;
    layer5_outputs(7540) <= a or b;
    layer5_outputs(7541) <= a;
    layer5_outputs(7542) <= a;
    layer5_outputs(7543) <= a;
    layer5_outputs(7544) <= b;
    layer5_outputs(7545) <= not b;
    layer5_outputs(7546) <= a xor b;
    layer5_outputs(7547) <= not b or a;
    layer5_outputs(7548) <= b and not a;
    layer5_outputs(7549) <= not b or a;
    layer5_outputs(7550) <= b;
    layer5_outputs(7551) <= a and not b;
    layer5_outputs(7552) <= b;
    layer5_outputs(7553) <= '1';
    layer5_outputs(7554) <= not a or b;
    layer5_outputs(7555) <= not a or b;
    layer5_outputs(7556) <= a or b;
    layer5_outputs(7557) <= a;
    layer5_outputs(7558) <= a or b;
    layer5_outputs(7559) <= a and b;
    layer5_outputs(7560) <= b;
    layer5_outputs(7561) <= not b;
    layer5_outputs(7562) <= not (a or b);
    layer5_outputs(7563) <= a and b;
    layer5_outputs(7564) <= not a;
    layer5_outputs(7565) <= not a;
    layer5_outputs(7566) <= not (a or b);
    layer5_outputs(7567) <= not a;
    layer5_outputs(7568) <= a;
    layer5_outputs(7569) <= not b or a;
    layer5_outputs(7570) <= not (a and b);
    layer5_outputs(7571) <= not a;
    layer5_outputs(7572) <= not (a xor b);
    layer5_outputs(7573) <= not a;
    layer5_outputs(7574) <= a;
    layer5_outputs(7575) <= not b or a;
    layer5_outputs(7576) <= not b;
    layer5_outputs(7577) <= a;
    layer5_outputs(7578) <= a;
    layer5_outputs(7579) <= a or b;
    layer5_outputs(7580) <= b and not a;
    layer5_outputs(7581) <= not b or a;
    layer5_outputs(7582) <= b;
    layer5_outputs(7583) <= not (a xor b);
    layer5_outputs(7584) <= not b;
    layer5_outputs(7585) <= not b;
    layer5_outputs(7586) <= a;
    layer5_outputs(7587) <= not (a and b);
    layer5_outputs(7588) <= not (a xor b);
    layer5_outputs(7589) <= a or b;
    layer5_outputs(7590) <= not b;
    layer5_outputs(7591) <= b;
    layer5_outputs(7592) <= not (a or b);
    layer5_outputs(7593) <= not (a xor b);
    layer5_outputs(7594) <= not b or a;
    layer5_outputs(7595) <= a;
    layer5_outputs(7596) <= not (a and b);
    layer5_outputs(7597) <= not b;
    layer5_outputs(7598) <= not b;
    layer5_outputs(7599) <= not (a or b);
    layer5_outputs(7600) <= a;
    layer5_outputs(7601) <= a xor b;
    layer5_outputs(7602) <= a xor b;
    layer5_outputs(7603) <= a;
    layer5_outputs(7604) <= not (a or b);
    layer5_outputs(7605) <= not b;
    layer5_outputs(7606) <= not b;
    layer5_outputs(7607) <= not (a xor b);
    layer5_outputs(7608) <= b and not a;
    layer5_outputs(7609) <= not b;
    layer5_outputs(7610) <= a xor b;
    layer5_outputs(7611) <= not a or b;
    layer5_outputs(7612) <= a;
    layer5_outputs(7613) <= b;
    layer5_outputs(7614) <= b;
    layer5_outputs(7615) <= not a;
    layer5_outputs(7616) <= not b;
    layer5_outputs(7617) <= not (a or b);
    layer5_outputs(7618) <= a and not b;
    layer5_outputs(7619) <= a;
    layer5_outputs(7620) <= a or b;
    layer5_outputs(7621) <= not a;
    layer5_outputs(7622) <= b and not a;
    layer5_outputs(7623) <= '0';
    layer5_outputs(7624) <= not b;
    layer5_outputs(7625) <= not a or b;
    layer5_outputs(7626) <= a xor b;
    layer5_outputs(7627) <= not a or b;
    layer5_outputs(7628) <= not b or a;
    layer5_outputs(7629) <= a or b;
    layer5_outputs(7630) <= b;
    layer5_outputs(7631) <= a xor b;
    layer5_outputs(7632) <= not a;
    layer5_outputs(7633) <= not b;
    layer5_outputs(7634) <= b;
    layer5_outputs(7635) <= not (a or b);
    layer5_outputs(7636) <= not b;
    layer5_outputs(7637) <= not (a xor b);
    layer5_outputs(7638) <= a and not b;
    layer5_outputs(7639) <= '1';
    layer5_outputs(7640) <= a xor b;
    layer5_outputs(7641) <= not b or a;
    layer5_outputs(7642) <= a;
    layer5_outputs(7643) <= not a;
    layer5_outputs(7644) <= a xor b;
    layer5_outputs(7645) <= b;
    layer5_outputs(7646) <= not b or a;
    layer5_outputs(7647) <= not b;
    layer5_outputs(7648) <= b;
    layer5_outputs(7649) <= not (a and b);
    layer5_outputs(7650) <= not b or a;
    layer5_outputs(7651) <= not b;
    layer5_outputs(7652) <= a;
    layer5_outputs(7653) <= b and not a;
    layer5_outputs(7654) <= not b or a;
    layer5_outputs(7655) <= not (a xor b);
    layer5_outputs(7656) <= b;
    layer5_outputs(7657) <= not (a and b);
    layer5_outputs(7658) <= not (a xor b);
    layer5_outputs(7659) <= a;
    layer5_outputs(7660) <= not (a and b);
    layer5_outputs(7661) <= not b;
    layer5_outputs(7662) <= not b;
    layer5_outputs(7663) <= not a;
    layer5_outputs(7664) <= not (a xor b);
    layer5_outputs(7665) <= b;
    layer5_outputs(7666) <= not (a xor b);
    layer5_outputs(7667) <= a or b;
    layer5_outputs(7668) <= a and not b;
    layer5_outputs(7669) <= not (a xor b);
    layer5_outputs(7670) <= a;
    layer5_outputs(7671) <= a xor b;
    layer5_outputs(7672) <= a;
    layer5_outputs(7673) <= not b or a;
    layer5_outputs(7674) <= a and not b;
    layer5_outputs(7675) <= a and b;
    layer5_outputs(7676) <= a;
    layer5_outputs(7677) <= b and not a;
    layer5_outputs(7678) <= a and not b;
    layer5_outputs(7679) <= not a or b;
    layer5_outputs(7680) <= a and not b;
    layer5_outputs(7681) <= '0';
    layer5_outputs(7682) <= a;
    layer5_outputs(7683) <= a or b;
    layer5_outputs(7684) <= b;
    layer5_outputs(7685) <= not a;
    layer5_outputs(7686) <= a xor b;
    layer5_outputs(7687) <= a and not b;
    layer5_outputs(7688) <= not (a or b);
    layer5_outputs(7689) <= b and not a;
    layer5_outputs(7690) <= not (a xor b);
    layer5_outputs(7691) <= not a;
    layer5_outputs(7692) <= not b or a;
    layer5_outputs(7693) <= a and not b;
    layer5_outputs(7694) <= b;
    layer5_outputs(7695) <= b and not a;
    layer5_outputs(7696) <= not b;
    layer5_outputs(7697) <= not a or b;
    layer5_outputs(7698) <= a or b;
    layer5_outputs(7699) <= b;
    layer5_outputs(7700) <= '0';
    layer5_outputs(7701) <= not a;
    layer5_outputs(7702) <= not (a xor b);
    layer5_outputs(7703) <= a or b;
    layer5_outputs(7704) <= not (a and b);
    layer5_outputs(7705) <= b and not a;
    layer5_outputs(7706) <= not a or b;
    layer5_outputs(7707) <= a;
    layer5_outputs(7708) <= b;
    layer5_outputs(7709) <= b and not a;
    layer5_outputs(7710) <= a;
    layer5_outputs(7711) <= a and not b;
    layer5_outputs(7712) <= a or b;
    layer5_outputs(7713) <= not b;
    layer5_outputs(7714) <= a or b;
    layer5_outputs(7715) <= b;
    layer5_outputs(7716) <= not a;
    layer5_outputs(7717) <= not b;
    layer5_outputs(7718) <= a;
    layer5_outputs(7719) <= a;
    layer5_outputs(7720) <= not (a xor b);
    layer5_outputs(7721) <= a or b;
    layer5_outputs(7722) <= '0';
    layer5_outputs(7723) <= a;
    layer5_outputs(7724) <= a xor b;
    layer5_outputs(7725) <= not b;
    layer5_outputs(7726) <= not (a or b);
    layer5_outputs(7727) <= a or b;
    layer5_outputs(7728) <= not a;
    layer5_outputs(7729) <= a;
    layer5_outputs(7730) <= not a;
    layer5_outputs(7731) <= a;
    layer5_outputs(7732) <= b;
    layer5_outputs(7733) <= a;
    layer5_outputs(7734) <= a and not b;
    layer5_outputs(7735) <= a and b;
    layer5_outputs(7736) <= not (a and b);
    layer5_outputs(7737) <= not b;
    layer5_outputs(7738) <= not a;
    layer5_outputs(7739) <= a and b;
    layer5_outputs(7740) <= not b;
    layer5_outputs(7741) <= a and not b;
    layer5_outputs(7742) <= b;
    layer5_outputs(7743) <= not a;
    layer5_outputs(7744) <= b;
    layer5_outputs(7745) <= b;
    layer5_outputs(7746) <= a and not b;
    layer5_outputs(7747) <= not b;
    layer5_outputs(7748) <= not b;
    layer5_outputs(7749) <= a;
    layer5_outputs(7750) <= not b or a;
    layer5_outputs(7751) <= a;
    layer5_outputs(7752) <= not b;
    layer5_outputs(7753) <= a;
    layer5_outputs(7754) <= a;
    layer5_outputs(7755) <= b;
    layer5_outputs(7756) <= a xor b;
    layer5_outputs(7757) <= '1';
    layer5_outputs(7758) <= a and not b;
    layer5_outputs(7759) <= b;
    layer5_outputs(7760) <= not (a or b);
    layer5_outputs(7761) <= a xor b;
    layer5_outputs(7762) <= b;
    layer5_outputs(7763) <= b and not a;
    layer5_outputs(7764) <= b and not a;
    layer5_outputs(7765) <= not a;
    layer5_outputs(7766) <= '1';
    layer5_outputs(7767) <= not a or b;
    layer5_outputs(7768) <= not b;
    layer5_outputs(7769) <= b;
    layer5_outputs(7770) <= not b;
    layer5_outputs(7771) <= not a;
    layer5_outputs(7772) <= not b;
    layer5_outputs(7773) <= '0';
    layer5_outputs(7774) <= not (a or b);
    layer5_outputs(7775) <= not a or b;
    layer5_outputs(7776) <= b and not a;
    layer5_outputs(7777) <= b and not a;
    layer5_outputs(7778) <= b;
    layer5_outputs(7779) <= a and b;
    layer5_outputs(7780) <= a or b;
    layer5_outputs(7781) <= not b;
    layer5_outputs(7782) <= a xor b;
    layer5_outputs(7783) <= not a;
    layer5_outputs(7784) <= '1';
    layer5_outputs(7785) <= not (a xor b);
    layer5_outputs(7786) <= not a;
    layer5_outputs(7787) <= a and not b;
    layer5_outputs(7788) <= b;
    layer5_outputs(7789) <= not (a xor b);
    layer5_outputs(7790) <= not a;
    layer5_outputs(7791) <= not a;
    layer5_outputs(7792) <= not (a or b);
    layer5_outputs(7793) <= not (a and b);
    layer5_outputs(7794) <= not a;
    layer5_outputs(7795) <= a;
    layer5_outputs(7796) <= a;
    layer5_outputs(7797) <= not a;
    layer5_outputs(7798) <= not b;
    layer5_outputs(7799) <= not a;
    layer5_outputs(7800) <= a;
    layer5_outputs(7801) <= not (a and b);
    layer5_outputs(7802) <= not a;
    layer5_outputs(7803) <= not a;
    layer5_outputs(7804) <= b;
    layer5_outputs(7805) <= a;
    layer5_outputs(7806) <= b and not a;
    layer5_outputs(7807) <= not a;
    layer5_outputs(7808) <= b;
    layer5_outputs(7809) <= b and not a;
    layer5_outputs(7810) <= not a;
    layer5_outputs(7811) <= a and b;
    layer5_outputs(7812) <= a;
    layer5_outputs(7813) <= not (a or b);
    layer5_outputs(7814) <= b;
    layer5_outputs(7815) <= not (a and b);
    layer5_outputs(7816) <= not a;
    layer5_outputs(7817) <= b;
    layer5_outputs(7818) <= a xor b;
    layer5_outputs(7819) <= '0';
    layer5_outputs(7820) <= a;
    layer5_outputs(7821) <= not (a xor b);
    layer5_outputs(7822) <= not b or a;
    layer5_outputs(7823) <= b;
    layer5_outputs(7824) <= a;
    layer5_outputs(7825) <= not a;
    layer5_outputs(7826) <= not (a or b);
    layer5_outputs(7827) <= b;
    layer5_outputs(7828) <= a and b;
    layer5_outputs(7829) <= a and not b;
    layer5_outputs(7830) <= b and not a;
    layer5_outputs(7831) <= a or b;
    layer5_outputs(7832) <= a or b;
    layer5_outputs(7833) <= b and not a;
    layer5_outputs(7834) <= '0';
    layer5_outputs(7835) <= not a;
    layer5_outputs(7836) <= b and not a;
    layer5_outputs(7837) <= not (a or b);
    layer5_outputs(7838) <= a;
    layer5_outputs(7839) <= not b or a;
    layer5_outputs(7840) <= not (a and b);
    layer5_outputs(7841) <= not a;
    layer5_outputs(7842) <= not (a or b);
    layer5_outputs(7843) <= a or b;
    layer5_outputs(7844) <= b;
    layer5_outputs(7845) <= not (a xor b);
    layer5_outputs(7846) <= not (a or b);
    layer5_outputs(7847) <= b and not a;
    layer5_outputs(7848) <= not b;
    layer5_outputs(7849) <= a;
    layer5_outputs(7850) <= not a;
    layer5_outputs(7851) <= a and b;
    layer5_outputs(7852) <= b;
    layer5_outputs(7853) <= not a;
    layer5_outputs(7854) <= not a;
    layer5_outputs(7855) <= not a;
    layer5_outputs(7856) <= '0';
    layer5_outputs(7857) <= not b;
    layer5_outputs(7858) <= a xor b;
    layer5_outputs(7859) <= not (a or b);
    layer5_outputs(7860) <= not b or a;
    layer5_outputs(7861) <= a and not b;
    layer5_outputs(7862) <= not b;
    layer5_outputs(7863) <= a xor b;
    layer5_outputs(7864) <= not b;
    layer5_outputs(7865) <= not (a and b);
    layer5_outputs(7866) <= not b;
    layer5_outputs(7867) <= a;
    layer5_outputs(7868) <= not (a and b);
    layer5_outputs(7869) <= not a;
    layer5_outputs(7870) <= not b;
    layer5_outputs(7871) <= b;
    layer5_outputs(7872) <= not b;
    layer5_outputs(7873) <= '1';
    layer5_outputs(7874) <= a or b;
    layer5_outputs(7875) <= a and b;
    layer5_outputs(7876) <= not b or a;
    layer5_outputs(7877) <= a;
    layer5_outputs(7878) <= not b;
    layer5_outputs(7879) <= not b;
    layer5_outputs(7880) <= a and not b;
    layer5_outputs(7881) <= not (a and b);
    layer5_outputs(7882) <= b and not a;
    layer5_outputs(7883) <= b and not a;
    layer5_outputs(7884) <= not b;
    layer5_outputs(7885) <= not (a and b);
    layer5_outputs(7886) <= a and b;
    layer5_outputs(7887) <= not a;
    layer5_outputs(7888) <= not b or a;
    layer5_outputs(7889) <= not a or b;
    layer5_outputs(7890) <= a xor b;
    layer5_outputs(7891) <= not a;
    layer5_outputs(7892) <= b;
    layer5_outputs(7893) <= not b;
    layer5_outputs(7894) <= not b;
    layer5_outputs(7895) <= b;
    layer5_outputs(7896) <= not (a or b);
    layer5_outputs(7897) <= a xor b;
    layer5_outputs(7898) <= a xor b;
    layer5_outputs(7899) <= not a;
    layer5_outputs(7900) <= not a;
    layer5_outputs(7901) <= not a;
    layer5_outputs(7902) <= not a;
    layer5_outputs(7903) <= not (a and b);
    layer5_outputs(7904) <= not a;
    layer5_outputs(7905) <= a xor b;
    layer5_outputs(7906) <= not b or a;
    layer5_outputs(7907) <= b;
    layer5_outputs(7908) <= not b;
    layer5_outputs(7909) <= not (a or b);
    layer5_outputs(7910) <= not (a or b);
    layer5_outputs(7911) <= not a;
    layer5_outputs(7912) <= b;
    layer5_outputs(7913) <= not (a and b);
    layer5_outputs(7914) <= not b;
    layer5_outputs(7915) <= not b;
    layer5_outputs(7916) <= '0';
    layer5_outputs(7917) <= '1';
    layer5_outputs(7918) <= not b;
    layer5_outputs(7919) <= not b;
    layer5_outputs(7920) <= a and b;
    layer5_outputs(7921) <= not a;
    layer5_outputs(7922) <= a and b;
    layer5_outputs(7923) <= a and not b;
    layer5_outputs(7924) <= not (a xor b);
    layer5_outputs(7925) <= not a;
    layer5_outputs(7926) <= '1';
    layer5_outputs(7927) <= not b;
    layer5_outputs(7928) <= a;
    layer5_outputs(7929) <= not b;
    layer5_outputs(7930) <= b and not a;
    layer5_outputs(7931) <= not b or a;
    layer5_outputs(7932) <= not (a or b);
    layer5_outputs(7933) <= not b;
    layer5_outputs(7934) <= b;
    layer5_outputs(7935) <= not b or a;
    layer5_outputs(7936) <= not b;
    layer5_outputs(7937) <= not a;
    layer5_outputs(7938) <= not b or a;
    layer5_outputs(7939) <= not b or a;
    layer5_outputs(7940) <= not (a and b);
    layer5_outputs(7941) <= not (a or b);
    layer5_outputs(7942) <= not (a or b);
    layer5_outputs(7943) <= b and not a;
    layer5_outputs(7944) <= not b;
    layer5_outputs(7945) <= a and not b;
    layer5_outputs(7946) <= not a;
    layer5_outputs(7947) <= a and b;
    layer5_outputs(7948) <= a or b;
    layer5_outputs(7949) <= not (a xor b);
    layer5_outputs(7950) <= a and not b;
    layer5_outputs(7951) <= a xor b;
    layer5_outputs(7952) <= not b;
    layer5_outputs(7953) <= not (a and b);
    layer5_outputs(7954) <= not (a xor b);
    layer5_outputs(7955) <= not (a and b);
    layer5_outputs(7956) <= a;
    layer5_outputs(7957) <= not a or b;
    layer5_outputs(7958) <= a xor b;
    layer5_outputs(7959) <= not (a or b);
    layer5_outputs(7960) <= not a or b;
    layer5_outputs(7961) <= not (a and b);
    layer5_outputs(7962) <= b and not a;
    layer5_outputs(7963) <= not a;
    layer5_outputs(7964) <= not a;
    layer5_outputs(7965) <= a and b;
    layer5_outputs(7966) <= '1';
    layer5_outputs(7967) <= a xor b;
    layer5_outputs(7968) <= b;
    layer5_outputs(7969) <= a;
    layer5_outputs(7970) <= a and b;
    layer5_outputs(7971) <= not (a or b);
    layer5_outputs(7972) <= a;
    layer5_outputs(7973) <= not b;
    layer5_outputs(7974) <= not a or b;
    layer5_outputs(7975) <= b;
    layer5_outputs(7976) <= b;
    layer5_outputs(7977) <= not (a xor b);
    layer5_outputs(7978) <= not a or b;
    layer5_outputs(7979) <= not b;
    layer5_outputs(7980) <= b;
    layer5_outputs(7981) <= a;
    layer5_outputs(7982) <= a;
    layer5_outputs(7983) <= not (a or b);
    layer5_outputs(7984) <= a or b;
    layer5_outputs(7985) <= a xor b;
    layer5_outputs(7986) <= a;
    layer5_outputs(7987) <= a and b;
    layer5_outputs(7988) <= a xor b;
    layer5_outputs(7989) <= not a;
    layer5_outputs(7990) <= not b or a;
    layer5_outputs(7991) <= not (a xor b);
    layer5_outputs(7992) <= a or b;
    layer5_outputs(7993) <= not b or a;
    layer5_outputs(7994) <= not b;
    layer5_outputs(7995) <= not a;
    layer5_outputs(7996) <= not a;
    layer5_outputs(7997) <= a;
    layer5_outputs(7998) <= not a;
    layer5_outputs(7999) <= not b;
    layer5_outputs(8000) <= not a;
    layer5_outputs(8001) <= not (a or b);
    layer5_outputs(8002) <= b and not a;
    layer5_outputs(8003) <= a or b;
    layer5_outputs(8004) <= not a;
    layer5_outputs(8005) <= b and not a;
    layer5_outputs(8006) <= a;
    layer5_outputs(8007) <= not (a xor b);
    layer5_outputs(8008) <= not b or a;
    layer5_outputs(8009) <= not b;
    layer5_outputs(8010) <= b and not a;
    layer5_outputs(8011) <= a;
    layer5_outputs(8012) <= a xor b;
    layer5_outputs(8013) <= not a;
    layer5_outputs(8014) <= b;
    layer5_outputs(8015) <= not (a or b);
    layer5_outputs(8016) <= b and not a;
    layer5_outputs(8017) <= not a or b;
    layer5_outputs(8018) <= a xor b;
    layer5_outputs(8019) <= not a;
    layer5_outputs(8020) <= b;
    layer5_outputs(8021) <= not b;
    layer5_outputs(8022) <= not (a xor b);
    layer5_outputs(8023) <= a and not b;
    layer5_outputs(8024) <= a and not b;
    layer5_outputs(8025) <= not (a xor b);
    layer5_outputs(8026) <= a;
    layer5_outputs(8027) <= not b;
    layer5_outputs(8028) <= a;
    layer5_outputs(8029) <= not (a and b);
    layer5_outputs(8030) <= not a;
    layer5_outputs(8031) <= a;
    layer5_outputs(8032) <= not (a and b);
    layer5_outputs(8033) <= not b or a;
    layer5_outputs(8034) <= not b;
    layer5_outputs(8035) <= not (a or b);
    layer5_outputs(8036) <= not b;
    layer5_outputs(8037) <= b;
    layer5_outputs(8038) <= a xor b;
    layer5_outputs(8039) <= not (a xor b);
    layer5_outputs(8040) <= not (a or b);
    layer5_outputs(8041) <= not (a xor b);
    layer5_outputs(8042) <= a;
    layer5_outputs(8043) <= not b or a;
    layer5_outputs(8044) <= not (a and b);
    layer5_outputs(8045) <= a or b;
    layer5_outputs(8046) <= not a;
    layer5_outputs(8047) <= not b or a;
    layer5_outputs(8048) <= b;
    layer5_outputs(8049) <= not b or a;
    layer5_outputs(8050) <= not b;
    layer5_outputs(8051) <= not b;
    layer5_outputs(8052) <= not b or a;
    layer5_outputs(8053) <= b and not a;
    layer5_outputs(8054) <= a or b;
    layer5_outputs(8055) <= a;
    layer5_outputs(8056) <= not a;
    layer5_outputs(8057) <= a xor b;
    layer5_outputs(8058) <= b and not a;
    layer5_outputs(8059) <= a;
    layer5_outputs(8060) <= not a;
    layer5_outputs(8061) <= b;
    layer5_outputs(8062) <= not a or b;
    layer5_outputs(8063) <= a;
    layer5_outputs(8064) <= a and not b;
    layer5_outputs(8065) <= b;
    layer5_outputs(8066) <= not b or a;
    layer5_outputs(8067) <= a and not b;
    layer5_outputs(8068) <= a;
    layer5_outputs(8069) <= not a or b;
    layer5_outputs(8070) <= not (a or b);
    layer5_outputs(8071) <= a xor b;
    layer5_outputs(8072) <= b and not a;
    layer5_outputs(8073) <= not b;
    layer5_outputs(8074) <= not b or a;
    layer5_outputs(8075) <= not a;
    layer5_outputs(8076) <= a and b;
    layer5_outputs(8077) <= a and b;
    layer5_outputs(8078) <= not (a xor b);
    layer5_outputs(8079) <= not b;
    layer5_outputs(8080) <= not (a and b);
    layer5_outputs(8081) <= not b;
    layer5_outputs(8082) <= b;
    layer5_outputs(8083) <= not (a xor b);
    layer5_outputs(8084) <= not b;
    layer5_outputs(8085) <= not a or b;
    layer5_outputs(8086) <= a xor b;
    layer5_outputs(8087) <= not a or b;
    layer5_outputs(8088) <= a;
    layer5_outputs(8089) <= not (a and b);
    layer5_outputs(8090) <= a xor b;
    layer5_outputs(8091) <= b;
    layer5_outputs(8092) <= a xor b;
    layer5_outputs(8093) <= b and not a;
    layer5_outputs(8094) <= a or b;
    layer5_outputs(8095) <= b;
    layer5_outputs(8096) <= a;
    layer5_outputs(8097) <= a and not b;
    layer5_outputs(8098) <= not a;
    layer5_outputs(8099) <= a and not b;
    layer5_outputs(8100) <= not b;
    layer5_outputs(8101) <= not b;
    layer5_outputs(8102) <= not (a and b);
    layer5_outputs(8103) <= b;
    layer5_outputs(8104) <= b;
    layer5_outputs(8105) <= a;
    layer5_outputs(8106) <= not a or b;
    layer5_outputs(8107) <= a;
    layer5_outputs(8108) <= not a;
    layer5_outputs(8109) <= '1';
    layer5_outputs(8110) <= not a;
    layer5_outputs(8111) <= a and not b;
    layer5_outputs(8112) <= a;
    layer5_outputs(8113) <= not (a xor b);
    layer5_outputs(8114) <= a and not b;
    layer5_outputs(8115) <= a;
    layer5_outputs(8116) <= a;
    layer5_outputs(8117) <= a;
    layer5_outputs(8118) <= a;
    layer5_outputs(8119) <= not (a and b);
    layer5_outputs(8120) <= not (a or b);
    layer5_outputs(8121) <= not b;
    layer5_outputs(8122) <= b;
    layer5_outputs(8123) <= a and b;
    layer5_outputs(8124) <= a;
    layer5_outputs(8125) <= not (a xor b);
    layer5_outputs(8126) <= not a;
    layer5_outputs(8127) <= b and not a;
    layer5_outputs(8128) <= a;
    layer5_outputs(8129) <= a or b;
    layer5_outputs(8130) <= '1';
    layer5_outputs(8131) <= a;
    layer5_outputs(8132) <= a;
    layer5_outputs(8133) <= b and not a;
    layer5_outputs(8134) <= b and not a;
    layer5_outputs(8135) <= not (a or b);
    layer5_outputs(8136) <= not b;
    layer5_outputs(8137) <= not a;
    layer5_outputs(8138) <= '1';
    layer5_outputs(8139) <= a;
    layer5_outputs(8140) <= a;
    layer5_outputs(8141) <= a and not b;
    layer5_outputs(8142) <= not a;
    layer5_outputs(8143) <= not b;
    layer5_outputs(8144) <= b;
    layer5_outputs(8145) <= not (a and b);
    layer5_outputs(8146) <= not b;
    layer5_outputs(8147) <= not a;
    layer5_outputs(8148) <= not b or a;
    layer5_outputs(8149) <= b and not a;
    layer5_outputs(8150) <= a;
    layer5_outputs(8151) <= a or b;
    layer5_outputs(8152) <= not (a and b);
    layer5_outputs(8153) <= not b;
    layer5_outputs(8154) <= not b or a;
    layer5_outputs(8155) <= not a;
    layer5_outputs(8156) <= a and b;
    layer5_outputs(8157) <= b;
    layer5_outputs(8158) <= not (a and b);
    layer5_outputs(8159) <= a;
    layer5_outputs(8160) <= not a;
    layer5_outputs(8161) <= b and not a;
    layer5_outputs(8162) <= a xor b;
    layer5_outputs(8163) <= a;
    layer5_outputs(8164) <= a;
    layer5_outputs(8165) <= not a or b;
    layer5_outputs(8166) <= not (a or b);
    layer5_outputs(8167) <= not b;
    layer5_outputs(8168) <= b and not a;
    layer5_outputs(8169) <= not (a or b);
    layer5_outputs(8170) <= not (a or b);
    layer5_outputs(8171) <= a;
    layer5_outputs(8172) <= not a or b;
    layer5_outputs(8173) <= not (a xor b);
    layer5_outputs(8174) <= b;
    layer5_outputs(8175) <= not b;
    layer5_outputs(8176) <= a and not b;
    layer5_outputs(8177) <= b and not a;
    layer5_outputs(8178) <= a;
    layer5_outputs(8179) <= a;
    layer5_outputs(8180) <= not (a or b);
    layer5_outputs(8181) <= a and b;
    layer5_outputs(8182) <= not a or b;
    layer5_outputs(8183) <= a;
    layer5_outputs(8184) <= a;
    layer5_outputs(8185) <= a and b;
    layer5_outputs(8186) <= a;
    layer5_outputs(8187) <= a and not b;
    layer5_outputs(8188) <= b;
    layer5_outputs(8189) <= a;
    layer5_outputs(8190) <= a and b;
    layer5_outputs(8191) <= not a;
    layer5_outputs(8192) <= '1';
    layer5_outputs(8193) <= a and b;
    layer5_outputs(8194) <= a;
    layer5_outputs(8195) <= a and b;
    layer5_outputs(8196) <= not b or a;
    layer5_outputs(8197) <= not b or a;
    layer5_outputs(8198) <= a and b;
    layer5_outputs(8199) <= not (a and b);
    layer5_outputs(8200) <= not (a or b);
    layer5_outputs(8201) <= a;
    layer5_outputs(8202) <= a and b;
    layer5_outputs(8203) <= not a;
    layer5_outputs(8204) <= not (a or b);
    layer5_outputs(8205) <= not a or b;
    layer5_outputs(8206) <= a;
    layer5_outputs(8207) <= b;
    layer5_outputs(8208) <= a and not b;
    layer5_outputs(8209) <= not a;
    layer5_outputs(8210) <= a xor b;
    layer5_outputs(8211) <= not a or b;
    layer5_outputs(8212) <= b and not a;
    layer5_outputs(8213) <= b and not a;
    layer5_outputs(8214) <= a;
    layer5_outputs(8215) <= not b;
    layer5_outputs(8216) <= not b;
    layer5_outputs(8217) <= not b;
    layer5_outputs(8218) <= a xor b;
    layer5_outputs(8219) <= a or b;
    layer5_outputs(8220) <= a;
    layer5_outputs(8221) <= b;
    layer5_outputs(8222) <= not b;
    layer5_outputs(8223) <= a and not b;
    layer5_outputs(8224) <= not (a xor b);
    layer5_outputs(8225) <= not (a and b);
    layer5_outputs(8226) <= a xor b;
    layer5_outputs(8227) <= b and not a;
    layer5_outputs(8228) <= a and b;
    layer5_outputs(8229) <= b;
    layer5_outputs(8230) <= not a;
    layer5_outputs(8231) <= a;
    layer5_outputs(8232) <= not (a xor b);
    layer5_outputs(8233) <= a xor b;
    layer5_outputs(8234) <= a xor b;
    layer5_outputs(8235) <= not b;
    layer5_outputs(8236) <= a and b;
    layer5_outputs(8237) <= not b;
    layer5_outputs(8238) <= not (a xor b);
    layer5_outputs(8239) <= not a;
    layer5_outputs(8240) <= a or b;
    layer5_outputs(8241) <= not a or b;
    layer5_outputs(8242) <= not a;
    layer5_outputs(8243) <= a;
    layer5_outputs(8244) <= not (a or b);
    layer5_outputs(8245) <= '0';
    layer5_outputs(8246) <= not a or b;
    layer5_outputs(8247) <= not b;
    layer5_outputs(8248) <= not (a xor b);
    layer5_outputs(8249) <= a;
    layer5_outputs(8250) <= not (a or b);
    layer5_outputs(8251) <= not a;
    layer5_outputs(8252) <= not b or a;
    layer5_outputs(8253) <= not a;
    layer5_outputs(8254) <= a xor b;
    layer5_outputs(8255) <= a or b;
    layer5_outputs(8256) <= not a or b;
    layer5_outputs(8257) <= a and not b;
    layer5_outputs(8258) <= a and not b;
    layer5_outputs(8259) <= b;
    layer5_outputs(8260) <= a;
    layer5_outputs(8261) <= a or b;
    layer5_outputs(8262) <= b;
    layer5_outputs(8263) <= a xor b;
    layer5_outputs(8264) <= not (a or b);
    layer5_outputs(8265) <= a or b;
    layer5_outputs(8266) <= not b or a;
    layer5_outputs(8267) <= b;
    layer5_outputs(8268) <= not a;
    layer5_outputs(8269) <= a or b;
    layer5_outputs(8270) <= not (a and b);
    layer5_outputs(8271) <= a xor b;
    layer5_outputs(8272) <= a xor b;
    layer5_outputs(8273) <= a;
    layer5_outputs(8274) <= not a;
    layer5_outputs(8275) <= a and b;
    layer5_outputs(8276) <= a xor b;
    layer5_outputs(8277) <= not a;
    layer5_outputs(8278) <= a and not b;
    layer5_outputs(8279) <= a and not b;
    layer5_outputs(8280) <= a or b;
    layer5_outputs(8281) <= not b or a;
    layer5_outputs(8282) <= not a;
    layer5_outputs(8283) <= a or b;
    layer5_outputs(8284) <= a xor b;
    layer5_outputs(8285) <= a;
    layer5_outputs(8286) <= b;
    layer5_outputs(8287) <= not b or a;
    layer5_outputs(8288) <= not (a and b);
    layer5_outputs(8289) <= not (a or b);
    layer5_outputs(8290) <= not (a or b);
    layer5_outputs(8291) <= not a;
    layer5_outputs(8292) <= b;
    layer5_outputs(8293) <= not b;
    layer5_outputs(8294) <= not (a and b);
    layer5_outputs(8295) <= '0';
    layer5_outputs(8296) <= b;
    layer5_outputs(8297) <= not b;
    layer5_outputs(8298) <= b;
    layer5_outputs(8299) <= not a;
    layer5_outputs(8300) <= a;
    layer5_outputs(8301) <= not a;
    layer5_outputs(8302) <= a xor b;
    layer5_outputs(8303) <= a xor b;
    layer5_outputs(8304) <= not b or a;
    layer5_outputs(8305) <= not (a or b);
    layer5_outputs(8306) <= a;
    layer5_outputs(8307) <= not b;
    layer5_outputs(8308) <= not (a xor b);
    layer5_outputs(8309) <= not (a or b);
    layer5_outputs(8310) <= not a or b;
    layer5_outputs(8311) <= a;
    layer5_outputs(8312) <= not a or b;
    layer5_outputs(8313) <= b;
    layer5_outputs(8314) <= not a;
    layer5_outputs(8315) <= '0';
    layer5_outputs(8316) <= a and not b;
    layer5_outputs(8317) <= a xor b;
    layer5_outputs(8318) <= not a;
    layer5_outputs(8319) <= a xor b;
    layer5_outputs(8320) <= not (a or b);
    layer5_outputs(8321) <= b;
    layer5_outputs(8322) <= not b;
    layer5_outputs(8323) <= a or b;
    layer5_outputs(8324) <= a xor b;
    layer5_outputs(8325) <= a xor b;
    layer5_outputs(8326) <= b;
    layer5_outputs(8327) <= not b or a;
    layer5_outputs(8328) <= not a;
    layer5_outputs(8329) <= b;
    layer5_outputs(8330) <= not (a xor b);
    layer5_outputs(8331) <= not b or a;
    layer5_outputs(8332) <= a xor b;
    layer5_outputs(8333) <= not a;
    layer5_outputs(8334) <= a or b;
    layer5_outputs(8335) <= not b;
    layer5_outputs(8336) <= a or b;
    layer5_outputs(8337) <= not a or b;
    layer5_outputs(8338) <= not a or b;
    layer5_outputs(8339) <= b;
    layer5_outputs(8340) <= '1';
    layer5_outputs(8341) <= b and not a;
    layer5_outputs(8342) <= b and not a;
    layer5_outputs(8343) <= b and not a;
    layer5_outputs(8344) <= a and b;
    layer5_outputs(8345) <= a and b;
    layer5_outputs(8346) <= a xor b;
    layer5_outputs(8347) <= a and not b;
    layer5_outputs(8348) <= not (a and b);
    layer5_outputs(8349) <= not (a and b);
    layer5_outputs(8350) <= a xor b;
    layer5_outputs(8351) <= b;
    layer5_outputs(8352) <= not (a and b);
    layer5_outputs(8353) <= not (a and b);
    layer5_outputs(8354) <= not b;
    layer5_outputs(8355) <= not (a xor b);
    layer5_outputs(8356) <= not (a and b);
    layer5_outputs(8357) <= b and not a;
    layer5_outputs(8358) <= a xor b;
    layer5_outputs(8359) <= b;
    layer5_outputs(8360) <= a and not b;
    layer5_outputs(8361) <= not (a xor b);
    layer5_outputs(8362) <= b and not a;
    layer5_outputs(8363) <= not (a or b);
    layer5_outputs(8364) <= not a;
    layer5_outputs(8365) <= not (a xor b);
    layer5_outputs(8366) <= b;
    layer5_outputs(8367) <= a;
    layer5_outputs(8368) <= not b;
    layer5_outputs(8369) <= not (a or b);
    layer5_outputs(8370) <= a;
    layer5_outputs(8371) <= not (a and b);
    layer5_outputs(8372) <= not (a and b);
    layer5_outputs(8373) <= b;
    layer5_outputs(8374) <= b;
    layer5_outputs(8375) <= a or b;
    layer5_outputs(8376) <= not (a and b);
    layer5_outputs(8377) <= a xor b;
    layer5_outputs(8378) <= a and b;
    layer5_outputs(8379) <= a;
    layer5_outputs(8380) <= not (a xor b);
    layer5_outputs(8381) <= not (a or b);
    layer5_outputs(8382) <= b;
    layer5_outputs(8383) <= b and not a;
    layer5_outputs(8384) <= a;
    layer5_outputs(8385) <= not b;
    layer5_outputs(8386) <= b and not a;
    layer5_outputs(8387) <= a and b;
    layer5_outputs(8388) <= not (a and b);
    layer5_outputs(8389) <= a;
    layer5_outputs(8390) <= not b;
    layer5_outputs(8391) <= not (a or b);
    layer5_outputs(8392) <= not a;
    layer5_outputs(8393) <= not b;
    layer5_outputs(8394) <= not (a or b);
    layer5_outputs(8395) <= not a;
    layer5_outputs(8396) <= not a;
    layer5_outputs(8397) <= b;
    layer5_outputs(8398) <= not b;
    layer5_outputs(8399) <= b;
    layer5_outputs(8400) <= not a;
    layer5_outputs(8401) <= '1';
    layer5_outputs(8402) <= not a or b;
    layer5_outputs(8403) <= not a;
    layer5_outputs(8404) <= b;
    layer5_outputs(8405) <= not (a xor b);
    layer5_outputs(8406) <= not (a xor b);
    layer5_outputs(8407) <= not b or a;
    layer5_outputs(8408) <= not a;
    layer5_outputs(8409) <= not (a and b);
    layer5_outputs(8410) <= not b;
    layer5_outputs(8411) <= not (a xor b);
    layer5_outputs(8412) <= a or b;
    layer5_outputs(8413) <= '0';
    layer5_outputs(8414) <= b;
    layer5_outputs(8415) <= b;
    layer5_outputs(8416) <= b;
    layer5_outputs(8417) <= b and not a;
    layer5_outputs(8418) <= a;
    layer5_outputs(8419) <= '0';
    layer5_outputs(8420) <= '0';
    layer5_outputs(8421) <= not (a and b);
    layer5_outputs(8422) <= not b;
    layer5_outputs(8423) <= a xor b;
    layer5_outputs(8424) <= b;
    layer5_outputs(8425) <= not (a xor b);
    layer5_outputs(8426) <= not (a xor b);
    layer5_outputs(8427) <= a xor b;
    layer5_outputs(8428) <= b;
    layer5_outputs(8429) <= not b or a;
    layer5_outputs(8430) <= not a;
    layer5_outputs(8431) <= not a;
    layer5_outputs(8432) <= b and not a;
    layer5_outputs(8433) <= b;
    layer5_outputs(8434) <= a and b;
    layer5_outputs(8435) <= b and not a;
    layer5_outputs(8436) <= not b or a;
    layer5_outputs(8437) <= b;
    layer5_outputs(8438) <= '0';
    layer5_outputs(8439) <= a xor b;
    layer5_outputs(8440) <= b and not a;
    layer5_outputs(8441) <= not a or b;
    layer5_outputs(8442) <= a and not b;
    layer5_outputs(8443) <= not b;
    layer5_outputs(8444) <= a and b;
    layer5_outputs(8445) <= not a;
    layer5_outputs(8446) <= b and not a;
    layer5_outputs(8447) <= a xor b;
    layer5_outputs(8448) <= not b;
    layer5_outputs(8449) <= not a or b;
    layer5_outputs(8450) <= not (a or b);
    layer5_outputs(8451) <= not (a or b);
    layer5_outputs(8452) <= not b;
    layer5_outputs(8453) <= not a;
    layer5_outputs(8454) <= not (a xor b);
    layer5_outputs(8455) <= b;
    layer5_outputs(8456) <= b;
    layer5_outputs(8457) <= not b;
    layer5_outputs(8458) <= not b or a;
    layer5_outputs(8459) <= a;
    layer5_outputs(8460) <= not b;
    layer5_outputs(8461) <= b;
    layer5_outputs(8462) <= not b;
    layer5_outputs(8463) <= a and b;
    layer5_outputs(8464) <= a and not b;
    layer5_outputs(8465) <= b;
    layer5_outputs(8466) <= a xor b;
    layer5_outputs(8467) <= a xor b;
    layer5_outputs(8468) <= a and b;
    layer5_outputs(8469) <= b;
    layer5_outputs(8470) <= not a or b;
    layer5_outputs(8471) <= not (a xor b);
    layer5_outputs(8472) <= b;
    layer5_outputs(8473) <= not a;
    layer5_outputs(8474) <= b;
    layer5_outputs(8475) <= b;
    layer5_outputs(8476) <= not (a or b);
    layer5_outputs(8477) <= not (a and b);
    layer5_outputs(8478) <= a;
    layer5_outputs(8479) <= a and b;
    layer5_outputs(8480) <= not (a xor b);
    layer5_outputs(8481) <= not b;
    layer5_outputs(8482) <= not (a and b);
    layer5_outputs(8483) <= not (a and b);
    layer5_outputs(8484) <= b;
    layer5_outputs(8485) <= not (a or b);
    layer5_outputs(8486) <= a;
    layer5_outputs(8487) <= not b or a;
    layer5_outputs(8488) <= b;
    layer5_outputs(8489) <= not b;
    layer5_outputs(8490) <= not a or b;
    layer5_outputs(8491) <= not (a or b);
    layer5_outputs(8492) <= not (a or b);
    layer5_outputs(8493) <= a and b;
    layer5_outputs(8494) <= b;
    layer5_outputs(8495) <= a and b;
    layer5_outputs(8496) <= not (a xor b);
    layer5_outputs(8497) <= not (a xor b);
    layer5_outputs(8498) <= not (a xor b);
    layer5_outputs(8499) <= not (a xor b);
    layer5_outputs(8500) <= not (a xor b);
    layer5_outputs(8501) <= a xor b;
    layer5_outputs(8502) <= not a or b;
    layer5_outputs(8503) <= not (a xor b);
    layer5_outputs(8504) <= not a;
    layer5_outputs(8505) <= not b;
    layer5_outputs(8506) <= b;
    layer5_outputs(8507) <= not (a or b);
    layer5_outputs(8508) <= a or b;
    layer5_outputs(8509) <= a and not b;
    layer5_outputs(8510) <= b;
    layer5_outputs(8511) <= not a or b;
    layer5_outputs(8512) <= not b or a;
    layer5_outputs(8513) <= b;
    layer5_outputs(8514) <= a and b;
    layer5_outputs(8515) <= b;
    layer5_outputs(8516) <= a;
    layer5_outputs(8517) <= a;
    layer5_outputs(8518) <= a;
    layer5_outputs(8519) <= not (a and b);
    layer5_outputs(8520) <= not b or a;
    layer5_outputs(8521) <= not a;
    layer5_outputs(8522) <= not (a or b);
    layer5_outputs(8523) <= not b;
    layer5_outputs(8524) <= not a or b;
    layer5_outputs(8525) <= a or b;
    layer5_outputs(8526) <= b and not a;
    layer5_outputs(8527) <= not (a and b);
    layer5_outputs(8528) <= not (a or b);
    layer5_outputs(8529) <= not b;
    layer5_outputs(8530) <= not b or a;
    layer5_outputs(8531) <= not b;
    layer5_outputs(8532) <= not b;
    layer5_outputs(8533) <= not b;
    layer5_outputs(8534) <= a;
    layer5_outputs(8535) <= a;
    layer5_outputs(8536) <= not (a and b);
    layer5_outputs(8537) <= not (a xor b);
    layer5_outputs(8538) <= a;
    layer5_outputs(8539) <= a and b;
    layer5_outputs(8540) <= b and not a;
    layer5_outputs(8541) <= not a;
    layer5_outputs(8542) <= not b or a;
    layer5_outputs(8543) <= not a or b;
    layer5_outputs(8544) <= not (a or b);
    layer5_outputs(8545) <= a and not b;
    layer5_outputs(8546) <= a;
    layer5_outputs(8547) <= '1';
    layer5_outputs(8548) <= a;
    layer5_outputs(8549) <= b and not a;
    layer5_outputs(8550) <= not a;
    layer5_outputs(8551) <= not a;
    layer5_outputs(8552) <= not b;
    layer5_outputs(8553) <= not (a xor b);
    layer5_outputs(8554) <= not b;
    layer5_outputs(8555) <= b;
    layer5_outputs(8556) <= not (a and b);
    layer5_outputs(8557) <= not (a and b);
    layer5_outputs(8558) <= not (a and b);
    layer5_outputs(8559) <= not (a and b);
    layer5_outputs(8560) <= a xor b;
    layer5_outputs(8561) <= a xor b;
    layer5_outputs(8562) <= a or b;
    layer5_outputs(8563) <= not (a or b);
    layer5_outputs(8564) <= not a;
    layer5_outputs(8565) <= b;
    layer5_outputs(8566) <= not a or b;
    layer5_outputs(8567) <= not a;
    layer5_outputs(8568) <= not a;
    layer5_outputs(8569) <= a;
    layer5_outputs(8570) <= a;
    layer5_outputs(8571) <= b;
    layer5_outputs(8572) <= not b;
    layer5_outputs(8573) <= a and b;
    layer5_outputs(8574) <= not (a and b);
    layer5_outputs(8575) <= not (a and b);
    layer5_outputs(8576) <= not a or b;
    layer5_outputs(8577) <= not a;
    layer5_outputs(8578) <= '1';
    layer5_outputs(8579) <= a;
    layer5_outputs(8580) <= not b or a;
    layer5_outputs(8581) <= not b or a;
    layer5_outputs(8582) <= not a;
    layer5_outputs(8583) <= a;
    layer5_outputs(8584) <= not (a and b);
    layer5_outputs(8585) <= a or b;
    layer5_outputs(8586) <= a;
    layer5_outputs(8587) <= a and b;
    layer5_outputs(8588) <= a;
    layer5_outputs(8589) <= b and not a;
    layer5_outputs(8590) <= a or b;
    layer5_outputs(8591) <= not b;
    layer5_outputs(8592) <= a;
    layer5_outputs(8593) <= not a;
    layer5_outputs(8594) <= a;
    layer5_outputs(8595) <= not b;
    layer5_outputs(8596) <= not b;
    layer5_outputs(8597) <= not (a and b);
    layer5_outputs(8598) <= a;
    layer5_outputs(8599) <= not (a xor b);
    layer5_outputs(8600) <= '0';
    layer5_outputs(8601) <= not (a or b);
    layer5_outputs(8602) <= a and b;
    layer5_outputs(8603) <= a;
    layer5_outputs(8604) <= b and not a;
    layer5_outputs(8605) <= b;
    layer5_outputs(8606) <= a;
    layer5_outputs(8607) <= a and not b;
    layer5_outputs(8608) <= not (a xor b);
    layer5_outputs(8609) <= not a or b;
    layer5_outputs(8610) <= not (a xor b);
    layer5_outputs(8611) <= a xor b;
    layer5_outputs(8612) <= not b;
    layer5_outputs(8613) <= a or b;
    layer5_outputs(8614) <= b and not a;
    layer5_outputs(8615) <= a or b;
    layer5_outputs(8616) <= a xor b;
    layer5_outputs(8617) <= b and not a;
    layer5_outputs(8618) <= b and not a;
    layer5_outputs(8619) <= not (a and b);
    layer5_outputs(8620) <= not (a and b);
    layer5_outputs(8621) <= b;
    layer5_outputs(8622) <= not b;
    layer5_outputs(8623) <= b;
    layer5_outputs(8624) <= not (a or b);
    layer5_outputs(8625) <= not a;
    layer5_outputs(8626) <= a;
    layer5_outputs(8627) <= b and not a;
    layer5_outputs(8628) <= b;
    layer5_outputs(8629) <= not (a or b);
    layer5_outputs(8630) <= not a;
    layer5_outputs(8631) <= not (a and b);
    layer5_outputs(8632) <= b;
    layer5_outputs(8633) <= not b;
    layer5_outputs(8634) <= not a;
    layer5_outputs(8635) <= not b;
    layer5_outputs(8636) <= b;
    layer5_outputs(8637) <= a;
    layer5_outputs(8638) <= not a;
    layer5_outputs(8639) <= a;
    layer5_outputs(8640) <= not (a and b);
    layer5_outputs(8641) <= not b;
    layer5_outputs(8642) <= a and not b;
    layer5_outputs(8643) <= a;
    layer5_outputs(8644) <= a;
    layer5_outputs(8645) <= a or b;
    layer5_outputs(8646) <= b;
    layer5_outputs(8647) <= b;
    layer5_outputs(8648) <= a and not b;
    layer5_outputs(8649) <= a or b;
    layer5_outputs(8650) <= b and not a;
    layer5_outputs(8651) <= b and not a;
    layer5_outputs(8652) <= b;
    layer5_outputs(8653) <= not a or b;
    layer5_outputs(8654) <= not a;
    layer5_outputs(8655) <= a xor b;
    layer5_outputs(8656) <= not (a or b);
    layer5_outputs(8657) <= not a;
    layer5_outputs(8658) <= a;
    layer5_outputs(8659) <= not a;
    layer5_outputs(8660) <= not (a xor b);
    layer5_outputs(8661) <= not (a xor b);
    layer5_outputs(8662) <= a and b;
    layer5_outputs(8663) <= '1';
    layer5_outputs(8664) <= a;
    layer5_outputs(8665) <= not a or b;
    layer5_outputs(8666) <= not b;
    layer5_outputs(8667) <= a;
    layer5_outputs(8668) <= a and not b;
    layer5_outputs(8669) <= a;
    layer5_outputs(8670) <= not b;
    layer5_outputs(8671) <= not (a xor b);
    layer5_outputs(8672) <= not (a or b);
    layer5_outputs(8673) <= a or b;
    layer5_outputs(8674) <= not (a and b);
    layer5_outputs(8675) <= not a;
    layer5_outputs(8676) <= b and not a;
    layer5_outputs(8677) <= not b;
    layer5_outputs(8678) <= b;
    layer5_outputs(8679) <= b;
    layer5_outputs(8680) <= a and not b;
    layer5_outputs(8681) <= a;
    layer5_outputs(8682) <= a xor b;
    layer5_outputs(8683) <= a or b;
    layer5_outputs(8684) <= a and not b;
    layer5_outputs(8685) <= a;
    layer5_outputs(8686) <= not b;
    layer5_outputs(8687) <= b;
    layer5_outputs(8688) <= not (a or b);
    layer5_outputs(8689) <= b;
    layer5_outputs(8690) <= b and not a;
    layer5_outputs(8691) <= not b;
    layer5_outputs(8692) <= not (a and b);
    layer5_outputs(8693) <= a or b;
    layer5_outputs(8694) <= a and b;
    layer5_outputs(8695) <= a;
    layer5_outputs(8696) <= a or b;
    layer5_outputs(8697) <= not a;
    layer5_outputs(8698) <= not b or a;
    layer5_outputs(8699) <= a and not b;
    layer5_outputs(8700) <= a;
    layer5_outputs(8701) <= not b;
    layer5_outputs(8702) <= not a or b;
    layer5_outputs(8703) <= not b;
    layer5_outputs(8704) <= '1';
    layer5_outputs(8705) <= not (a or b);
    layer5_outputs(8706) <= not a;
    layer5_outputs(8707) <= b;
    layer5_outputs(8708) <= not b or a;
    layer5_outputs(8709) <= not a or b;
    layer5_outputs(8710) <= a;
    layer5_outputs(8711) <= a or b;
    layer5_outputs(8712) <= b;
    layer5_outputs(8713) <= not b;
    layer5_outputs(8714) <= not a;
    layer5_outputs(8715) <= not (a xor b);
    layer5_outputs(8716) <= b;
    layer5_outputs(8717) <= a;
    layer5_outputs(8718) <= a and not b;
    layer5_outputs(8719) <= not b;
    layer5_outputs(8720) <= not a;
    layer5_outputs(8721) <= not (a and b);
    layer5_outputs(8722) <= a;
    layer5_outputs(8723) <= a and not b;
    layer5_outputs(8724) <= a or b;
    layer5_outputs(8725) <= not (a and b);
    layer5_outputs(8726) <= a and not b;
    layer5_outputs(8727) <= a;
    layer5_outputs(8728) <= not (a and b);
    layer5_outputs(8729) <= not (a xor b);
    layer5_outputs(8730) <= not (a xor b);
    layer5_outputs(8731) <= b;
    layer5_outputs(8732) <= a xor b;
    layer5_outputs(8733) <= b;
    layer5_outputs(8734) <= a or b;
    layer5_outputs(8735) <= not a;
    layer5_outputs(8736) <= not (a xor b);
    layer5_outputs(8737) <= a;
    layer5_outputs(8738) <= not b;
    layer5_outputs(8739) <= not b or a;
    layer5_outputs(8740) <= not a;
    layer5_outputs(8741) <= b and not a;
    layer5_outputs(8742) <= a and not b;
    layer5_outputs(8743) <= a;
    layer5_outputs(8744) <= a;
    layer5_outputs(8745) <= not (a xor b);
    layer5_outputs(8746) <= not a;
    layer5_outputs(8747) <= not a or b;
    layer5_outputs(8748) <= '1';
    layer5_outputs(8749) <= not (a xor b);
    layer5_outputs(8750) <= a or b;
    layer5_outputs(8751) <= a;
    layer5_outputs(8752) <= b;
    layer5_outputs(8753) <= not a;
    layer5_outputs(8754) <= a or b;
    layer5_outputs(8755) <= b;
    layer5_outputs(8756) <= not b;
    layer5_outputs(8757) <= not a;
    layer5_outputs(8758) <= a;
    layer5_outputs(8759) <= not a;
    layer5_outputs(8760) <= '0';
    layer5_outputs(8761) <= a or b;
    layer5_outputs(8762) <= not a or b;
    layer5_outputs(8763) <= b and not a;
    layer5_outputs(8764) <= b;
    layer5_outputs(8765) <= not (a or b);
    layer5_outputs(8766) <= not b or a;
    layer5_outputs(8767) <= not (a or b);
    layer5_outputs(8768) <= not (a xor b);
    layer5_outputs(8769) <= '0';
    layer5_outputs(8770) <= b;
    layer5_outputs(8771) <= not a or b;
    layer5_outputs(8772) <= a and not b;
    layer5_outputs(8773) <= b;
    layer5_outputs(8774) <= '0';
    layer5_outputs(8775) <= a;
    layer5_outputs(8776) <= a and not b;
    layer5_outputs(8777) <= a and not b;
    layer5_outputs(8778) <= not b or a;
    layer5_outputs(8779) <= not b;
    layer5_outputs(8780) <= a;
    layer5_outputs(8781) <= not a;
    layer5_outputs(8782) <= not b;
    layer5_outputs(8783) <= not (a or b);
    layer5_outputs(8784) <= not (a xor b);
    layer5_outputs(8785) <= a;
    layer5_outputs(8786) <= '0';
    layer5_outputs(8787) <= a xor b;
    layer5_outputs(8788) <= not (a xor b);
    layer5_outputs(8789) <= not b or a;
    layer5_outputs(8790) <= not b;
    layer5_outputs(8791) <= a or b;
    layer5_outputs(8792) <= not a or b;
    layer5_outputs(8793) <= not b or a;
    layer5_outputs(8794) <= b;
    layer5_outputs(8795) <= not b;
    layer5_outputs(8796) <= not b or a;
    layer5_outputs(8797) <= b;
    layer5_outputs(8798) <= a or b;
    layer5_outputs(8799) <= not (a and b);
    layer5_outputs(8800) <= not a;
    layer5_outputs(8801) <= not (a xor b);
    layer5_outputs(8802) <= a and not b;
    layer5_outputs(8803) <= not (a or b);
    layer5_outputs(8804) <= b;
    layer5_outputs(8805) <= not b or a;
    layer5_outputs(8806) <= not b;
    layer5_outputs(8807) <= a or b;
    layer5_outputs(8808) <= not a;
    layer5_outputs(8809) <= not b;
    layer5_outputs(8810) <= not (a or b);
    layer5_outputs(8811) <= not b or a;
    layer5_outputs(8812) <= a and b;
    layer5_outputs(8813) <= a;
    layer5_outputs(8814) <= b;
    layer5_outputs(8815) <= not a or b;
    layer5_outputs(8816) <= b;
    layer5_outputs(8817) <= not (a or b);
    layer5_outputs(8818) <= not b;
    layer5_outputs(8819) <= not b or a;
    layer5_outputs(8820) <= b;
    layer5_outputs(8821) <= b;
    layer5_outputs(8822) <= '0';
    layer5_outputs(8823) <= not (a or b);
    layer5_outputs(8824) <= not (a xor b);
    layer5_outputs(8825) <= not (a xor b);
    layer5_outputs(8826) <= a;
    layer5_outputs(8827) <= not (a xor b);
    layer5_outputs(8828) <= not b or a;
    layer5_outputs(8829) <= not (a xor b);
    layer5_outputs(8830) <= not b;
    layer5_outputs(8831) <= not (a xor b);
    layer5_outputs(8832) <= not (a or b);
    layer5_outputs(8833) <= not a;
    layer5_outputs(8834) <= a;
    layer5_outputs(8835) <= a;
    layer5_outputs(8836) <= not a or b;
    layer5_outputs(8837) <= not a;
    layer5_outputs(8838) <= a and b;
    layer5_outputs(8839) <= a and b;
    layer5_outputs(8840) <= a;
    layer5_outputs(8841) <= a;
    layer5_outputs(8842) <= a xor b;
    layer5_outputs(8843) <= not a or b;
    layer5_outputs(8844) <= not (a xor b);
    layer5_outputs(8845) <= not b;
    layer5_outputs(8846) <= not b;
    layer5_outputs(8847) <= not (a and b);
    layer5_outputs(8848) <= a or b;
    layer5_outputs(8849) <= not b or a;
    layer5_outputs(8850) <= not a or b;
    layer5_outputs(8851) <= not b;
    layer5_outputs(8852) <= a or b;
    layer5_outputs(8853) <= b;
    layer5_outputs(8854) <= not a;
    layer5_outputs(8855) <= a and b;
    layer5_outputs(8856) <= not (a or b);
    layer5_outputs(8857) <= a and not b;
    layer5_outputs(8858) <= a;
    layer5_outputs(8859) <= not b;
    layer5_outputs(8860) <= not a;
    layer5_outputs(8861) <= '1';
    layer5_outputs(8862) <= not (a and b);
    layer5_outputs(8863) <= b;
    layer5_outputs(8864) <= not a;
    layer5_outputs(8865) <= not a or b;
    layer5_outputs(8866) <= b;
    layer5_outputs(8867) <= a;
    layer5_outputs(8868) <= b;
    layer5_outputs(8869) <= '0';
    layer5_outputs(8870) <= not b;
    layer5_outputs(8871) <= b;
    layer5_outputs(8872) <= not b;
    layer5_outputs(8873) <= b and not a;
    layer5_outputs(8874) <= a and b;
    layer5_outputs(8875) <= not a or b;
    layer5_outputs(8876) <= b;
    layer5_outputs(8877) <= not a;
    layer5_outputs(8878) <= a and b;
    layer5_outputs(8879) <= b;
    layer5_outputs(8880) <= not b;
    layer5_outputs(8881) <= not b;
    layer5_outputs(8882) <= a;
    layer5_outputs(8883) <= a and not b;
    layer5_outputs(8884) <= a or b;
    layer5_outputs(8885) <= not a;
    layer5_outputs(8886) <= a;
    layer5_outputs(8887) <= a and not b;
    layer5_outputs(8888) <= '0';
    layer5_outputs(8889) <= a;
    layer5_outputs(8890) <= a or b;
    layer5_outputs(8891) <= not (a xor b);
    layer5_outputs(8892) <= b;
    layer5_outputs(8893) <= not a;
    layer5_outputs(8894) <= a or b;
    layer5_outputs(8895) <= not (a and b);
    layer5_outputs(8896) <= not a;
    layer5_outputs(8897) <= b;
    layer5_outputs(8898) <= b;
    layer5_outputs(8899) <= a;
    layer5_outputs(8900) <= b;
    layer5_outputs(8901) <= a or b;
    layer5_outputs(8902) <= not (a or b);
    layer5_outputs(8903) <= not b;
    layer5_outputs(8904) <= a and b;
    layer5_outputs(8905) <= not a;
    layer5_outputs(8906) <= a and not b;
    layer5_outputs(8907) <= a or b;
    layer5_outputs(8908) <= a;
    layer5_outputs(8909) <= not b or a;
    layer5_outputs(8910) <= a or b;
    layer5_outputs(8911) <= not a or b;
    layer5_outputs(8912) <= not b;
    layer5_outputs(8913) <= a xor b;
    layer5_outputs(8914) <= b;
    layer5_outputs(8915) <= a and b;
    layer5_outputs(8916) <= not a;
    layer5_outputs(8917) <= b and not a;
    layer5_outputs(8918) <= a and b;
    layer5_outputs(8919) <= not (a or b);
    layer5_outputs(8920) <= a or b;
    layer5_outputs(8921) <= b and not a;
    layer5_outputs(8922) <= a and b;
    layer5_outputs(8923) <= not a or b;
    layer5_outputs(8924) <= not (a or b);
    layer5_outputs(8925) <= a;
    layer5_outputs(8926) <= not b or a;
    layer5_outputs(8927) <= '1';
    layer5_outputs(8928) <= b;
    layer5_outputs(8929) <= not a or b;
    layer5_outputs(8930) <= not (a and b);
    layer5_outputs(8931) <= not b or a;
    layer5_outputs(8932) <= not a or b;
    layer5_outputs(8933) <= b;
    layer5_outputs(8934) <= not (a xor b);
    layer5_outputs(8935) <= a;
    layer5_outputs(8936) <= not b or a;
    layer5_outputs(8937) <= not (a or b);
    layer5_outputs(8938) <= not b or a;
    layer5_outputs(8939) <= b;
    layer5_outputs(8940) <= not (a xor b);
    layer5_outputs(8941) <= a and not b;
    layer5_outputs(8942) <= b;
    layer5_outputs(8943) <= not a;
    layer5_outputs(8944) <= not b;
    layer5_outputs(8945) <= not (a xor b);
    layer5_outputs(8946) <= a;
    layer5_outputs(8947) <= b;
    layer5_outputs(8948) <= '1';
    layer5_outputs(8949) <= not (a xor b);
    layer5_outputs(8950) <= b and not a;
    layer5_outputs(8951) <= b and not a;
    layer5_outputs(8952) <= a and not b;
    layer5_outputs(8953) <= a;
    layer5_outputs(8954) <= a or b;
    layer5_outputs(8955) <= not b;
    layer5_outputs(8956) <= not b or a;
    layer5_outputs(8957) <= not b;
    layer5_outputs(8958) <= not b;
    layer5_outputs(8959) <= b;
    layer5_outputs(8960) <= a xor b;
    layer5_outputs(8961) <= a xor b;
    layer5_outputs(8962) <= a and not b;
    layer5_outputs(8963) <= a xor b;
    layer5_outputs(8964) <= not a;
    layer5_outputs(8965) <= not (a and b);
    layer5_outputs(8966) <= a or b;
    layer5_outputs(8967) <= a;
    layer5_outputs(8968) <= not a;
    layer5_outputs(8969) <= a and not b;
    layer5_outputs(8970) <= not (a and b);
    layer5_outputs(8971) <= a or b;
    layer5_outputs(8972) <= not a;
    layer5_outputs(8973) <= b and not a;
    layer5_outputs(8974) <= a xor b;
    layer5_outputs(8975) <= a and not b;
    layer5_outputs(8976) <= not b or a;
    layer5_outputs(8977) <= b;
    layer5_outputs(8978) <= a;
    layer5_outputs(8979) <= b;
    layer5_outputs(8980) <= b;
    layer5_outputs(8981) <= not b;
    layer5_outputs(8982) <= not b;
    layer5_outputs(8983) <= b;
    layer5_outputs(8984) <= not a;
    layer5_outputs(8985) <= not a or b;
    layer5_outputs(8986) <= not b;
    layer5_outputs(8987) <= not (a and b);
    layer5_outputs(8988) <= not (a xor b);
    layer5_outputs(8989) <= a and not b;
    layer5_outputs(8990) <= not a;
    layer5_outputs(8991) <= a xor b;
    layer5_outputs(8992) <= b and not a;
    layer5_outputs(8993) <= not a or b;
    layer5_outputs(8994) <= a;
    layer5_outputs(8995) <= a or b;
    layer5_outputs(8996) <= b;
    layer5_outputs(8997) <= not (a or b);
    layer5_outputs(8998) <= a and b;
    layer5_outputs(8999) <= not (a xor b);
    layer5_outputs(9000) <= not b or a;
    layer5_outputs(9001) <= a;
    layer5_outputs(9002) <= not a;
    layer5_outputs(9003) <= b;
    layer5_outputs(9004) <= not a;
    layer5_outputs(9005) <= a;
    layer5_outputs(9006) <= not (a xor b);
    layer5_outputs(9007) <= not a or b;
    layer5_outputs(9008) <= not (a or b);
    layer5_outputs(9009) <= not (a or b);
    layer5_outputs(9010) <= not a;
    layer5_outputs(9011) <= not b or a;
    layer5_outputs(9012) <= b;
    layer5_outputs(9013) <= a;
    layer5_outputs(9014) <= a and not b;
    layer5_outputs(9015) <= not (a xor b);
    layer5_outputs(9016) <= a or b;
    layer5_outputs(9017) <= a xor b;
    layer5_outputs(9018) <= a;
    layer5_outputs(9019) <= b and not a;
    layer5_outputs(9020) <= a and b;
    layer5_outputs(9021) <= a and b;
    layer5_outputs(9022) <= not (a xor b);
    layer5_outputs(9023) <= not a;
    layer5_outputs(9024) <= not a or b;
    layer5_outputs(9025) <= not (a or b);
    layer5_outputs(9026) <= a or b;
    layer5_outputs(9027) <= not b or a;
    layer5_outputs(9028) <= not b;
    layer5_outputs(9029) <= a xor b;
    layer5_outputs(9030) <= not b or a;
    layer5_outputs(9031) <= not b or a;
    layer5_outputs(9032) <= b;
    layer5_outputs(9033) <= a xor b;
    layer5_outputs(9034) <= not b;
    layer5_outputs(9035) <= a or b;
    layer5_outputs(9036) <= not a or b;
    layer5_outputs(9037) <= a;
    layer5_outputs(9038) <= not b or a;
    layer5_outputs(9039) <= a xor b;
    layer5_outputs(9040) <= b and not a;
    layer5_outputs(9041) <= not (a or b);
    layer5_outputs(9042) <= not b or a;
    layer5_outputs(9043) <= a or b;
    layer5_outputs(9044) <= not b;
    layer5_outputs(9045) <= not b;
    layer5_outputs(9046) <= not (a and b);
    layer5_outputs(9047) <= not b;
    layer5_outputs(9048) <= not a;
    layer5_outputs(9049) <= a or b;
    layer5_outputs(9050) <= a xor b;
    layer5_outputs(9051) <= b;
    layer5_outputs(9052) <= not (a xor b);
    layer5_outputs(9053) <= a;
    layer5_outputs(9054) <= not (a or b);
    layer5_outputs(9055) <= not a;
    layer5_outputs(9056) <= a and b;
    layer5_outputs(9057) <= a;
    layer5_outputs(9058) <= a and not b;
    layer5_outputs(9059) <= not (a xor b);
    layer5_outputs(9060) <= not a;
    layer5_outputs(9061) <= a or b;
    layer5_outputs(9062) <= not b;
    layer5_outputs(9063) <= not (a xor b);
    layer5_outputs(9064) <= a xor b;
    layer5_outputs(9065) <= a;
    layer5_outputs(9066) <= not a;
    layer5_outputs(9067) <= not a;
    layer5_outputs(9068) <= a and not b;
    layer5_outputs(9069) <= a;
    layer5_outputs(9070) <= not (a and b);
    layer5_outputs(9071) <= not a or b;
    layer5_outputs(9072) <= '1';
    layer5_outputs(9073) <= not (a and b);
    layer5_outputs(9074) <= not (a and b);
    layer5_outputs(9075) <= a and b;
    layer5_outputs(9076) <= not b;
    layer5_outputs(9077) <= a xor b;
    layer5_outputs(9078) <= not a;
    layer5_outputs(9079) <= b and not a;
    layer5_outputs(9080) <= not a;
    layer5_outputs(9081) <= a or b;
    layer5_outputs(9082) <= not (a xor b);
    layer5_outputs(9083) <= not (a and b);
    layer5_outputs(9084) <= '0';
    layer5_outputs(9085) <= not b or a;
    layer5_outputs(9086) <= a;
    layer5_outputs(9087) <= b;
    layer5_outputs(9088) <= a;
    layer5_outputs(9089) <= a and b;
    layer5_outputs(9090) <= not (a xor b);
    layer5_outputs(9091) <= a xor b;
    layer5_outputs(9092) <= not b or a;
    layer5_outputs(9093) <= not b or a;
    layer5_outputs(9094) <= a xor b;
    layer5_outputs(9095) <= a;
    layer5_outputs(9096) <= a;
    layer5_outputs(9097) <= not a;
    layer5_outputs(9098) <= not (a xor b);
    layer5_outputs(9099) <= a and not b;
    layer5_outputs(9100) <= a xor b;
    layer5_outputs(9101) <= a and not b;
    layer5_outputs(9102) <= a;
    layer5_outputs(9103) <= not (a xor b);
    layer5_outputs(9104) <= a;
    layer5_outputs(9105) <= a xor b;
    layer5_outputs(9106) <= b;
    layer5_outputs(9107) <= b;
    layer5_outputs(9108) <= not (a and b);
    layer5_outputs(9109) <= not a;
    layer5_outputs(9110) <= b and not a;
    layer5_outputs(9111) <= b;
    layer5_outputs(9112) <= not a;
    layer5_outputs(9113) <= not b or a;
    layer5_outputs(9114) <= not b;
    layer5_outputs(9115) <= not (a or b);
    layer5_outputs(9116) <= not a;
    layer5_outputs(9117) <= not (a or b);
    layer5_outputs(9118) <= not (a and b);
    layer5_outputs(9119) <= a and not b;
    layer5_outputs(9120) <= a;
    layer5_outputs(9121) <= not (a and b);
    layer5_outputs(9122) <= not (a and b);
    layer5_outputs(9123) <= not b;
    layer5_outputs(9124) <= not b;
    layer5_outputs(9125) <= b;
    layer5_outputs(9126) <= a;
    layer5_outputs(9127) <= not b or a;
    layer5_outputs(9128) <= not (a and b);
    layer5_outputs(9129) <= not (a xor b);
    layer5_outputs(9130) <= not b;
    layer5_outputs(9131) <= b and not a;
    layer5_outputs(9132) <= a and b;
    layer5_outputs(9133) <= not b;
    layer5_outputs(9134) <= not (a or b);
    layer5_outputs(9135) <= a and b;
    layer5_outputs(9136) <= not a or b;
    layer5_outputs(9137) <= a;
    layer5_outputs(9138) <= not b;
    layer5_outputs(9139) <= not (a and b);
    layer5_outputs(9140) <= not (a or b);
    layer5_outputs(9141) <= a xor b;
    layer5_outputs(9142) <= a xor b;
    layer5_outputs(9143) <= not (a and b);
    layer5_outputs(9144) <= a;
    layer5_outputs(9145) <= not b;
    layer5_outputs(9146) <= not b;
    layer5_outputs(9147) <= a and not b;
    layer5_outputs(9148) <= a;
    layer5_outputs(9149) <= not b or a;
    layer5_outputs(9150) <= a xor b;
    layer5_outputs(9151) <= a and b;
    layer5_outputs(9152) <= a;
    layer5_outputs(9153) <= '0';
    layer5_outputs(9154) <= '0';
    layer5_outputs(9155) <= not a;
    layer5_outputs(9156) <= b;
    layer5_outputs(9157) <= not a or b;
    layer5_outputs(9158) <= not b;
    layer5_outputs(9159) <= a;
    layer5_outputs(9160) <= not a or b;
    layer5_outputs(9161) <= a and b;
    layer5_outputs(9162) <= b;
    layer5_outputs(9163) <= b;
    layer5_outputs(9164) <= not a or b;
    layer5_outputs(9165) <= not (a xor b);
    layer5_outputs(9166) <= b;
    layer5_outputs(9167) <= a;
    layer5_outputs(9168) <= not b;
    layer5_outputs(9169) <= a or b;
    layer5_outputs(9170) <= not (a and b);
    layer5_outputs(9171) <= a;
    layer5_outputs(9172) <= not a or b;
    layer5_outputs(9173) <= not a;
    layer5_outputs(9174) <= not b;
    layer5_outputs(9175) <= a or b;
    layer5_outputs(9176) <= not (a or b);
    layer5_outputs(9177) <= a xor b;
    layer5_outputs(9178) <= a xor b;
    layer5_outputs(9179) <= a and not b;
    layer5_outputs(9180) <= a and not b;
    layer5_outputs(9181) <= a xor b;
    layer5_outputs(9182) <= not (a or b);
    layer5_outputs(9183) <= b and not a;
    layer5_outputs(9184) <= not (a xor b);
    layer5_outputs(9185) <= a xor b;
    layer5_outputs(9186) <= not b or a;
    layer5_outputs(9187) <= not a;
    layer5_outputs(9188) <= a and b;
    layer5_outputs(9189) <= a xor b;
    layer5_outputs(9190) <= not (a and b);
    layer5_outputs(9191) <= a or b;
    layer5_outputs(9192) <= not b;
    layer5_outputs(9193) <= a and b;
    layer5_outputs(9194) <= a;
    layer5_outputs(9195) <= not b or a;
    layer5_outputs(9196) <= not a;
    layer5_outputs(9197) <= a xor b;
    layer5_outputs(9198) <= a;
    layer5_outputs(9199) <= not b;
    layer5_outputs(9200) <= a;
    layer5_outputs(9201) <= not (a xor b);
    layer5_outputs(9202) <= a;
    layer5_outputs(9203) <= a or b;
    layer5_outputs(9204) <= a;
    layer5_outputs(9205) <= b and not a;
    layer5_outputs(9206) <= a and b;
    layer5_outputs(9207) <= a and b;
    layer5_outputs(9208) <= not a;
    layer5_outputs(9209) <= a or b;
    layer5_outputs(9210) <= a;
    layer5_outputs(9211) <= a and not b;
    layer5_outputs(9212) <= not b;
    layer5_outputs(9213) <= not b or a;
    layer5_outputs(9214) <= a;
    layer5_outputs(9215) <= a or b;
    layer5_outputs(9216) <= not a;
    layer5_outputs(9217) <= a;
    layer5_outputs(9218) <= not b or a;
    layer5_outputs(9219) <= b;
    layer5_outputs(9220) <= b;
    layer5_outputs(9221) <= not b;
    layer5_outputs(9222) <= a or b;
    layer5_outputs(9223) <= a or b;
    layer5_outputs(9224) <= a and not b;
    layer5_outputs(9225) <= a;
    layer5_outputs(9226) <= not b;
    layer5_outputs(9227) <= not (a xor b);
    layer5_outputs(9228) <= not b or a;
    layer5_outputs(9229) <= a and b;
    layer5_outputs(9230) <= a;
    layer5_outputs(9231) <= not b or a;
    layer5_outputs(9232) <= not a;
    layer5_outputs(9233) <= not (a or b);
    layer5_outputs(9234) <= not b;
    layer5_outputs(9235) <= b and not a;
    layer5_outputs(9236) <= a;
    layer5_outputs(9237) <= not (a or b);
    layer5_outputs(9238) <= not (a or b);
    layer5_outputs(9239) <= a;
    layer5_outputs(9240) <= a or b;
    layer5_outputs(9241) <= a;
    layer5_outputs(9242) <= not a;
    layer5_outputs(9243) <= a;
    layer5_outputs(9244) <= b;
    layer5_outputs(9245) <= not (a or b);
    layer5_outputs(9246) <= a;
    layer5_outputs(9247) <= not (a or b);
    layer5_outputs(9248) <= a and not b;
    layer5_outputs(9249) <= a;
    layer5_outputs(9250) <= '0';
    layer5_outputs(9251) <= not (a and b);
    layer5_outputs(9252) <= not a;
    layer5_outputs(9253) <= not a;
    layer5_outputs(9254) <= b;
    layer5_outputs(9255) <= not b;
    layer5_outputs(9256) <= a;
    layer5_outputs(9257) <= b;
    layer5_outputs(9258) <= a xor b;
    layer5_outputs(9259) <= not b;
    layer5_outputs(9260) <= not (a and b);
    layer5_outputs(9261) <= b;
    layer5_outputs(9262) <= not b;
    layer5_outputs(9263) <= a and b;
    layer5_outputs(9264) <= not (a or b);
    layer5_outputs(9265) <= not b or a;
    layer5_outputs(9266) <= a or b;
    layer5_outputs(9267) <= a;
    layer5_outputs(9268) <= not (a xor b);
    layer5_outputs(9269) <= a;
    layer5_outputs(9270) <= not b;
    layer5_outputs(9271) <= a and not b;
    layer5_outputs(9272) <= not b or a;
    layer5_outputs(9273) <= not b;
    layer5_outputs(9274) <= b;
    layer5_outputs(9275) <= not a or b;
    layer5_outputs(9276) <= not (a and b);
    layer5_outputs(9277) <= not a or b;
    layer5_outputs(9278) <= not b or a;
    layer5_outputs(9279) <= b;
    layer5_outputs(9280) <= a or b;
    layer5_outputs(9281) <= a or b;
    layer5_outputs(9282) <= not a;
    layer5_outputs(9283) <= not a;
    layer5_outputs(9284) <= not b;
    layer5_outputs(9285) <= b;
    layer5_outputs(9286) <= not a or b;
    layer5_outputs(9287) <= not a;
    layer5_outputs(9288) <= not a;
    layer5_outputs(9289) <= not b;
    layer5_outputs(9290) <= a and not b;
    layer5_outputs(9291) <= not (a and b);
    layer5_outputs(9292) <= b;
    layer5_outputs(9293) <= not a or b;
    layer5_outputs(9294) <= not b;
    layer5_outputs(9295) <= b;
    layer5_outputs(9296) <= b;
    layer5_outputs(9297) <= not b or a;
    layer5_outputs(9298) <= not a;
    layer5_outputs(9299) <= a and not b;
    layer5_outputs(9300) <= not a or b;
    layer5_outputs(9301) <= a;
    layer5_outputs(9302) <= not (a and b);
    layer5_outputs(9303) <= not a or b;
    layer5_outputs(9304) <= not (a and b);
    layer5_outputs(9305) <= a;
    layer5_outputs(9306) <= not a;
    layer5_outputs(9307) <= a xor b;
    layer5_outputs(9308) <= not (a xor b);
    layer5_outputs(9309) <= not (a or b);
    layer5_outputs(9310) <= not b;
    layer5_outputs(9311) <= b and not a;
    layer5_outputs(9312) <= a and b;
    layer5_outputs(9313) <= a;
    layer5_outputs(9314) <= not b;
    layer5_outputs(9315) <= not b or a;
    layer5_outputs(9316) <= not b;
    layer5_outputs(9317) <= a and b;
    layer5_outputs(9318) <= a or b;
    layer5_outputs(9319) <= not b or a;
    layer5_outputs(9320) <= b and not a;
    layer5_outputs(9321) <= not a or b;
    layer5_outputs(9322) <= b;
    layer5_outputs(9323) <= not a;
    layer5_outputs(9324) <= not b;
    layer5_outputs(9325) <= not a or b;
    layer5_outputs(9326) <= not b;
    layer5_outputs(9327) <= b;
    layer5_outputs(9328) <= not b;
    layer5_outputs(9329) <= not a;
    layer5_outputs(9330) <= not (a xor b);
    layer5_outputs(9331) <= not b;
    layer5_outputs(9332) <= b;
    layer5_outputs(9333) <= not a;
    layer5_outputs(9334) <= not a;
    layer5_outputs(9335) <= a or b;
    layer5_outputs(9336) <= a and b;
    layer5_outputs(9337) <= not (a or b);
    layer5_outputs(9338) <= a or b;
    layer5_outputs(9339) <= b;
    layer5_outputs(9340) <= a and b;
    layer5_outputs(9341) <= not (a or b);
    layer5_outputs(9342) <= a;
    layer5_outputs(9343) <= not a or b;
    layer5_outputs(9344) <= not a;
    layer5_outputs(9345) <= not a;
    layer5_outputs(9346) <= not b or a;
    layer5_outputs(9347) <= b;
    layer5_outputs(9348) <= a;
    layer5_outputs(9349) <= not b;
    layer5_outputs(9350) <= b;
    layer5_outputs(9351) <= b;
    layer5_outputs(9352) <= not (a or b);
    layer5_outputs(9353) <= b;
    layer5_outputs(9354) <= not (a and b);
    layer5_outputs(9355) <= b;
    layer5_outputs(9356) <= not b;
    layer5_outputs(9357) <= not b;
    layer5_outputs(9358) <= not a or b;
    layer5_outputs(9359) <= a or b;
    layer5_outputs(9360) <= a xor b;
    layer5_outputs(9361) <= not (a and b);
    layer5_outputs(9362) <= a;
    layer5_outputs(9363) <= a xor b;
    layer5_outputs(9364) <= not a;
    layer5_outputs(9365) <= a and not b;
    layer5_outputs(9366) <= not a;
    layer5_outputs(9367) <= a;
    layer5_outputs(9368) <= not a;
    layer5_outputs(9369) <= a;
    layer5_outputs(9370) <= not a;
    layer5_outputs(9371) <= not b or a;
    layer5_outputs(9372) <= b;
    layer5_outputs(9373) <= not (a and b);
    layer5_outputs(9374) <= not a;
    layer5_outputs(9375) <= b and not a;
    layer5_outputs(9376) <= not (a xor b);
    layer5_outputs(9377) <= a xor b;
    layer5_outputs(9378) <= not (a or b);
    layer5_outputs(9379) <= '1';
    layer5_outputs(9380) <= b and not a;
    layer5_outputs(9381) <= a xor b;
    layer5_outputs(9382) <= a;
    layer5_outputs(9383) <= b and not a;
    layer5_outputs(9384) <= not (a and b);
    layer5_outputs(9385) <= not (a xor b);
    layer5_outputs(9386) <= b;
    layer5_outputs(9387) <= not a;
    layer5_outputs(9388) <= a and not b;
    layer5_outputs(9389) <= not b or a;
    layer5_outputs(9390) <= not a;
    layer5_outputs(9391) <= b;
    layer5_outputs(9392) <= not (a xor b);
    layer5_outputs(9393) <= a and not b;
    layer5_outputs(9394) <= not b;
    layer5_outputs(9395) <= a;
    layer5_outputs(9396) <= a and b;
    layer5_outputs(9397) <= a and not b;
    layer5_outputs(9398) <= not a;
    layer5_outputs(9399) <= b;
    layer5_outputs(9400) <= a;
    layer5_outputs(9401) <= not (a or b);
    layer5_outputs(9402) <= b;
    layer5_outputs(9403) <= a and not b;
    layer5_outputs(9404) <= not a;
    layer5_outputs(9405) <= b and not a;
    layer5_outputs(9406) <= b and not a;
    layer5_outputs(9407) <= not (a xor b);
    layer5_outputs(9408) <= b;
    layer5_outputs(9409) <= not b;
    layer5_outputs(9410) <= b;
    layer5_outputs(9411) <= a;
    layer5_outputs(9412) <= a xor b;
    layer5_outputs(9413) <= b;
    layer5_outputs(9414) <= not (a xor b);
    layer5_outputs(9415) <= b;
    layer5_outputs(9416) <= not (a and b);
    layer5_outputs(9417) <= not (a and b);
    layer5_outputs(9418) <= a;
    layer5_outputs(9419) <= a;
    layer5_outputs(9420) <= not a or b;
    layer5_outputs(9421) <= not a;
    layer5_outputs(9422) <= not (a xor b);
    layer5_outputs(9423) <= not a or b;
    layer5_outputs(9424) <= a;
    layer5_outputs(9425) <= '0';
    layer5_outputs(9426) <= a and b;
    layer5_outputs(9427) <= a xor b;
    layer5_outputs(9428) <= not (a or b);
    layer5_outputs(9429) <= b;
    layer5_outputs(9430) <= not (a and b);
    layer5_outputs(9431) <= not (a and b);
    layer5_outputs(9432) <= not b;
    layer5_outputs(9433) <= not (a and b);
    layer5_outputs(9434) <= not a;
    layer5_outputs(9435) <= a;
    layer5_outputs(9436) <= a and not b;
    layer5_outputs(9437) <= not b or a;
    layer5_outputs(9438) <= a;
    layer5_outputs(9439) <= not (a or b);
    layer5_outputs(9440) <= not b or a;
    layer5_outputs(9441) <= a;
    layer5_outputs(9442) <= a and b;
    layer5_outputs(9443) <= b and not a;
    layer5_outputs(9444) <= not a;
    layer5_outputs(9445) <= not b or a;
    layer5_outputs(9446) <= not b;
    layer5_outputs(9447) <= not b;
    layer5_outputs(9448) <= b;
    layer5_outputs(9449) <= a xor b;
    layer5_outputs(9450) <= not a;
    layer5_outputs(9451) <= not (a xor b);
    layer5_outputs(9452) <= not b or a;
    layer5_outputs(9453) <= a or b;
    layer5_outputs(9454) <= a and not b;
    layer5_outputs(9455) <= not b;
    layer5_outputs(9456) <= not b or a;
    layer5_outputs(9457) <= not a;
    layer5_outputs(9458) <= a xor b;
    layer5_outputs(9459) <= not a;
    layer5_outputs(9460) <= a and not b;
    layer5_outputs(9461) <= a and not b;
    layer5_outputs(9462) <= b;
    layer5_outputs(9463) <= not b;
    layer5_outputs(9464) <= not (a xor b);
    layer5_outputs(9465) <= a or b;
    layer5_outputs(9466) <= not (a xor b);
    layer5_outputs(9467) <= b;
    layer5_outputs(9468) <= a and b;
    layer5_outputs(9469) <= a or b;
    layer5_outputs(9470) <= b and not a;
    layer5_outputs(9471) <= not b or a;
    layer5_outputs(9472) <= b and not a;
    layer5_outputs(9473) <= a and b;
    layer5_outputs(9474) <= not (a and b);
    layer5_outputs(9475) <= not (a or b);
    layer5_outputs(9476) <= b and not a;
    layer5_outputs(9477) <= not a;
    layer5_outputs(9478) <= not a;
    layer5_outputs(9479) <= not (a xor b);
    layer5_outputs(9480) <= not (a and b);
    layer5_outputs(9481) <= not (a xor b);
    layer5_outputs(9482) <= not b;
    layer5_outputs(9483) <= b and not a;
    layer5_outputs(9484) <= b and not a;
    layer5_outputs(9485) <= a;
    layer5_outputs(9486) <= a and not b;
    layer5_outputs(9487) <= b;
    layer5_outputs(9488) <= a and not b;
    layer5_outputs(9489) <= a;
    layer5_outputs(9490) <= b and not a;
    layer5_outputs(9491) <= a;
    layer5_outputs(9492) <= b and not a;
    layer5_outputs(9493) <= b;
    layer5_outputs(9494) <= not b or a;
    layer5_outputs(9495) <= a;
    layer5_outputs(9496) <= a xor b;
    layer5_outputs(9497) <= not (a xor b);
    layer5_outputs(9498) <= a and not b;
    layer5_outputs(9499) <= b;
    layer5_outputs(9500) <= not b or a;
    layer5_outputs(9501) <= a xor b;
    layer5_outputs(9502) <= not a;
    layer5_outputs(9503) <= b and not a;
    layer5_outputs(9504) <= not a or b;
    layer5_outputs(9505) <= a and b;
    layer5_outputs(9506) <= not b;
    layer5_outputs(9507) <= '0';
    layer5_outputs(9508) <= a and not b;
    layer5_outputs(9509) <= not (a and b);
    layer5_outputs(9510) <= a or b;
    layer5_outputs(9511) <= b;
    layer5_outputs(9512) <= a or b;
    layer5_outputs(9513) <= a xor b;
    layer5_outputs(9514) <= a or b;
    layer5_outputs(9515) <= not (a xor b);
    layer5_outputs(9516) <= not (a and b);
    layer5_outputs(9517) <= not (a or b);
    layer5_outputs(9518) <= a and b;
    layer5_outputs(9519) <= not a or b;
    layer5_outputs(9520) <= a xor b;
    layer5_outputs(9521) <= b;
    layer5_outputs(9522) <= a and b;
    layer5_outputs(9523) <= a xor b;
    layer5_outputs(9524) <= a and b;
    layer5_outputs(9525) <= a;
    layer5_outputs(9526) <= a and b;
    layer5_outputs(9527) <= a and b;
    layer5_outputs(9528) <= not b or a;
    layer5_outputs(9529) <= b and not a;
    layer5_outputs(9530) <= a and b;
    layer5_outputs(9531) <= not b;
    layer5_outputs(9532) <= b;
    layer5_outputs(9533) <= a and not b;
    layer5_outputs(9534) <= not (a and b);
    layer5_outputs(9535) <= not (a and b);
    layer5_outputs(9536) <= not (a xor b);
    layer5_outputs(9537) <= a;
    layer5_outputs(9538) <= b;
    layer5_outputs(9539) <= '0';
    layer5_outputs(9540) <= a xor b;
    layer5_outputs(9541) <= a xor b;
    layer5_outputs(9542) <= not (a or b);
    layer5_outputs(9543) <= a xor b;
    layer5_outputs(9544) <= b;
    layer5_outputs(9545) <= a;
    layer5_outputs(9546) <= a;
    layer5_outputs(9547) <= not b;
    layer5_outputs(9548) <= not b;
    layer5_outputs(9549) <= b;
    layer5_outputs(9550) <= not (a xor b);
    layer5_outputs(9551) <= b;
    layer5_outputs(9552) <= not b;
    layer5_outputs(9553) <= not a or b;
    layer5_outputs(9554) <= not a;
    layer5_outputs(9555) <= a or b;
    layer5_outputs(9556) <= a xor b;
    layer5_outputs(9557) <= not b;
    layer5_outputs(9558) <= not (a or b);
    layer5_outputs(9559) <= not a or b;
    layer5_outputs(9560) <= b and not a;
    layer5_outputs(9561) <= a;
    layer5_outputs(9562) <= b and not a;
    layer5_outputs(9563) <= a;
    layer5_outputs(9564) <= not b or a;
    layer5_outputs(9565) <= not (a xor b);
    layer5_outputs(9566) <= not b or a;
    layer5_outputs(9567) <= a and not b;
    layer5_outputs(9568) <= b and not a;
    layer5_outputs(9569) <= a or b;
    layer5_outputs(9570) <= b;
    layer5_outputs(9571) <= a and not b;
    layer5_outputs(9572) <= not a;
    layer5_outputs(9573) <= b and not a;
    layer5_outputs(9574) <= not b;
    layer5_outputs(9575) <= a xor b;
    layer5_outputs(9576) <= not (a and b);
    layer5_outputs(9577) <= '0';
    layer5_outputs(9578) <= not b;
    layer5_outputs(9579) <= not (a or b);
    layer5_outputs(9580) <= not b;
    layer5_outputs(9581) <= not (a and b);
    layer5_outputs(9582) <= not a;
    layer5_outputs(9583) <= not (a and b);
    layer5_outputs(9584) <= a xor b;
    layer5_outputs(9585) <= a and not b;
    layer5_outputs(9586) <= a or b;
    layer5_outputs(9587) <= not a;
    layer5_outputs(9588) <= a or b;
    layer5_outputs(9589) <= not (a xor b);
    layer5_outputs(9590) <= a and b;
    layer5_outputs(9591) <= not a;
    layer5_outputs(9592) <= not (a and b);
    layer5_outputs(9593) <= a and b;
    layer5_outputs(9594) <= not (a xor b);
    layer5_outputs(9595) <= a;
    layer5_outputs(9596) <= b and not a;
    layer5_outputs(9597) <= b;
    layer5_outputs(9598) <= b;
    layer5_outputs(9599) <= a xor b;
    layer5_outputs(9600) <= not a;
    layer5_outputs(9601) <= not a or b;
    layer5_outputs(9602) <= not a or b;
    layer5_outputs(9603) <= not b or a;
    layer5_outputs(9604) <= not b or a;
    layer5_outputs(9605) <= not (a xor b);
    layer5_outputs(9606) <= a and b;
    layer5_outputs(9607) <= b;
    layer5_outputs(9608) <= a and b;
    layer5_outputs(9609) <= not b;
    layer5_outputs(9610) <= a;
    layer5_outputs(9611) <= b and not a;
    layer5_outputs(9612) <= a or b;
    layer5_outputs(9613) <= a or b;
    layer5_outputs(9614) <= a and not b;
    layer5_outputs(9615) <= not a or b;
    layer5_outputs(9616) <= not b;
    layer5_outputs(9617) <= a and not b;
    layer5_outputs(9618) <= a;
    layer5_outputs(9619) <= a;
    layer5_outputs(9620) <= a and not b;
    layer5_outputs(9621) <= a or b;
    layer5_outputs(9622) <= a;
    layer5_outputs(9623) <= not a;
    layer5_outputs(9624) <= not b;
    layer5_outputs(9625) <= a xor b;
    layer5_outputs(9626) <= a xor b;
    layer5_outputs(9627) <= a;
    layer5_outputs(9628) <= a and b;
    layer5_outputs(9629) <= a xor b;
    layer5_outputs(9630) <= not (a or b);
    layer5_outputs(9631) <= not (a or b);
    layer5_outputs(9632) <= a;
    layer5_outputs(9633) <= b and not a;
    layer5_outputs(9634) <= a xor b;
    layer5_outputs(9635) <= b and not a;
    layer5_outputs(9636) <= b;
    layer5_outputs(9637) <= '1';
    layer5_outputs(9638) <= b;
    layer5_outputs(9639) <= not a;
    layer5_outputs(9640) <= not b;
    layer5_outputs(9641) <= a and b;
    layer5_outputs(9642) <= not (a xor b);
    layer5_outputs(9643) <= not a or b;
    layer5_outputs(9644) <= not b;
    layer5_outputs(9645) <= not b;
    layer5_outputs(9646) <= b;
    layer5_outputs(9647) <= '1';
    layer5_outputs(9648) <= not b;
    layer5_outputs(9649) <= a;
    layer5_outputs(9650) <= not (a and b);
    layer5_outputs(9651) <= b;
    layer5_outputs(9652) <= not a;
    layer5_outputs(9653) <= not a;
    layer5_outputs(9654) <= a;
    layer5_outputs(9655) <= not b;
    layer5_outputs(9656) <= '0';
    layer5_outputs(9657) <= a;
    layer5_outputs(9658) <= a or b;
    layer5_outputs(9659) <= not a;
    layer5_outputs(9660) <= b;
    layer5_outputs(9661) <= not b;
    layer5_outputs(9662) <= a and b;
    layer5_outputs(9663) <= b;
    layer5_outputs(9664) <= b and not a;
    layer5_outputs(9665) <= a and b;
    layer5_outputs(9666) <= '1';
    layer5_outputs(9667) <= not b or a;
    layer5_outputs(9668) <= not b;
    layer5_outputs(9669) <= a and not b;
    layer5_outputs(9670) <= not (a xor b);
    layer5_outputs(9671) <= not a or b;
    layer5_outputs(9672) <= a and b;
    layer5_outputs(9673) <= a and not b;
    layer5_outputs(9674) <= not (a xor b);
    layer5_outputs(9675) <= not a or b;
    layer5_outputs(9676) <= a and not b;
    layer5_outputs(9677) <= not (a and b);
    layer5_outputs(9678) <= not b;
    layer5_outputs(9679) <= a;
    layer5_outputs(9680) <= b;
    layer5_outputs(9681) <= not b or a;
    layer5_outputs(9682) <= not b;
    layer5_outputs(9683) <= not b;
    layer5_outputs(9684) <= not (a xor b);
    layer5_outputs(9685) <= a and b;
    layer5_outputs(9686) <= a;
    layer5_outputs(9687) <= a;
    layer5_outputs(9688) <= not b;
    layer5_outputs(9689) <= b;
    layer5_outputs(9690) <= not a or b;
    layer5_outputs(9691) <= b and not a;
    layer5_outputs(9692) <= b;
    layer5_outputs(9693) <= not (a and b);
    layer5_outputs(9694) <= not (a or b);
    layer5_outputs(9695) <= not (a xor b);
    layer5_outputs(9696) <= a and not b;
    layer5_outputs(9697) <= not a;
    layer5_outputs(9698) <= b and not a;
    layer5_outputs(9699) <= b;
    layer5_outputs(9700) <= not a;
    layer5_outputs(9701) <= not (a or b);
    layer5_outputs(9702) <= not b;
    layer5_outputs(9703) <= not a;
    layer5_outputs(9704) <= b;
    layer5_outputs(9705) <= a xor b;
    layer5_outputs(9706) <= not (a and b);
    layer5_outputs(9707) <= not b;
    layer5_outputs(9708) <= a or b;
    layer5_outputs(9709) <= not b;
    layer5_outputs(9710) <= not a;
    layer5_outputs(9711) <= a xor b;
    layer5_outputs(9712) <= b and not a;
    layer5_outputs(9713) <= a;
    layer5_outputs(9714) <= b;
    layer5_outputs(9715) <= not (a xor b);
    layer5_outputs(9716) <= not a;
    layer5_outputs(9717) <= b;
    layer5_outputs(9718) <= a and b;
    layer5_outputs(9719) <= not a;
    layer5_outputs(9720) <= not a;
    layer5_outputs(9721) <= b and not a;
    layer5_outputs(9722) <= not b;
    layer5_outputs(9723) <= a xor b;
    layer5_outputs(9724) <= not a;
    layer5_outputs(9725) <= b;
    layer5_outputs(9726) <= not b or a;
    layer5_outputs(9727) <= '1';
    layer5_outputs(9728) <= b and not a;
    layer5_outputs(9729) <= not b or a;
    layer5_outputs(9730) <= a;
    layer5_outputs(9731) <= a xor b;
    layer5_outputs(9732) <= a;
    layer5_outputs(9733) <= a and not b;
    layer5_outputs(9734) <= a or b;
    layer5_outputs(9735) <= not b;
    layer5_outputs(9736) <= not (a xor b);
    layer5_outputs(9737) <= a or b;
    layer5_outputs(9738) <= a and not b;
    layer5_outputs(9739) <= a;
    layer5_outputs(9740) <= a;
    layer5_outputs(9741) <= a xor b;
    layer5_outputs(9742) <= not (a and b);
    layer5_outputs(9743) <= not a;
    layer5_outputs(9744) <= b and not a;
    layer5_outputs(9745) <= a and not b;
    layer5_outputs(9746) <= not a;
    layer5_outputs(9747) <= not b or a;
    layer5_outputs(9748) <= a xor b;
    layer5_outputs(9749) <= a and not b;
    layer5_outputs(9750) <= b;
    layer5_outputs(9751) <= a xor b;
    layer5_outputs(9752) <= not (a xor b);
    layer5_outputs(9753) <= not b or a;
    layer5_outputs(9754) <= not a or b;
    layer5_outputs(9755) <= not b or a;
    layer5_outputs(9756) <= b;
    layer5_outputs(9757) <= a;
    layer5_outputs(9758) <= not a;
    layer5_outputs(9759) <= a and b;
    layer5_outputs(9760) <= not b;
    layer5_outputs(9761) <= not a;
    layer5_outputs(9762) <= b;
    layer5_outputs(9763) <= b and not a;
    layer5_outputs(9764) <= '1';
    layer5_outputs(9765) <= not a;
    layer5_outputs(9766) <= not (a and b);
    layer5_outputs(9767) <= a and not b;
    layer5_outputs(9768) <= not b;
    layer5_outputs(9769) <= not b;
    layer5_outputs(9770) <= a and b;
    layer5_outputs(9771) <= not (a and b);
    layer5_outputs(9772) <= a;
    layer5_outputs(9773) <= a xor b;
    layer5_outputs(9774) <= not b;
    layer5_outputs(9775) <= a xor b;
    layer5_outputs(9776) <= a or b;
    layer5_outputs(9777) <= not (a xor b);
    layer5_outputs(9778) <= a and b;
    layer5_outputs(9779) <= not a;
    layer5_outputs(9780) <= not a or b;
    layer5_outputs(9781) <= a or b;
    layer5_outputs(9782) <= b;
    layer5_outputs(9783) <= b and not a;
    layer5_outputs(9784) <= a and not b;
    layer5_outputs(9785) <= not a or b;
    layer5_outputs(9786) <= a xor b;
    layer5_outputs(9787) <= a xor b;
    layer5_outputs(9788) <= a and b;
    layer5_outputs(9789) <= not b or a;
    layer5_outputs(9790) <= a xor b;
    layer5_outputs(9791) <= b and not a;
    layer5_outputs(9792) <= b;
    layer5_outputs(9793) <= '1';
    layer5_outputs(9794) <= not (a and b);
    layer5_outputs(9795) <= a and not b;
    layer5_outputs(9796) <= not a;
    layer5_outputs(9797) <= not b;
    layer5_outputs(9798) <= a;
    layer5_outputs(9799) <= not (a and b);
    layer5_outputs(9800) <= not (a xor b);
    layer5_outputs(9801) <= not a or b;
    layer5_outputs(9802) <= b;
    layer5_outputs(9803) <= a;
    layer5_outputs(9804) <= not b;
    layer5_outputs(9805) <= a or b;
    layer5_outputs(9806) <= a;
    layer5_outputs(9807) <= a xor b;
    layer5_outputs(9808) <= not b;
    layer5_outputs(9809) <= not a;
    layer5_outputs(9810) <= a xor b;
    layer5_outputs(9811) <= not (a or b);
    layer5_outputs(9812) <= b;
    layer5_outputs(9813) <= a or b;
    layer5_outputs(9814) <= not b or a;
    layer5_outputs(9815) <= b;
    layer5_outputs(9816) <= a xor b;
    layer5_outputs(9817) <= a and not b;
    layer5_outputs(9818) <= a xor b;
    layer5_outputs(9819) <= a;
    layer5_outputs(9820) <= a xor b;
    layer5_outputs(9821) <= a and b;
    layer5_outputs(9822) <= b;
    layer5_outputs(9823) <= a or b;
    layer5_outputs(9824) <= not (a and b);
    layer5_outputs(9825) <= not b;
    layer5_outputs(9826) <= not b;
    layer5_outputs(9827) <= b;
    layer5_outputs(9828) <= a;
    layer5_outputs(9829) <= not (a xor b);
    layer5_outputs(9830) <= b;
    layer5_outputs(9831) <= not b or a;
    layer5_outputs(9832) <= a and b;
    layer5_outputs(9833) <= not (a and b);
    layer5_outputs(9834) <= not b or a;
    layer5_outputs(9835) <= '0';
    layer5_outputs(9836) <= not a;
    layer5_outputs(9837) <= a and b;
    layer5_outputs(9838) <= not a;
    layer5_outputs(9839) <= a;
    layer5_outputs(9840) <= not a;
    layer5_outputs(9841) <= not b;
    layer5_outputs(9842) <= b;
    layer5_outputs(9843) <= not a;
    layer5_outputs(9844) <= a and b;
    layer5_outputs(9845) <= not (a xor b);
    layer5_outputs(9846) <= a and not b;
    layer5_outputs(9847) <= not (a and b);
    layer5_outputs(9848) <= not b;
    layer5_outputs(9849) <= not b or a;
    layer5_outputs(9850) <= a;
    layer5_outputs(9851) <= not b or a;
    layer5_outputs(9852) <= not b;
    layer5_outputs(9853) <= not a or b;
    layer5_outputs(9854) <= a xor b;
    layer5_outputs(9855) <= a;
    layer5_outputs(9856) <= '1';
    layer5_outputs(9857) <= a;
    layer5_outputs(9858) <= a xor b;
    layer5_outputs(9859) <= not a;
    layer5_outputs(9860) <= not (a and b);
    layer5_outputs(9861) <= not (a or b);
    layer5_outputs(9862) <= not a;
    layer5_outputs(9863) <= '0';
    layer5_outputs(9864) <= a xor b;
    layer5_outputs(9865) <= not b or a;
    layer5_outputs(9866) <= b;
    layer5_outputs(9867) <= a;
    layer5_outputs(9868) <= not (a xor b);
    layer5_outputs(9869) <= a;
    layer5_outputs(9870) <= a and b;
    layer5_outputs(9871) <= not a;
    layer5_outputs(9872) <= b;
    layer5_outputs(9873) <= not (a and b);
    layer5_outputs(9874) <= not a or b;
    layer5_outputs(9875) <= not b;
    layer5_outputs(9876) <= not (a xor b);
    layer5_outputs(9877) <= a xor b;
    layer5_outputs(9878) <= not b;
    layer5_outputs(9879) <= a or b;
    layer5_outputs(9880) <= not a;
    layer5_outputs(9881) <= a or b;
    layer5_outputs(9882) <= a and not b;
    layer5_outputs(9883) <= not (a or b);
    layer5_outputs(9884) <= not b;
    layer5_outputs(9885) <= a;
    layer5_outputs(9886) <= not b;
    layer5_outputs(9887) <= not a;
    layer5_outputs(9888) <= b and not a;
    layer5_outputs(9889) <= not a or b;
    layer5_outputs(9890) <= a and b;
    layer5_outputs(9891) <= not (a xor b);
    layer5_outputs(9892) <= a and b;
    layer5_outputs(9893) <= a;
    layer5_outputs(9894) <= b;
    layer5_outputs(9895) <= a and b;
    layer5_outputs(9896) <= b;
    layer5_outputs(9897) <= b and not a;
    layer5_outputs(9898) <= not a;
    layer5_outputs(9899) <= not a;
    layer5_outputs(9900) <= not (a and b);
    layer5_outputs(9901) <= not b;
    layer5_outputs(9902) <= '0';
    layer5_outputs(9903) <= a and b;
    layer5_outputs(9904) <= not b;
    layer5_outputs(9905) <= a and b;
    layer5_outputs(9906) <= a xor b;
    layer5_outputs(9907) <= b;
    layer5_outputs(9908) <= not a;
    layer5_outputs(9909) <= a and b;
    layer5_outputs(9910) <= not b or a;
    layer5_outputs(9911) <= a and not b;
    layer5_outputs(9912) <= not a or b;
    layer5_outputs(9913) <= not b;
    layer5_outputs(9914) <= a xor b;
    layer5_outputs(9915) <= '1';
    layer5_outputs(9916) <= a and b;
    layer5_outputs(9917) <= a and b;
    layer5_outputs(9918) <= a xor b;
    layer5_outputs(9919) <= not b or a;
    layer5_outputs(9920) <= not a;
    layer5_outputs(9921) <= not b or a;
    layer5_outputs(9922) <= a or b;
    layer5_outputs(9923) <= a and b;
    layer5_outputs(9924) <= not (a xor b);
    layer5_outputs(9925) <= '0';
    layer5_outputs(9926) <= not a;
    layer5_outputs(9927) <= not (a or b);
    layer5_outputs(9928) <= a or b;
    layer5_outputs(9929) <= not b or a;
    layer5_outputs(9930) <= not (a and b);
    layer5_outputs(9931) <= b;
    layer5_outputs(9932) <= not a;
    layer5_outputs(9933) <= b and not a;
    layer5_outputs(9934) <= not a;
    layer5_outputs(9935) <= b and not a;
    layer5_outputs(9936) <= a xor b;
    layer5_outputs(9937) <= '1';
    layer5_outputs(9938) <= b;
    layer5_outputs(9939) <= b;
    layer5_outputs(9940) <= not b;
    layer5_outputs(9941) <= not (a and b);
    layer5_outputs(9942) <= not (a or b);
    layer5_outputs(9943) <= not a or b;
    layer5_outputs(9944) <= not b;
    layer5_outputs(9945) <= not a or b;
    layer5_outputs(9946) <= a and b;
    layer5_outputs(9947) <= not (a or b);
    layer5_outputs(9948) <= not (a or b);
    layer5_outputs(9949) <= a and not b;
    layer5_outputs(9950) <= not (a and b);
    layer5_outputs(9951) <= a;
    layer5_outputs(9952) <= '0';
    layer5_outputs(9953) <= not b or a;
    layer5_outputs(9954) <= not b;
    layer5_outputs(9955) <= a xor b;
    layer5_outputs(9956) <= not a;
    layer5_outputs(9957) <= a and not b;
    layer5_outputs(9958) <= a and b;
    layer5_outputs(9959) <= a or b;
    layer5_outputs(9960) <= not b;
    layer5_outputs(9961) <= a and b;
    layer5_outputs(9962) <= a;
    layer5_outputs(9963) <= not b;
    layer5_outputs(9964) <= a or b;
    layer5_outputs(9965) <= a or b;
    layer5_outputs(9966) <= a and b;
    layer5_outputs(9967) <= b;
    layer5_outputs(9968) <= a and not b;
    layer5_outputs(9969) <= b and not a;
    layer5_outputs(9970) <= a;
    layer5_outputs(9971) <= not b;
    layer5_outputs(9972) <= b;
    layer5_outputs(9973) <= a or b;
    layer5_outputs(9974) <= b;
    layer5_outputs(9975) <= a xor b;
    layer5_outputs(9976) <= a and not b;
    layer5_outputs(9977) <= a xor b;
    layer5_outputs(9978) <= '0';
    layer5_outputs(9979) <= not a;
    layer5_outputs(9980) <= b;
    layer5_outputs(9981) <= b;
    layer5_outputs(9982) <= not b;
    layer5_outputs(9983) <= b;
    layer5_outputs(9984) <= not a;
    layer5_outputs(9985) <= not b;
    layer5_outputs(9986) <= not a;
    layer5_outputs(9987) <= a and b;
    layer5_outputs(9988) <= b;
    layer5_outputs(9989) <= '1';
    layer5_outputs(9990) <= b;
    layer5_outputs(9991) <= a and b;
    layer5_outputs(9992) <= not a;
    layer5_outputs(9993) <= not b or a;
    layer5_outputs(9994) <= not (a and b);
    layer5_outputs(9995) <= a or b;
    layer5_outputs(9996) <= not b or a;
    layer5_outputs(9997) <= not a;
    layer5_outputs(9998) <= not b;
    layer5_outputs(9999) <= b;
    layer5_outputs(10000) <= a;
    layer5_outputs(10001) <= not a;
    layer5_outputs(10002) <= b;
    layer5_outputs(10003) <= b;
    layer5_outputs(10004) <= b and not a;
    layer5_outputs(10005) <= not (a and b);
    layer5_outputs(10006) <= not a;
    layer5_outputs(10007) <= not b;
    layer5_outputs(10008) <= a or b;
    layer5_outputs(10009) <= not b;
    layer5_outputs(10010) <= not a or b;
    layer5_outputs(10011) <= b;
    layer5_outputs(10012) <= not a;
    layer5_outputs(10013) <= not (a xor b);
    layer5_outputs(10014) <= not (a and b);
    layer5_outputs(10015) <= a or b;
    layer5_outputs(10016) <= not a;
    layer5_outputs(10017) <= not (a and b);
    layer5_outputs(10018) <= not a;
    layer5_outputs(10019) <= not b;
    layer5_outputs(10020) <= b and not a;
    layer5_outputs(10021) <= not b;
    layer5_outputs(10022) <= not (a and b);
    layer5_outputs(10023) <= not (a or b);
    layer5_outputs(10024) <= b;
    layer5_outputs(10025) <= not b or a;
    layer5_outputs(10026) <= a or b;
    layer5_outputs(10027) <= not b;
    layer5_outputs(10028) <= a;
    layer5_outputs(10029) <= not (a xor b);
    layer5_outputs(10030) <= not a or b;
    layer5_outputs(10031) <= not b;
    layer5_outputs(10032) <= not (a xor b);
    layer5_outputs(10033) <= b;
    layer5_outputs(10034) <= not a;
    layer5_outputs(10035) <= a;
    layer5_outputs(10036) <= b and not a;
    layer5_outputs(10037) <= not (a xor b);
    layer5_outputs(10038) <= b;
    layer5_outputs(10039) <= not b;
    layer5_outputs(10040) <= not b or a;
    layer5_outputs(10041) <= '0';
    layer5_outputs(10042) <= a;
    layer5_outputs(10043) <= a;
    layer5_outputs(10044) <= not (a xor b);
    layer5_outputs(10045) <= not b;
    layer5_outputs(10046) <= not a or b;
    layer5_outputs(10047) <= not (a xor b);
    layer5_outputs(10048) <= not a or b;
    layer5_outputs(10049) <= b;
    layer5_outputs(10050) <= a;
    layer5_outputs(10051) <= not a;
    layer5_outputs(10052) <= not (a xor b);
    layer5_outputs(10053) <= a or b;
    layer5_outputs(10054) <= a and b;
    layer5_outputs(10055) <= not a;
    layer5_outputs(10056) <= a;
    layer5_outputs(10057) <= a and not b;
    layer5_outputs(10058) <= a;
    layer5_outputs(10059) <= not b;
    layer5_outputs(10060) <= not a;
    layer5_outputs(10061) <= a xor b;
    layer5_outputs(10062) <= a and b;
    layer5_outputs(10063) <= b;
    layer5_outputs(10064) <= a xor b;
    layer5_outputs(10065) <= a;
    layer5_outputs(10066) <= b;
    layer5_outputs(10067) <= b;
    layer5_outputs(10068) <= not a;
    layer5_outputs(10069) <= b;
    layer5_outputs(10070) <= a and not b;
    layer5_outputs(10071) <= not (a or b);
    layer5_outputs(10072) <= not b;
    layer5_outputs(10073) <= a or b;
    layer5_outputs(10074) <= not a;
    layer5_outputs(10075) <= a;
    layer5_outputs(10076) <= a xor b;
    layer5_outputs(10077) <= not (a xor b);
    layer5_outputs(10078) <= a and b;
    layer5_outputs(10079) <= a and not b;
    layer5_outputs(10080) <= b;
    layer5_outputs(10081) <= b;
    layer5_outputs(10082) <= a and not b;
    layer5_outputs(10083) <= not (a xor b);
    layer5_outputs(10084) <= a;
    layer5_outputs(10085) <= not (a and b);
    layer5_outputs(10086) <= not b;
    layer5_outputs(10087) <= not a or b;
    layer5_outputs(10088) <= a and not b;
    layer5_outputs(10089) <= not (a and b);
    layer5_outputs(10090) <= not a;
    layer5_outputs(10091) <= a and b;
    layer5_outputs(10092) <= a;
    layer5_outputs(10093) <= not (a or b);
    layer5_outputs(10094) <= a and not b;
    layer5_outputs(10095) <= not (a and b);
    layer5_outputs(10096) <= not a or b;
    layer5_outputs(10097) <= '0';
    layer5_outputs(10098) <= not b or a;
    layer5_outputs(10099) <= not (a or b);
    layer5_outputs(10100) <= not (a and b);
    layer5_outputs(10101) <= not a;
    layer5_outputs(10102) <= a;
    layer5_outputs(10103) <= not a;
    layer5_outputs(10104) <= a and not b;
    layer5_outputs(10105) <= not b;
    layer5_outputs(10106) <= not (a xor b);
    layer5_outputs(10107) <= not a;
    layer5_outputs(10108) <= not a;
    layer5_outputs(10109) <= not a;
    layer5_outputs(10110) <= not b;
    layer5_outputs(10111) <= not a;
    layer5_outputs(10112) <= b;
    layer5_outputs(10113) <= not a or b;
    layer5_outputs(10114) <= not a;
    layer5_outputs(10115) <= not b or a;
    layer5_outputs(10116) <= not b or a;
    layer5_outputs(10117) <= not b or a;
    layer5_outputs(10118) <= a and b;
    layer5_outputs(10119) <= not a;
    layer5_outputs(10120) <= not a or b;
    layer5_outputs(10121) <= not a;
    layer5_outputs(10122) <= a and b;
    layer5_outputs(10123) <= b;
    layer5_outputs(10124) <= not (a or b);
    layer5_outputs(10125) <= not (a or b);
    layer5_outputs(10126) <= not (a and b);
    layer5_outputs(10127) <= a or b;
    layer5_outputs(10128) <= a;
    layer5_outputs(10129) <= not (a xor b);
    layer5_outputs(10130) <= not a;
    layer5_outputs(10131) <= not (a or b);
    layer5_outputs(10132) <= a;
    layer5_outputs(10133) <= not b or a;
    layer5_outputs(10134) <= not (a xor b);
    layer5_outputs(10135) <= not a;
    layer5_outputs(10136) <= a;
    layer5_outputs(10137) <= b;
    layer5_outputs(10138) <= not b;
    layer5_outputs(10139) <= not b;
    layer5_outputs(10140) <= not (a xor b);
    layer5_outputs(10141) <= not a;
    layer5_outputs(10142) <= not a;
    layer5_outputs(10143) <= not a;
    layer5_outputs(10144) <= a and b;
    layer5_outputs(10145) <= b;
    layer5_outputs(10146) <= a;
    layer5_outputs(10147) <= not b;
    layer5_outputs(10148) <= b and not a;
    layer5_outputs(10149) <= not b;
    layer5_outputs(10150) <= not b or a;
    layer5_outputs(10151) <= not b or a;
    layer5_outputs(10152) <= a and b;
    layer5_outputs(10153) <= b;
    layer5_outputs(10154) <= a and not b;
    layer5_outputs(10155) <= not (a or b);
    layer5_outputs(10156) <= b;
    layer5_outputs(10157) <= not b or a;
    layer5_outputs(10158) <= not a;
    layer5_outputs(10159) <= a;
    layer5_outputs(10160) <= not (a xor b);
    layer5_outputs(10161) <= b;
    layer5_outputs(10162) <= b and not a;
    layer5_outputs(10163) <= a xor b;
    layer5_outputs(10164) <= a and b;
    layer5_outputs(10165) <= a;
    layer5_outputs(10166) <= b;
    layer5_outputs(10167) <= not a or b;
    layer5_outputs(10168) <= a or b;
    layer5_outputs(10169) <= a;
    layer5_outputs(10170) <= not a;
    layer5_outputs(10171) <= not a;
    layer5_outputs(10172) <= not b;
    layer5_outputs(10173) <= a;
    layer5_outputs(10174) <= b;
    layer5_outputs(10175) <= b;
    layer5_outputs(10176) <= a and b;
    layer5_outputs(10177) <= b and not a;
    layer5_outputs(10178) <= b;
    layer5_outputs(10179) <= not b;
    layer5_outputs(10180) <= b;
    layer5_outputs(10181) <= a;
    layer5_outputs(10182) <= not b;
    layer5_outputs(10183) <= b;
    layer5_outputs(10184) <= not a or b;
    layer5_outputs(10185) <= not (a or b);
    layer5_outputs(10186) <= b and not a;
    layer5_outputs(10187) <= a and b;
    layer5_outputs(10188) <= a;
    layer5_outputs(10189) <= a;
    layer5_outputs(10190) <= not (a or b);
    layer5_outputs(10191) <= not b;
    layer5_outputs(10192) <= b;
    layer5_outputs(10193) <= not a;
    layer5_outputs(10194) <= not a or b;
    layer5_outputs(10195) <= a xor b;
    layer5_outputs(10196) <= '1';
    layer5_outputs(10197) <= not (a or b);
    layer5_outputs(10198) <= a and not b;
    layer5_outputs(10199) <= b and not a;
    layer5_outputs(10200) <= a xor b;
    layer5_outputs(10201) <= not a;
    layer5_outputs(10202) <= a xor b;
    layer5_outputs(10203) <= not b or a;
    layer5_outputs(10204) <= '0';
    layer5_outputs(10205) <= a xor b;
    layer5_outputs(10206) <= not a or b;
    layer5_outputs(10207) <= a;
    layer5_outputs(10208) <= not b;
    layer5_outputs(10209) <= b;
    layer5_outputs(10210) <= a and not b;
    layer5_outputs(10211) <= b;
    layer5_outputs(10212) <= a xor b;
    layer5_outputs(10213) <= not b or a;
    layer5_outputs(10214) <= not a;
    layer5_outputs(10215) <= not a;
    layer5_outputs(10216) <= a;
    layer5_outputs(10217) <= not (a or b);
    layer5_outputs(10218) <= not a;
    layer5_outputs(10219) <= not (a xor b);
    layer5_outputs(10220) <= not b;
    layer5_outputs(10221) <= not (a or b);
    layer5_outputs(10222) <= a and not b;
    layer5_outputs(10223) <= b;
    layer5_outputs(10224) <= a and not b;
    layer5_outputs(10225) <= not b or a;
    layer5_outputs(10226) <= a;
    layer5_outputs(10227) <= not (a and b);
    layer5_outputs(10228) <= not a;
    layer5_outputs(10229) <= not b;
    layer5_outputs(10230) <= a;
    layer5_outputs(10231) <= not a;
    layer5_outputs(10232) <= a xor b;
    layer5_outputs(10233) <= b;
    layer5_outputs(10234) <= a;
    layer5_outputs(10235) <= b and not a;
    layer5_outputs(10236) <= a and not b;
    layer5_outputs(10237) <= not a;
    layer5_outputs(10238) <= a xor b;
    layer5_outputs(10239) <= a;
    layer6_outputs(0) <= not b;
    layer6_outputs(1) <= a and b;
    layer6_outputs(2) <= not b;
    layer6_outputs(3) <= not a;
    layer6_outputs(4) <= a;
    layer6_outputs(5) <= b;
    layer6_outputs(6) <= a xor b;
    layer6_outputs(7) <= a xor b;
    layer6_outputs(8) <= a and not b;
    layer6_outputs(9) <= not (a xor b);
    layer6_outputs(10) <= not b;
    layer6_outputs(11) <= b;
    layer6_outputs(12) <= a and not b;
    layer6_outputs(13) <= a and not b;
    layer6_outputs(14) <= a;
    layer6_outputs(15) <= not b;
    layer6_outputs(16) <= not b;
    layer6_outputs(17) <= not (a and b);
    layer6_outputs(18) <= not (a xor b);
    layer6_outputs(19) <= not b or a;
    layer6_outputs(20) <= a;
    layer6_outputs(21) <= not b;
    layer6_outputs(22) <= b;
    layer6_outputs(23) <= not (a xor b);
    layer6_outputs(24) <= not a;
    layer6_outputs(25) <= not b;
    layer6_outputs(26) <= not a;
    layer6_outputs(27) <= not a;
    layer6_outputs(28) <= b;
    layer6_outputs(29) <= not a;
    layer6_outputs(30) <= b and not a;
    layer6_outputs(31) <= not b;
    layer6_outputs(32) <= a xor b;
    layer6_outputs(33) <= a xor b;
    layer6_outputs(34) <= a;
    layer6_outputs(35) <= a;
    layer6_outputs(36) <= not a;
    layer6_outputs(37) <= not a;
    layer6_outputs(38) <= a;
    layer6_outputs(39) <= not (a xor b);
    layer6_outputs(40) <= a or b;
    layer6_outputs(41) <= a;
    layer6_outputs(42) <= not a;
    layer6_outputs(43) <= not a or b;
    layer6_outputs(44) <= not a;
    layer6_outputs(45) <= not (a xor b);
    layer6_outputs(46) <= not b;
    layer6_outputs(47) <= a;
    layer6_outputs(48) <= a;
    layer6_outputs(49) <= not b;
    layer6_outputs(50) <= a and not b;
    layer6_outputs(51) <= b;
    layer6_outputs(52) <= a xor b;
    layer6_outputs(53) <= not a;
    layer6_outputs(54) <= a xor b;
    layer6_outputs(55) <= b;
    layer6_outputs(56) <= '0';
    layer6_outputs(57) <= not b;
    layer6_outputs(58) <= a;
    layer6_outputs(59) <= not b;
    layer6_outputs(60) <= a or b;
    layer6_outputs(61) <= not (a or b);
    layer6_outputs(62) <= b;
    layer6_outputs(63) <= a or b;
    layer6_outputs(64) <= a xor b;
    layer6_outputs(65) <= b;
    layer6_outputs(66) <= not a;
    layer6_outputs(67) <= b and not a;
    layer6_outputs(68) <= a and not b;
    layer6_outputs(69) <= b;
    layer6_outputs(70) <= not (a or b);
    layer6_outputs(71) <= not (a or b);
    layer6_outputs(72) <= not b;
    layer6_outputs(73) <= not b;
    layer6_outputs(74) <= a xor b;
    layer6_outputs(75) <= b;
    layer6_outputs(76) <= not a;
    layer6_outputs(77) <= not a or b;
    layer6_outputs(78) <= a;
    layer6_outputs(79) <= not (a xor b);
    layer6_outputs(80) <= b;
    layer6_outputs(81) <= not (a and b);
    layer6_outputs(82) <= not a;
    layer6_outputs(83) <= not a;
    layer6_outputs(84) <= a;
    layer6_outputs(85) <= b;
    layer6_outputs(86) <= not a;
    layer6_outputs(87) <= a and not b;
    layer6_outputs(88) <= not b;
    layer6_outputs(89) <= a;
    layer6_outputs(90) <= a and b;
    layer6_outputs(91) <= b;
    layer6_outputs(92) <= not b;
    layer6_outputs(93) <= not a;
    layer6_outputs(94) <= not a;
    layer6_outputs(95) <= b;
    layer6_outputs(96) <= a;
    layer6_outputs(97) <= a;
    layer6_outputs(98) <= a xor b;
    layer6_outputs(99) <= not b;
    layer6_outputs(100) <= not (a and b);
    layer6_outputs(101) <= not b;
    layer6_outputs(102) <= b;
    layer6_outputs(103) <= not b;
    layer6_outputs(104) <= not (a or b);
    layer6_outputs(105) <= not b;
    layer6_outputs(106) <= b;
    layer6_outputs(107) <= not (a xor b);
    layer6_outputs(108) <= a;
    layer6_outputs(109) <= not b;
    layer6_outputs(110) <= a;
    layer6_outputs(111) <= a and not b;
    layer6_outputs(112) <= not (a xor b);
    layer6_outputs(113) <= b;
    layer6_outputs(114) <= not (a xor b);
    layer6_outputs(115) <= a;
    layer6_outputs(116) <= a xor b;
    layer6_outputs(117) <= a and not b;
    layer6_outputs(118) <= b;
    layer6_outputs(119) <= a or b;
    layer6_outputs(120) <= a or b;
    layer6_outputs(121) <= not a;
    layer6_outputs(122) <= not a;
    layer6_outputs(123) <= a;
    layer6_outputs(124) <= a xor b;
    layer6_outputs(125) <= not a;
    layer6_outputs(126) <= a;
    layer6_outputs(127) <= not b or a;
    layer6_outputs(128) <= not a or b;
    layer6_outputs(129) <= a and not b;
    layer6_outputs(130) <= not (a xor b);
    layer6_outputs(131) <= a;
    layer6_outputs(132) <= not (a xor b);
    layer6_outputs(133) <= a and not b;
    layer6_outputs(134) <= not a or b;
    layer6_outputs(135) <= a and b;
    layer6_outputs(136) <= not a;
    layer6_outputs(137) <= not (a or b);
    layer6_outputs(138) <= a and not b;
    layer6_outputs(139) <= not a or b;
    layer6_outputs(140) <= not (a xor b);
    layer6_outputs(141) <= a or b;
    layer6_outputs(142) <= not b;
    layer6_outputs(143) <= b;
    layer6_outputs(144) <= b and not a;
    layer6_outputs(145) <= b;
    layer6_outputs(146) <= a and b;
    layer6_outputs(147) <= not (a xor b);
    layer6_outputs(148) <= not b;
    layer6_outputs(149) <= not b or a;
    layer6_outputs(150) <= not a;
    layer6_outputs(151) <= not b;
    layer6_outputs(152) <= not b;
    layer6_outputs(153) <= not b;
    layer6_outputs(154) <= a or b;
    layer6_outputs(155) <= a and b;
    layer6_outputs(156) <= a and not b;
    layer6_outputs(157) <= not a or b;
    layer6_outputs(158) <= '1';
    layer6_outputs(159) <= b and not a;
    layer6_outputs(160) <= not (a xor b);
    layer6_outputs(161) <= not b or a;
    layer6_outputs(162) <= not (a xor b);
    layer6_outputs(163) <= a and not b;
    layer6_outputs(164) <= a;
    layer6_outputs(165) <= a or b;
    layer6_outputs(166) <= not b;
    layer6_outputs(167) <= not b or a;
    layer6_outputs(168) <= not (a xor b);
    layer6_outputs(169) <= not (a or b);
    layer6_outputs(170) <= a or b;
    layer6_outputs(171) <= a and b;
    layer6_outputs(172) <= not (a xor b);
    layer6_outputs(173) <= a and not b;
    layer6_outputs(174) <= not a or b;
    layer6_outputs(175) <= a and b;
    layer6_outputs(176) <= a and b;
    layer6_outputs(177) <= a and b;
    layer6_outputs(178) <= a;
    layer6_outputs(179) <= a;
    layer6_outputs(180) <= not a;
    layer6_outputs(181) <= b and not a;
    layer6_outputs(182) <= not a;
    layer6_outputs(183) <= not b or a;
    layer6_outputs(184) <= a and b;
    layer6_outputs(185) <= a xor b;
    layer6_outputs(186) <= not a;
    layer6_outputs(187) <= b;
    layer6_outputs(188) <= a and not b;
    layer6_outputs(189) <= not (a xor b);
    layer6_outputs(190) <= a xor b;
    layer6_outputs(191) <= not a or b;
    layer6_outputs(192) <= not a or b;
    layer6_outputs(193) <= not a or b;
    layer6_outputs(194) <= not b;
    layer6_outputs(195) <= a xor b;
    layer6_outputs(196) <= a xor b;
    layer6_outputs(197) <= a;
    layer6_outputs(198) <= a and not b;
    layer6_outputs(199) <= not (a or b);
    layer6_outputs(200) <= a;
    layer6_outputs(201) <= b and not a;
    layer6_outputs(202) <= a;
    layer6_outputs(203) <= not (a and b);
    layer6_outputs(204) <= not b;
    layer6_outputs(205) <= not (a and b);
    layer6_outputs(206) <= b and not a;
    layer6_outputs(207) <= a and b;
    layer6_outputs(208) <= not b;
    layer6_outputs(209) <= not (a and b);
    layer6_outputs(210) <= a xor b;
    layer6_outputs(211) <= a or b;
    layer6_outputs(212) <= a xor b;
    layer6_outputs(213) <= a or b;
    layer6_outputs(214) <= a and b;
    layer6_outputs(215) <= not b;
    layer6_outputs(216) <= a;
    layer6_outputs(217) <= a xor b;
    layer6_outputs(218) <= not a;
    layer6_outputs(219) <= b and not a;
    layer6_outputs(220) <= b;
    layer6_outputs(221) <= not b or a;
    layer6_outputs(222) <= a xor b;
    layer6_outputs(223) <= b;
    layer6_outputs(224) <= a or b;
    layer6_outputs(225) <= not b;
    layer6_outputs(226) <= not (a xor b);
    layer6_outputs(227) <= a xor b;
    layer6_outputs(228) <= not a;
    layer6_outputs(229) <= a;
    layer6_outputs(230) <= b and not a;
    layer6_outputs(231) <= not (a and b);
    layer6_outputs(232) <= a;
    layer6_outputs(233) <= a xor b;
    layer6_outputs(234) <= a;
    layer6_outputs(235) <= not b or a;
    layer6_outputs(236) <= a;
    layer6_outputs(237) <= a xor b;
    layer6_outputs(238) <= b;
    layer6_outputs(239) <= not b;
    layer6_outputs(240) <= a and not b;
    layer6_outputs(241) <= b;
    layer6_outputs(242) <= not (a or b);
    layer6_outputs(243) <= not (a xor b);
    layer6_outputs(244) <= not b;
    layer6_outputs(245) <= not (a or b);
    layer6_outputs(246) <= a and not b;
    layer6_outputs(247) <= not (a xor b);
    layer6_outputs(248) <= b and not a;
    layer6_outputs(249) <= a and not b;
    layer6_outputs(250) <= a and not b;
    layer6_outputs(251) <= a and b;
    layer6_outputs(252) <= not b or a;
    layer6_outputs(253) <= not a;
    layer6_outputs(254) <= a;
    layer6_outputs(255) <= not a or b;
    layer6_outputs(256) <= b;
    layer6_outputs(257) <= not (a xor b);
    layer6_outputs(258) <= not a;
    layer6_outputs(259) <= not a;
    layer6_outputs(260) <= b;
    layer6_outputs(261) <= b;
    layer6_outputs(262) <= a and not b;
    layer6_outputs(263) <= not a or b;
    layer6_outputs(264) <= a;
    layer6_outputs(265) <= not a;
    layer6_outputs(266) <= not b;
    layer6_outputs(267) <= not a;
    layer6_outputs(268) <= a xor b;
    layer6_outputs(269) <= not a;
    layer6_outputs(270) <= a or b;
    layer6_outputs(271) <= not a;
    layer6_outputs(272) <= a and not b;
    layer6_outputs(273) <= not b or a;
    layer6_outputs(274) <= a or b;
    layer6_outputs(275) <= a and not b;
    layer6_outputs(276) <= a or b;
    layer6_outputs(277) <= a;
    layer6_outputs(278) <= a xor b;
    layer6_outputs(279) <= b;
    layer6_outputs(280) <= a;
    layer6_outputs(281) <= b;
    layer6_outputs(282) <= a;
    layer6_outputs(283) <= not b or a;
    layer6_outputs(284) <= a;
    layer6_outputs(285) <= a or b;
    layer6_outputs(286) <= not (a and b);
    layer6_outputs(287) <= b;
    layer6_outputs(288) <= b;
    layer6_outputs(289) <= not (a xor b);
    layer6_outputs(290) <= a;
    layer6_outputs(291) <= not b;
    layer6_outputs(292) <= a;
    layer6_outputs(293) <= not a or b;
    layer6_outputs(294) <= not (a and b);
    layer6_outputs(295) <= b;
    layer6_outputs(296) <= a or b;
    layer6_outputs(297) <= a;
    layer6_outputs(298) <= b and not a;
    layer6_outputs(299) <= not (a xor b);
    layer6_outputs(300) <= not (a and b);
    layer6_outputs(301) <= '1';
    layer6_outputs(302) <= not b;
    layer6_outputs(303) <= not a;
    layer6_outputs(304) <= not (a and b);
    layer6_outputs(305) <= not a;
    layer6_outputs(306) <= a or b;
    layer6_outputs(307) <= not a;
    layer6_outputs(308) <= a;
    layer6_outputs(309) <= b;
    layer6_outputs(310) <= not b;
    layer6_outputs(311) <= not (a xor b);
    layer6_outputs(312) <= b;
    layer6_outputs(313) <= a xor b;
    layer6_outputs(314) <= not a;
    layer6_outputs(315) <= not a;
    layer6_outputs(316) <= a xor b;
    layer6_outputs(317) <= not b;
    layer6_outputs(318) <= a xor b;
    layer6_outputs(319) <= not (a xor b);
    layer6_outputs(320) <= a and not b;
    layer6_outputs(321) <= not a or b;
    layer6_outputs(322) <= a;
    layer6_outputs(323) <= b;
    layer6_outputs(324) <= b and not a;
    layer6_outputs(325) <= b and not a;
    layer6_outputs(326) <= not (a xor b);
    layer6_outputs(327) <= not (a xor b);
    layer6_outputs(328) <= a xor b;
    layer6_outputs(329) <= not b;
    layer6_outputs(330) <= a;
    layer6_outputs(331) <= not (a xor b);
    layer6_outputs(332) <= not b or a;
    layer6_outputs(333) <= b and not a;
    layer6_outputs(334) <= not (a or b);
    layer6_outputs(335) <= b;
    layer6_outputs(336) <= not a;
    layer6_outputs(337) <= not b;
    layer6_outputs(338) <= a and not b;
    layer6_outputs(339) <= not b;
    layer6_outputs(340) <= a;
    layer6_outputs(341) <= not (a xor b);
    layer6_outputs(342) <= a and b;
    layer6_outputs(343) <= not a or b;
    layer6_outputs(344) <= a and not b;
    layer6_outputs(345) <= a or b;
    layer6_outputs(346) <= not (a or b);
    layer6_outputs(347) <= a;
    layer6_outputs(348) <= not (a or b);
    layer6_outputs(349) <= not a;
    layer6_outputs(350) <= not (a xor b);
    layer6_outputs(351) <= a xor b;
    layer6_outputs(352) <= not a or b;
    layer6_outputs(353) <= b;
    layer6_outputs(354) <= a;
    layer6_outputs(355) <= not a;
    layer6_outputs(356) <= a;
    layer6_outputs(357) <= a xor b;
    layer6_outputs(358) <= not (a xor b);
    layer6_outputs(359) <= not a;
    layer6_outputs(360) <= a xor b;
    layer6_outputs(361) <= a;
    layer6_outputs(362) <= b;
    layer6_outputs(363) <= a or b;
    layer6_outputs(364) <= not a or b;
    layer6_outputs(365) <= b;
    layer6_outputs(366) <= not b;
    layer6_outputs(367) <= a xor b;
    layer6_outputs(368) <= a and b;
    layer6_outputs(369) <= not b or a;
    layer6_outputs(370) <= not (a xor b);
    layer6_outputs(371) <= b;
    layer6_outputs(372) <= a and b;
    layer6_outputs(373) <= a and b;
    layer6_outputs(374) <= a;
    layer6_outputs(375) <= b and not a;
    layer6_outputs(376) <= not a;
    layer6_outputs(377) <= a;
    layer6_outputs(378) <= b;
    layer6_outputs(379) <= a xor b;
    layer6_outputs(380) <= a;
    layer6_outputs(381) <= a or b;
    layer6_outputs(382) <= a;
    layer6_outputs(383) <= a or b;
    layer6_outputs(384) <= b;
    layer6_outputs(385) <= b and not a;
    layer6_outputs(386) <= not a;
    layer6_outputs(387) <= not (a xor b);
    layer6_outputs(388) <= not (a xor b);
    layer6_outputs(389) <= not (a or b);
    layer6_outputs(390) <= a;
    layer6_outputs(391) <= a;
    layer6_outputs(392) <= not a or b;
    layer6_outputs(393) <= '1';
    layer6_outputs(394) <= a and b;
    layer6_outputs(395) <= not b;
    layer6_outputs(396) <= not (a or b);
    layer6_outputs(397) <= a or b;
    layer6_outputs(398) <= a and not b;
    layer6_outputs(399) <= not a;
    layer6_outputs(400) <= not b;
    layer6_outputs(401) <= a or b;
    layer6_outputs(402) <= not (a xor b);
    layer6_outputs(403) <= a;
    layer6_outputs(404) <= b and not a;
    layer6_outputs(405) <= not (a xor b);
    layer6_outputs(406) <= a or b;
    layer6_outputs(407) <= a;
    layer6_outputs(408) <= not (a xor b);
    layer6_outputs(409) <= a or b;
    layer6_outputs(410) <= a xor b;
    layer6_outputs(411) <= not b;
    layer6_outputs(412) <= a or b;
    layer6_outputs(413) <= not (a xor b);
    layer6_outputs(414) <= not (a or b);
    layer6_outputs(415) <= not a;
    layer6_outputs(416) <= a and not b;
    layer6_outputs(417) <= a or b;
    layer6_outputs(418) <= not (a or b);
    layer6_outputs(419) <= a and b;
    layer6_outputs(420) <= a;
    layer6_outputs(421) <= not (a or b);
    layer6_outputs(422) <= not b or a;
    layer6_outputs(423) <= not (a and b);
    layer6_outputs(424) <= a xor b;
    layer6_outputs(425) <= not b;
    layer6_outputs(426) <= b and not a;
    layer6_outputs(427) <= a xor b;
    layer6_outputs(428) <= not (a or b);
    layer6_outputs(429) <= a xor b;
    layer6_outputs(430) <= not a or b;
    layer6_outputs(431) <= '1';
    layer6_outputs(432) <= not a;
    layer6_outputs(433) <= b and not a;
    layer6_outputs(434) <= not a;
    layer6_outputs(435) <= not a;
    layer6_outputs(436) <= not (a or b);
    layer6_outputs(437) <= not b;
    layer6_outputs(438) <= not (a xor b);
    layer6_outputs(439) <= b;
    layer6_outputs(440) <= a;
    layer6_outputs(441) <= b;
    layer6_outputs(442) <= not a;
    layer6_outputs(443) <= not (a and b);
    layer6_outputs(444) <= not (a and b);
    layer6_outputs(445) <= b;
    layer6_outputs(446) <= a;
    layer6_outputs(447) <= a;
    layer6_outputs(448) <= a and b;
    layer6_outputs(449) <= a and b;
    layer6_outputs(450) <= b and not a;
    layer6_outputs(451) <= not b;
    layer6_outputs(452) <= a;
    layer6_outputs(453) <= b;
    layer6_outputs(454) <= a xor b;
    layer6_outputs(455) <= a xor b;
    layer6_outputs(456) <= not (a xor b);
    layer6_outputs(457) <= b;
    layer6_outputs(458) <= not a;
    layer6_outputs(459) <= not a;
    layer6_outputs(460) <= not b;
    layer6_outputs(461) <= not (a xor b);
    layer6_outputs(462) <= a;
    layer6_outputs(463) <= not a;
    layer6_outputs(464) <= a or b;
    layer6_outputs(465) <= not (a or b);
    layer6_outputs(466) <= b and not a;
    layer6_outputs(467) <= not b or a;
    layer6_outputs(468) <= not a;
    layer6_outputs(469) <= not b;
    layer6_outputs(470) <= a;
    layer6_outputs(471) <= not b;
    layer6_outputs(472) <= not (a xor b);
    layer6_outputs(473) <= b;
    layer6_outputs(474) <= b;
    layer6_outputs(475) <= '0';
    layer6_outputs(476) <= not (a xor b);
    layer6_outputs(477) <= a xor b;
    layer6_outputs(478) <= not (a and b);
    layer6_outputs(479) <= not b;
    layer6_outputs(480) <= not a;
    layer6_outputs(481) <= not b or a;
    layer6_outputs(482) <= not b;
    layer6_outputs(483) <= a;
    layer6_outputs(484) <= not (a or b);
    layer6_outputs(485) <= not (a or b);
    layer6_outputs(486) <= a or b;
    layer6_outputs(487) <= not (a xor b);
    layer6_outputs(488) <= not b;
    layer6_outputs(489) <= a or b;
    layer6_outputs(490) <= a and b;
    layer6_outputs(491) <= a xor b;
    layer6_outputs(492) <= not b;
    layer6_outputs(493) <= not (a and b);
    layer6_outputs(494) <= b and not a;
    layer6_outputs(495) <= not a or b;
    layer6_outputs(496) <= not a;
    layer6_outputs(497) <= not b;
    layer6_outputs(498) <= a or b;
    layer6_outputs(499) <= not b or a;
    layer6_outputs(500) <= not b;
    layer6_outputs(501) <= not (a and b);
    layer6_outputs(502) <= '0';
    layer6_outputs(503) <= a or b;
    layer6_outputs(504) <= not (a and b);
    layer6_outputs(505) <= b;
    layer6_outputs(506) <= a and b;
    layer6_outputs(507) <= not b;
    layer6_outputs(508) <= b;
    layer6_outputs(509) <= '0';
    layer6_outputs(510) <= b;
    layer6_outputs(511) <= a;
    layer6_outputs(512) <= b;
    layer6_outputs(513) <= not (a xor b);
    layer6_outputs(514) <= not (a or b);
    layer6_outputs(515) <= not (a and b);
    layer6_outputs(516) <= not a;
    layer6_outputs(517) <= not (a or b);
    layer6_outputs(518) <= a;
    layer6_outputs(519) <= '1';
    layer6_outputs(520) <= not (a and b);
    layer6_outputs(521) <= a;
    layer6_outputs(522) <= a and not b;
    layer6_outputs(523) <= not (a and b);
    layer6_outputs(524) <= a xor b;
    layer6_outputs(525) <= not (a and b);
    layer6_outputs(526) <= a;
    layer6_outputs(527) <= not b or a;
    layer6_outputs(528) <= a and b;
    layer6_outputs(529) <= a;
    layer6_outputs(530) <= not b;
    layer6_outputs(531) <= not (a xor b);
    layer6_outputs(532) <= not (a xor b);
    layer6_outputs(533) <= not a;
    layer6_outputs(534) <= not b;
    layer6_outputs(535) <= not b;
    layer6_outputs(536) <= a and b;
    layer6_outputs(537) <= not (a and b);
    layer6_outputs(538) <= a;
    layer6_outputs(539) <= a;
    layer6_outputs(540) <= a and b;
    layer6_outputs(541) <= a xor b;
    layer6_outputs(542) <= not (a or b);
    layer6_outputs(543) <= not a;
    layer6_outputs(544) <= a;
    layer6_outputs(545) <= not b;
    layer6_outputs(546) <= a;
    layer6_outputs(547) <= not a;
    layer6_outputs(548) <= not b;
    layer6_outputs(549) <= b;
    layer6_outputs(550) <= not a or b;
    layer6_outputs(551) <= not (a xor b);
    layer6_outputs(552) <= not b;
    layer6_outputs(553) <= not (a xor b);
    layer6_outputs(554) <= not (a xor b);
    layer6_outputs(555) <= not (a xor b);
    layer6_outputs(556) <= not (a or b);
    layer6_outputs(557) <= not (a or b);
    layer6_outputs(558) <= b and not a;
    layer6_outputs(559) <= not a;
    layer6_outputs(560) <= a;
    layer6_outputs(561) <= not (a xor b);
    layer6_outputs(562) <= not b;
    layer6_outputs(563) <= a xor b;
    layer6_outputs(564) <= a xor b;
    layer6_outputs(565) <= not a;
    layer6_outputs(566) <= a xor b;
    layer6_outputs(567) <= not (a and b);
    layer6_outputs(568) <= not b or a;
    layer6_outputs(569) <= not b;
    layer6_outputs(570) <= a and b;
    layer6_outputs(571) <= b;
    layer6_outputs(572) <= not (a and b);
    layer6_outputs(573) <= a;
    layer6_outputs(574) <= not a;
    layer6_outputs(575) <= not (a or b);
    layer6_outputs(576) <= a and not b;
    layer6_outputs(577) <= not b;
    layer6_outputs(578) <= b;
    layer6_outputs(579) <= a;
    layer6_outputs(580) <= not b;
    layer6_outputs(581) <= not (a and b);
    layer6_outputs(582) <= not (a xor b);
    layer6_outputs(583) <= b;
    layer6_outputs(584) <= not (a and b);
    layer6_outputs(585) <= a or b;
    layer6_outputs(586) <= not b;
    layer6_outputs(587) <= not a;
    layer6_outputs(588) <= not (a xor b);
    layer6_outputs(589) <= not a or b;
    layer6_outputs(590) <= a;
    layer6_outputs(591) <= a or b;
    layer6_outputs(592) <= b;
    layer6_outputs(593) <= not b;
    layer6_outputs(594) <= b;
    layer6_outputs(595) <= not a;
    layer6_outputs(596) <= not b or a;
    layer6_outputs(597) <= not b;
    layer6_outputs(598) <= b;
    layer6_outputs(599) <= b;
    layer6_outputs(600) <= not (a xor b);
    layer6_outputs(601) <= a;
    layer6_outputs(602) <= a xor b;
    layer6_outputs(603) <= b;
    layer6_outputs(604) <= b and not a;
    layer6_outputs(605) <= not b;
    layer6_outputs(606) <= b and not a;
    layer6_outputs(607) <= b;
    layer6_outputs(608) <= a and not b;
    layer6_outputs(609) <= not (a and b);
    layer6_outputs(610) <= not b;
    layer6_outputs(611) <= not a;
    layer6_outputs(612) <= a and not b;
    layer6_outputs(613) <= a or b;
    layer6_outputs(614) <= b and not a;
    layer6_outputs(615) <= not b;
    layer6_outputs(616) <= not a;
    layer6_outputs(617) <= not a;
    layer6_outputs(618) <= not (a or b);
    layer6_outputs(619) <= not b;
    layer6_outputs(620) <= not b;
    layer6_outputs(621) <= a;
    layer6_outputs(622) <= a;
    layer6_outputs(623) <= not a;
    layer6_outputs(624) <= a and not b;
    layer6_outputs(625) <= b;
    layer6_outputs(626) <= a xor b;
    layer6_outputs(627) <= not (a or b);
    layer6_outputs(628) <= a xor b;
    layer6_outputs(629) <= a xor b;
    layer6_outputs(630) <= b;
    layer6_outputs(631) <= a and b;
    layer6_outputs(632) <= a and not b;
    layer6_outputs(633) <= not a;
    layer6_outputs(634) <= a and not b;
    layer6_outputs(635) <= not (a and b);
    layer6_outputs(636) <= b;
    layer6_outputs(637) <= not b;
    layer6_outputs(638) <= a xor b;
    layer6_outputs(639) <= not b or a;
    layer6_outputs(640) <= a and b;
    layer6_outputs(641) <= a;
    layer6_outputs(642) <= b and not a;
    layer6_outputs(643) <= not (a and b);
    layer6_outputs(644) <= not a;
    layer6_outputs(645) <= a;
    layer6_outputs(646) <= not a;
    layer6_outputs(647) <= not (a or b);
    layer6_outputs(648) <= a xor b;
    layer6_outputs(649) <= a xor b;
    layer6_outputs(650) <= b;
    layer6_outputs(651) <= not (a xor b);
    layer6_outputs(652) <= a xor b;
    layer6_outputs(653) <= b;
    layer6_outputs(654) <= not (a and b);
    layer6_outputs(655) <= not (a or b);
    layer6_outputs(656) <= not (a xor b);
    layer6_outputs(657) <= not b;
    layer6_outputs(658) <= a or b;
    layer6_outputs(659) <= not a or b;
    layer6_outputs(660) <= not (a or b);
    layer6_outputs(661) <= not a or b;
    layer6_outputs(662) <= a xor b;
    layer6_outputs(663) <= not (a xor b);
    layer6_outputs(664) <= b;
    layer6_outputs(665) <= not b or a;
    layer6_outputs(666) <= '1';
    layer6_outputs(667) <= not a;
    layer6_outputs(668) <= a xor b;
    layer6_outputs(669) <= not b;
    layer6_outputs(670) <= b;
    layer6_outputs(671) <= not a or b;
    layer6_outputs(672) <= not b;
    layer6_outputs(673) <= a;
    layer6_outputs(674) <= not a or b;
    layer6_outputs(675) <= not (a xor b);
    layer6_outputs(676) <= a and not b;
    layer6_outputs(677) <= not a or b;
    layer6_outputs(678) <= b;
    layer6_outputs(679) <= a xor b;
    layer6_outputs(680) <= not b or a;
    layer6_outputs(681) <= not (a or b);
    layer6_outputs(682) <= a;
    layer6_outputs(683) <= not b;
    layer6_outputs(684) <= a;
    layer6_outputs(685) <= a;
    layer6_outputs(686) <= not (a or b);
    layer6_outputs(687) <= not a;
    layer6_outputs(688) <= not (a xor b);
    layer6_outputs(689) <= a xor b;
    layer6_outputs(690) <= b;
    layer6_outputs(691) <= a and not b;
    layer6_outputs(692) <= a xor b;
    layer6_outputs(693) <= not a or b;
    layer6_outputs(694) <= a;
    layer6_outputs(695) <= a xor b;
    layer6_outputs(696) <= a;
    layer6_outputs(697) <= not (a xor b);
    layer6_outputs(698) <= a;
    layer6_outputs(699) <= not (a xor b);
    layer6_outputs(700) <= b and not a;
    layer6_outputs(701) <= b;
    layer6_outputs(702) <= not b;
    layer6_outputs(703) <= not b or a;
    layer6_outputs(704) <= a and b;
    layer6_outputs(705) <= a;
    layer6_outputs(706) <= not b;
    layer6_outputs(707) <= not a;
    layer6_outputs(708) <= a and not b;
    layer6_outputs(709) <= not b;
    layer6_outputs(710) <= b;
    layer6_outputs(711) <= not b;
    layer6_outputs(712) <= not (a xor b);
    layer6_outputs(713) <= a xor b;
    layer6_outputs(714) <= not b or a;
    layer6_outputs(715) <= not (a and b);
    layer6_outputs(716) <= not a or b;
    layer6_outputs(717) <= not (a and b);
    layer6_outputs(718) <= not b;
    layer6_outputs(719) <= not b;
    layer6_outputs(720) <= a and not b;
    layer6_outputs(721) <= not (a xor b);
    layer6_outputs(722) <= not b;
    layer6_outputs(723) <= b;
    layer6_outputs(724) <= a;
    layer6_outputs(725) <= not a;
    layer6_outputs(726) <= not (a and b);
    layer6_outputs(727) <= b;
    layer6_outputs(728) <= not a;
    layer6_outputs(729) <= a xor b;
    layer6_outputs(730) <= a and b;
    layer6_outputs(731) <= not b;
    layer6_outputs(732) <= a xor b;
    layer6_outputs(733) <= a and b;
    layer6_outputs(734) <= a or b;
    layer6_outputs(735) <= not a;
    layer6_outputs(736) <= a or b;
    layer6_outputs(737) <= a;
    layer6_outputs(738) <= not (a or b);
    layer6_outputs(739) <= a;
    layer6_outputs(740) <= b;
    layer6_outputs(741) <= a;
    layer6_outputs(742) <= not a;
    layer6_outputs(743) <= a or b;
    layer6_outputs(744) <= a;
    layer6_outputs(745) <= not a;
    layer6_outputs(746) <= not (a or b);
    layer6_outputs(747) <= not a;
    layer6_outputs(748) <= not (a and b);
    layer6_outputs(749) <= not a;
    layer6_outputs(750) <= a or b;
    layer6_outputs(751) <= not (a or b);
    layer6_outputs(752) <= a xor b;
    layer6_outputs(753) <= not a;
    layer6_outputs(754) <= b;
    layer6_outputs(755) <= not a or b;
    layer6_outputs(756) <= a or b;
    layer6_outputs(757) <= a;
    layer6_outputs(758) <= a and b;
    layer6_outputs(759) <= a or b;
    layer6_outputs(760) <= not (a or b);
    layer6_outputs(761) <= a and not b;
    layer6_outputs(762) <= a and not b;
    layer6_outputs(763) <= a xor b;
    layer6_outputs(764) <= not b or a;
    layer6_outputs(765) <= a;
    layer6_outputs(766) <= a;
    layer6_outputs(767) <= b;
    layer6_outputs(768) <= not a;
    layer6_outputs(769) <= not b or a;
    layer6_outputs(770) <= b;
    layer6_outputs(771) <= a xor b;
    layer6_outputs(772) <= not (a xor b);
    layer6_outputs(773) <= b;
    layer6_outputs(774) <= a xor b;
    layer6_outputs(775) <= not (a xor b);
    layer6_outputs(776) <= not a;
    layer6_outputs(777) <= a and b;
    layer6_outputs(778) <= a;
    layer6_outputs(779) <= not b;
    layer6_outputs(780) <= b;
    layer6_outputs(781) <= not a;
    layer6_outputs(782) <= not b;
    layer6_outputs(783) <= a xor b;
    layer6_outputs(784) <= not (a xor b);
    layer6_outputs(785) <= b;
    layer6_outputs(786) <= not (a and b);
    layer6_outputs(787) <= not a;
    layer6_outputs(788) <= not a or b;
    layer6_outputs(789) <= not (a or b);
    layer6_outputs(790) <= not b;
    layer6_outputs(791) <= b and not a;
    layer6_outputs(792) <= a;
    layer6_outputs(793) <= a xor b;
    layer6_outputs(794) <= b;
    layer6_outputs(795) <= b;
    layer6_outputs(796) <= b;
    layer6_outputs(797) <= not a;
    layer6_outputs(798) <= a xor b;
    layer6_outputs(799) <= b;
    layer6_outputs(800) <= not a;
    layer6_outputs(801) <= not b;
    layer6_outputs(802) <= not a;
    layer6_outputs(803) <= not (a xor b);
    layer6_outputs(804) <= a;
    layer6_outputs(805) <= not (a or b);
    layer6_outputs(806) <= not b;
    layer6_outputs(807) <= not (a xor b);
    layer6_outputs(808) <= b and not a;
    layer6_outputs(809) <= a or b;
    layer6_outputs(810) <= not (a and b);
    layer6_outputs(811) <= not b;
    layer6_outputs(812) <= not b;
    layer6_outputs(813) <= a or b;
    layer6_outputs(814) <= a xor b;
    layer6_outputs(815) <= not b;
    layer6_outputs(816) <= not (a or b);
    layer6_outputs(817) <= a or b;
    layer6_outputs(818) <= a or b;
    layer6_outputs(819) <= not (a or b);
    layer6_outputs(820) <= a;
    layer6_outputs(821) <= not b;
    layer6_outputs(822) <= b;
    layer6_outputs(823) <= not (a and b);
    layer6_outputs(824) <= b and not a;
    layer6_outputs(825) <= b and not a;
    layer6_outputs(826) <= a or b;
    layer6_outputs(827) <= not b or a;
    layer6_outputs(828) <= a and not b;
    layer6_outputs(829) <= b;
    layer6_outputs(830) <= a and b;
    layer6_outputs(831) <= a or b;
    layer6_outputs(832) <= a and b;
    layer6_outputs(833) <= a and b;
    layer6_outputs(834) <= not (a or b);
    layer6_outputs(835) <= a;
    layer6_outputs(836) <= not (a xor b);
    layer6_outputs(837) <= a;
    layer6_outputs(838) <= a;
    layer6_outputs(839) <= not (a xor b);
    layer6_outputs(840) <= not b;
    layer6_outputs(841) <= b;
    layer6_outputs(842) <= not b;
    layer6_outputs(843) <= a and b;
    layer6_outputs(844) <= b;
    layer6_outputs(845) <= b and not a;
    layer6_outputs(846) <= a;
    layer6_outputs(847) <= not a;
    layer6_outputs(848) <= not a;
    layer6_outputs(849) <= a;
    layer6_outputs(850) <= a xor b;
    layer6_outputs(851) <= not b;
    layer6_outputs(852) <= not a or b;
    layer6_outputs(853) <= a and not b;
    layer6_outputs(854) <= a or b;
    layer6_outputs(855) <= not a or b;
    layer6_outputs(856) <= a and not b;
    layer6_outputs(857) <= a;
    layer6_outputs(858) <= not a or b;
    layer6_outputs(859) <= not a;
    layer6_outputs(860) <= a xor b;
    layer6_outputs(861) <= a xor b;
    layer6_outputs(862) <= b;
    layer6_outputs(863) <= b;
    layer6_outputs(864) <= not a;
    layer6_outputs(865) <= not b or a;
    layer6_outputs(866) <= not a or b;
    layer6_outputs(867) <= not b;
    layer6_outputs(868) <= a;
    layer6_outputs(869) <= a;
    layer6_outputs(870) <= not (a and b);
    layer6_outputs(871) <= not (a xor b);
    layer6_outputs(872) <= '0';
    layer6_outputs(873) <= not b or a;
    layer6_outputs(874) <= b;
    layer6_outputs(875) <= not (a and b);
    layer6_outputs(876) <= a;
    layer6_outputs(877) <= not a;
    layer6_outputs(878) <= not b or a;
    layer6_outputs(879) <= not b;
    layer6_outputs(880) <= a or b;
    layer6_outputs(881) <= a;
    layer6_outputs(882) <= not a;
    layer6_outputs(883) <= not b;
    layer6_outputs(884) <= b;
    layer6_outputs(885) <= not a;
    layer6_outputs(886) <= a;
    layer6_outputs(887) <= not a;
    layer6_outputs(888) <= not b or a;
    layer6_outputs(889) <= a;
    layer6_outputs(890) <= a and not b;
    layer6_outputs(891) <= not a;
    layer6_outputs(892) <= b;
    layer6_outputs(893) <= not (a xor b);
    layer6_outputs(894) <= not b;
    layer6_outputs(895) <= a or b;
    layer6_outputs(896) <= b;
    layer6_outputs(897) <= a;
    layer6_outputs(898) <= a xor b;
    layer6_outputs(899) <= not b;
    layer6_outputs(900) <= not (a xor b);
    layer6_outputs(901) <= b and not a;
    layer6_outputs(902) <= not (a xor b);
    layer6_outputs(903) <= a;
    layer6_outputs(904) <= a;
    layer6_outputs(905) <= a xor b;
    layer6_outputs(906) <= not (a xor b);
    layer6_outputs(907) <= a;
    layer6_outputs(908) <= a;
    layer6_outputs(909) <= not a;
    layer6_outputs(910) <= a;
    layer6_outputs(911) <= not a;
    layer6_outputs(912) <= a xor b;
    layer6_outputs(913) <= not (a xor b);
    layer6_outputs(914) <= a xor b;
    layer6_outputs(915) <= not (a and b);
    layer6_outputs(916) <= not a;
    layer6_outputs(917) <= not a or b;
    layer6_outputs(918) <= not (a xor b);
    layer6_outputs(919) <= b;
    layer6_outputs(920) <= a;
    layer6_outputs(921) <= not a;
    layer6_outputs(922) <= not b or a;
    layer6_outputs(923) <= a;
    layer6_outputs(924) <= a;
    layer6_outputs(925) <= not a;
    layer6_outputs(926) <= not a or b;
    layer6_outputs(927) <= '0';
    layer6_outputs(928) <= a;
    layer6_outputs(929) <= not a;
    layer6_outputs(930) <= a;
    layer6_outputs(931) <= not b or a;
    layer6_outputs(932) <= a and b;
    layer6_outputs(933) <= b and not a;
    layer6_outputs(934) <= not (a xor b);
    layer6_outputs(935) <= b;
    layer6_outputs(936) <= b;
    layer6_outputs(937) <= not b;
    layer6_outputs(938) <= not b;
    layer6_outputs(939) <= a xor b;
    layer6_outputs(940) <= not a;
    layer6_outputs(941) <= not b;
    layer6_outputs(942) <= a and not b;
    layer6_outputs(943) <= not (a or b);
    layer6_outputs(944) <= a and not b;
    layer6_outputs(945) <= not a;
    layer6_outputs(946) <= a or b;
    layer6_outputs(947) <= not (a or b);
    layer6_outputs(948) <= not a or b;
    layer6_outputs(949) <= not b;
    layer6_outputs(950) <= not a;
    layer6_outputs(951) <= a and not b;
    layer6_outputs(952) <= a;
    layer6_outputs(953) <= not b;
    layer6_outputs(954) <= a xor b;
    layer6_outputs(955) <= not a;
    layer6_outputs(956) <= not (a xor b);
    layer6_outputs(957) <= a and b;
    layer6_outputs(958) <= not (a xor b);
    layer6_outputs(959) <= not (a and b);
    layer6_outputs(960) <= not b;
    layer6_outputs(961) <= a;
    layer6_outputs(962) <= a and b;
    layer6_outputs(963) <= b;
    layer6_outputs(964) <= not a;
    layer6_outputs(965) <= a;
    layer6_outputs(966) <= a xor b;
    layer6_outputs(967) <= not b;
    layer6_outputs(968) <= not (a xor b);
    layer6_outputs(969) <= a;
    layer6_outputs(970) <= not a;
    layer6_outputs(971) <= not (a xor b);
    layer6_outputs(972) <= not (a xor b);
    layer6_outputs(973) <= not b;
    layer6_outputs(974) <= not a or b;
    layer6_outputs(975) <= not b;
    layer6_outputs(976) <= not (a or b);
    layer6_outputs(977) <= not b;
    layer6_outputs(978) <= a;
    layer6_outputs(979) <= b;
    layer6_outputs(980) <= a;
    layer6_outputs(981) <= not a or b;
    layer6_outputs(982) <= b;
    layer6_outputs(983) <= not (a xor b);
    layer6_outputs(984) <= a;
    layer6_outputs(985) <= a or b;
    layer6_outputs(986) <= a and not b;
    layer6_outputs(987) <= b;
    layer6_outputs(988) <= b and not a;
    layer6_outputs(989) <= a;
    layer6_outputs(990) <= not (a xor b);
    layer6_outputs(991) <= a and not b;
    layer6_outputs(992) <= a and not b;
    layer6_outputs(993) <= not b;
    layer6_outputs(994) <= not a;
    layer6_outputs(995) <= a;
    layer6_outputs(996) <= b;
    layer6_outputs(997) <= a xor b;
    layer6_outputs(998) <= not a or b;
    layer6_outputs(999) <= a;
    layer6_outputs(1000) <= a;
    layer6_outputs(1001) <= not a;
    layer6_outputs(1002) <= not b or a;
    layer6_outputs(1003) <= a;
    layer6_outputs(1004) <= not a;
    layer6_outputs(1005) <= not (a xor b);
    layer6_outputs(1006) <= not (a xor b);
    layer6_outputs(1007) <= a;
    layer6_outputs(1008) <= not b;
    layer6_outputs(1009) <= a;
    layer6_outputs(1010) <= a and not b;
    layer6_outputs(1011) <= a;
    layer6_outputs(1012) <= not b or a;
    layer6_outputs(1013) <= not (a xor b);
    layer6_outputs(1014) <= not a or b;
    layer6_outputs(1015) <= a;
    layer6_outputs(1016) <= a;
    layer6_outputs(1017) <= not a;
    layer6_outputs(1018) <= not a;
    layer6_outputs(1019) <= a or b;
    layer6_outputs(1020) <= b and not a;
    layer6_outputs(1021) <= not b;
    layer6_outputs(1022) <= not a or b;
    layer6_outputs(1023) <= not (a xor b);
    layer6_outputs(1024) <= not a;
    layer6_outputs(1025) <= b and not a;
    layer6_outputs(1026) <= a or b;
    layer6_outputs(1027) <= a xor b;
    layer6_outputs(1028) <= a xor b;
    layer6_outputs(1029) <= a and not b;
    layer6_outputs(1030) <= b and not a;
    layer6_outputs(1031) <= not a;
    layer6_outputs(1032) <= a;
    layer6_outputs(1033) <= b;
    layer6_outputs(1034) <= not b;
    layer6_outputs(1035) <= b and not a;
    layer6_outputs(1036) <= not (a and b);
    layer6_outputs(1037) <= not b or a;
    layer6_outputs(1038) <= a;
    layer6_outputs(1039) <= b and not a;
    layer6_outputs(1040) <= b and not a;
    layer6_outputs(1041) <= not a or b;
    layer6_outputs(1042) <= b;
    layer6_outputs(1043) <= not a;
    layer6_outputs(1044) <= a;
    layer6_outputs(1045) <= not a;
    layer6_outputs(1046) <= not a or b;
    layer6_outputs(1047) <= not a;
    layer6_outputs(1048) <= not a or b;
    layer6_outputs(1049) <= a xor b;
    layer6_outputs(1050) <= a xor b;
    layer6_outputs(1051) <= b and not a;
    layer6_outputs(1052) <= a xor b;
    layer6_outputs(1053) <= not (a xor b);
    layer6_outputs(1054) <= not (a xor b);
    layer6_outputs(1055) <= not a;
    layer6_outputs(1056) <= a or b;
    layer6_outputs(1057) <= not b;
    layer6_outputs(1058) <= b;
    layer6_outputs(1059) <= not a;
    layer6_outputs(1060) <= not (a xor b);
    layer6_outputs(1061) <= a;
    layer6_outputs(1062) <= b;
    layer6_outputs(1063) <= a;
    layer6_outputs(1064) <= a xor b;
    layer6_outputs(1065) <= a;
    layer6_outputs(1066) <= a or b;
    layer6_outputs(1067) <= a;
    layer6_outputs(1068) <= not b;
    layer6_outputs(1069) <= a xor b;
    layer6_outputs(1070) <= not b;
    layer6_outputs(1071) <= not (a xor b);
    layer6_outputs(1072) <= a xor b;
    layer6_outputs(1073) <= a xor b;
    layer6_outputs(1074) <= a xor b;
    layer6_outputs(1075) <= not a;
    layer6_outputs(1076) <= not b;
    layer6_outputs(1077) <= a xor b;
    layer6_outputs(1078) <= b;
    layer6_outputs(1079) <= not (a xor b);
    layer6_outputs(1080) <= not b or a;
    layer6_outputs(1081) <= not b;
    layer6_outputs(1082) <= a;
    layer6_outputs(1083) <= not (a or b);
    layer6_outputs(1084) <= a xor b;
    layer6_outputs(1085) <= not a;
    layer6_outputs(1086) <= a or b;
    layer6_outputs(1087) <= not b;
    layer6_outputs(1088) <= not b or a;
    layer6_outputs(1089) <= a;
    layer6_outputs(1090) <= not (a xor b);
    layer6_outputs(1091) <= a;
    layer6_outputs(1092) <= b;
    layer6_outputs(1093) <= a xor b;
    layer6_outputs(1094) <= b;
    layer6_outputs(1095) <= '0';
    layer6_outputs(1096) <= not a or b;
    layer6_outputs(1097) <= not b;
    layer6_outputs(1098) <= not b;
    layer6_outputs(1099) <= b;
    layer6_outputs(1100) <= b;
    layer6_outputs(1101) <= not a;
    layer6_outputs(1102) <= not (a and b);
    layer6_outputs(1103) <= not b or a;
    layer6_outputs(1104) <= not (a and b);
    layer6_outputs(1105) <= b and not a;
    layer6_outputs(1106) <= not a or b;
    layer6_outputs(1107) <= not (a or b);
    layer6_outputs(1108) <= b;
    layer6_outputs(1109) <= a xor b;
    layer6_outputs(1110) <= a xor b;
    layer6_outputs(1111) <= not (a xor b);
    layer6_outputs(1112) <= a;
    layer6_outputs(1113) <= b;
    layer6_outputs(1114) <= b;
    layer6_outputs(1115) <= b;
    layer6_outputs(1116) <= b;
    layer6_outputs(1117) <= a or b;
    layer6_outputs(1118) <= b;
    layer6_outputs(1119) <= not b;
    layer6_outputs(1120) <= not (a xor b);
    layer6_outputs(1121) <= not (a or b);
    layer6_outputs(1122) <= not (a xor b);
    layer6_outputs(1123) <= a and b;
    layer6_outputs(1124) <= not (a xor b);
    layer6_outputs(1125) <= a;
    layer6_outputs(1126) <= b;
    layer6_outputs(1127) <= not (a xor b);
    layer6_outputs(1128) <= a or b;
    layer6_outputs(1129) <= not (a xor b);
    layer6_outputs(1130) <= not a;
    layer6_outputs(1131) <= not a;
    layer6_outputs(1132) <= not (a and b);
    layer6_outputs(1133) <= b;
    layer6_outputs(1134) <= not b;
    layer6_outputs(1135) <= not a;
    layer6_outputs(1136) <= not (a xor b);
    layer6_outputs(1137) <= not a;
    layer6_outputs(1138) <= a;
    layer6_outputs(1139) <= not (a xor b);
    layer6_outputs(1140) <= b;
    layer6_outputs(1141) <= not a;
    layer6_outputs(1142) <= '0';
    layer6_outputs(1143) <= b and not a;
    layer6_outputs(1144) <= a xor b;
    layer6_outputs(1145) <= a or b;
    layer6_outputs(1146) <= not b;
    layer6_outputs(1147) <= b;
    layer6_outputs(1148) <= a;
    layer6_outputs(1149) <= not b;
    layer6_outputs(1150) <= a;
    layer6_outputs(1151) <= not a;
    layer6_outputs(1152) <= a and b;
    layer6_outputs(1153) <= b and not a;
    layer6_outputs(1154) <= not (a or b);
    layer6_outputs(1155) <= not b;
    layer6_outputs(1156) <= b;
    layer6_outputs(1157) <= b;
    layer6_outputs(1158) <= not (a or b);
    layer6_outputs(1159) <= a xor b;
    layer6_outputs(1160) <= b;
    layer6_outputs(1161) <= b;
    layer6_outputs(1162) <= not b;
    layer6_outputs(1163) <= not (a and b);
    layer6_outputs(1164) <= b;
    layer6_outputs(1165) <= not (a and b);
    layer6_outputs(1166) <= not b;
    layer6_outputs(1167) <= a;
    layer6_outputs(1168) <= not a;
    layer6_outputs(1169) <= b and not a;
    layer6_outputs(1170) <= not (a or b);
    layer6_outputs(1171) <= not (a or b);
    layer6_outputs(1172) <= a xor b;
    layer6_outputs(1173) <= not b;
    layer6_outputs(1174) <= not a;
    layer6_outputs(1175) <= a;
    layer6_outputs(1176) <= not b or a;
    layer6_outputs(1177) <= not (a or b);
    layer6_outputs(1178) <= not a;
    layer6_outputs(1179) <= a xor b;
    layer6_outputs(1180) <= a and not b;
    layer6_outputs(1181) <= not a;
    layer6_outputs(1182) <= b;
    layer6_outputs(1183) <= not a;
    layer6_outputs(1184) <= not b;
    layer6_outputs(1185) <= not b;
    layer6_outputs(1186) <= a or b;
    layer6_outputs(1187) <= not (a and b);
    layer6_outputs(1188) <= a xor b;
    layer6_outputs(1189) <= b;
    layer6_outputs(1190) <= not a;
    layer6_outputs(1191) <= not a;
    layer6_outputs(1192) <= not a or b;
    layer6_outputs(1193) <= not b or a;
    layer6_outputs(1194) <= not (a and b);
    layer6_outputs(1195) <= b;
    layer6_outputs(1196) <= a xor b;
    layer6_outputs(1197) <= a;
    layer6_outputs(1198) <= not (a xor b);
    layer6_outputs(1199) <= not a;
    layer6_outputs(1200) <= not b;
    layer6_outputs(1201) <= not (a xor b);
    layer6_outputs(1202) <= not b;
    layer6_outputs(1203) <= not (a or b);
    layer6_outputs(1204) <= b and not a;
    layer6_outputs(1205) <= not (a or b);
    layer6_outputs(1206) <= not a;
    layer6_outputs(1207) <= b;
    layer6_outputs(1208) <= '1';
    layer6_outputs(1209) <= not b or a;
    layer6_outputs(1210) <= not (a or b);
    layer6_outputs(1211) <= b;
    layer6_outputs(1212) <= a xor b;
    layer6_outputs(1213) <= a xor b;
    layer6_outputs(1214) <= not b;
    layer6_outputs(1215) <= not (a or b);
    layer6_outputs(1216) <= not a;
    layer6_outputs(1217) <= not (a or b);
    layer6_outputs(1218) <= a and not b;
    layer6_outputs(1219) <= a and b;
    layer6_outputs(1220) <= a or b;
    layer6_outputs(1221) <= a;
    layer6_outputs(1222) <= a and not b;
    layer6_outputs(1223) <= not (a xor b);
    layer6_outputs(1224) <= b;
    layer6_outputs(1225) <= a or b;
    layer6_outputs(1226) <= a;
    layer6_outputs(1227) <= b;
    layer6_outputs(1228) <= b and not a;
    layer6_outputs(1229) <= not a;
    layer6_outputs(1230) <= b;
    layer6_outputs(1231) <= not b or a;
    layer6_outputs(1232) <= b;
    layer6_outputs(1233) <= not b or a;
    layer6_outputs(1234) <= b and not a;
    layer6_outputs(1235) <= b;
    layer6_outputs(1236) <= not a;
    layer6_outputs(1237) <= not (a xor b);
    layer6_outputs(1238) <= a xor b;
    layer6_outputs(1239) <= not b or a;
    layer6_outputs(1240) <= not (a xor b);
    layer6_outputs(1241) <= not (a xor b);
    layer6_outputs(1242) <= b and not a;
    layer6_outputs(1243) <= not a;
    layer6_outputs(1244) <= a;
    layer6_outputs(1245) <= a or b;
    layer6_outputs(1246) <= not (a or b);
    layer6_outputs(1247) <= not b;
    layer6_outputs(1248) <= a;
    layer6_outputs(1249) <= not a;
    layer6_outputs(1250) <= not (a xor b);
    layer6_outputs(1251) <= not b;
    layer6_outputs(1252) <= not b;
    layer6_outputs(1253) <= a or b;
    layer6_outputs(1254) <= not (a xor b);
    layer6_outputs(1255) <= not a;
    layer6_outputs(1256) <= not b;
    layer6_outputs(1257) <= a xor b;
    layer6_outputs(1258) <= a or b;
    layer6_outputs(1259) <= not (a xor b);
    layer6_outputs(1260) <= b and not a;
    layer6_outputs(1261) <= not b or a;
    layer6_outputs(1262) <= not (a or b);
    layer6_outputs(1263) <= not a;
    layer6_outputs(1264) <= not a;
    layer6_outputs(1265) <= a or b;
    layer6_outputs(1266) <= a;
    layer6_outputs(1267) <= not b or a;
    layer6_outputs(1268) <= a;
    layer6_outputs(1269) <= b and not a;
    layer6_outputs(1270) <= not a or b;
    layer6_outputs(1271) <= not b or a;
    layer6_outputs(1272) <= not (a and b);
    layer6_outputs(1273) <= a and b;
    layer6_outputs(1274) <= not (a and b);
    layer6_outputs(1275) <= not b;
    layer6_outputs(1276) <= a and b;
    layer6_outputs(1277) <= not b;
    layer6_outputs(1278) <= a xor b;
    layer6_outputs(1279) <= not b or a;
    layer6_outputs(1280) <= a or b;
    layer6_outputs(1281) <= a and not b;
    layer6_outputs(1282) <= a and b;
    layer6_outputs(1283) <= not b;
    layer6_outputs(1284) <= not b;
    layer6_outputs(1285) <= a and b;
    layer6_outputs(1286) <= not (a or b);
    layer6_outputs(1287) <= a;
    layer6_outputs(1288) <= not b;
    layer6_outputs(1289) <= a and b;
    layer6_outputs(1290) <= a;
    layer6_outputs(1291) <= b;
    layer6_outputs(1292) <= a and b;
    layer6_outputs(1293) <= a;
    layer6_outputs(1294) <= b and not a;
    layer6_outputs(1295) <= not a;
    layer6_outputs(1296) <= not (a xor b);
    layer6_outputs(1297) <= not a or b;
    layer6_outputs(1298) <= not a;
    layer6_outputs(1299) <= a and b;
    layer6_outputs(1300) <= not b;
    layer6_outputs(1301) <= not (a xor b);
    layer6_outputs(1302) <= a;
    layer6_outputs(1303) <= a and b;
    layer6_outputs(1304) <= a xor b;
    layer6_outputs(1305) <= b;
    layer6_outputs(1306) <= a;
    layer6_outputs(1307) <= not b;
    layer6_outputs(1308) <= b;
    layer6_outputs(1309) <= b and not a;
    layer6_outputs(1310) <= not (a xor b);
    layer6_outputs(1311) <= a or b;
    layer6_outputs(1312) <= a or b;
    layer6_outputs(1313) <= not (a xor b);
    layer6_outputs(1314) <= a xor b;
    layer6_outputs(1315) <= a xor b;
    layer6_outputs(1316) <= not (a xor b);
    layer6_outputs(1317) <= b;
    layer6_outputs(1318) <= not a;
    layer6_outputs(1319) <= not (a and b);
    layer6_outputs(1320) <= a xor b;
    layer6_outputs(1321) <= not a;
    layer6_outputs(1322) <= a xor b;
    layer6_outputs(1323) <= not (a and b);
    layer6_outputs(1324) <= a xor b;
    layer6_outputs(1325) <= a and not b;
    layer6_outputs(1326) <= not a;
    layer6_outputs(1327) <= not a;
    layer6_outputs(1328) <= a;
    layer6_outputs(1329) <= b;
    layer6_outputs(1330) <= not a;
    layer6_outputs(1331) <= a xor b;
    layer6_outputs(1332) <= b and not a;
    layer6_outputs(1333) <= not a;
    layer6_outputs(1334) <= a and b;
    layer6_outputs(1335) <= b;
    layer6_outputs(1336) <= not (a xor b);
    layer6_outputs(1337) <= not (a xor b);
    layer6_outputs(1338) <= not a;
    layer6_outputs(1339) <= not b or a;
    layer6_outputs(1340) <= a;
    layer6_outputs(1341) <= a;
    layer6_outputs(1342) <= a;
    layer6_outputs(1343) <= a;
    layer6_outputs(1344) <= not (a or b);
    layer6_outputs(1345) <= not a or b;
    layer6_outputs(1346) <= not a or b;
    layer6_outputs(1347) <= a and not b;
    layer6_outputs(1348) <= a xor b;
    layer6_outputs(1349) <= not b;
    layer6_outputs(1350) <= not (a and b);
    layer6_outputs(1351) <= b;
    layer6_outputs(1352) <= not b;
    layer6_outputs(1353) <= a and not b;
    layer6_outputs(1354) <= not b or a;
    layer6_outputs(1355) <= b;
    layer6_outputs(1356) <= not (a xor b);
    layer6_outputs(1357) <= b;
    layer6_outputs(1358) <= b;
    layer6_outputs(1359) <= a xor b;
    layer6_outputs(1360) <= not (a and b);
    layer6_outputs(1361) <= not a;
    layer6_outputs(1362) <= not (a or b);
    layer6_outputs(1363) <= a;
    layer6_outputs(1364) <= a or b;
    layer6_outputs(1365) <= not b;
    layer6_outputs(1366) <= not (a and b);
    layer6_outputs(1367) <= not a;
    layer6_outputs(1368) <= not a;
    layer6_outputs(1369) <= b;
    layer6_outputs(1370) <= b;
    layer6_outputs(1371) <= a and not b;
    layer6_outputs(1372) <= not a;
    layer6_outputs(1373) <= a and not b;
    layer6_outputs(1374) <= a;
    layer6_outputs(1375) <= not b;
    layer6_outputs(1376) <= not a;
    layer6_outputs(1377) <= b;
    layer6_outputs(1378) <= not b or a;
    layer6_outputs(1379) <= a and not b;
    layer6_outputs(1380) <= not a;
    layer6_outputs(1381) <= not a or b;
    layer6_outputs(1382) <= not (a xor b);
    layer6_outputs(1383) <= not a or b;
    layer6_outputs(1384) <= b;
    layer6_outputs(1385) <= not (a or b);
    layer6_outputs(1386) <= not a;
    layer6_outputs(1387) <= not (a and b);
    layer6_outputs(1388) <= a;
    layer6_outputs(1389) <= a xor b;
    layer6_outputs(1390) <= not b;
    layer6_outputs(1391) <= not a;
    layer6_outputs(1392) <= not b;
    layer6_outputs(1393) <= not a or b;
    layer6_outputs(1394) <= a or b;
    layer6_outputs(1395) <= a xor b;
    layer6_outputs(1396) <= not b or a;
    layer6_outputs(1397) <= a or b;
    layer6_outputs(1398) <= b;
    layer6_outputs(1399) <= a;
    layer6_outputs(1400) <= not a;
    layer6_outputs(1401) <= a xor b;
    layer6_outputs(1402) <= a;
    layer6_outputs(1403) <= a xor b;
    layer6_outputs(1404) <= not b or a;
    layer6_outputs(1405) <= a xor b;
    layer6_outputs(1406) <= a;
    layer6_outputs(1407) <= a xor b;
    layer6_outputs(1408) <= not (a and b);
    layer6_outputs(1409) <= a and not b;
    layer6_outputs(1410) <= not a;
    layer6_outputs(1411) <= not a;
    layer6_outputs(1412) <= b;
    layer6_outputs(1413) <= a xor b;
    layer6_outputs(1414) <= not b;
    layer6_outputs(1415) <= not (a xor b);
    layer6_outputs(1416) <= not a;
    layer6_outputs(1417) <= a xor b;
    layer6_outputs(1418) <= not (a and b);
    layer6_outputs(1419) <= '0';
    layer6_outputs(1420) <= a;
    layer6_outputs(1421) <= b;
    layer6_outputs(1422) <= a xor b;
    layer6_outputs(1423) <= b;
    layer6_outputs(1424) <= b and not a;
    layer6_outputs(1425) <= not (a or b);
    layer6_outputs(1426) <= b;
    layer6_outputs(1427) <= not a;
    layer6_outputs(1428) <= a xor b;
    layer6_outputs(1429) <= not b;
    layer6_outputs(1430) <= a xor b;
    layer6_outputs(1431) <= not (a and b);
    layer6_outputs(1432) <= a xor b;
    layer6_outputs(1433) <= not b;
    layer6_outputs(1434) <= not a or b;
    layer6_outputs(1435) <= not b;
    layer6_outputs(1436) <= a xor b;
    layer6_outputs(1437) <= not (a xor b);
    layer6_outputs(1438) <= a;
    layer6_outputs(1439) <= not (a xor b);
    layer6_outputs(1440) <= not a;
    layer6_outputs(1441) <= not (a and b);
    layer6_outputs(1442) <= not (a and b);
    layer6_outputs(1443) <= a xor b;
    layer6_outputs(1444) <= not b;
    layer6_outputs(1445) <= a xor b;
    layer6_outputs(1446) <= b and not a;
    layer6_outputs(1447) <= not (a and b);
    layer6_outputs(1448) <= a;
    layer6_outputs(1449) <= not a;
    layer6_outputs(1450) <= not a;
    layer6_outputs(1451) <= not b;
    layer6_outputs(1452) <= b;
    layer6_outputs(1453) <= a;
    layer6_outputs(1454) <= a or b;
    layer6_outputs(1455) <= not b;
    layer6_outputs(1456) <= not (a and b);
    layer6_outputs(1457) <= not b;
    layer6_outputs(1458) <= b;
    layer6_outputs(1459) <= not a or b;
    layer6_outputs(1460) <= a;
    layer6_outputs(1461) <= not (a xor b);
    layer6_outputs(1462) <= not b;
    layer6_outputs(1463) <= not a or b;
    layer6_outputs(1464) <= not (a xor b);
    layer6_outputs(1465) <= not a;
    layer6_outputs(1466) <= not (a or b);
    layer6_outputs(1467) <= a xor b;
    layer6_outputs(1468) <= not b;
    layer6_outputs(1469) <= not a;
    layer6_outputs(1470) <= a xor b;
    layer6_outputs(1471) <= not (a and b);
    layer6_outputs(1472) <= a and b;
    layer6_outputs(1473) <= not (a and b);
    layer6_outputs(1474) <= a and not b;
    layer6_outputs(1475) <= b;
    layer6_outputs(1476) <= a and b;
    layer6_outputs(1477) <= b;
    layer6_outputs(1478) <= not (a and b);
    layer6_outputs(1479) <= b;
    layer6_outputs(1480) <= a and b;
    layer6_outputs(1481) <= b and not a;
    layer6_outputs(1482) <= not a;
    layer6_outputs(1483) <= a and not b;
    layer6_outputs(1484) <= not (a xor b);
    layer6_outputs(1485) <= not a;
    layer6_outputs(1486) <= b;
    layer6_outputs(1487) <= a xor b;
    layer6_outputs(1488) <= b;
    layer6_outputs(1489) <= not a;
    layer6_outputs(1490) <= not (a xor b);
    layer6_outputs(1491) <= not b;
    layer6_outputs(1492) <= a and b;
    layer6_outputs(1493) <= b and not a;
    layer6_outputs(1494) <= not (a and b);
    layer6_outputs(1495) <= not (a or b);
    layer6_outputs(1496) <= a;
    layer6_outputs(1497) <= not (a xor b);
    layer6_outputs(1498) <= a and not b;
    layer6_outputs(1499) <= not b;
    layer6_outputs(1500) <= not (a xor b);
    layer6_outputs(1501) <= '1';
    layer6_outputs(1502) <= not b;
    layer6_outputs(1503) <= a;
    layer6_outputs(1504) <= a or b;
    layer6_outputs(1505) <= not a;
    layer6_outputs(1506) <= b;
    layer6_outputs(1507) <= not (a or b);
    layer6_outputs(1508) <= b and not a;
    layer6_outputs(1509) <= not b;
    layer6_outputs(1510) <= not a;
    layer6_outputs(1511) <= a;
    layer6_outputs(1512) <= b and not a;
    layer6_outputs(1513) <= not (a xor b);
    layer6_outputs(1514) <= not (a xor b);
    layer6_outputs(1515) <= not a;
    layer6_outputs(1516) <= b and not a;
    layer6_outputs(1517) <= not a;
    layer6_outputs(1518) <= not b;
    layer6_outputs(1519) <= b;
    layer6_outputs(1520) <= a;
    layer6_outputs(1521) <= not (a xor b);
    layer6_outputs(1522) <= a;
    layer6_outputs(1523) <= a and not b;
    layer6_outputs(1524) <= a and b;
    layer6_outputs(1525) <= not a;
    layer6_outputs(1526) <= a or b;
    layer6_outputs(1527) <= not a;
    layer6_outputs(1528) <= not a or b;
    layer6_outputs(1529) <= a;
    layer6_outputs(1530) <= a;
    layer6_outputs(1531) <= not (a xor b);
    layer6_outputs(1532) <= not a;
    layer6_outputs(1533) <= a or b;
    layer6_outputs(1534) <= '1';
    layer6_outputs(1535) <= a;
    layer6_outputs(1536) <= a;
    layer6_outputs(1537) <= not a;
    layer6_outputs(1538) <= a and b;
    layer6_outputs(1539) <= not (a xor b);
    layer6_outputs(1540) <= b;
    layer6_outputs(1541) <= a xor b;
    layer6_outputs(1542) <= a xor b;
    layer6_outputs(1543) <= a xor b;
    layer6_outputs(1544) <= a xor b;
    layer6_outputs(1545) <= a or b;
    layer6_outputs(1546) <= not a;
    layer6_outputs(1547) <= not b or a;
    layer6_outputs(1548) <= not (a xor b);
    layer6_outputs(1549) <= b and not a;
    layer6_outputs(1550) <= a or b;
    layer6_outputs(1551) <= not a;
    layer6_outputs(1552) <= b;
    layer6_outputs(1553) <= not b or a;
    layer6_outputs(1554) <= not a;
    layer6_outputs(1555) <= a;
    layer6_outputs(1556) <= b;
    layer6_outputs(1557) <= b;
    layer6_outputs(1558) <= a and b;
    layer6_outputs(1559) <= a xor b;
    layer6_outputs(1560) <= not (a or b);
    layer6_outputs(1561) <= not a;
    layer6_outputs(1562) <= not a;
    layer6_outputs(1563) <= not b;
    layer6_outputs(1564) <= b;
    layer6_outputs(1565) <= not b or a;
    layer6_outputs(1566) <= not (a and b);
    layer6_outputs(1567) <= not a;
    layer6_outputs(1568) <= a;
    layer6_outputs(1569) <= not (a or b);
    layer6_outputs(1570) <= not b;
    layer6_outputs(1571) <= not (a xor b);
    layer6_outputs(1572) <= not b or a;
    layer6_outputs(1573) <= not a;
    layer6_outputs(1574) <= not a;
    layer6_outputs(1575) <= b;
    layer6_outputs(1576) <= a;
    layer6_outputs(1577) <= a xor b;
    layer6_outputs(1578) <= not b;
    layer6_outputs(1579) <= b;
    layer6_outputs(1580) <= a and b;
    layer6_outputs(1581) <= a;
    layer6_outputs(1582) <= not b;
    layer6_outputs(1583) <= not (a and b);
    layer6_outputs(1584) <= a;
    layer6_outputs(1585) <= not a;
    layer6_outputs(1586) <= not b or a;
    layer6_outputs(1587) <= not a;
    layer6_outputs(1588) <= not a;
    layer6_outputs(1589) <= not b or a;
    layer6_outputs(1590) <= not b;
    layer6_outputs(1591) <= b and not a;
    layer6_outputs(1592) <= b;
    layer6_outputs(1593) <= not a;
    layer6_outputs(1594) <= not b;
    layer6_outputs(1595) <= a xor b;
    layer6_outputs(1596) <= not a;
    layer6_outputs(1597) <= b and not a;
    layer6_outputs(1598) <= not (a and b);
    layer6_outputs(1599) <= b and not a;
    layer6_outputs(1600) <= a;
    layer6_outputs(1601) <= a;
    layer6_outputs(1602) <= not (a or b);
    layer6_outputs(1603) <= not b;
    layer6_outputs(1604) <= not a;
    layer6_outputs(1605) <= not (a xor b);
    layer6_outputs(1606) <= not (a xor b);
    layer6_outputs(1607) <= b and not a;
    layer6_outputs(1608) <= not b;
    layer6_outputs(1609) <= b;
    layer6_outputs(1610) <= not b;
    layer6_outputs(1611) <= b;
    layer6_outputs(1612) <= not a or b;
    layer6_outputs(1613) <= not a;
    layer6_outputs(1614) <= not a;
    layer6_outputs(1615) <= not (a or b);
    layer6_outputs(1616) <= b and not a;
    layer6_outputs(1617) <= b;
    layer6_outputs(1618) <= a xor b;
    layer6_outputs(1619) <= not b;
    layer6_outputs(1620) <= not (a xor b);
    layer6_outputs(1621) <= not b or a;
    layer6_outputs(1622) <= not (a and b);
    layer6_outputs(1623) <= not (a xor b);
    layer6_outputs(1624) <= not b;
    layer6_outputs(1625) <= not b;
    layer6_outputs(1626) <= b and not a;
    layer6_outputs(1627) <= a xor b;
    layer6_outputs(1628) <= a and b;
    layer6_outputs(1629) <= a or b;
    layer6_outputs(1630) <= a;
    layer6_outputs(1631) <= a;
    layer6_outputs(1632) <= a and b;
    layer6_outputs(1633) <= not (a xor b);
    layer6_outputs(1634) <= not (a xor b);
    layer6_outputs(1635) <= not a;
    layer6_outputs(1636) <= a xor b;
    layer6_outputs(1637) <= b and not a;
    layer6_outputs(1638) <= a and not b;
    layer6_outputs(1639) <= not (a or b);
    layer6_outputs(1640) <= b;
    layer6_outputs(1641) <= a;
    layer6_outputs(1642) <= not (a and b);
    layer6_outputs(1643) <= not a or b;
    layer6_outputs(1644) <= a;
    layer6_outputs(1645) <= a xor b;
    layer6_outputs(1646) <= not b;
    layer6_outputs(1647) <= not (a xor b);
    layer6_outputs(1648) <= not a;
    layer6_outputs(1649) <= a;
    layer6_outputs(1650) <= not a;
    layer6_outputs(1651) <= not b;
    layer6_outputs(1652) <= not (a and b);
    layer6_outputs(1653) <= not b;
    layer6_outputs(1654) <= a and not b;
    layer6_outputs(1655) <= a xor b;
    layer6_outputs(1656) <= not a;
    layer6_outputs(1657) <= not (a xor b);
    layer6_outputs(1658) <= not b or a;
    layer6_outputs(1659) <= b and not a;
    layer6_outputs(1660) <= b;
    layer6_outputs(1661) <= not a;
    layer6_outputs(1662) <= not a;
    layer6_outputs(1663) <= a;
    layer6_outputs(1664) <= not b;
    layer6_outputs(1665) <= a;
    layer6_outputs(1666) <= not a;
    layer6_outputs(1667) <= not a;
    layer6_outputs(1668) <= b;
    layer6_outputs(1669) <= b and not a;
    layer6_outputs(1670) <= not (a or b);
    layer6_outputs(1671) <= not a;
    layer6_outputs(1672) <= a and not b;
    layer6_outputs(1673) <= b;
    layer6_outputs(1674) <= not b;
    layer6_outputs(1675) <= a xor b;
    layer6_outputs(1676) <= a;
    layer6_outputs(1677) <= not (a xor b);
    layer6_outputs(1678) <= b;
    layer6_outputs(1679) <= a xor b;
    layer6_outputs(1680) <= b;
    layer6_outputs(1681) <= not a;
    layer6_outputs(1682) <= a xor b;
    layer6_outputs(1683) <= b and not a;
    layer6_outputs(1684) <= a or b;
    layer6_outputs(1685) <= a or b;
    layer6_outputs(1686) <= a;
    layer6_outputs(1687) <= not b;
    layer6_outputs(1688) <= not (a xor b);
    layer6_outputs(1689) <= a and not b;
    layer6_outputs(1690) <= not (a xor b);
    layer6_outputs(1691) <= not b;
    layer6_outputs(1692) <= a xor b;
    layer6_outputs(1693) <= a xor b;
    layer6_outputs(1694) <= b and not a;
    layer6_outputs(1695) <= not (a xor b);
    layer6_outputs(1696) <= a and b;
    layer6_outputs(1697) <= a xor b;
    layer6_outputs(1698) <= a or b;
    layer6_outputs(1699) <= a;
    layer6_outputs(1700) <= not a;
    layer6_outputs(1701) <= a and b;
    layer6_outputs(1702) <= not b;
    layer6_outputs(1703) <= not b;
    layer6_outputs(1704) <= a xor b;
    layer6_outputs(1705) <= not b;
    layer6_outputs(1706) <= not b;
    layer6_outputs(1707) <= a xor b;
    layer6_outputs(1708) <= not (a xor b);
    layer6_outputs(1709) <= not b;
    layer6_outputs(1710) <= a;
    layer6_outputs(1711) <= not (a xor b);
    layer6_outputs(1712) <= not (a xor b);
    layer6_outputs(1713) <= a xor b;
    layer6_outputs(1714) <= a;
    layer6_outputs(1715) <= not b;
    layer6_outputs(1716) <= a and not b;
    layer6_outputs(1717) <= not b;
    layer6_outputs(1718) <= a xor b;
    layer6_outputs(1719) <= '0';
    layer6_outputs(1720) <= b;
    layer6_outputs(1721) <= not a;
    layer6_outputs(1722) <= b and not a;
    layer6_outputs(1723) <= not b or a;
    layer6_outputs(1724) <= a;
    layer6_outputs(1725) <= not b;
    layer6_outputs(1726) <= a xor b;
    layer6_outputs(1727) <= a;
    layer6_outputs(1728) <= a xor b;
    layer6_outputs(1729) <= b;
    layer6_outputs(1730) <= not b;
    layer6_outputs(1731) <= not a or b;
    layer6_outputs(1732) <= not a or b;
    layer6_outputs(1733) <= not b or a;
    layer6_outputs(1734) <= not a;
    layer6_outputs(1735) <= not b;
    layer6_outputs(1736) <= a;
    layer6_outputs(1737) <= a;
    layer6_outputs(1738) <= a;
    layer6_outputs(1739) <= a;
    layer6_outputs(1740) <= a;
    layer6_outputs(1741) <= a and not b;
    layer6_outputs(1742) <= not (a xor b);
    layer6_outputs(1743) <= not b;
    layer6_outputs(1744) <= not b;
    layer6_outputs(1745) <= not (a or b);
    layer6_outputs(1746) <= not b or a;
    layer6_outputs(1747) <= not a;
    layer6_outputs(1748) <= not a;
    layer6_outputs(1749) <= a xor b;
    layer6_outputs(1750) <= not (a or b);
    layer6_outputs(1751) <= a;
    layer6_outputs(1752) <= not a;
    layer6_outputs(1753) <= a;
    layer6_outputs(1754) <= a xor b;
    layer6_outputs(1755) <= not (a or b);
    layer6_outputs(1756) <= a xor b;
    layer6_outputs(1757) <= not b;
    layer6_outputs(1758) <= a;
    layer6_outputs(1759) <= not a;
    layer6_outputs(1760) <= a or b;
    layer6_outputs(1761) <= a xor b;
    layer6_outputs(1762) <= b;
    layer6_outputs(1763) <= a xor b;
    layer6_outputs(1764) <= a xor b;
    layer6_outputs(1765) <= not (a xor b);
    layer6_outputs(1766) <= b;
    layer6_outputs(1767) <= not a;
    layer6_outputs(1768) <= b;
    layer6_outputs(1769) <= a;
    layer6_outputs(1770) <= not (a xor b);
    layer6_outputs(1771) <= not b or a;
    layer6_outputs(1772) <= a xor b;
    layer6_outputs(1773) <= not a;
    layer6_outputs(1774) <= not b;
    layer6_outputs(1775) <= a;
    layer6_outputs(1776) <= not a;
    layer6_outputs(1777) <= not b;
    layer6_outputs(1778) <= not a;
    layer6_outputs(1779) <= a xor b;
    layer6_outputs(1780) <= a xor b;
    layer6_outputs(1781) <= not (a xor b);
    layer6_outputs(1782) <= not b;
    layer6_outputs(1783) <= not (a xor b);
    layer6_outputs(1784) <= not a;
    layer6_outputs(1785) <= b and not a;
    layer6_outputs(1786) <= not b;
    layer6_outputs(1787) <= not a or b;
    layer6_outputs(1788) <= a xor b;
    layer6_outputs(1789) <= b;
    layer6_outputs(1790) <= not b;
    layer6_outputs(1791) <= not a or b;
    layer6_outputs(1792) <= not (a xor b);
    layer6_outputs(1793) <= not (a xor b);
    layer6_outputs(1794) <= a and not b;
    layer6_outputs(1795) <= a xor b;
    layer6_outputs(1796) <= not a;
    layer6_outputs(1797) <= not b or a;
    layer6_outputs(1798) <= not a;
    layer6_outputs(1799) <= a;
    layer6_outputs(1800) <= b;
    layer6_outputs(1801) <= not (a xor b);
    layer6_outputs(1802) <= a and not b;
    layer6_outputs(1803) <= a or b;
    layer6_outputs(1804) <= a xor b;
    layer6_outputs(1805) <= a;
    layer6_outputs(1806) <= not a;
    layer6_outputs(1807) <= a;
    layer6_outputs(1808) <= not b or a;
    layer6_outputs(1809) <= a and b;
    layer6_outputs(1810) <= not a or b;
    layer6_outputs(1811) <= b;
    layer6_outputs(1812) <= b;
    layer6_outputs(1813) <= a xor b;
    layer6_outputs(1814) <= a xor b;
    layer6_outputs(1815) <= b;
    layer6_outputs(1816) <= a;
    layer6_outputs(1817) <= not b or a;
    layer6_outputs(1818) <= a xor b;
    layer6_outputs(1819) <= b and not a;
    layer6_outputs(1820) <= not (a and b);
    layer6_outputs(1821) <= a;
    layer6_outputs(1822) <= not a or b;
    layer6_outputs(1823) <= not a;
    layer6_outputs(1824) <= b;
    layer6_outputs(1825) <= a xor b;
    layer6_outputs(1826) <= a;
    layer6_outputs(1827) <= a and b;
    layer6_outputs(1828) <= not a or b;
    layer6_outputs(1829) <= b;
    layer6_outputs(1830) <= not (a and b);
    layer6_outputs(1831) <= a and not b;
    layer6_outputs(1832) <= not a;
    layer6_outputs(1833) <= not a;
    layer6_outputs(1834) <= a and not b;
    layer6_outputs(1835) <= not (a and b);
    layer6_outputs(1836) <= a xor b;
    layer6_outputs(1837) <= a xor b;
    layer6_outputs(1838) <= not b or a;
    layer6_outputs(1839) <= not (a xor b);
    layer6_outputs(1840) <= not a;
    layer6_outputs(1841) <= not (a xor b);
    layer6_outputs(1842) <= a and not b;
    layer6_outputs(1843) <= not a;
    layer6_outputs(1844) <= not (a xor b);
    layer6_outputs(1845) <= not (a or b);
    layer6_outputs(1846) <= a or b;
    layer6_outputs(1847) <= not b or a;
    layer6_outputs(1848) <= b and not a;
    layer6_outputs(1849) <= not (a and b);
    layer6_outputs(1850) <= a;
    layer6_outputs(1851) <= not b or a;
    layer6_outputs(1852) <= not (a xor b);
    layer6_outputs(1853) <= b;
    layer6_outputs(1854) <= not (a xor b);
    layer6_outputs(1855) <= b;
    layer6_outputs(1856) <= not a;
    layer6_outputs(1857) <= not b;
    layer6_outputs(1858) <= not (a xor b);
    layer6_outputs(1859) <= not a;
    layer6_outputs(1860) <= a and not b;
    layer6_outputs(1861) <= b;
    layer6_outputs(1862) <= b;
    layer6_outputs(1863) <= not a or b;
    layer6_outputs(1864) <= not (a xor b);
    layer6_outputs(1865) <= b and not a;
    layer6_outputs(1866) <= not a;
    layer6_outputs(1867) <= not (a and b);
    layer6_outputs(1868) <= not b;
    layer6_outputs(1869) <= a;
    layer6_outputs(1870) <= a;
    layer6_outputs(1871) <= b and not a;
    layer6_outputs(1872) <= not a;
    layer6_outputs(1873) <= not b;
    layer6_outputs(1874) <= a or b;
    layer6_outputs(1875) <= a xor b;
    layer6_outputs(1876) <= not (a and b);
    layer6_outputs(1877) <= a and not b;
    layer6_outputs(1878) <= not a;
    layer6_outputs(1879) <= not b or a;
    layer6_outputs(1880) <= a and not b;
    layer6_outputs(1881) <= a and not b;
    layer6_outputs(1882) <= a and b;
    layer6_outputs(1883) <= not a;
    layer6_outputs(1884) <= a xor b;
    layer6_outputs(1885) <= not a or b;
    layer6_outputs(1886) <= b and not a;
    layer6_outputs(1887) <= b;
    layer6_outputs(1888) <= not b;
    layer6_outputs(1889) <= a and b;
    layer6_outputs(1890) <= not a;
    layer6_outputs(1891) <= not (a or b);
    layer6_outputs(1892) <= not b;
    layer6_outputs(1893) <= a or b;
    layer6_outputs(1894) <= not (a and b);
    layer6_outputs(1895) <= not a;
    layer6_outputs(1896) <= a and not b;
    layer6_outputs(1897) <= not (a xor b);
    layer6_outputs(1898) <= not (a xor b);
    layer6_outputs(1899) <= b;
    layer6_outputs(1900) <= not (a xor b);
    layer6_outputs(1901) <= not b;
    layer6_outputs(1902) <= not b or a;
    layer6_outputs(1903) <= not a or b;
    layer6_outputs(1904) <= not b or a;
    layer6_outputs(1905) <= b;
    layer6_outputs(1906) <= a xor b;
    layer6_outputs(1907) <= not (a and b);
    layer6_outputs(1908) <= not b or a;
    layer6_outputs(1909) <= not a;
    layer6_outputs(1910) <= a;
    layer6_outputs(1911) <= not (a and b);
    layer6_outputs(1912) <= a xor b;
    layer6_outputs(1913) <= a;
    layer6_outputs(1914) <= b;
    layer6_outputs(1915) <= a and not b;
    layer6_outputs(1916) <= not (a or b);
    layer6_outputs(1917) <= b;
    layer6_outputs(1918) <= not (a or b);
    layer6_outputs(1919) <= a;
    layer6_outputs(1920) <= not a;
    layer6_outputs(1921) <= not b;
    layer6_outputs(1922) <= b;
    layer6_outputs(1923) <= a;
    layer6_outputs(1924) <= not a;
    layer6_outputs(1925) <= b and not a;
    layer6_outputs(1926) <= a;
    layer6_outputs(1927) <= not b or a;
    layer6_outputs(1928) <= not (a xor b);
    layer6_outputs(1929) <= a xor b;
    layer6_outputs(1930) <= not b;
    layer6_outputs(1931) <= not a;
    layer6_outputs(1932) <= not (a xor b);
    layer6_outputs(1933) <= not (a and b);
    layer6_outputs(1934) <= b and not a;
    layer6_outputs(1935) <= b and not a;
    layer6_outputs(1936) <= not (a xor b);
    layer6_outputs(1937) <= not a;
    layer6_outputs(1938) <= a xor b;
    layer6_outputs(1939) <= a xor b;
    layer6_outputs(1940) <= not a;
    layer6_outputs(1941) <= a and b;
    layer6_outputs(1942) <= not a;
    layer6_outputs(1943) <= not b or a;
    layer6_outputs(1944) <= not a;
    layer6_outputs(1945) <= b;
    layer6_outputs(1946) <= not (a xor b);
    layer6_outputs(1947) <= not b or a;
    layer6_outputs(1948) <= '0';
    layer6_outputs(1949) <= not b or a;
    layer6_outputs(1950) <= b;
    layer6_outputs(1951) <= not (a or b);
    layer6_outputs(1952) <= not (a and b);
    layer6_outputs(1953) <= a xor b;
    layer6_outputs(1954) <= b;
    layer6_outputs(1955) <= a;
    layer6_outputs(1956) <= not (a or b);
    layer6_outputs(1957) <= not a;
    layer6_outputs(1958) <= a;
    layer6_outputs(1959) <= not b;
    layer6_outputs(1960) <= a and b;
    layer6_outputs(1961) <= a or b;
    layer6_outputs(1962) <= a or b;
    layer6_outputs(1963) <= not b;
    layer6_outputs(1964) <= a;
    layer6_outputs(1965) <= not a or b;
    layer6_outputs(1966) <= a and not b;
    layer6_outputs(1967) <= a or b;
    layer6_outputs(1968) <= not a;
    layer6_outputs(1969) <= not b or a;
    layer6_outputs(1970) <= a;
    layer6_outputs(1971) <= not a;
    layer6_outputs(1972) <= a;
    layer6_outputs(1973) <= a;
    layer6_outputs(1974) <= a or b;
    layer6_outputs(1975) <= b and not a;
    layer6_outputs(1976) <= '1';
    layer6_outputs(1977) <= a and not b;
    layer6_outputs(1978) <= a and not b;
    layer6_outputs(1979) <= a xor b;
    layer6_outputs(1980) <= not (a and b);
    layer6_outputs(1981) <= not a;
    layer6_outputs(1982) <= a and b;
    layer6_outputs(1983) <= not (a and b);
    layer6_outputs(1984) <= not a;
    layer6_outputs(1985) <= b;
    layer6_outputs(1986) <= a and not b;
    layer6_outputs(1987) <= a;
    layer6_outputs(1988) <= b;
    layer6_outputs(1989) <= not a;
    layer6_outputs(1990) <= a and not b;
    layer6_outputs(1991) <= not (a and b);
    layer6_outputs(1992) <= not b;
    layer6_outputs(1993) <= a xor b;
    layer6_outputs(1994) <= not a;
    layer6_outputs(1995) <= not a or b;
    layer6_outputs(1996) <= not a;
    layer6_outputs(1997) <= b and not a;
    layer6_outputs(1998) <= a xor b;
    layer6_outputs(1999) <= a;
    layer6_outputs(2000) <= b;
    layer6_outputs(2001) <= not b or a;
    layer6_outputs(2002) <= not b or a;
    layer6_outputs(2003) <= a;
    layer6_outputs(2004) <= not (a xor b);
    layer6_outputs(2005) <= not a or b;
    layer6_outputs(2006) <= a;
    layer6_outputs(2007) <= not b;
    layer6_outputs(2008) <= not a;
    layer6_outputs(2009) <= a xor b;
    layer6_outputs(2010) <= a;
    layer6_outputs(2011) <= a xor b;
    layer6_outputs(2012) <= not b or a;
    layer6_outputs(2013) <= a;
    layer6_outputs(2014) <= a or b;
    layer6_outputs(2015) <= not a;
    layer6_outputs(2016) <= not b;
    layer6_outputs(2017) <= a;
    layer6_outputs(2018) <= b;
    layer6_outputs(2019) <= not (a xor b);
    layer6_outputs(2020) <= not (a or b);
    layer6_outputs(2021) <= a and b;
    layer6_outputs(2022) <= not (a and b);
    layer6_outputs(2023) <= not (a and b);
    layer6_outputs(2024) <= b;
    layer6_outputs(2025) <= a or b;
    layer6_outputs(2026) <= a or b;
    layer6_outputs(2027) <= a xor b;
    layer6_outputs(2028) <= not b or a;
    layer6_outputs(2029) <= a xor b;
    layer6_outputs(2030) <= b;
    layer6_outputs(2031) <= b and not a;
    layer6_outputs(2032) <= not a or b;
    layer6_outputs(2033) <= not (a xor b);
    layer6_outputs(2034) <= a xor b;
    layer6_outputs(2035) <= a xor b;
    layer6_outputs(2036) <= b;
    layer6_outputs(2037) <= not (a or b);
    layer6_outputs(2038) <= not b or a;
    layer6_outputs(2039) <= b;
    layer6_outputs(2040) <= a xor b;
    layer6_outputs(2041) <= not b or a;
    layer6_outputs(2042) <= a xor b;
    layer6_outputs(2043) <= a xor b;
    layer6_outputs(2044) <= a;
    layer6_outputs(2045) <= not (a and b);
    layer6_outputs(2046) <= a and b;
    layer6_outputs(2047) <= not (a and b);
    layer6_outputs(2048) <= a;
    layer6_outputs(2049) <= b;
    layer6_outputs(2050) <= b;
    layer6_outputs(2051) <= not b or a;
    layer6_outputs(2052) <= not b;
    layer6_outputs(2053) <= not b;
    layer6_outputs(2054) <= a or b;
    layer6_outputs(2055) <= not a;
    layer6_outputs(2056) <= a or b;
    layer6_outputs(2057) <= not b;
    layer6_outputs(2058) <= a xor b;
    layer6_outputs(2059) <= a;
    layer6_outputs(2060) <= not b;
    layer6_outputs(2061) <= a and b;
    layer6_outputs(2062) <= not a;
    layer6_outputs(2063) <= not (a and b);
    layer6_outputs(2064) <= b;
    layer6_outputs(2065) <= a or b;
    layer6_outputs(2066) <= a or b;
    layer6_outputs(2067) <= not a or b;
    layer6_outputs(2068) <= not (a and b);
    layer6_outputs(2069) <= b;
    layer6_outputs(2070) <= not (a xor b);
    layer6_outputs(2071) <= not (a and b);
    layer6_outputs(2072) <= not a;
    layer6_outputs(2073) <= not b or a;
    layer6_outputs(2074) <= not b;
    layer6_outputs(2075) <= a or b;
    layer6_outputs(2076) <= a;
    layer6_outputs(2077) <= b and not a;
    layer6_outputs(2078) <= a xor b;
    layer6_outputs(2079) <= not a;
    layer6_outputs(2080) <= not b;
    layer6_outputs(2081) <= not b;
    layer6_outputs(2082) <= not b or a;
    layer6_outputs(2083) <= b;
    layer6_outputs(2084) <= a or b;
    layer6_outputs(2085) <= not a or b;
    layer6_outputs(2086) <= not (a or b);
    layer6_outputs(2087) <= not (a xor b);
    layer6_outputs(2088) <= not (a or b);
    layer6_outputs(2089) <= not a;
    layer6_outputs(2090) <= a;
    layer6_outputs(2091) <= a and not b;
    layer6_outputs(2092) <= not a;
    layer6_outputs(2093) <= not b;
    layer6_outputs(2094) <= not a;
    layer6_outputs(2095) <= a xor b;
    layer6_outputs(2096) <= not b;
    layer6_outputs(2097) <= not (a or b);
    layer6_outputs(2098) <= b and not a;
    layer6_outputs(2099) <= b;
    layer6_outputs(2100) <= a or b;
    layer6_outputs(2101) <= not b;
    layer6_outputs(2102) <= not a;
    layer6_outputs(2103) <= a xor b;
    layer6_outputs(2104) <= a xor b;
    layer6_outputs(2105) <= not b or a;
    layer6_outputs(2106) <= not a;
    layer6_outputs(2107) <= not b;
    layer6_outputs(2108) <= b and not a;
    layer6_outputs(2109) <= a;
    layer6_outputs(2110) <= not (a and b);
    layer6_outputs(2111) <= not (a and b);
    layer6_outputs(2112) <= a;
    layer6_outputs(2113) <= not b;
    layer6_outputs(2114) <= not (a xor b);
    layer6_outputs(2115) <= not a or b;
    layer6_outputs(2116) <= a;
    layer6_outputs(2117) <= a or b;
    layer6_outputs(2118) <= b;
    layer6_outputs(2119) <= not (a xor b);
    layer6_outputs(2120) <= b;
    layer6_outputs(2121) <= not (a xor b);
    layer6_outputs(2122) <= not (a and b);
    layer6_outputs(2123) <= a or b;
    layer6_outputs(2124) <= not (a xor b);
    layer6_outputs(2125) <= b;
    layer6_outputs(2126) <= not a;
    layer6_outputs(2127) <= not b;
    layer6_outputs(2128) <= a xor b;
    layer6_outputs(2129) <= a;
    layer6_outputs(2130) <= b;
    layer6_outputs(2131) <= a and b;
    layer6_outputs(2132) <= not b;
    layer6_outputs(2133) <= b and not a;
    layer6_outputs(2134) <= b and not a;
    layer6_outputs(2135) <= not a or b;
    layer6_outputs(2136) <= b;
    layer6_outputs(2137) <= not a;
    layer6_outputs(2138) <= not (a xor b);
    layer6_outputs(2139) <= not b or a;
    layer6_outputs(2140) <= a and b;
    layer6_outputs(2141) <= a;
    layer6_outputs(2142) <= not b;
    layer6_outputs(2143) <= not b or a;
    layer6_outputs(2144) <= a xor b;
    layer6_outputs(2145) <= a and not b;
    layer6_outputs(2146) <= '0';
    layer6_outputs(2147) <= b;
    layer6_outputs(2148) <= b;
    layer6_outputs(2149) <= a and b;
    layer6_outputs(2150) <= '0';
    layer6_outputs(2151) <= b and not a;
    layer6_outputs(2152) <= not (a and b);
    layer6_outputs(2153) <= a xor b;
    layer6_outputs(2154) <= b;
    layer6_outputs(2155) <= not a;
    layer6_outputs(2156) <= not b or a;
    layer6_outputs(2157) <= not b;
    layer6_outputs(2158) <= a and b;
    layer6_outputs(2159) <= a;
    layer6_outputs(2160) <= b and not a;
    layer6_outputs(2161) <= b;
    layer6_outputs(2162) <= a;
    layer6_outputs(2163) <= a;
    layer6_outputs(2164) <= not (a xor b);
    layer6_outputs(2165) <= not a;
    layer6_outputs(2166) <= a;
    layer6_outputs(2167) <= '1';
    layer6_outputs(2168) <= a xor b;
    layer6_outputs(2169) <= not (a and b);
    layer6_outputs(2170) <= not b or a;
    layer6_outputs(2171) <= not (a xor b);
    layer6_outputs(2172) <= a and not b;
    layer6_outputs(2173) <= not b;
    layer6_outputs(2174) <= b;
    layer6_outputs(2175) <= a and b;
    layer6_outputs(2176) <= a;
    layer6_outputs(2177) <= a xor b;
    layer6_outputs(2178) <= a and b;
    layer6_outputs(2179) <= a and b;
    layer6_outputs(2180) <= not b;
    layer6_outputs(2181) <= a;
    layer6_outputs(2182) <= b;
    layer6_outputs(2183) <= b;
    layer6_outputs(2184) <= not (a xor b);
    layer6_outputs(2185) <= a xor b;
    layer6_outputs(2186) <= a;
    layer6_outputs(2187) <= not a;
    layer6_outputs(2188) <= not a;
    layer6_outputs(2189) <= a or b;
    layer6_outputs(2190) <= a xor b;
    layer6_outputs(2191) <= not a or b;
    layer6_outputs(2192) <= not b;
    layer6_outputs(2193) <= a or b;
    layer6_outputs(2194) <= not a;
    layer6_outputs(2195) <= a;
    layer6_outputs(2196) <= not a;
    layer6_outputs(2197) <= a and b;
    layer6_outputs(2198) <= a;
    layer6_outputs(2199) <= not (a xor b);
    layer6_outputs(2200) <= not a;
    layer6_outputs(2201) <= a xor b;
    layer6_outputs(2202) <= not b;
    layer6_outputs(2203) <= b and not a;
    layer6_outputs(2204) <= not (a and b);
    layer6_outputs(2205) <= not (a xor b);
    layer6_outputs(2206) <= not (a xor b);
    layer6_outputs(2207) <= a or b;
    layer6_outputs(2208) <= a;
    layer6_outputs(2209) <= a and not b;
    layer6_outputs(2210) <= not a;
    layer6_outputs(2211) <= not a;
    layer6_outputs(2212) <= not (a and b);
    layer6_outputs(2213) <= a xor b;
    layer6_outputs(2214) <= b;
    layer6_outputs(2215) <= not a;
    layer6_outputs(2216) <= a;
    layer6_outputs(2217) <= not a or b;
    layer6_outputs(2218) <= not a;
    layer6_outputs(2219) <= a;
    layer6_outputs(2220) <= not a;
    layer6_outputs(2221) <= a and b;
    layer6_outputs(2222) <= a and b;
    layer6_outputs(2223) <= b;
    layer6_outputs(2224) <= not b;
    layer6_outputs(2225) <= not a;
    layer6_outputs(2226) <= not b;
    layer6_outputs(2227) <= not (a and b);
    layer6_outputs(2228) <= not b;
    layer6_outputs(2229) <= a xor b;
    layer6_outputs(2230) <= a;
    layer6_outputs(2231) <= not a;
    layer6_outputs(2232) <= not b;
    layer6_outputs(2233) <= not (a xor b);
    layer6_outputs(2234) <= not a;
    layer6_outputs(2235) <= not a;
    layer6_outputs(2236) <= not (a or b);
    layer6_outputs(2237) <= a xor b;
    layer6_outputs(2238) <= b;
    layer6_outputs(2239) <= a xor b;
    layer6_outputs(2240) <= a;
    layer6_outputs(2241) <= not (a and b);
    layer6_outputs(2242) <= a xor b;
    layer6_outputs(2243) <= b and not a;
    layer6_outputs(2244) <= not a;
    layer6_outputs(2245) <= a xor b;
    layer6_outputs(2246) <= b;
    layer6_outputs(2247) <= not (a xor b);
    layer6_outputs(2248) <= not b;
    layer6_outputs(2249) <= not (a or b);
    layer6_outputs(2250) <= not (a xor b);
    layer6_outputs(2251) <= not (a xor b);
    layer6_outputs(2252) <= a and b;
    layer6_outputs(2253) <= not a or b;
    layer6_outputs(2254) <= not b or a;
    layer6_outputs(2255) <= not (a or b);
    layer6_outputs(2256) <= not a;
    layer6_outputs(2257) <= not (a or b);
    layer6_outputs(2258) <= not b;
    layer6_outputs(2259) <= not b or a;
    layer6_outputs(2260) <= not b;
    layer6_outputs(2261) <= not a;
    layer6_outputs(2262) <= a xor b;
    layer6_outputs(2263) <= a or b;
    layer6_outputs(2264) <= not a or b;
    layer6_outputs(2265) <= not (a or b);
    layer6_outputs(2266) <= not (a or b);
    layer6_outputs(2267) <= not b;
    layer6_outputs(2268) <= a and not b;
    layer6_outputs(2269) <= not (a xor b);
    layer6_outputs(2270) <= a;
    layer6_outputs(2271) <= a and not b;
    layer6_outputs(2272) <= not a;
    layer6_outputs(2273) <= a and not b;
    layer6_outputs(2274) <= not b;
    layer6_outputs(2275) <= b;
    layer6_outputs(2276) <= not (a xor b);
    layer6_outputs(2277) <= not b;
    layer6_outputs(2278) <= a;
    layer6_outputs(2279) <= a;
    layer6_outputs(2280) <= not b or a;
    layer6_outputs(2281) <= b and not a;
    layer6_outputs(2282) <= a or b;
    layer6_outputs(2283) <= not b;
    layer6_outputs(2284) <= not a;
    layer6_outputs(2285) <= not a;
    layer6_outputs(2286) <= not (a and b);
    layer6_outputs(2287) <= not b;
    layer6_outputs(2288) <= a xor b;
    layer6_outputs(2289) <= not a;
    layer6_outputs(2290) <= not b;
    layer6_outputs(2291) <= not b;
    layer6_outputs(2292) <= a or b;
    layer6_outputs(2293) <= '0';
    layer6_outputs(2294) <= not b;
    layer6_outputs(2295) <= not a or b;
    layer6_outputs(2296) <= a;
    layer6_outputs(2297) <= a and not b;
    layer6_outputs(2298) <= b and not a;
    layer6_outputs(2299) <= a and b;
    layer6_outputs(2300) <= not a or b;
    layer6_outputs(2301) <= a xor b;
    layer6_outputs(2302) <= not b;
    layer6_outputs(2303) <= not b;
    layer6_outputs(2304) <= a;
    layer6_outputs(2305) <= not a;
    layer6_outputs(2306) <= a and not b;
    layer6_outputs(2307) <= a;
    layer6_outputs(2308) <= a xor b;
    layer6_outputs(2309) <= not b;
    layer6_outputs(2310) <= not a or b;
    layer6_outputs(2311) <= not (a or b);
    layer6_outputs(2312) <= not a;
    layer6_outputs(2313) <= a and b;
    layer6_outputs(2314) <= not (a xor b);
    layer6_outputs(2315) <= not b or a;
    layer6_outputs(2316) <= a;
    layer6_outputs(2317) <= b and not a;
    layer6_outputs(2318) <= not (a or b);
    layer6_outputs(2319) <= not (a or b);
    layer6_outputs(2320) <= not a;
    layer6_outputs(2321) <= not b;
    layer6_outputs(2322) <= not a;
    layer6_outputs(2323) <= b and not a;
    layer6_outputs(2324) <= a;
    layer6_outputs(2325) <= a;
    layer6_outputs(2326) <= not b;
    layer6_outputs(2327) <= a;
    layer6_outputs(2328) <= a;
    layer6_outputs(2329) <= a and b;
    layer6_outputs(2330) <= b;
    layer6_outputs(2331) <= not a;
    layer6_outputs(2332) <= b;
    layer6_outputs(2333) <= not a;
    layer6_outputs(2334) <= a;
    layer6_outputs(2335) <= b and not a;
    layer6_outputs(2336) <= not a or b;
    layer6_outputs(2337) <= a;
    layer6_outputs(2338) <= a;
    layer6_outputs(2339) <= a xor b;
    layer6_outputs(2340) <= a;
    layer6_outputs(2341) <= b;
    layer6_outputs(2342) <= not b;
    layer6_outputs(2343) <= not a or b;
    layer6_outputs(2344) <= a and not b;
    layer6_outputs(2345) <= not b;
    layer6_outputs(2346) <= not b;
    layer6_outputs(2347) <= not b;
    layer6_outputs(2348) <= b and not a;
    layer6_outputs(2349) <= not a;
    layer6_outputs(2350) <= not a;
    layer6_outputs(2351) <= not b;
    layer6_outputs(2352) <= '0';
    layer6_outputs(2353) <= not a or b;
    layer6_outputs(2354) <= b;
    layer6_outputs(2355) <= a and b;
    layer6_outputs(2356) <= not a or b;
    layer6_outputs(2357) <= b;
    layer6_outputs(2358) <= a;
    layer6_outputs(2359) <= not b;
    layer6_outputs(2360) <= not b;
    layer6_outputs(2361) <= a xor b;
    layer6_outputs(2362) <= not (a xor b);
    layer6_outputs(2363) <= a;
    layer6_outputs(2364) <= not (a xor b);
    layer6_outputs(2365) <= not b;
    layer6_outputs(2366) <= not (a xor b);
    layer6_outputs(2367) <= '0';
    layer6_outputs(2368) <= not a;
    layer6_outputs(2369) <= a and not b;
    layer6_outputs(2370) <= not b;
    layer6_outputs(2371) <= a and not b;
    layer6_outputs(2372) <= not (a xor b);
    layer6_outputs(2373) <= not b;
    layer6_outputs(2374) <= a;
    layer6_outputs(2375) <= a and b;
    layer6_outputs(2376) <= a xor b;
    layer6_outputs(2377) <= b;
    layer6_outputs(2378) <= a;
    layer6_outputs(2379) <= not (a xor b);
    layer6_outputs(2380) <= not (a xor b);
    layer6_outputs(2381) <= a and b;
    layer6_outputs(2382) <= a and b;
    layer6_outputs(2383) <= b;
    layer6_outputs(2384) <= a;
    layer6_outputs(2385) <= a;
    layer6_outputs(2386) <= not (a xor b);
    layer6_outputs(2387) <= not b;
    layer6_outputs(2388) <= b;
    layer6_outputs(2389) <= b;
    layer6_outputs(2390) <= not b or a;
    layer6_outputs(2391) <= not a;
    layer6_outputs(2392) <= a;
    layer6_outputs(2393) <= b and not a;
    layer6_outputs(2394) <= a;
    layer6_outputs(2395) <= not b;
    layer6_outputs(2396) <= a;
    layer6_outputs(2397) <= a;
    layer6_outputs(2398) <= not (a or b);
    layer6_outputs(2399) <= not b;
    layer6_outputs(2400) <= not b or a;
    layer6_outputs(2401) <= b;
    layer6_outputs(2402) <= '1';
    layer6_outputs(2403) <= a;
    layer6_outputs(2404) <= a;
    layer6_outputs(2405) <= a or b;
    layer6_outputs(2406) <= a xor b;
    layer6_outputs(2407) <= b and not a;
    layer6_outputs(2408) <= a and b;
    layer6_outputs(2409) <= a or b;
    layer6_outputs(2410) <= not b;
    layer6_outputs(2411) <= not (a or b);
    layer6_outputs(2412) <= not a;
    layer6_outputs(2413) <= b;
    layer6_outputs(2414) <= not (a and b);
    layer6_outputs(2415) <= not b;
    layer6_outputs(2416) <= a and b;
    layer6_outputs(2417) <= a;
    layer6_outputs(2418) <= not (a and b);
    layer6_outputs(2419) <= a;
    layer6_outputs(2420) <= not a;
    layer6_outputs(2421) <= a or b;
    layer6_outputs(2422) <= a;
    layer6_outputs(2423) <= a and not b;
    layer6_outputs(2424) <= not (a or b);
    layer6_outputs(2425) <= a xor b;
    layer6_outputs(2426) <= b;
    layer6_outputs(2427) <= a;
    layer6_outputs(2428) <= not a;
    layer6_outputs(2429) <= not a or b;
    layer6_outputs(2430) <= a and not b;
    layer6_outputs(2431) <= not b or a;
    layer6_outputs(2432) <= a and not b;
    layer6_outputs(2433) <= not a;
    layer6_outputs(2434) <= not (a xor b);
    layer6_outputs(2435) <= a;
    layer6_outputs(2436) <= not a;
    layer6_outputs(2437) <= not b or a;
    layer6_outputs(2438) <= a;
    layer6_outputs(2439) <= not b or a;
    layer6_outputs(2440) <= not b or a;
    layer6_outputs(2441) <= not (a xor b);
    layer6_outputs(2442) <= not (a and b);
    layer6_outputs(2443) <= b and not a;
    layer6_outputs(2444) <= a xor b;
    layer6_outputs(2445) <= b and not a;
    layer6_outputs(2446) <= a;
    layer6_outputs(2447) <= a and not b;
    layer6_outputs(2448) <= not (a xor b);
    layer6_outputs(2449) <= a and b;
    layer6_outputs(2450) <= a and b;
    layer6_outputs(2451) <= a or b;
    layer6_outputs(2452) <= b and not a;
    layer6_outputs(2453) <= a xor b;
    layer6_outputs(2454) <= a xor b;
    layer6_outputs(2455) <= not a;
    layer6_outputs(2456) <= not (a xor b);
    layer6_outputs(2457) <= not a;
    layer6_outputs(2458) <= not a;
    layer6_outputs(2459) <= a or b;
    layer6_outputs(2460) <= not a;
    layer6_outputs(2461) <= not b;
    layer6_outputs(2462) <= b;
    layer6_outputs(2463) <= b;
    layer6_outputs(2464) <= not b;
    layer6_outputs(2465) <= '0';
    layer6_outputs(2466) <= a;
    layer6_outputs(2467) <= not (a xor b);
    layer6_outputs(2468) <= not a;
    layer6_outputs(2469) <= b;
    layer6_outputs(2470) <= b and not a;
    layer6_outputs(2471) <= a xor b;
    layer6_outputs(2472) <= b;
    layer6_outputs(2473) <= a and b;
    layer6_outputs(2474) <= not (a and b);
    layer6_outputs(2475) <= not a;
    layer6_outputs(2476) <= a and not b;
    layer6_outputs(2477) <= not b;
    layer6_outputs(2478) <= a;
    layer6_outputs(2479) <= a and not b;
    layer6_outputs(2480) <= b;
    layer6_outputs(2481) <= not a or b;
    layer6_outputs(2482) <= b;
    layer6_outputs(2483) <= a;
    layer6_outputs(2484) <= not a;
    layer6_outputs(2485) <= not (a and b);
    layer6_outputs(2486) <= b and not a;
    layer6_outputs(2487) <= a or b;
    layer6_outputs(2488) <= not (a xor b);
    layer6_outputs(2489) <= not a;
    layer6_outputs(2490) <= b and not a;
    layer6_outputs(2491) <= not a;
    layer6_outputs(2492) <= not (a xor b);
    layer6_outputs(2493) <= a;
    layer6_outputs(2494) <= not a;
    layer6_outputs(2495) <= '0';
    layer6_outputs(2496) <= not a;
    layer6_outputs(2497) <= b and not a;
    layer6_outputs(2498) <= not (a or b);
    layer6_outputs(2499) <= not a;
    layer6_outputs(2500) <= not b or a;
    layer6_outputs(2501) <= a or b;
    layer6_outputs(2502) <= not a or b;
    layer6_outputs(2503) <= not a or b;
    layer6_outputs(2504) <= not a;
    layer6_outputs(2505) <= not a;
    layer6_outputs(2506) <= not (a xor b);
    layer6_outputs(2507) <= not (a xor b);
    layer6_outputs(2508) <= not (a xor b);
    layer6_outputs(2509) <= not a;
    layer6_outputs(2510) <= a xor b;
    layer6_outputs(2511) <= not a or b;
    layer6_outputs(2512) <= '0';
    layer6_outputs(2513) <= not (a or b);
    layer6_outputs(2514) <= not b;
    layer6_outputs(2515) <= not a;
    layer6_outputs(2516) <= a;
    layer6_outputs(2517) <= a xor b;
    layer6_outputs(2518) <= b;
    layer6_outputs(2519) <= not (a and b);
    layer6_outputs(2520) <= not b or a;
    layer6_outputs(2521) <= not a or b;
    layer6_outputs(2522) <= a;
    layer6_outputs(2523) <= not a;
    layer6_outputs(2524) <= not (a xor b);
    layer6_outputs(2525) <= b;
    layer6_outputs(2526) <= not b;
    layer6_outputs(2527) <= a;
    layer6_outputs(2528) <= not (a xor b);
    layer6_outputs(2529) <= not b or a;
    layer6_outputs(2530) <= a or b;
    layer6_outputs(2531) <= not (a or b);
    layer6_outputs(2532) <= b;
    layer6_outputs(2533) <= a;
    layer6_outputs(2534) <= not (a or b);
    layer6_outputs(2535) <= not (a xor b);
    layer6_outputs(2536) <= a xor b;
    layer6_outputs(2537) <= a xor b;
    layer6_outputs(2538) <= a;
    layer6_outputs(2539) <= not (a or b);
    layer6_outputs(2540) <= not a;
    layer6_outputs(2541) <= not b;
    layer6_outputs(2542) <= not a;
    layer6_outputs(2543) <= not (a or b);
    layer6_outputs(2544) <= a xor b;
    layer6_outputs(2545) <= a or b;
    layer6_outputs(2546) <= not b;
    layer6_outputs(2547) <= not a or b;
    layer6_outputs(2548) <= not (a or b);
    layer6_outputs(2549) <= a;
    layer6_outputs(2550) <= a;
    layer6_outputs(2551) <= not a;
    layer6_outputs(2552) <= not b;
    layer6_outputs(2553) <= not a;
    layer6_outputs(2554) <= a or b;
    layer6_outputs(2555) <= a xor b;
    layer6_outputs(2556) <= not (a xor b);
    layer6_outputs(2557) <= b;
    layer6_outputs(2558) <= a and not b;
    layer6_outputs(2559) <= not b;
    layer6_outputs(2560) <= not (a or b);
    layer6_outputs(2561) <= not b or a;
    layer6_outputs(2562) <= b;
    layer6_outputs(2563) <= a and b;
    layer6_outputs(2564) <= a xor b;
    layer6_outputs(2565) <= b;
    layer6_outputs(2566) <= not (a xor b);
    layer6_outputs(2567) <= a xor b;
    layer6_outputs(2568) <= a xor b;
    layer6_outputs(2569) <= a or b;
    layer6_outputs(2570) <= '1';
    layer6_outputs(2571) <= not a;
    layer6_outputs(2572) <= not (a or b);
    layer6_outputs(2573) <= not b;
    layer6_outputs(2574) <= a xor b;
    layer6_outputs(2575) <= not b;
    layer6_outputs(2576) <= not (a and b);
    layer6_outputs(2577) <= b;
    layer6_outputs(2578) <= not a or b;
    layer6_outputs(2579) <= a and b;
    layer6_outputs(2580) <= a or b;
    layer6_outputs(2581) <= not a;
    layer6_outputs(2582) <= b;
    layer6_outputs(2583) <= not a;
    layer6_outputs(2584) <= a or b;
    layer6_outputs(2585) <= a;
    layer6_outputs(2586) <= '0';
    layer6_outputs(2587) <= not a;
    layer6_outputs(2588) <= not a;
    layer6_outputs(2589) <= a;
    layer6_outputs(2590) <= not a;
    layer6_outputs(2591) <= not b;
    layer6_outputs(2592) <= a and b;
    layer6_outputs(2593) <= a and not b;
    layer6_outputs(2594) <= '1';
    layer6_outputs(2595) <= not (a xor b);
    layer6_outputs(2596) <= a and not b;
    layer6_outputs(2597) <= not b or a;
    layer6_outputs(2598) <= not (a or b);
    layer6_outputs(2599) <= a;
    layer6_outputs(2600) <= a;
    layer6_outputs(2601) <= a xor b;
    layer6_outputs(2602) <= not b;
    layer6_outputs(2603) <= not (a xor b);
    layer6_outputs(2604) <= not b;
    layer6_outputs(2605) <= a xor b;
    layer6_outputs(2606) <= a;
    layer6_outputs(2607) <= b and not a;
    layer6_outputs(2608) <= a and b;
    layer6_outputs(2609) <= b;
    layer6_outputs(2610) <= a;
    layer6_outputs(2611) <= not b;
    layer6_outputs(2612) <= not a or b;
    layer6_outputs(2613) <= not b;
    layer6_outputs(2614) <= b;
    layer6_outputs(2615) <= not (a xor b);
    layer6_outputs(2616) <= not b;
    layer6_outputs(2617) <= b;
    layer6_outputs(2618) <= not b or a;
    layer6_outputs(2619) <= not a;
    layer6_outputs(2620) <= not (a xor b);
    layer6_outputs(2621) <= not a;
    layer6_outputs(2622) <= a;
    layer6_outputs(2623) <= a;
    layer6_outputs(2624) <= not a;
    layer6_outputs(2625) <= a and not b;
    layer6_outputs(2626) <= not a;
    layer6_outputs(2627) <= not (a xor b);
    layer6_outputs(2628) <= a xor b;
    layer6_outputs(2629) <= not b;
    layer6_outputs(2630) <= a;
    layer6_outputs(2631) <= not (a xor b);
    layer6_outputs(2632) <= not a;
    layer6_outputs(2633) <= not b;
    layer6_outputs(2634) <= a;
    layer6_outputs(2635) <= a and b;
    layer6_outputs(2636) <= a or b;
    layer6_outputs(2637) <= b and not a;
    layer6_outputs(2638) <= not a or b;
    layer6_outputs(2639) <= not (a and b);
    layer6_outputs(2640) <= '1';
    layer6_outputs(2641) <= not a or b;
    layer6_outputs(2642) <= a xor b;
    layer6_outputs(2643) <= not (a xor b);
    layer6_outputs(2644) <= not a or b;
    layer6_outputs(2645) <= not b;
    layer6_outputs(2646) <= a xor b;
    layer6_outputs(2647) <= a;
    layer6_outputs(2648) <= not a or b;
    layer6_outputs(2649) <= a xor b;
    layer6_outputs(2650) <= a and not b;
    layer6_outputs(2651) <= a xor b;
    layer6_outputs(2652) <= not (a and b);
    layer6_outputs(2653) <= not b or a;
    layer6_outputs(2654) <= not (a xor b);
    layer6_outputs(2655) <= b;
    layer6_outputs(2656) <= a xor b;
    layer6_outputs(2657) <= not (a or b);
    layer6_outputs(2658) <= b and not a;
    layer6_outputs(2659) <= b;
    layer6_outputs(2660) <= not (a xor b);
    layer6_outputs(2661) <= not a or b;
    layer6_outputs(2662) <= not b;
    layer6_outputs(2663) <= a;
    layer6_outputs(2664) <= a xor b;
    layer6_outputs(2665) <= b;
    layer6_outputs(2666) <= a xor b;
    layer6_outputs(2667) <= not (a xor b);
    layer6_outputs(2668) <= not b;
    layer6_outputs(2669) <= not b;
    layer6_outputs(2670) <= not (a or b);
    layer6_outputs(2671) <= a;
    layer6_outputs(2672) <= not a or b;
    layer6_outputs(2673) <= a xor b;
    layer6_outputs(2674) <= a and b;
    layer6_outputs(2675) <= b;
    layer6_outputs(2676) <= not b;
    layer6_outputs(2677) <= not (a xor b);
    layer6_outputs(2678) <= a and b;
    layer6_outputs(2679) <= a and b;
    layer6_outputs(2680) <= a;
    layer6_outputs(2681) <= b and not a;
    layer6_outputs(2682) <= b and not a;
    layer6_outputs(2683) <= not (a or b);
    layer6_outputs(2684) <= a;
    layer6_outputs(2685) <= a and not b;
    layer6_outputs(2686) <= a;
    layer6_outputs(2687) <= b;
    layer6_outputs(2688) <= not a;
    layer6_outputs(2689) <= a or b;
    layer6_outputs(2690) <= b;
    layer6_outputs(2691) <= a;
    layer6_outputs(2692) <= not (a xor b);
    layer6_outputs(2693) <= not a or b;
    layer6_outputs(2694) <= a or b;
    layer6_outputs(2695) <= not (a or b);
    layer6_outputs(2696) <= a;
    layer6_outputs(2697) <= not (a and b);
    layer6_outputs(2698) <= not (a and b);
    layer6_outputs(2699) <= a or b;
    layer6_outputs(2700) <= b and not a;
    layer6_outputs(2701) <= not b;
    layer6_outputs(2702) <= a xor b;
    layer6_outputs(2703) <= b and not a;
    layer6_outputs(2704) <= not a;
    layer6_outputs(2705) <= a xor b;
    layer6_outputs(2706) <= a xor b;
    layer6_outputs(2707) <= '0';
    layer6_outputs(2708) <= not (a or b);
    layer6_outputs(2709) <= a;
    layer6_outputs(2710) <= a or b;
    layer6_outputs(2711) <= b;
    layer6_outputs(2712) <= not (a or b);
    layer6_outputs(2713) <= not b;
    layer6_outputs(2714) <= b;
    layer6_outputs(2715) <= b;
    layer6_outputs(2716) <= not (a xor b);
    layer6_outputs(2717) <= a and not b;
    layer6_outputs(2718) <= a xor b;
    layer6_outputs(2719) <= a xor b;
    layer6_outputs(2720) <= not b;
    layer6_outputs(2721) <= a or b;
    layer6_outputs(2722) <= not a;
    layer6_outputs(2723) <= not a;
    layer6_outputs(2724) <= not a;
    layer6_outputs(2725) <= not a;
    layer6_outputs(2726) <= a xor b;
    layer6_outputs(2727) <= not b;
    layer6_outputs(2728) <= not a or b;
    layer6_outputs(2729) <= a xor b;
    layer6_outputs(2730) <= '1';
    layer6_outputs(2731) <= a;
    layer6_outputs(2732) <= not a;
    layer6_outputs(2733) <= not (a or b);
    layer6_outputs(2734) <= b;
    layer6_outputs(2735) <= not (a xor b);
    layer6_outputs(2736) <= a;
    layer6_outputs(2737) <= a;
    layer6_outputs(2738) <= not (a and b);
    layer6_outputs(2739) <= not a;
    layer6_outputs(2740) <= not a;
    layer6_outputs(2741) <= a;
    layer6_outputs(2742) <= not (a and b);
    layer6_outputs(2743) <= a xor b;
    layer6_outputs(2744) <= b;
    layer6_outputs(2745) <= a and b;
    layer6_outputs(2746) <= b;
    layer6_outputs(2747) <= a and b;
    layer6_outputs(2748) <= a xor b;
    layer6_outputs(2749) <= b;
    layer6_outputs(2750) <= b and not a;
    layer6_outputs(2751) <= not (a and b);
    layer6_outputs(2752) <= b;
    layer6_outputs(2753) <= a xor b;
    layer6_outputs(2754) <= b and not a;
    layer6_outputs(2755) <= a and b;
    layer6_outputs(2756) <= b and not a;
    layer6_outputs(2757) <= a xor b;
    layer6_outputs(2758) <= a;
    layer6_outputs(2759) <= a;
    layer6_outputs(2760) <= a;
    layer6_outputs(2761) <= a;
    layer6_outputs(2762) <= b;
    layer6_outputs(2763) <= not b;
    layer6_outputs(2764) <= not (a xor b);
    layer6_outputs(2765) <= not a or b;
    layer6_outputs(2766) <= b;
    layer6_outputs(2767) <= b and not a;
    layer6_outputs(2768) <= not b;
    layer6_outputs(2769) <= not (a and b);
    layer6_outputs(2770) <= '1';
    layer6_outputs(2771) <= not a;
    layer6_outputs(2772) <= a and not b;
    layer6_outputs(2773) <= b;
    layer6_outputs(2774) <= a and not b;
    layer6_outputs(2775) <= not a;
    layer6_outputs(2776) <= a and b;
    layer6_outputs(2777) <= a;
    layer6_outputs(2778) <= not (a or b);
    layer6_outputs(2779) <= not a;
    layer6_outputs(2780) <= '1';
    layer6_outputs(2781) <= a and b;
    layer6_outputs(2782) <= a and b;
    layer6_outputs(2783) <= not (a and b);
    layer6_outputs(2784) <= b and not a;
    layer6_outputs(2785) <= not a or b;
    layer6_outputs(2786) <= not (a xor b);
    layer6_outputs(2787) <= not a;
    layer6_outputs(2788) <= '0';
    layer6_outputs(2789) <= a and b;
    layer6_outputs(2790) <= not a or b;
    layer6_outputs(2791) <= not b or a;
    layer6_outputs(2792) <= b;
    layer6_outputs(2793) <= not b;
    layer6_outputs(2794) <= not a or b;
    layer6_outputs(2795) <= a xor b;
    layer6_outputs(2796) <= a and b;
    layer6_outputs(2797) <= not a;
    layer6_outputs(2798) <= not (a or b);
    layer6_outputs(2799) <= not (a or b);
    layer6_outputs(2800) <= a and b;
    layer6_outputs(2801) <= a xor b;
    layer6_outputs(2802) <= not a or b;
    layer6_outputs(2803) <= not b;
    layer6_outputs(2804) <= not a;
    layer6_outputs(2805) <= not (a xor b);
    layer6_outputs(2806) <= not a;
    layer6_outputs(2807) <= a and b;
    layer6_outputs(2808) <= b;
    layer6_outputs(2809) <= not a;
    layer6_outputs(2810) <= a and b;
    layer6_outputs(2811) <= a and b;
    layer6_outputs(2812) <= a or b;
    layer6_outputs(2813) <= b and not a;
    layer6_outputs(2814) <= a xor b;
    layer6_outputs(2815) <= a xor b;
    layer6_outputs(2816) <= not a;
    layer6_outputs(2817) <= not b;
    layer6_outputs(2818) <= a or b;
    layer6_outputs(2819) <= not (a xor b);
    layer6_outputs(2820) <= a and b;
    layer6_outputs(2821) <= not (a xor b);
    layer6_outputs(2822) <= not a;
    layer6_outputs(2823) <= a;
    layer6_outputs(2824) <= a and not b;
    layer6_outputs(2825) <= not b or a;
    layer6_outputs(2826) <= not b;
    layer6_outputs(2827) <= not (a and b);
    layer6_outputs(2828) <= b;
    layer6_outputs(2829) <= not a;
    layer6_outputs(2830) <= a and not b;
    layer6_outputs(2831) <= not b or a;
    layer6_outputs(2832) <= not a;
    layer6_outputs(2833) <= not (a xor b);
    layer6_outputs(2834) <= not a;
    layer6_outputs(2835) <= not a or b;
    layer6_outputs(2836) <= a and b;
    layer6_outputs(2837) <= a xor b;
    layer6_outputs(2838) <= not b or a;
    layer6_outputs(2839) <= not (a and b);
    layer6_outputs(2840) <= not a;
    layer6_outputs(2841) <= a;
    layer6_outputs(2842) <= not (a xor b);
    layer6_outputs(2843) <= not a;
    layer6_outputs(2844) <= b;
    layer6_outputs(2845) <= a and not b;
    layer6_outputs(2846) <= not (a or b);
    layer6_outputs(2847) <= not a;
    layer6_outputs(2848) <= a;
    layer6_outputs(2849) <= not b;
    layer6_outputs(2850) <= not a;
    layer6_outputs(2851) <= not a or b;
    layer6_outputs(2852) <= a;
    layer6_outputs(2853) <= a and b;
    layer6_outputs(2854) <= a or b;
    layer6_outputs(2855) <= not (a xor b);
    layer6_outputs(2856) <= not b;
    layer6_outputs(2857) <= not b;
    layer6_outputs(2858) <= b;
    layer6_outputs(2859) <= a;
    layer6_outputs(2860) <= not (a xor b);
    layer6_outputs(2861) <= not b;
    layer6_outputs(2862) <= a and not b;
    layer6_outputs(2863) <= not (a xor b);
    layer6_outputs(2864) <= a xor b;
    layer6_outputs(2865) <= not b or a;
    layer6_outputs(2866) <= not (a or b);
    layer6_outputs(2867) <= not (a and b);
    layer6_outputs(2868) <= not a or b;
    layer6_outputs(2869) <= not (a xor b);
    layer6_outputs(2870) <= not b;
    layer6_outputs(2871) <= b;
    layer6_outputs(2872) <= not (a and b);
    layer6_outputs(2873) <= not (a xor b);
    layer6_outputs(2874) <= a;
    layer6_outputs(2875) <= a;
    layer6_outputs(2876) <= not a;
    layer6_outputs(2877) <= not (a xor b);
    layer6_outputs(2878) <= not a;
    layer6_outputs(2879) <= a xor b;
    layer6_outputs(2880) <= not (a xor b);
    layer6_outputs(2881) <= not b or a;
    layer6_outputs(2882) <= a and not b;
    layer6_outputs(2883) <= b;
    layer6_outputs(2884) <= not a;
    layer6_outputs(2885) <= not (a xor b);
    layer6_outputs(2886) <= a;
    layer6_outputs(2887) <= not a;
    layer6_outputs(2888) <= not (a and b);
    layer6_outputs(2889) <= b;
    layer6_outputs(2890) <= a;
    layer6_outputs(2891) <= not (a xor b);
    layer6_outputs(2892) <= a;
    layer6_outputs(2893) <= not b;
    layer6_outputs(2894) <= a xor b;
    layer6_outputs(2895) <= not a or b;
    layer6_outputs(2896) <= b;
    layer6_outputs(2897) <= not (a and b);
    layer6_outputs(2898) <= not (a or b);
    layer6_outputs(2899) <= not (a xor b);
    layer6_outputs(2900) <= a xor b;
    layer6_outputs(2901) <= a and b;
    layer6_outputs(2902) <= not a;
    layer6_outputs(2903) <= b and not a;
    layer6_outputs(2904) <= not b;
    layer6_outputs(2905) <= b and not a;
    layer6_outputs(2906) <= not (a or b);
    layer6_outputs(2907) <= not (a or b);
    layer6_outputs(2908) <= not b;
    layer6_outputs(2909) <= not b;
    layer6_outputs(2910) <= b;
    layer6_outputs(2911) <= b;
    layer6_outputs(2912) <= b and not a;
    layer6_outputs(2913) <= not (a or b);
    layer6_outputs(2914) <= a;
    layer6_outputs(2915) <= a xor b;
    layer6_outputs(2916) <= not a or b;
    layer6_outputs(2917) <= not (a and b);
    layer6_outputs(2918) <= not b;
    layer6_outputs(2919) <= not (a xor b);
    layer6_outputs(2920) <= b;
    layer6_outputs(2921) <= a;
    layer6_outputs(2922) <= not (a xor b);
    layer6_outputs(2923) <= a or b;
    layer6_outputs(2924) <= not (a and b);
    layer6_outputs(2925) <= not b;
    layer6_outputs(2926) <= not b or a;
    layer6_outputs(2927) <= a;
    layer6_outputs(2928) <= not b or a;
    layer6_outputs(2929) <= not a or b;
    layer6_outputs(2930) <= not a;
    layer6_outputs(2931) <= a and not b;
    layer6_outputs(2932) <= a and b;
    layer6_outputs(2933) <= '0';
    layer6_outputs(2934) <= not b;
    layer6_outputs(2935) <= b;
    layer6_outputs(2936) <= not (a or b);
    layer6_outputs(2937) <= not a;
    layer6_outputs(2938) <= not (a xor b);
    layer6_outputs(2939) <= not (a and b);
    layer6_outputs(2940) <= not (a xor b);
    layer6_outputs(2941) <= b;
    layer6_outputs(2942) <= b;
    layer6_outputs(2943) <= not (a and b);
    layer6_outputs(2944) <= b;
    layer6_outputs(2945) <= b;
    layer6_outputs(2946) <= not b or a;
    layer6_outputs(2947) <= a;
    layer6_outputs(2948) <= not a;
    layer6_outputs(2949) <= b and not a;
    layer6_outputs(2950) <= not a;
    layer6_outputs(2951) <= a;
    layer6_outputs(2952) <= a xor b;
    layer6_outputs(2953) <= b and not a;
    layer6_outputs(2954) <= not a;
    layer6_outputs(2955) <= b;
    layer6_outputs(2956) <= not b;
    layer6_outputs(2957) <= b;
    layer6_outputs(2958) <= not (a and b);
    layer6_outputs(2959) <= a and not b;
    layer6_outputs(2960) <= a;
    layer6_outputs(2961) <= not a or b;
    layer6_outputs(2962) <= a xor b;
    layer6_outputs(2963) <= b;
    layer6_outputs(2964) <= a or b;
    layer6_outputs(2965) <= not (a xor b);
    layer6_outputs(2966) <= not a or b;
    layer6_outputs(2967) <= b and not a;
    layer6_outputs(2968) <= b;
    layer6_outputs(2969) <= b and not a;
    layer6_outputs(2970) <= a;
    layer6_outputs(2971) <= not b;
    layer6_outputs(2972) <= not (a or b);
    layer6_outputs(2973) <= not b;
    layer6_outputs(2974) <= b;
    layer6_outputs(2975) <= a xor b;
    layer6_outputs(2976) <= not b;
    layer6_outputs(2977) <= not b;
    layer6_outputs(2978) <= a xor b;
    layer6_outputs(2979) <= a and b;
    layer6_outputs(2980) <= a and not b;
    layer6_outputs(2981) <= not (a xor b);
    layer6_outputs(2982) <= a;
    layer6_outputs(2983) <= a;
    layer6_outputs(2984) <= a;
    layer6_outputs(2985) <= a and b;
    layer6_outputs(2986) <= not (a and b);
    layer6_outputs(2987) <= not a;
    layer6_outputs(2988) <= b and not a;
    layer6_outputs(2989) <= b and not a;
    layer6_outputs(2990) <= not (a and b);
    layer6_outputs(2991) <= not b or a;
    layer6_outputs(2992) <= a;
    layer6_outputs(2993) <= a xor b;
    layer6_outputs(2994) <= not a;
    layer6_outputs(2995) <= a;
    layer6_outputs(2996) <= a xor b;
    layer6_outputs(2997) <= a xor b;
    layer6_outputs(2998) <= a or b;
    layer6_outputs(2999) <= not b;
    layer6_outputs(3000) <= not a;
    layer6_outputs(3001) <= not a;
    layer6_outputs(3002) <= not a;
    layer6_outputs(3003) <= not a or b;
    layer6_outputs(3004) <= a xor b;
    layer6_outputs(3005) <= not b;
    layer6_outputs(3006) <= b and not a;
    layer6_outputs(3007) <= not a or b;
    layer6_outputs(3008) <= not b;
    layer6_outputs(3009) <= a;
    layer6_outputs(3010) <= not a;
    layer6_outputs(3011) <= not a;
    layer6_outputs(3012) <= a xor b;
    layer6_outputs(3013) <= a and b;
    layer6_outputs(3014) <= a or b;
    layer6_outputs(3015) <= not b;
    layer6_outputs(3016) <= b and not a;
    layer6_outputs(3017) <= not a;
    layer6_outputs(3018) <= not (a or b);
    layer6_outputs(3019) <= a;
    layer6_outputs(3020) <= not b;
    layer6_outputs(3021) <= b;
    layer6_outputs(3022) <= not (a and b);
    layer6_outputs(3023) <= not b;
    layer6_outputs(3024) <= not a;
    layer6_outputs(3025) <= a or b;
    layer6_outputs(3026) <= b and not a;
    layer6_outputs(3027) <= not (a and b);
    layer6_outputs(3028) <= a;
    layer6_outputs(3029) <= not (a xor b);
    layer6_outputs(3030) <= not b;
    layer6_outputs(3031) <= a xor b;
    layer6_outputs(3032) <= a;
    layer6_outputs(3033) <= a or b;
    layer6_outputs(3034) <= not a or b;
    layer6_outputs(3035) <= not (a xor b);
    layer6_outputs(3036) <= b;
    layer6_outputs(3037) <= b;
    layer6_outputs(3038) <= not (a xor b);
    layer6_outputs(3039) <= b;
    layer6_outputs(3040) <= a and not b;
    layer6_outputs(3041) <= a;
    layer6_outputs(3042) <= a;
    layer6_outputs(3043) <= not a;
    layer6_outputs(3044) <= not b;
    layer6_outputs(3045) <= a;
    layer6_outputs(3046) <= a or b;
    layer6_outputs(3047) <= b;
    layer6_outputs(3048) <= not b;
    layer6_outputs(3049) <= not (a and b);
    layer6_outputs(3050) <= a;
    layer6_outputs(3051) <= b;
    layer6_outputs(3052) <= not (a or b);
    layer6_outputs(3053) <= not (a or b);
    layer6_outputs(3054) <= not (a or b);
    layer6_outputs(3055) <= not b or a;
    layer6_outputs(3056) <= a;
    layer6_outputs(3057) <= not (a xor b);
    layer6_outputs(3058) <= not (a and b);
    layer6_outputs(3059) <= not b;
    layer6_outputs(3060) <= not a or b;
    layer6_outputs(3061) <= a xor b;
    layer6_outputs(3062) <= not (a and b);
    layer6_outputs(3063) <= not b;
    layer6_outputs(3064) <= a;
    layer6_outputs(3065) <= not b or a;
    layer6_outputs(3066) <= not b;
    layer6_outputs(3067) <= not (a xor b);
    layer6_outputs(3068) <= not (a xor b);
    layer6_outputs(3069) <= not b;
    layer6_outputs(3070) <= b;
    layer6_outputs(3071) <= a;
    layer6_outputs(3072) <= a;
    layer6_outputs(3073) <= b;
    layer6_outputs(3074) <= b and not a;
    layer6_outputs(3075) <= a and not b;
    layer6_outputs(3076) <= not b;
    layer6_outputs(3077) <= b;
    layer6_outputs(3078) <= not a;
    layer6_outputs(3079) <= not (a and b);
    layer6_outputs(3080) <= not (a and b);
    layer6_outputs(3081) <= not (a and b);
    layer6_outputs(3082) <= a xor b;
    layer6_outputs(3083) <= a;
    layer6_outputs(3084) <= a xor b;
    layer6_outputs(3085) <= not b;
    layer6_outputs(3086) <= a xor b;
    layer6_outputs(3087) <= a and b;
    layer6_outputs(3088) <= a xor b;
    layer6_outputs(3089) <= b;
    layer6_outputs(3090) <= a and b;
    layer6_outputs(3091) <= b and not a;
    layer6_outputs(3092) <= a;
    layer6_outputs(3093) <= a and not b;
    layer6_outputs(3094) <= not (a and b);
    layer6_outputs(3095) <= not a or b;
    layer6_outputs(3096) <= '0';
    layer6_outputs(3097) <= a and not b;
    layer6_outputs(3098) <= b;
    layer6_outputs(3099) <= b;
    layer6_outputs(3100) <= b;
    layer6_outputs(3101) <= a xor b;
    layer6_outputs(3102) <= a;
    layer6_outputs(3103) <= a xor b;
    layer6_outputs(3104) <= b;
    layer6_outputs(3105) <= b;
    layer6_outputs(3106) <= not b;
    layer6_outputs(3107) <= a xor b;
    layer6_outputs(3108) <= a and not b;
    layer6_outputs(3109) <= a xor b;
    layer6_outputs(3110) <= a and b;
    layer6_outputs(3111) <= not a;
    layer6_outputs(3112) <= a and b;
    layer6_outputs(3113) <= a and not b;
    layer6_outputs(3114) <= not b;
    layer6_outputs(3115) <= not (a xor b);
    layer6_outputs(3116) <= not b or a;
    layer6_outputs(3117) <= not a or b;
    layer6_outputs(3118) <= a or b;
    layer6_outputs(3119) <= b and not a;
    layer6_outputs(3120) <= not (a or b);
    layer6_outputs(3121) <= not b;
    layer6_outputs(3122) <= a and not b;
    layer6_outputs(3123) <= not (a xor b);
    layer6_outputs(3124) <= a and b;
    layer6_outputs(3125) <= a xor b;
    layer6_outputs(3126) <= a;
    layer6_outputs(3127) <= not (a and b);
    layer6_outputs(3128) <= a and not b;
    layer6_outputs(3129) <= a;
    layer6_outputs(3130) <= not (a xor b);
    layer6_outputs(3131) <= b;
    layer6_outputs(3132) <= a;
    layer6_outputs(3133) <= a and b;
    layer6_outputs(3134) <= not (a xor b);
    layer6_outputs(3135) <= a;
    layer6_outputs(3136) <= not b;
    layer6_outputs(3137) <= b;
    layer6_outputs(3138) <= a;
    layer6_outputs(3139) <= a;
    layer6_outputs(3140) <= a and not b;
    layer6_outputs(3141) <= not (a xor b);
    layer6_outputs(3142) <= not a or b;
    layer6_outputs(3143) <= b;
    layer6_outputs(3144) <= not b;
    layer6_outputs(3145) <= not (a xor b);
    layer6_outputs(3146) <= not (a xor b);
    layer6_outputs(3147) <= b;
    layer6_outputs(3148) <= not (a or b);
    layer6_outputs(3149) <= a;
    layer6_outputs(3150) <= not a;
    layer6_outputs(3151) <= not a or b;
    layer6_outputs(3152) <= a or b;
    layer6_outputs(3153) <= not b;
    layer6_outputs(3154) <= not (a xor b);
    layer6_outputs(3155) <= a;
    layer6_outputs(3156) <= a;
    layer6_outputs(3157) <= a or b;
    layer6_outputs(3158) <= not (a xor b);
    layer6_outputs(3159) <= not (a and b);
    layer6_outputs(3160) <= a and not b;
    layer6_outputs(3161) <= a and b;
    layer6_outputs(3162) <= a xor b;
    layer6_outputs(3163) <= a and b;
    layer6_outputs(3164) <= not (a xor b);
    layer6_outputs(3165) <= not (a and b);
    layer6_outputs(3166) <= b and not a;
    layer6_outputs(3167) <= not a;
    layer6_outputs(3168) <= a;
    layer6_outputs(3169) <= a;
    layer6_outputs(3170) <= not b;
    layer6_outputs(3171) <= not (a xor b);
    layer6_outputs(3172) <= not (a xor b);
    layer6_outputs(3173) <= not a or b;
    layer6_outputs(3174) <= a;
    layer6_outputs(3175) <= '1';
    layer6_outputs(3176) <= a and b;
    layer6_outputs(3177) <= a and b;
    layer6_outputs(3178) <= a or b;
    layer6_outputs(3179) <= a;
    layer6_outputs(3180) <= not (a xor b);
    layer6_outputs(3181) <= not b;
    layer6_outputs(3182) <= not (a and b);
    layer6_outputs(3183) <= not a;
    layer6_outputs(3184) <= b and not a;
    layer6_outputs(3185) <= not b;
    layer6_outputs(3186) <= not a;
    layer6_outputs(3187) <= not a or b;
    layer6_outputs(3188) <= not (a xor b);
    layer6_outputs(3189) <= b;
    layer6_outputs(3190) <= a xor b;
    layer6_outputs(3191) <= not (a or b);
    layer6_outputs(3192) <= not (a and b);
    layer6_outputs(3193) <= a or b;
    layer6_outputs(3194) <= not (a xor b);
    layer6_outputs(3195) <= a xor b;
    layer6_outputs(3196) <= b;
    layer6_outputs(3197) <= not (a or b);
    layer6_outputs(3198) <= not a;
    layer6_outputs(3199) <= a and b;
    layer6_outputs(3200) <= a;
    layer6_outputs(3201) <= a;
    layer6_outputs(3202) <= not (a xor b);
    layer6_outputs(3203) <= a or b;
    layer6_outputs(3204) <= b;
    layer6_outputs(3205) <= a or b;
    layer6_outputs(3206) <= not b or a;
    layer6_outputs(3207) <= not b;
    layer6_outputs(3208) <= not b;
    layer6_outputs(3209) <= not b;
    layer6_outputs(3210) <= a or b;
    layer6_outputs(3211) <= a;
    layer6_outputs(3212) <= a xor b;
    layer6_outputs(3213) <= not (a and b);
    layer6_outputs(3214) <= b and not a;
    layer6_outputs(3215) <= b and not a;
    layer6_outputs(3216) <= a;
    layer6_outputs(3217) <= not b;
    layer6_outputs(3218) <= not b;
    layer6_outputs(3219) <= a;
    layer6_outputs(3220) <= not b;
    layer6_outputs(3221) <= not a or b;
    layer6_outputs(3222) <= not a or b;
    layer6_outputs(3223) <= a;
    layer6_outputs(3224) <= a xor b;
    layer6_outputs(3225) <= b;
    layer6_outputs(3226) <= not (a xor b);
    layer6_outputs(3227) <= a and b;
    layer6_outputs(3228) <= a;
    layer6_outputs(3229) <= not a;
    layer6_outputs(3230) <= a and not b;
    layer6_outputs(3231) <= a;
    layer6_outputs(3232) <= a xor b;
    layer6_outputs(3233) <= not a;
    layer6_outputs(3234) <= not b;
    layer6_outputs(3235) <= a xor b;
    layer6_outputs(3236) <= a or b;
    layer6_outputs(3237) <= not b or a;
    layer6_outputs(3238) <= b and not a;
    layer6_outputs(3239) <= a and b;
    layer6_outputs(3240) <= not a;
    layer6_outputs(3241) <= b and not a;
    layer6_outputs(3242) <= not (a xor b);
    layer6_outputs(3243) <= a;
    layer6_outputs(3244) <= a and b;
    layer6_outputs(3245) <= a and b;
    layer6_outputs(3246) <= not a;
    layer6_outputs(3247) <= not b;
    layer6_outputs(3248) <= not (a and b);
    layer6_outputs(3249) <= not b;
    layer6_outputs(3250) <= not b;
    layer6_outputs(3251) <= not a or b;
    layer6_outputs(3252) <= not (a xor b);
    layer6_outputs(3253) <= not (a or b);
    layer6_outputs(3254) <= b and not a;
    layer6_outputs(3255) <= not a;
    layer6_outputs(3256) <= not (a xor b);
    layer6_outputs(3257) <= not (a or b);
    layer6_outputs(3258) <= not (a and b);
    layer6_outputs(3259) <= a or b;
    layer6_outputs(3260) <= a xor b;
    layer6_outputs(3261) <= not (a and b);
    layer6_outputs(3262) <= not b;
    layer6_outputs(3263) <= '1';
    layer6_outputs(3264) <= a;
    layer6_outputs(3265) <= not a;
    layer6_outputs(3266) <= a xor b;
    layer6_outputs(3267) <= not a or b;
    layer6_outputs(3268) <= not a;
    layer6_outputs(3269) <= a and b;
    layer6_outputs(3270) <= not b or a;
    layer6_outputs(3271) <= a;
    layer6_outputs(3272) <= not b or a;
    layer6_outputs(3273) <= a;
    layer6_outputs(3274) <= not (a xor b);
    layer6_outputs(3275) <= not a;
    layer6_outputs(3276) <= b;
    layer6_outputs(3277) <= not b or a;
    layer6_outputs(3278) <= not (a xor b);
    layer6_outputs(3279) <= b;
    layer6_outputs(3280) <= a or b;
    layer6_outputs(3281) <= not b;
    layer6_outputs(3282) <= not b;
    layer6_outputs(3283) <= a xor b;
    layer6_outputs(3284) <= a and not b;
    layer6_outputs(3285) <= not (a and b);
    layer6_outputs(3286) <= not b or a;
    layer6_outputs(3287) <= not a;
    layer6_outputs(3288) <= a;
    layer6_outputs(3289) <= not (a xor b);
    layer6_outputs(3290) <= not (a xor b);
    layer6_outputs(3291) <= a and b;
    layer6_outputs(3292) <= b;
    layer6_outputs(3293) <= not a;
    layer6_outputs(3294) <= not b;
    layer6_outputs(3295) <= not b or a;
    layer6_outputs(3296) <= a and b;
    layer6_outputs(3297) <= not (a and b);
    layer6_outputs(3298) <= a;
    layer6_outputs(3299) <= not a;
    layer6_outputs(3300) <= not b or a;
    layer6_outputs(3301) <= not a or b;
    layer6_outputs(3302) <= a xor b;
    layer6_outputs(3303) <= not (a xor b);
    layer6_outputs(3304) <= a;
    layer6_outputs(3305) <= not (a or b);
    layer6_outputs(3306) <= b;
    layer6_outputs(3307) <= not (a and b);
    layer6_outputs(3308) <= not b;
    layer6_outputs(3309) <= not b;
    layer6_outputs(3310) <= not b;
    layer6_outputs(3311) <= not (a or b);
    layer6_outputs(3312) <= a;
    layer6_outputs(3313) <= not a;
    layer6_outputs(3314) <= b;
    layer6_outputs(3315) <= not b or a;
    layer6_outputs(3316) <= not a;
    layer6_outputs(3317) <= not (a and b);
    layer6_outputs(3318) <= not a or b;
    layer6_outputs(3319) <= a xor b;
    layer6_outputs(3320) <= a xor b;
    layer6_outputs(3321) <= not a;
    layer6_outputs(3322) <= not (a xor b);
    layer6_outputs(3323) <= not b or a;
    layer6_outputs(3324) <= b and not a;
    layer6_outputs(3325) <= not b or a;
    layer6_outputs(3326) <= not (a and b);
    layer6_outputs(3327) <= a and b;
    layer6_outputs(3328) <= not b;
    layer6_outputs(3329) <= not (a xor b);
    layer6_outputs(3330) <= not b;
    layer6_outputs(3331) <= a;
    layer6_outputs(3332) <= a xor b;
    layer6_outputs(3333) <= a;
    layer6_outputs(3334) <= not a;
    layer6_outputs(3335) <= a xor b;
    layer6_outputs(3336) <= not (a xor b);
    layer6_outputs(3337) <= a;
    layer6_outputs(3338) <= b;
    layer6_outputs(3339) <= a and b;
    layer6_outputs(3340) <= b;
    layer6_outputs(3341) <= a or b;
    layer6_outputs(3342) <= not (a and b);
    layer6_outputs(3343) <= a xor b;
    layer6_outputs(3344) <= not (a xor b);
    layer6_outputs(3345) <= b;
    layer6_outputs(3346) <= not b or a;
    layer6_outputs(3347) <= b;
    layer6_outputs(3348) <= '0';
    layer6_outputs(3349) <= not b or a;
    layer6_outputs(3350) <= a;
    layer6_outputs(3351) <= not b;
    layer6_outputs(3352) <= not b;
    layer6_outputs(3353) <= b and not a;
    layer6_outputs(3354) <= a and not b;
    layer6_outputs(3355) <= a;
    layer6_outputs(3356) <= a;
    layer6_outputs(3357) <= b;
    layer6_outputs(3358) <= not (a and b);
    layer6_outputs(3359) <= b;
    layer6_outputs(3360) <= not b or a;
    layer6_outputs(3361) <= a;
    layer6_outputs(3362) <= a;
    layer6_outputs(3363) <= a;
    layer6_outputs(3364) <= a xor b;
    layer6_outputs(3365) <= a;
    layer6_outputs(3366) <= not (a or b);
    layer6_outputs(3367) <= a xor b;
    layer6_outputs(3368) <= b;
    layer6_outputs(3369) <= a or b;
    layer6_outputs(3370) <= not (a and b);
    layer6_outputs(3371) <= b;
    layer6_outputs(3372) <= a and b;
    layer6_outputs(3373) <= not (a xor b);
    layer6_outputs(3374) <= not a;
    layer6_outputs(3375) <= a xor b;
    layer6_outputs(3376) <= not b;
    layer6_outputs(3377) <= not (a or b);
    layer6_outputs(3378) <= a and not b;
    layer6_outputs(3379) <= not a or b;
    layer6_outputs(3380) <= a xor b;
    layer6_outputs(3381) <= b;
    layer6_outputs(3382) <= not a;
    layer6_outputs(3383) <= not a;
    layer6_outputs(3384) <= not (a xor b);
    layer6_outputs(3385) <= not (a and b);
    layer6_outputs(3386) <= b;
    layer6_outputs(3387) <= b;
    layer6_outputs(3388) <= not (a xor b);
    layer6_outputs(3389) <= a or b;
    layer6_outputs(3390) <= not (a xor b);
    layer6_outputs(3391) <= not a;
    layer6_outputs(3392) <= b;
    layer6_outputs(3393) <= a and not b;
    layer6_outputs(3394) <= not a;
    layer6_outputs(3395) <= not (a and b);
    layer6_outputs(3396) <= not a or b;
    layer6_outputs(3397) <= a xor b;
    layer6_outputs(3398) <= a;
    layer6_outputs(3399) <= not a or b;
    layer6_outputs(3400) <= not (a and b);
    layer6_outputs(3401) <= not b;
    layer6_outputs(3402) <= a xor b;
    layer6_outputs(3403) <= b;
    layer6_outputs(3404) <= a;
    layer6_outputs(3405) <= not (a and b);
    layer6_outputs(3406) <= not (a or b);
    layer6_outputs(3407) <= not b or a;
    layer6_outputs(3408) <= b and not a;
    layer6_outputs(3409) <= b;
    layer6_outputs(3410) <= a xor b;
    layer6_outputs(3411) <= b and not a;
    layer6_outputs(3412) <= not (a xor b);
    layer6_outputs(3413) <= b;
    layer6_outputs(3414) <= not (a or b);
    layer6_outputs(3415) <= not b;
    layer6_outputs(3416) <= a and b;
    layer6_outputs(3417) <= a and b;
    layer6_outputs(3418) <= not b;
    layer6_outputs(3419) <= b and not a;
    layer6_outputs(3420) <= b and not a;
    layer6_outputs(3421) <= not a;
    layer6_outputs(3422) <= a;
    layer6_outputs(3423) <= a;
    layer6_outputs(3424) <= b;
    layer6_outputs(3425) <= not (a xor b);
    layer6_outputs(3426) <= a or b;
    layer6_outputs(3427) <= a xor b;
    layer6_outputs(3428) <= b;
    layer6_outputs(3429) <= b;
    layer6_outputs(3430) <= a xor b;
    layer6_outputs(3431) <= a;
    layer6_outputs(3432) <= a and not b;
    layer6_outputs(3433) <= not (a and b);
    layer6_outputs(3434) <= not a;
    layer6_outputs(3435) <= b;
    layer6_outputs(3436) <= not a;
    layer6_outputs(3437) <= not b;
    layer6_outputs(3438) <= not (a and b);
    layer6_outputs(3439) <= not b or a;
    layer6_outputs(3440) <= not a;
    layer6_outputs(3441) <= a;
    layer6_outputs(3442) <= not (a xor b);
    layer6_outputs(3443) <= b;
    layer6_outputs(3444) <= a;
    layer6_outputs(3445) <= not b;
    layer6_outputs(3446) <= b;
    layer6_outputs(3447) <= not a or b;
    layer6_outputs(3448) <= not b or a;
    layer6_outputs(3449) <= not (a xor b);
    layer6_outputs(3450) <= a;
    layer6_outputs(3451) <= a xor b;
    layer6_outputs(3452) <= b;
    layer6_outputs(3453) <= not (a or b);
    layer6_outputs(3454) <= a xor b;
    layer6_outputs(3455) <= not a;
    layer6_outputs(3456) <= '1';
    layer6_outputs(3457) <= not (a xor b);
    layer6_outputs(3458) <= a;
    layer6_outputs(3459) <= not b;
    layer6_outputs(3460) <= not b;
    layer6_outputs(3461) <= b;
    layer6_outputs(3462) <= b;
    layer6_outputs(3463) <= a xor b;
    layer6_outputs(3464) <= not (a xor b);
    layer6_outputs(3465) <= not (a or b);
    layer6_outputs(3466) <= not a;
    layer6_outputs(3467) <= b and not a;
    layer6_outputs(3468) <= a;
    layer6_outputs(3469) <= not b;
    layer6_outputs(3470) <= not b;
    layer6_outputs(3471) <= not a;
    layer6_outputs(3472) <= not b;
    layer6_outputs(3473) <= not b;
    layer6_outputs(3474) <= a xor b;
    layer6_outputs(3475) <= not a;
    layer6_outputs(3476) <= a;
    layer6_outputs(3477) <= not a;
    layer6_outputs(3478) <= b;
    layer6_outputs(3479) <= a;
    layer6_outputs(3480) <= not b or a;
    layer6_outputs(3481) <= not (a xor b);
    layer6_outputs(3482) <= a;
    layer6_outputs(3483) <= a;
    layer6_outputs(3484) <= a;
    layer6_outputs(3485) <= b;
    layer6_outputs(3486) <= '0';
    layer6_outputs(3487) <= a and not b;
    layer6_outputs(3488) <= not (a xor b);
    layer6_outputs(3489) <= not a or b;
    layer6_outputs(3490) <= not (a and b);
    layer6_outputs(3491) <= a;
    layer6_outputs(3492) <= b;
    layer6_outputs(3493) <= a;
    layer6_outputs(3494) <= a;
    layer6_outputs(3495) <= not (a or b);
    layer6_outputs(3496) <= b and not a;
    layer6_outputs(3497) <= '1';
    layer6_outputs(3498) <= not (a xor b);
    layer6_outputs(3499) <= a and b;
    layer6_outputs(3500) <= b;
    layer6_outputs(3501) <= not a;
    layer6_outputs(3502) <= not (a xor b);
    layer6_outputs(3503) <= a xor b;
    layer6_outputs(3504) <= a;
    layer6_outputs(3505) <= a;
    layer6_outputs(3506) <= a;
    layer6_outputs(3507) <= not (a or b);
    layer6_outputs(3508) <= a and b;
    layer6_outputs(3509) <= a and b;
    layer6_outputs(3510) <= not (a xor b);
    layer6_outputs(3511) <= not (a and b);
    layer6_outputs(3512) <= b;
    layer6_outputs(3513) <= not a;
    layer6_outputs(3514) <= not (a and b);
    layer6_outputs(3515) <= a;
    layer6_outputs(3516) <= b and not a;
    layer6_outputs(3517) <= a and b;
    layer6_outputs(3518) <= not b;
    layer6_outputs(3519) <= b;
    layer6_outputs(3520) <= a;
    layer6_outputs(3521) <= a xor b;
    layer6_outputs(3522) <= not (a or b);
    layer6_outputs(3523) <= not (a xor b);
    layer6_outputs(3524) <= not b;
    layer6_outputs(3525) <= a;
    layer6_outputs(3526) <= a xor b;
    layer6_outputs(3527) <= a;
    layer6_outputs(3528) <= not (a xor b);
    layer6_outputs(3529) <= not b or a;
    layer6_outputs(3530) <= b;
    layer6_outputs(3531) <= not (a or b);
    layer6_outputs(3532) <= b and not a;
    layer6_outputs(3533) <= not (a and b);
    layer6_outputs(3534) <= not b;
    layer6_outputs(3535) <= not (a xor b);
    layer6_outputs(3536) <= a xor b;
    layer6_outputs(3537) <= a;
    layer6_outputs(3538) <= a xor b;
    layer6_outputs(3539) <= a xor b;
    layer6_outputs(3540) <= not b;
    layer6_outputs(3541) <= not a or b;
    layer6_outputs(3542) <= a and not b;
    layer6_outputs(3543) <= not b;
    layer6_outputs(3544) <= not (a and b);
    layer6_outputs(3545) <= not b or a;
    layer6_outputs(3546) <= b;
    layer6_outputs(3547) <= a xor b;
    layer6_outputs(3548) <= a;
    layer6_outputs(3549) <= not a;
    layer6_outputs(3550) <= a and b;
    layer6_outputs(3551) <= not b;
    layer6_outputs(3552) <= b and not a;
    layer6_outputs(3553) <= not b;
    layer6_outputs(3554) <= '1';
    layer6_outputs(3555) <= not a;
    layer6_outputs(3556) <= a;
    layer6_outputs(3557) <= b;
    layer6_outputs(3558) <= a or b;
    layer6_outputs(3559) <= b;
    layer6_outputs(3560) <= not (a xor b);
    layer6_outputs(3561) <= a xor b;
    layer6_outputs(3562) <= a and not b;
    layer6_outputs(3563) <= b;
    layer6_outputs(3564) <= not a;
    layer6_outputs(3565) <= a xor b;
    layer6_outputs(3566) <= a or b;
    layer6_outputs(3567) <= b;
    layer6_outputs(3568) <= b and not a;
    layer6_outputs(3569) <= not (a or b);
    layer6_outputs(3570) <= not b;
    layer6_outputs(3571) <= not a;
    layer6_outputs(3572) <= not a;
    layer6_outputs(3573) <= not (a xor b);
    layer6_outputs(3574) <= b;
    layer6_outputs(3575) <= a;
    layer6_outputs(3576) <= a;
    layer6_outputs(3577) <= b and not a;
    layer6_outputs(3578) <= a xor b;
    layer6_outputs(3579) <= not (a xor b);
    layer6_outputs(3580) <= not (a and b);
    layer6_outputs(3581) <= not (a xor b);
    layer6_outputs(3582) <= '1';
    layer6_outputs(3583) <= not b;
    layer6_outputs(3584) <= b and not a;
    layer6_outputs(3585) <= not b;
    layer6_outputs(3586) <= b;
    layer6_outputs(3587) <= a and b;
    layer6_outputs(3588) <= not a;
    layer6_outputs(3589) <= b and not a;
    layer6_outputs(3590) <= a and not b;
    layer6_outputs(3591) <= a and not b;
    layer6_outputs(3592) <= not b;
    layer6_outputs(3593) <= not (a xor b);
    layer6_outputs(3594) <= not (a xor b);
    layer6_outputs(3595) <= not b;
    layer6_outputs(3596) <= a;
    layer6_outputs(3597) <= not (a xor b);
    layer6_outputs(3598) <= a and b;
    layer6_outputs(3599) <= a or b;
    layer6_outputs(3600) <= a;
    layer6_outputs(3601) <= a;
    layer6_outputs(3602) <= not a;
    layer6_outputs(3603) <= '0';
    layer6_outputs(3604) <= not a or b;
    layer6_outputs(3605) <= not b;
    layer6_outputs(3606) <= a;
    layer6_outputs(3607) <= not b;
    layer6_outputs(3608) <= not a;
    layer6_outputs(3609) <= not b;
    layer6_outputs(3610) <= b and not a;
    layer6_outputs(3611) <= not a;
    layer6_outputs(3612) <= not a or b;
    layer6_outputs(3613) <= a;
    layer6_outputs(3614) <= not a;
    layer6_outputs(3615) <= not b or a;
    layer6_outputs(3616) <= not b;
    layer6_outputs(3617) <= not a;
    layer6_outputs(3618) <= '1';
    layer6_outputs(3619) <= a and b;
    layer6_outputs(3620) <= a;
    layer6_outputs(3621) <= a and not b;
    layer6_outputs(3622) <= not (a or b);
    layer6_outputs(3623) <= not (a or b);
    layer6_outputs(3624) <= not b;
    layer6_outputs(3625) <= not (a xor b);
    layer6_outputs(3626) <= a and not b;
    layer6_outputs(3627) <= b;
    layer6_outputs(3628) <= b;
    layer6_outputs(3629) <= a;
    layer6_outputs(3630) <= a;
    layer6_outputs(3631) <= a xor b;
    layer6_outputs(3632) <= not a or b;
    layer6_outputs(3633) <= not (a xor b);
    layer6_outputs(3634) <= a xor b;
    layer6_outputs(3635) <= a or b;
    layer6_outputs(3636) <= a or b;
    layer6_outputs(3637) <= not a;
    layer6_outputs(3638) <= not b;
    layer6_outputs(3639) <= a xor b;
    layer6_outputs(3640) <= a xor b;
    layer6_outputs(3641) <= a;
    layer6_outputs(3642) <= not a;
    layer6_outputs(3643) <= a xor b;
    layer6_outputs(3644) <= a and not b;
    layer6_outputs(3645) <= a and not b;
    layer6_outputs(3646) <= b;
    layer6_outputs(3647) <= not (a xor b);
    layer6_outputs(3648) <= not b or a;
    layer6_outputs(3649) <= b;
    layer6_outputs(3650) <= not b;
    layer6_outputs(3651) <= '1';
    layer6_outputs(3652) <= not (a or b);
    layer6_outputs(3653) <= a;
    layer6_outputs(3654) <= not b or a;
    layer6_outputs(3655) <= a and b;
    layer6_outputs(3656) <= b;
    layer6_outputs(3657) <= not b;
    layer6_outputs(3658) <= not (a or b);
    layer6_outputs(3659) <= not b;
    layer6_outputs(3660) <= not a or b;
    layer6_outputs(3661) <= not b or a;
    layer6_outputs(3662) <= not (a or b);
    layer6_outputs(3663) <= not b;
    layer6_outputs(3664) <= not (a xor b);
    layer6_outputs(3665) <= a;
    layer6_outputs(3666) <= not (a and b);
    layer6_outputs(3667) <= a;
    layer6_outputs(3668) <= a xor b;
    layer6_outputs(3669) <= b and not a;
    layer6_outputs(3670) <= not (a or b);
    layer6_outputs(3671) <= b;
    layer6_outputs(3672) <= a xor b;
    layer6_outputs(3673) <= b;
    layer6_outputs(3674) <= b;
    layer6_outputs(3675) <= not (a or b);
    layer6_outputs(3676) <= not a or b;
    layer6_outputs(3677) <= not (a or b);
    layer6_outputs(3678) <= not b or a;
    layer6_outputs(3679) <= not b;
    layer6_outputs(3680) <= a;
    layer6_outputs(3681) <= not a or b;
    layer6_outputs(3682) <= a or b;
    layer6_outputs(3683) <= not (a xor b);
    layer6_outputs(3684) <= not a or b;
    layer6_outputs(3685) <= '0';
    layer6_outputs(3686) <= b;
    layer6_outputs(3687) <= b;
    layer6_outputs(3688) <= b;
    layer6_outputs(3689) <= not b;
    layer6_outputs(3690) <= not (a or b);
    layer6_outputs(3691) <= a xor b;
    layer6_outputs(3692) <= a;
    layer6_outputs(3693) <= a xor b;
    layer6_outputs(3694) <= not (a xor b);
    layer6_outputs(3695) <= not a;
    layer6_outputs(3696) <= not (a xor b);
    layer6_outputs(3697) <= a;
    layer6_outputs(3698) <= b;
    layer6_outputs(3699) <= not b or a;
    layer6_outputs(3700) <= a xor b;
    layer6_outputs(3701) <= a;
    layer6_outputs(3702) <= not b;
    layer6_outputs(3703) <= a or b;
    layer6_outputs(3704) <= a;
    layer6_outputs(3705) <= b;
    layer6_outputs(3706) <= b;
    layer6_outputs(3707) <= b;
    layer6_outputs(3708) <= a;
    layer6_outputs(3709) <= a;
    layer6_outputs(3710) <= b;
    layer6_outputs(3711) <= not a;
    layer6_outputs(3712) <= not b;
    layer6_outputs(3713) <= b;
    layer6_outputs(3714) <= '0';
    layer6_outputs(3715) <= b and not a;
    layer6_outputs(3716) <= not b or a;
    layer6_outputs(3717) <= not a;
    layer6_outputs(3718) <= a;
    layer6_outputs(3719) <= not (a and b);
    layer6_outputs(3720) <= b and not a;
    layer6_outputs(3721) <= a and not b;
    layer6_outputs(3722) <= a xor b;
    layer6_outputs(3723) <= not (a xor b);
    layer6_outputs(3724) <= b and not a;
    layer6_outputs(3725) <= not (a xor b);
    layer6_outputs(3726) <= not (a or b);
    layer6_outputs(3727) <= not b;
    layer6_outputs(3728) <= b and not a;
    layer6_outputs(3729) <= b;
    layer6_outputs(3730) <= b;
    layer6_outputs(3731) <= not b;
    layer6_outputs(3732) <= a;
    layer6_outputs(3733) <= b;
    layer6_outputs(3734) <= b;
    layer6_outputs(3735) <= not b;
    layer6_outputs(3736) <= not a;
    layer6_outputs(3737) <= a and not b;
    layer6_outputs(3738) <= not (a and b);
    layer6_outputs(3739) <= a xor b;
    layer6_outputs(3740) <= not a;
    layer6_outputs(3741) <= not (a xor b);
    layer6_outputs(3742) <= b and not a;
    layer6_outputs(3743) <= b;
    layer6_outputs(3744) <= not a;
    layer6_outputs(3745) <= b;
    layer6_outputs(3746) <= a xor b;
    layer6_outputs(3747) <= not a;
    layer6_outputs(3748) <= not (a and b);
    layer6_outputs(3749) <= a;
    layer6_outputs(3750) <= b and not a;
    layer6_outputs(3751) <= not b;
    layer6_outputs(3752) <= not (a or b);
    layer6_outputs(3753) <= a;
    layer6_outputs(3754) <= not a;
    layer6_outputs(3755) <= not (a xor b);
    layer6_outputs(3756) <= not (a xor b);
    layer6_outputs(3757) <= a;
    layer6_outputs(3758) <= not a;
    layer6_outputs(3759) <= a;
    layer6_outputs(3760) <= not b or a;
    layer6_outputs(3761) <= b;
    layer6_outputs(3762) <= not (a xor b);
    layer6_outputs(3763) <= a and not b;
    layer6_outputs(3764) <= b;
    layer6_outputs(3765) <= a;
    layer6_outputs(3766) <= a or b;
    layer6_outputs(3767) <= not b or a;
    layer6_outputs(3768) <= a and b;
    layer6_outputs(3769) <= not b or a;
    layer6_outputs(3770) <= a or b;
    layer6_outputs(3771) <= not a;
    layer6_outputs(3772) <= a xor b;
    layer6_outputs(3773) <= a;
    layer6_outputs(3774) <= b;
    layer6_outputs(3775) <= not b;
    layer6_outputs(3776) <= a xor b;
    layer6_outputs(3777) <= not a;
    layer6_outputs(3778) <= b;
    layer6_outputs(3779) <= a;
    layer6_outputs(3780) <= not a;
    layer6_outputs(3781) <= not a;
    layer6_outputs(3782) <= a;
    layer6_outputs(3783) <= a and not b;
    layer6_outputs(3784) <= a or b;
    layer6_outputs(3785) <= not (a or b);
    layer6_outputs(3786) <= not (a or b);
    layer6_outputs(3787) <= a;
    layer6_outputs(3788) <= not a;
    layer6_outputs(3789) <= not (a and b);
    layer6_outputs(3790) <= not a;
    layer6_outputs(3791) <= not (a xor b);
    layer6_outputs(3792) <= a and not b;
    layer6_outputs(3793) <= not (a and b);
    layer6_outputs(3794) <= not a;
    layer6_outputs(3795) <= not b;
    layer6_outputs(3796) <= a and not b;
    layer6_outputs(3797) <= '0';
    layer6_outputs(3798) <= '0';
    layer6_outputs(3799) <= a;
    layer6_outputs(3800) <= b;
    layer6_outputs(3801) <= a;
    layer6_outputs(3802) <= a and b;
    layer6_outputs(3803) <= b;
    layer6_outputs(3804) <= b and not a;
    layer6_outputs(3805) <= a and b;
    layer6_outputs(3806) <= a;
    layer6_outputs(3807) <= not a or b;
    layer6_outputs(3808) <= not a or b;
    layer6_outputs(3809) <= b;
    layer6_outputs(3810) <= not b or a;
    layer6_outputs(3811) <= not (a or b);
    layer6_outputs(3812) <= not a;
    layer6_outputs(3813) <= b;
    layer6_outputs(3814) <= not b or a;
    layer6_outputs(3815) <= not (a and b);
    layer6_outputs(3816) <= b;
    layer6_outputs(3817) <= not b;
    layer6_outputs(3818) <= b;
    layer6_outputs(3819) <= not b;
    layer6_outputs(3820) <= not (a and b);
    layer6_outputs(3821) <= not (a or b);
    layer6_outputs(3822) <= a xor b;
    layer6_outputs(3823) <= a and b;
    layer6_outputs(3824) <= a and b;
    layer6_outputs(3825) <= not (a xor b);
    layer6_outputs(3826) <= a xor b;
    layer6_outputs(3827) <= not b or a;
    layer6_outputs(3828) <= not b;
    layer6_outputs(3829) <= a xor b;
    layer6_outputs(3830) <= not b;
    layer6_outputs(3831) <= a;
    layer6_outputs(3832) <= not a;
    layer6_outputs(3833) <= a xor b;
    layer6_outputs(3834) <= b;
    layer6_outputs(3835) <= not (a or b);
    layer6_outputs(3836) <= not (a and b);
    layer6_outputs(3837) <= not a;
    layer6_outputs(3838) <= not b;
    layer6_outputs(3839) <= not b or a;
    layer6_outputs(3840) <= not b or a;
    layer6_outputs(3841) <= a and b;
    layer6_outputs(3842) <= a or b;
    layer6_outputs(3843) <= a and b;
    layer6_outputs(3844) <= not (a xor b);
    layer6_outputs(3845) <= not b;
    layer6_outputs(3846) <= not b or a;
    layer6_outputs(3847) <= not (a and b);
    layer6_outputs(3848) <= not b;
    layer6_outputs(3849) <= not (a xor b);
    layer6_outputs(3850) <= not b;
    layer6_outputs(3851) <= not b;
    layer6_outputs(3852) <= not (a or b);
    layer6_outputs(3853) <= a and not b;
    layer6_outputs(3854) <= not (a xor b);
    layer6_outputs(3855) <= not b;
    layer6_outputs(3856) <= b and not a;
    layer6_outputs(3857) <= a;
    layer6_outputs(3858) <= not a;
    layer6_outputs(3859) <= a and not b;
    layer6_outputs(3860) <= a and b;
    layer6_outputs(3861) <= a xor b;
    layer6_outputs(3862) <= not (a xor b);
    layer6_outputs(3863) <= a xor b;
    layer6_outputs(3864) <= a and not b;
    layer6_outputs(3865) <= a;
    layer6_outputs(3866) <= not (a xor b);
    layer6_outputs(3867) <= a and not b;
    layer6_outputs(3868) <= b;
    layer6_outputs(3869) <= not (a or b);
    layer6_outputs(3870) <= a;
    layer6_outputs(3871) <= not b;
    layer6_outputs(3872) <= a or b;
    layer6_outputs(3873) <= a xor b;
    layer6_outputs(3874) <= not (a and b);
    layer6_outputs(3875) <= a and not b;
    layer6_outputs(3876) <= not a;
    layer6_outputs(3877) <= a and b;
    layer6_outputs(3878) <= not a;
    layer6_outputs(3879) <= not (a or b);
    layer6_outputs(3880) <= not (a xor b);
    layer6_outputs(3881) <= b;
    layer6_outputs(3882) <= not a;
    layer6_outputs(3883) <= not b;
    layer6_outputs(3884) <= b;
    layer6_outputs(3885) <= not (a xor b);
    layer6_outputs(3886) <= not (a and b);
    layer6_outputs(3887) <= a xor b;
    layer6_outputs(3888) <= b;
    layer6_outputs(3889) <= a xor b;
    layer6_outputs(3890) <= a xor b;
    layer6_outputs(3891) <= not a or b;
    layer6_outputs(3892) <= not b or a;
    layer6_outputs(3893) <= a;
    layer6_outputs(3894) <= b;
    layer6_outputs(3895) <= b;
    layer6_outputs(3896) <= b;
    layer6_outputs(3897) <= b;
    layer6_outputs(3898) <= a;
    layer6_outputs(3899) <= a or b;
    layer6_outputs(3900) <= not b;
    layer6_outputs(3901) <= not (a xor b);
    layer6_outputs(3902) <= a or b;
    layer6_outputs(3903) <= not b or a;
    layer6_outputs(3904) <= a;
    layer6_outputs(3905) <= b;
    layer6_outputs(3906) <= b;
    layer6_outputs(3907) <= not a or b;
    layer6_outputs(3908) <= a or b;
    layer6_outputs(3909) <= a;
    layer6_outputs(3910) <= not b;
    layer6_outputs(3911) <= a;
    layer6_outputs(3912) <= a xor b;
    layer6_outputs(3913) <= not b;
    layer6_outputs(3914) <= a xor b;
    layer6_outputs(3915) <= a xor b;
    layer6_outputs(3916) <= b and not a;
    layer6_outputs(3917) <= not b;
    layer6_outputs(3918) <= not (a or b);
    layer6_outputs(3919) <= b and not a;
    layer6_outputs(3920) <= not a;
    layer6_outputs(3921) <= a xor b;
    layer6_outputs(3922) <= not a;
    layer6_outputs(3923) <= not b or a;
    layer6_outputs(3924) <= a or b;
    layer6_outputs(3925) <= not b;
    layer6_outputs(3926) <= not b;
    layer6_outputs(3927) <= not (a xor b);
    layer6_outputs(3928) <= a;
    layer6_outputs(3929) <= b;
    layer6_outputs(3930) <= not b or a;
    layer6_outputs(3931) <= a;
    layer6_outputs(3932) <= a;
    layer6_outputs(3933) <= a;
    layer6_outputs(3934) <= not a or b;
    layer6_outputs(3935) <= not a;
    layer6_outputs(3936) <= b and not a;
    layer6_outputs(3937) <= not b;
    layer6_outputs(3938) <= a xor b;
    layer6_outputs(3939) <= not b;
    layer6_outputs(3940) <= not (a or b);
    layer6_outputs(3941) <= not b;
    layer6_outputs(3942) <= a xor b;
    layer6_outputs(3943) <= not (a xor b);
    layer6_outputs(3944) <= not a or b;
    layer6_outputs(3945) <= a xor b;
    layer6_outputs(3946) <= a or b;
    layer6_outputs(3947) <= a;
    layer6_outputs(3948) <= a;
    layer6_outputs(3949) <= not b;
    layer6_outputs(3950) <= a xor b;
    layer6_outputs(3951) <= a;
    layer6_outputs(3952) <= not (a xor b);
    layer6_outputs(3953) <= '0';
    layer6_outputs(3954) <= not (a xor b);
    layer6_outputs(3955) <= b and not a;
    layer6_outputs(3956) <= a and b;
    layer6_outputs(3957) <= a and not b;
    layer6_outputs(3958) <= a and b;
    layer6_outputs(3959) <= not b;
    layer6_outputs(3960) <= not (a or b);
    layer6_outputs(3961) <= not b;
    layer6_outputs(3962) <= a;
    layer6_outputs(3963) <= not a;
    layer6_outputs(3964) <= not b;
    layer6_outputs(3965) <= a and b;
    layer6_outputs(3966) <= a or b;
    layer6_outputs(3967) <= a and not b;
    layer6_outputs(3968) <= not b;
    layer6_outputs(3969) <= not a or b;
    layer6_outputs(3970) <= not b;
    layer6_outputs(3971) <= b;
    layer6_outputs(3972) <= a and not b;
    layer6_outputs(3973) <= not b;
    layer6_outputs(3974) <= not a;
    layer6_outputs(3975) <= a xor b;
    layer6_outputs(3976) <= not (a xor b);
    layer6_outputs(3977) <= not a or b;
    layer6_outputs(3978) <= not (a or b);
    layer6_outputs(3979) <= not b;
    layer6_outputs(3980) <= not b or a;
    layer6_outputs(3981) <= not a;
    layer6_outputs(3982) <= a;
    layer6_outputs(3983) <= not a or b;
    layer6_outputs(3984) <= a;
    layer6_outputs(3985) <= b;
    layer6_outputs(3986) <= a and not b;
    layer6_outputs(3987) <= not (a xor b);
    layer6_outputs(3988) <= '1';
    layer6_outputs(3989) <= a xor b;
    layer6_outputs(3990) <= not (a and b);
    layer6_outputs(3991) <= not b;
    layer6_outputs(3992) <= not b;
    layer6_outputs(3993) <= a or b;
    layer6_outputs(3994) <= not b;
    layer6_outputs(3995) <= not b;
    layer6_outputs(3996) <= not b or a;
    layer6_outputs(3997) <= a or b;
    layer6_outputs(3998) <= not a;
    layer6_outputs(3999) <= not (a and b);
    layer6_outputs(4000) <= not b or a;
    layer6_outputs(4001) <= not b;
    layer6_outputs(4002) <= not (a xor b);
    layer6_outputs(4003) <= not a;
    layer6_outputs(4004) <= not (a and b);
    layer6_outputs(4005) <= a and b;
    layer6_outputs(4006) <= a xor b;
    layer6_outputs(4007) <= not (a xor b);
    layer6_outputs(4008) <= a or b;
    layer6_outputs(4009) <= not a;
    layer6_outputs(4010) <= not (a or b);
    layer6_outputs(4011) <= not a;
    layer6_outputs(4012) <= not (a xor b);
    layer6_outputs(4013) <= not (a xor b);
    layer6_outputs(4014) <= b and not a;
    layer6_outputs(4015) <= not b or a;
    layer6_outputs(4016) <= a and not b;
    layer6_outputs(4017) <= not a;
    layer6_outputs(4018) <= not (a and b);
    layer6_outputs(4019) <= not (a and b);
    layer6_outputs(4020) <= not a;
    layer6_outputs(4021) <= b;
    layer6_outputs(4022) <= a;
    layer6_outputs(4023) <= not (a xor b);
    layer6_outputs(4024) <= not (a or b);
    layer6_outputs(4025) <= b;
    layer6_outputs(4026) <= not a;
    layer6_outputs(4027) <= not b;
    layer6_outputs(4028) <= b and not a;
    layer6_outputs(4029) <= not b;
    layer6_outputs(4030) <= not (a xor b);
    layer6_outputs(4031) <= b and not a;
    layer6_outputs(4032) <= not a or b;
    layer6_outputs(4033) <= a and b;
    layer6_outputs(4034) <= b and not a;
    layer6_outputs(4035) <= a xor b;
    layer6_outputs(4036) <= not a;
    layer6_outputs(4037) <= b and not a;
    layer6_outputs(4038) <= not a or b;
    layer6_outputs(4039) <= a and not b;
    layer6_outputs(4040) <= not a;
    layer6_outputs(4041) <= not (a and b);
    layer6_outputs(4042) <= a xor b;
    layer6_outputs(4043) <= a and not b;
    layer6_outputs(4044) <= not b;
    layer6_outputs(4045) <= a xor b;
    layer6_outputs(4046) <= not (a xor b);
    layer6_outputs(4047) <= b;
    layer6_outputs(4048) <= not a;
    layer6_outputs(4049) <= not (a and b);
    layer6_outputs(4050) <= not b or a;
    layer6_outputs(4051) <= a and not b;
    layer6_outputs(4052) <= not (a xor b);
    layer6_outputs(4053) <= a and b;
    layer6_outputs(4054) <= a;
    layer6_outputs(4055) <= not b;
    layer6_outputs(4056) <= not a;
    layer6_outputs(4057) <= a;
    layer6_outputs(4058) <= not b;
    layer6_outputs(4059) <= not (a and b);
    layer6_outputs(4060) <= a;
    layer6_outputs(4061) <= b;
    layer6_outputs(4062) <= not (a or b);
    layer6_outputs(4063) <= b;
    layer6_outputs(4064) <= not a;
    layer6_outputs(4065) <= a xor b;
    layer6_outputs(4066) <= a;
    layer6_outputs(4067) <= b;
    layer6_outputs(4068) <= b;
    layer6_outputs(4069) <= not (a and b);
    layer6_outputs(4070) <= a xor b;
    layer6_outputs(4071) <= a and not b;
    layer6_outputs(4072) <= a;
    layer6_outputs(4073) <= b;
    layer6_outputs(4074) <= not (a xor b);
    layer6_outputs(4075) <= not a or b;
    layer6_outputs(4076) <= b;
    layer6_outputs(4077) <= not b;
    layer6_outputs(4078) <= not (a xor b);
    layer6_outputs(4079) <= not b;
    layer6_outputs(4080) <= b;
    layer6_outputs(4081) <= not a;
    layer6_outputs(4082) <= not (a xor b);
    layer6_outputs(4083) <= not (a xor b);
    layer6_outputs(4084) <= a and b;
    layer6_outputs(4085) <= a and b;
    layer6_outputs(4086) <= a xor b;
    layer6_outputs(4087) <= a and b;
    layer6_outputs(4088) <= b;
    layer6_outputs(4089) <= a xor b;
    layer6_outputs(4090) <= not (a and b);
    layer6_outputs(4091) <= a xor b;
    layer6_outputs(4092) <= not a or b;
    layer6_outputs(4093) <= not (a and b);
    layer6_outputs(4094) <= a;
    layer6_outputs(4095) <= a xor b;
    layer6_outputs(4096) <= a and b;
    layer6_outputs(4097) <= a xor b;
    layer6_outputs(4098) <= a xor b;
    layer6_outputs(4099) <= a;
    layer6_outputs(4100) <= not b;
    layer6_outputs(4101) <= a xor b;
    layer6_outputs(4102) <= not a or b;
    layer6_outputs(4103) <= not b or a;
    layer6_outputs(4104) <= not b or a;
    layer6_outputs(4105) <= a xor b;
    layer6_outputs(4106) <= a and not b;
    layer6_outputs(4107) <= a and b;
    layer6_outputs(4108) <= a and b;
    layer6_outputs(4109) <= a and b;
    layer6_outputs(4110) <= not (a xor b);
    layer6_outputs(4111) <= not b;
    layer6_outputs(4112) <= not a;
    layer6_outputs(4113) <= not b or a;
    layer6_outputs(4114) <= a;
    layer6_outputs(4115) <= b;
    layer6_outputs(4116) <= a and not b;
    layer6_outputs(4117) <= a and b;
    layer6_outputs(4118) <= not (a xor b);
    layer6_outputs(4119) <= not (a xor b);
    layer6_outputs(4120) <= a and not b;
    layer6_outputs(4121) <= not (a and b);
    layer6_outputs(4122) <= a xor b;
    layer6_outputs(4123) <= not (a xor b);
    layer6_outputs(4124) <= not b;
    layer6_outputs(4125) <= not a;
    layer6_outputs(4126) <= a;
    layer6_outputs(4127) <= a and not b;
    layer6_outputs(4128) <= a and b;
    layer6_outputs(4129) <= a;
    layer6_outputs(4130) <= not b;
    layer6_outputs(4131) <= b;
    layer6_outputs(4132) <= not b or a;
    layer6_outputs(4133) <= b;
    layer6_outputs(4134) <= not (a xor b);
    layer6_outputs(4135) <= not b or a;
    layer6_outputs(4136) <= b and not a;
    layer6_outputs(4137) <= not (a xor b);
    layer6_outputs(4138) <= not (a or b);
    layer6_outputs(4139) <= a xor b;
    layer6_outputs(4140) <= a and not b;
    layer6_outputs(4141) <= not (a xor b);
    layer6_outputs(4142) <= a;
    layer6_outputs(4143) <= not (a xor b);
    layer6_outputs(4144) <= not a;
    layer6_outputs(4145) <= not a or b;
    layer6_outputs(4146) <= not (a and b);
    layer6_outputs(4147) <= not (a xor b);
    layer6_outputs(4148) <= not b;
    layer6_outputs(4149) <= a;
    layer6_outputs(4150) <= not (a xor b);
    layer6_outputs(4151) <= not a;
    layer6_outputs(4152) <= not b or a;
    layer6_outputs(4153) <= b;
    layer6_outputs(4154) <= a or b;
    layer6_outputs(4155) <= a;
    layer6_outputs(4156) <= not (a and b);
    layer6_outputs(4157) <= not (a and b);
    layer6_outputs(4158) <= b and not a;
    layer6_outputs(4159) <= a xor b;
    layer6_outputs(4160) <= a xor b;
    layer6_outputs(4161) <= a xor b;
    layer6_outputs(4162) <= not a;
    layer6_outputs(4163) <= not a;
    layer6_outputs(4164) <= a xor b;
    layer6_outputs(4165) <= not b;
    layer6_outputs(4166) <= a or b;
    layer6_outputs(4167) <= a;
    layer6_outputs(4168) <= not (a and b);
    layer6_outputs(4169) <= '0';
    layer6_outputs(4170) <= not a;
    layer6_outputs(4171) <= not a or b;
    layer6_outputs(4172) <= a;
    layer6_outputs(4173) <= not a;
    layer6_outputs(4174) <= not a;
    layer6_outputs(4175) <= a and not b;
    layer6_outputs(4176) <= not b;
    layer6_outputs(4177) <= a or b;
    layer6_outputs(4178) <= a and b;
    layer6_outputs(4179) <= not b;
    layer6_outputs(4180) <= not b;
    layer6_outputs(4181) <= not b or a;
    layer6_outputs(4182) <= b and not a;
    layer6_outputs(4183) <= not (a xor b);
    layer6_outputs(4184) <= a xor b;
    layer6_outputs(4185) <= b;
    layer6_outputs(4186) <= a;
    layer6_outputs(4187) <= not b or a;
    layer6_outputs(4188) <= not a;
    layer6_outputs(4189) <= b;
    layer6_outputs(4190) <= not a or b;
    layer6_outputs(4191) <= a;
    layer6_outputs(4192) <= not a or b;
    layer6_outputs(4193) <= not a;
    layer6_outputs(4194) <= b;
    layer6_outputs(4195) <= a and not b;
    layer6_outputs(4196) <= not (a xor b);
    layer6_outputs(4197) <= b;
    layer6_outputs(4198) <= a;
    layer6_outputs(4199) <= not (a or b);
    layer6_outputs(4200) <= not b or a;
    layer6_outputs(4201) <= not b;
    layer6_outputs(4202) <= not a or b;
    layer6_outputs(4203) <= not (a or b);
    layer6_outputs(4204) <= b and not a;
    layer6_outputs(4205) <= a;
    layer6_outputs(4206) <= not (a or b);
    layer6_outputs(4207) <= not a;
    layer6_outputs(4208) <= b;
    layer6_outputs(4209) <= not (a xor b);
    layer6_outputs(4210) <= not (a xor b);
    layer6_outputs(4211) <= a or b;
    layer6_outputs(4212) <= not (a xor b);
    layer6_outputs(4213) <= b and not a;
    layer6_outputs(4214) <= b and not a;
    layer6_outputs(4215) <= not b;
    layer6_outputs(4216) <= a or b;
    layer6_outputs(4217) <= a xor b;
    layer6_outputs(4218) <= a xor b;
    layer6_outputs(4219) <= a xor b;
    layer6_outputs(4220) <= a;
    layer6_outputs(4221) <= not b or a;
    layer6_outputs(4222) <= not b;
    layer6_outputs(4223) <= a or b;
    layer6_outputs(4224) <= not a;
    layer6_outputs(4225) <= b;
    layer6_outputs(4226) <= not a or b;
    layer6_outputs(4227) <= not b or a;
    layer6_outputs(4228) <= a xor b;
    layer6_outputs(4229) <= b;
    layer6_outputs(4230) <= not a;
    layer6_outputs(4231) <= not b or a;
    layer6_outputs(4232) <= b and not a;
    layer6_outputs(4233) <= b;
    layer6_outputs(4234) <= not b;
    layer6_outputs(4235) <= not (a xor b);
    layer6_outputs(4236) <= not (a or b);
    layer6_outputs(4237) <= a;
    layer6_outputs(4238) <= not (a xor b);
    layer6_outputs(4239) <= not (a xor b);
    layer6_outputs(4240) <= not (a or b);
    layer6_outputs(4241) <= not (a xor b);
    layer6_outputs(4242) <= a and not b;
    layer6_outputs(4243) <= a or b;
    layer6_outputs(4244) <= not (a xor b);
    layer6_outputs(4245) <= a or b;
    layer6_outputs(4246) <= a and b;
    layer6_outputs(4247) <= a xor b;
    layer6_outputs(4248) <= b;
    layer6_outputs(4249) <= b;
    layer6_outputs(4250) <= not (a and b);
    layer6_outputs(4251) <= b;
    layer6_outputs(4252) <= a xor b;
    layer6_outputs(4253) <= a;
    layer6_outputs(4254) <= not (a xor b);
    layer6_outputs(4255) <= a or b;
    layer6_outputs(4256) <= b;
    layer6_outputs(4257) <= not (a xor b);
    layer6_outputs(4258) <= b and not a;
    layer6_outputs(4259) <= not (a and b);
    layer6_outputs(4260) <= not b or a;
    layer6_outputs(4261) <= not b;
    layer6_outputs(4262) <= not (a or b);
    layer6_outputs(4263) <= a or b;
    layer6_outputs(4264) <= a;
    layer6_outputs(4265) <= a and not b;
    layer6_outputs(4266) <= a;
    layer6_outputs(4267) <= not a;
    layer6_outputs(4268) <= not b;
    layer6_outputs(4269) <= a and b;
    layer6_outputs(4270) <= a xor b;
    layer6_outputs(4271) <= not a or b;
    layer6_outputs(4272) <= not b;
    layer6_outputs(4273) <= not (a and b);
    layer6_outputs(4274) <= not a;
    layer6_outputs(4275) <= a;
    layer6_outputs(4276) <= b;
    layer6_outputs(4277) <= b;
    layer6_outputs(4278) <= not (a and b);
    layer6_outputs(4279) <= not b or a;
    layer6_outputs(4280) <= not (a and b);
    layer6_outputs(4281) <= not b;
    layer6_outputs(4282) <= a;
    layer6_outputs(4283) <= b;
    layer6_outputs(4284) <= not a;
    layer6_outputs(4285) <= not (a xor b);
    layer6_outputs(4286) <= a;
    layer6_outputs(4287) <= not b;
    layer6_outputs(4288) <= b;
    layer6_outputs(4289) <= not (a or b);
    layer6_outputs(4290) <= not (a xor b);
    layer6_outputs(4291) <= not a;
    layer6_outputs(4292) <= not a;
    layer6_outputs(4293) <= a and b;
    layer6_outputs(4294) <= not (a xor b);
    layer6_outputs(4295) <= not (a or b);
    layer6_outputs(4296) <= b and not a;
    layer6_outputs(4297) <= a and not b;
    layer6_outputs(4298) <= a;
    layer6_outputs(4299) <= b;
    layer6_outputs(4300) <= not (a or b);
    layer6_outputs(4301) <= not a;
    layer6_outputs(4302) <= not a;
    layer6_outputs(4303) <= not a or b;
    layer6_outputs(4304) <= not (a xor b);
    layer6_outputs(4305) <= not (a or b);
    layer6_outputs(4306) <= '1';
    layer6_outputs(4307) <= a xor b;
    layer6_outputs(4308) <= a xor b;
    layer6_outputs(4309) <= not (a and b);
    layer6_outputs(4310) <= a;
    layer6_outputs(4311) <= not a;
    layer6_outputs(4312) <= '0';
    layer6_outputs(4313) <= not a;
    layer6_outputs(4314) <= a;
    layer6_outputs(4315) <= a xor b;
    layer6_outputs(4316) <= not b or a;
    layer6_outputs(4317) <= not a;
    layer6_outputs(4318) <= not (a and b);
    layer6_outputs(4319) <= not b;
    layer6_outputs(4320) <= b and not a;
    layer6_outputs(4321) <= b;
    layer6_outputs(4322) <= b;
    layer6_outputs(4323) <= not b;
    layer6_outputs(4324) <= b;
    layer6_outputs(4325) <= a;
    layer6_outputs(4326) <= a;
    layer6_outputs(4327) <= a and not b;
    layer6_outputs(4328) <= not b;
    layer6_outputs(4329) <= not a or b;
    layer6_outputs(4330) <= not b or a;
    layer6_outputs(4331) <= not (a or b);
    layer6_outputs(4332) <= a xor b;
    layer6_outputs(4333) <= a xor b;
    layer6_outputs(4334) <= b;
    layer6_outputs(4335) <= not (a and b);
    layer6_outputs(4336) <= a xor b;
    layer6_outputs(4337) <= b;
    layer6_outputs(4338) <= not a;
    layer6_outputs(4339) <= a;
    layer6_outputs(4340) <= a;
    layer6_outputs(4341) <= b;
    layer6_outputs(4342) <= not a or b;
    layer6_outputs(4343) <= a xor b;
    layer6_outputs(4344) <= a and not b;
    layer6_outputs(4345) <= not a or b;
    layer6_outputs(4346) <= b;
    layer6_outputs(4347) <= not b;
    layer6_outputs(4348) <= not b;
    layer6_outputs(4349) <= a;
    layer6_outputs(4350) <= not b;
    layer6_outputs(4351) <= not a;
    layer6_outputs(4352) <= a;
    layer6_outputs(4353) <= a;
    layer6_outputs(4354) <= a and b;
    layer6_outputs(4355) <= a;
    layer6_outputs(4356) <= b;
    layer6_outputs(4357) <= a xor b;
    layer6_outputs(4358) <= not (a xor b);
    layer6_outputs(4359) <= not a or b;
    layer6_outputs(4360) <= not a or b;
    layer6_outputs(4361) <= a and not b;
    layer6_outputs(4362) <= a xor b;
    layer6_outputs(4363) <= a;
    layer6_outputs(4364) <= a xor b;
    layer6_outputs(4365) <= not a;
    layer6_outputs(4366) <= a;
    layer6_outputs(4367) <= b and not a;
    layer6_outputs(4368) <= a;
    layer6_outputs(4369) <= a;
    layer6_outputs(4370) <= a and b;
    layer6_outputs(4371) <= not b;
    layer6_outputs(4372) <= '0';
    layer6_outputs(4373) <= not (a xor b);
    layer6_outputs(4374) <= not (a xor b);
    layer6_outputs(4375) <= not (a xor b);
    layer6_outputs(4376) <= not b or a;
    layer6_outputs(4377) <= not (a xor b);
    layer6_outputs(4378) <= b;
    layer6_outputs(4379) <= not b or a;
    layer6_outputs(4380) <= a xor b;
    layer6_outputs(4381) <= not (a xor b);
    layer6_outputs(4382) <= a xor b;
    layer6_outputs(4383) <= not b;
    layer6_outputs(4384) <= a and b;
    layer6_outputs(4385) <= b;
    layer6_outputs(4386) <= a;
    layer6_outputs(4387) <= not a;
    layer6_outputs(4388) <= a and not b;
    layer6_outputs(4389) <= not b;
    layer6_outputs(4390) <= b;
    layer6_outputs(4391) <= not (a or b);
    layer6_outputs(4392) <= not a;
    layer6_outputs(4393) <= b;
    layer6_outputs(4394) <= not (a xor b);
    layer6_outputs(4395) <= a or b;
    layer6_outputs(4396) <= a xor b;
    layer6_outputs(4397) <= not a;
    layer6_outputs(4398) <= a or b;
    layer6_outputs(4399) <= a xor b;
    layer6_outputs(4400) <= not (a or b);
    layer6_outputs(4401) <= b;
    layer6_outputs(4402) <= b;
    layer6_outputs(4403) <= b;
    layer6_outputs(4404) <= b;
    layer6_outputs(4405) <= not a;
    layer6_outputs(4406) <= not b;
    layer6_outputs(4407) <= not (a xor b);
    layer6_outputs(4408) <= a and b;
    layer6_outputs(4409) <= a and not b;
    layer6_outputs(4410) <= not (a xor b);
    layer6_outputs(4411) <= a;
    layer6_outputs(4412) <= b and not a;
    layer6_outputs(4413) <= not a;
    layer6_outputs(4414) <= not (a xor b);
    layer6_outputs(4415) <= a and b;
    layer6_outputs(4416) <= a;
    layer6_outputs(4417) <= not b or a;
    layer6_outputs(4418) <= not b;
    layer6_outputs(4419) <= not b;
    layer6_outputs(4420) <= a;
    layer6_outputs(4421) <= b;
    layer6_outputs(4422) <= not b or a;
    layer6_outputs(4423) <= a xor b;
    layer6_outputs(4424) <= a xor b;
    layer6_outputs(4425) <= a or b;
    layer6_outputs(4426) <= not a;
    layer6_outputs(4427) <= not a;
    layer6_outputs(4428) <= a xor b;
    layer6_outputs(4429) <= a;
    layer6_outputs(4430) <= a or b;
    layer6_outputs(4431) <= not a;
    layer6_outputs(4432) <= not (a or b);
    layer6_outputs(4433) <= not b;
    layer6_outputs(4434) <= a and b;
    layer6_outputs(4435) <= not b or a;
    layer6_outputs(4436) <= b;
    layer6_outputs(4437) <= not (a xor b);
    layer6_outputs(4438) <= a;
    layer6_outputs(4439) <= not (a xor b);
    layer6_outputs(4440) <= a;
    layer6_outputs(4441) <= '0';
    layer6_outputs(4442) <= not b or a;
    layer6_outputs(4443) <= not (a xor b);
    layer6_outputs(4444) <= b;
    layer6_outputs(4445) <= a and b;
    layer6_outputs(4446) <= not a;
    layer6_outputs(4447) <= not (a and b);
    layer6_outputs(4448) <= not b;
    layer6_outputs(4449) <= a;
    layer6_outputs(4450) <= b and not a;
    layer6_outputs(4451) <= b;
    layer6_outputs(4452) <= a and not b;
    layer6_outputs(4453) <= a;
    layer6_outputs(4454) <= a xor b;
    layer6_outputs(4455) <= not (a and b);
    layer6_outputs(4456) <= a;
    layer6_outputs(4457) <= not b;
    layer6_outputs(4458) <= a xor b;
    layer6_outputs(4459) <= not b or a;
    layer6_outputs(4460) <= b;
    layer6_outputs(4461) <= b;
    layer6_outputs(4462) <= a;
    layer6_outputs(4463) <= a xor b;
    layer6_outputs(4464) <= not b or a;
    layer6_outputs(4465) <= a and b;
    layer6_outputs(4466) <= b;
    layer6_outputs(4467) <= a xor b;
    layer6_outputs(4468) <= a;
    layer6_outputs(4469) <= a xor b;
    layer6_outputs(4470) <= a and not b;
    layer6_outputs(4471) <= not b;
    layer6_outputs(4472) <= a or b;
    layer6_outputs(4473) <= a;
    layer6_outputs(4474) <= b;
    layer6_outputs(4475) <= '0';
    layer6_outputs(4476) <= not b;
    layer6_outputs(4477) <= b;
    layer6_outputs(4478) <= a;
    layer6_outputs(4479) <= a xor b;
    layer6_outputs(4480) <= not a;
    layer6_outputs(4481) <= a and not b;
    layer6_outputs(4482) <= not b;
    layer6_outputs(4483) <= not (a xor b);
    layer6_outputs(4484) <= not (a or b);
    layer6_outputs(4485) <= a xor b;
    layer6_outputs(4486) <= a;
    layer6_outputs(4487) <= not a;
    layer6_outputs(4488) <= not a;
    layer6_outputs(4489) <= a xor b;
    layer6_outputs(4490) <= not b;
    layer6_outputs(4491) <= a and b;
    layer6_outputs(4492) <= b;
    layer6_outputs(4493) <= not b;
    layer6_outputs(4494) <= a and b;
    layer6_outputs(4495) <= not (a xor b);
    layer6_outputs(4496) <= b;
    layer6_outputs(4497) <= not b;
    layer6_outputs(4498) <= a;
    layer6_outputs(4499) <= b and not a;
    layer6_outputs(4500) <= a;
    layer6_outputs(4501) <= a;
    layer6_outputs(4502) <= not b;
    layer6_outputs(4503) <= not (a xor b);
    layer6_outputs(4504) <= b;
    layer6_outputs(4505) <= not a;
    layer6_outputs(4506) <= b and not a;
    layer6_outputs(4507) <= not a or b;
    layer6_outputs(4508) <= not b;
    layer6_outputs(4509) <= not (a or b);
    layer6_outputs(4510) <= a xor b;
    layer6_outputs(4511) <= b and not a;
    layer6_outputs(4512) <= a xor b;
    layer6_outputs(4513) <= a;
    layer6_outputs(4514) <= a;
    layer6_outputs(4515) <= a or b;
    layer6_outputs(4516) <= not b;
    layer6_outputs(4517) <= not (a and b);
    layer6_outputs(4518) <= a;
    layer6_outputs(4519) <= a and not b;
    layer6_outputs(4520) <= b and not a;
    layer6_outputs(4521) <= b;
    layer6_outputs(4522) <= not a;
    layer6_outputs(4523) <= not a;
    layer6_outputs(4524) <= not b;
    layer6_outputs(4525) <= not b or a;
    layer6_outputs(4526) <= not b or a;
    layer6_outputs(4527) <= a;
    layer6_outputs(4528) <= not (a and b);
    layer6_outputs(4529) <= b;
    layer6_outputs(4530) <= a or b;
    layer6_outputs(4531) <= not a or b;
    layer6_outputs(4532) <= b;
    layer6_outputs(4533) <= not b;
    layer6_outputs(4534) <= not (a and b);
    layer6_outputs(4535) <= not b;
    layer6_outputs(4536) <= not b;
    layer6_outputs(4537) <= b;
    layer6_outputs(4538) <= b;
    layer6_outputs(4539) <= a xor b;
    layer6_outputs(4540) <= not a;
    layer6_outputs(4541) <= not b;
    layer6_outputs(4542) <= a xor b;
    layer6_outputs(4543) <= a and b;
    layer6_outputs(4544) <= a;
    layer6_outputs(4545) <= a;
    layer6_outputs(4546) <= not b;
    layer6_outputs(4547) <= b;
    layer6_outputs(4548) <= '1';
    layer6_outputs(4549) <= a;
    layer6_outputs(4550) <= not (a xor b);
    layer6_outputs(4551) <= a xor b;
    layer6_outputs(4552) <= not (a and b);
    layer6_outputs(4553) <= a xor b;
    layer6_outputs(4554) <= a or b;
    layer6_outputs(4555) <= a xor b;
    layer6_outputs(4556) <= not b;
    layer6_outputs(4557) <= b;
    layer6_outputs(4558) <= not a;
    layer6_outputs(4559) <= a;
    layer6_outputs(4560) <= not (a or b);
    layer6_outputs(4561) <= not (a and b);
    layer6_outputs(4562) <= not a;
    layer6_outputs(4563) <= not (a xor b);
    layer6_outputs(4564) <= b and not a;
    layer6_outputs(4565) <= a and not b;
    layer6_outputs(4566) <= not b or a;
    layer6_outputs(4567) <= b;
    layer6_outputs(4568) <= b;
    layer6_outputs(4569) <= a xor b;
    layer6_outputs(4570) <= not b;
    layer6_outputs(4571) <= a;
    layer6_outputs(4572) <= not a or b;
    layer6_outputs(4573) <= b;
    layer6_outputs(4574) <= not (a xor b);
    layer6_outputs(4575) <= b;
    layer6_outputs(4576) <= b and not a;
    layer6_outputs(4577) <= b;
    layer6_outputs(4578) <= '1';
    layer6_outputs(4579) <= b;
    layer6_outputs(4580) <= not a;
    layer6_outputs(4581) <= a and not b;
    layer6_outputs(4582) <= not a;
    layer6_outputs(4583) <= not (a xor b);
    layer6_outputs(4584) <= not b;
    layer6_outputs(4585) <= not b or a;
    layer6_outputs(4586) <= not b or a;
    layer6_outputs(4587) <= not a;
    layer6_outputs(4588) <= b;
    layer6_outputs(4589) <= not b or a;
    layer6_outputs(4590) <= not (a xor b);
    layer6_outputs(4591) <= not a;
    layer6_outputs(4592) <= a xor b;
    layer6_outputs(4593) <= not a;
    layer6_outputs(4594) <= a xor b;
    layer6_outputs(4595) <= not a;
    layer6_outputs(4596) <= not b;
    layer6_outputs(4597) <= a xor b;
    layer6_outputs(4598) <= not a;
    layer6_outputs(4599) <= b and not a;
    layer6_outputs(4600) <= not a;
    layer6_outputs(4601) <= not a or b;
    layer6_outputs(4602) <= a or b;
    layer6_outputs(4603) <= a or b;
    layer6_outputs(4604) <= not a;
    layer6_outputs(4605) <= not a;
    layer6_outputs(4606) <= not a;
    layer6_outputs(4607) <= not a;
    layer6_outputs(4608) <= not a or b;
    layer6_outputs(4609) <= not b;
    layer6_outputs(4610) <= b;
    layer6_outputs(4611) <= not b or a;
    layer6_outputs(4612) <= a xor b;
    layer6_outputs(4613) <= a xor b;
    layer6_outputs(4614) <= not b;
    layer6_outputs(4615) <= a;
    layer6_outputs(4616) <= a;
    layer6_outputs(4617) <= not (a and b);
    layer6_outputs(4618) <= not (a and b);
    layer6_outputs(4619) <= not (a xor b);
    layer6_outputs(4620) <= not (a and b);
    layer6_outputs(4621) <= a and not b;
    layer6_outputs(4622) <= a;
    layer6_outputs(4623) <= a or b;
    layer6_outputs(4624) <= not b;
    layer6_outputs(4625) <= a xor b;
    layer6_outputs(4626) <= b;
    layer6_outputs(4627) <= a;
    layer6_outputs(4628) <= a xor b;
    layer6_outputs(4629) <= not b;
    layer6_outputs(4630) <= a;
    layer6_outputs(4631) <= b;
    layer6_outputs(4632) <= a or b;
    layer6_outputs(4633) <= not (a xor b);
    layer6_outputs(4634) <= a xor b;
    layer6_outputs(4635) <= not a;
    layer6_outputs(4636) <= b;
    layer6_outputs(4637) <= a;
    layer6_outputs(4638) <= not b;
    layer6_outputs(4639) <= not (a xor b);
    layer6_outputs(4640) <= not (a and b);
    layer6_outputs(4641) <= not (a or b);
    layer6_outputs(4642) <= not (a or b);
    layer6_outputs(4643) <= a xor b;
    layer6_outputs(4644) <= not a or b;
    layer6_outputs(4645) <= not (a or b);
    layer6_outputs(4646) <= not (a and b);
    layer6_outputs(4647) <= a;
    layer6_outputs(4648) <= a;
    layer6_outputs(4649) <= not (a or b);
    layer6_outputs(4650) <= a or b;
    layer6_outputs(4651) <= not b;
    layer6_outputs(4652) <= a and b;
    layer6_outputs(4653) <= a;
    layer6_outputs(4654) <= a and not b;
    layer6_outputs(4655) <= '1';
    layer6_outputs(4656) <= b and not a;
    layer6_outputs(4657) <= not b;
    layer6_outputs(4658) <= b and not a;
    layer6_outputs(4659) <= not (a or b);
    layer6_outputs(4660) <= not a or b;
    layer6_outputs(4661) <= a xor b;
    layer6_outputs(4662) <= a and b;
    layer6_outputs(4663) <= not b;
    layer6_outputs(4664) <= not a;
    layer6_outputs(4665) <= b;
    layer6_outputs(4666) <= a;
    layer6_outputs(4667) <= b;
    layer6_outputs(4668) <= a and b;
    layer6_outputs(4669) <= not b;
    layer6_outputs(4670) <= not (a xor b);
    layer6_outputs(4671) <= a;
    layer6_outputs(4672) <= not a or b;
    layer6_outputs(4673) <= not b or a;
    layer6_outputs(4674) <= a and not b;
    layer6_outputs(4675) <= not (a xor b);
    layer6_outputs(4676) <= b;
    layer6_outputs(4677) <= b;
    layer6_outputs(4678) <= not a;
    layer6_outputs(4679) <= a and b;
    layer6_outputs(4680) <= a;
    layer6_outputs(4681) <= b and not a;
    layer6_outputs(4682) <= a xor b;
    layer6_outputs(4683) <= not (a xor b);
    layer6_outputs(4684) <= not (a xor b);
    layer6_outputs(4685) <= not b;
    layer6_outputs(4686) <= not (a xor b);
    layer6_outputs(4687) <= a;
    layer6_outputs(4688) <= not b;
    layer6_outputs(4689) <= b;
    layer6_outputs(4690) <= not b;
    layer6_outputs(4691) <= not (a xor b);
    layer6_outputs(4692) <= b and not a;
    layer6_outputs(4693) <= a;
    layer6_outputs(4694) <= a and not b;
    layer6_outputs(4695) <= a xor b;
    layer6_outputs(4696) <= b;
    layer6_outputs(4697) <= b and not a;
    layer6_outputs(4698) <= a;
    layer6_outputs(4699) <= not (a xor b);
    layer6_outputs(4700) <= not a;
    layer6_outputs(4701) <= not b;
    layer6_outputs(4702) <= not a or b;
    layer6_outputs(4703) <= not a;
    layer6_outputs(4704) <= not (a xor b);
    layer6_outputs(4705) <= a xor b;
    layer6_outputs(4706) <= a xor b;
    layer6_outputs(4707) <= a xor b;
    layer6_outputs(4708) <= not b;
    layer6_outputs(4709) <= a;
    layer6_outputs(4710) <= not a or b;
    layer6_outputs(4711) <= a or b;
    layer6_outputs(4712) <= b;
    layer6_outputs(4713) <= not (a or b);
    layer6_outputs(4714) <= not a or b;
    layer6_outputs(4715) <= not (a or b);
    layer6_outputs(4716) <= a;
    layer6_outputs(4717) <= not b;
    layer6_outputs(4718) <= a or b;
    layer6_outputs(4719) <= b and not a;
    layer6_outputs(4720) <= not a;
    layer6_outputs(4721) <= a;
    layer6_outputs(4722) <= not (a xor b);
    layer6_outputs(4723) <= not b;
    layer6_outputs(4724) <= not b;
    layer6_outputs(4725) <= a;
    layer6_outputs(4726) <= b and not a;
    layer6_outputs(4727) <= not b or a;
    layer6_outputs(4728) <= not a;
    layer6_outputs(4729) <= not b or a;
    layer6_outputs(4730) <= b;
    layer6_outputs(4731) <= not (a or b);
    layer6_outputs(4732) <= not (a xor b);
    layer6_outputs(4733) <= a and b;
    layer6_outputs(4734) <= a and b;
    layer6_outputs(4735) <= a and b;
    layer6_outputs(4736) <= not b or a;
    layer6_outputs(4737) <= a xor b;
    layer6_outputs(4738) <= not b or a;
    layer6_outputs(4739) <= a;
    layer6_outputs(4740) <= not b or a;
    layer6_outputs(4741) <= a and b;
    layer6_outputs(4742) <= a;
    layer6_outputs(4743) <= not b or a;
    layer6_outputs(4744) <= a;
    layer6_outputs(4745) <= not (a xor b);
    layer6_outputs(4746) <= b;
    layer6_outputs(4747) <= a xor b;
    layer6_outputs(4748) <= a xor b;
    layer6_outputs(4749) <= not b;
    layer6_outputs(4750) <= b;
    layer6_outputs(4751) <= a and b;
    layer6_outputs(4752) <= not b or a;
    layer6_outputs(4753) <= a;
    layer6_outputs(4754) <= not b or a;
    layer6_outputs(4755) <= not b or a;
    layer6_outputs(4756) <= not b;
    layer6_outputs(4757) <= b;
    layer6_outputs(4758) <= a xor b;
    layer6_outputs(4759) <= a xor b;
    layer6_outputs(4760) <= not b;
    layer6_outputs(4761) <= not b;
    layer6_outputs(4762) <= a xor b;
    layer6_outputs(4763) <= b;
    layer6_outputs(4764) <= a;
    layer6_outputs(4765) <= not b;
    layer6_outputs(4766) <= not a or b;
    layer6_outputs(4767) <= a;
    layer6_outputs(4768) <= not (a xor b);
    layer6_outputs(4769) <= b;
    layer6_outputs(4770) <= not b;
    layer6_outputs(4771) <= not a or b;
    layer6_outputs(4772) <= b;
    layer6_outputs(4773) <= a or b;
    layer6_outputs(4774) <= not a;
    layer6_outputs(4775) <= a or b;
    layer6_outputs(4776) <= b;
    layer6_outputs(4777) <= not (a and b);
    layer6_outputs(4778) <= a or b;
    layer6_outputs(4779) <= not (a xor b);
    layer6_outputs(4780) <= not b or a;
    layer6_outputs(4781) <= b and not a;
    layer6_outputs(4782) <= a and b;
    layer6_outputs(4783) <= not b;
    layer6_outputs(4784) <= not (a and b);
    layer6_outputs(4785) <= a and b;
    layer6_outputs(4786) <= not b;
    layer6_outputs(4787) <= a;
    layer6_outputs(4788) <= not (a xor b);
    layer6_outputs(4789) <= not a;
    layer6_outputs(4790) <= not b or a;
    layer6_outputs(4791) <= b;
    layer6_outputs(4792) <= a;
    layer6_outputs(4793) <= b and not a;
    layer6_outputs(4794) <= a and b;
    layer6_outputs(4795) <= not a;
    layer6_outputs(4796) <= b and not a;
    layer6_outputs(4797) <= a xor b;
    layer6_outputs(4798) <= not (a xor b);
    layer6_outputs(4799) <= not (a xor b);
    layer6_outputs(4800) <= b and not a;
    layer6_outputs(4801) <= not b;
    layer6_outputs(4802) <= b;
    layer6_outputs(4803) <= a and not b;
    layer6_outputs(4804) <= a and b;
    layer6_outputs(4805) <= not a;
    layer6_outputs(4806) <= not a or b;
    layer6_outputs(4807) <= not b;
    layer6_outputs(4808) <= a xor b;
    layer6_outputs(4809) <= not a;
    layer6_outputs(4810) <= not a;
    layer6_outputs(4811) <= b;
    layer6_outputs(4812) <= b;
    layer6_outputs(4813) <= not (a xor b);
    layer6_outputs(4814) <= b;
    layer6_outputs(4815) <= not a or b;
    layer6_outputs(4816) <= a and not b;
    layer6_outputs(4817) <= not b;
    layer6_outputs(4818) <= b and not a;
    layer6_outputs(4819) <= a or b;
    layer6_outputs(4820) <= a;
    layer6_outputs(4821) <= b;
    layer6_outputs(4822) <= not (a and b);
    layer6_outputs(4823) <= a xor b;
    layer6_outputs(4824) <= b and not a;
    layer6_outputs(4825) <= b;
    layer6_outputs(4826) <= not (a xor b);
    layer6_outputs(4827) <= not b;
    layer6_outputs(4828) <= not (a xor b);
    layer6_outputs(4829) <= b and not a;
    layer6_outputs(4830) <= not a;
    layer6_outputs(4831) <= a and not b;
    layer6_outputs(4832) <= not b;
    layer6_outputs(4833) <= a and not b;
    layer6_outputs(4834) <= a;
    layer6_outputs(4835) <= a;
    layer6_outputs(4836) <= b;
    layer6_outputs(4837) <= b;
    layer6_outputs(4838) <= not (a xor b);
    layer6_outputs(4839) <= a;
    layer6_outputs(4840) <= not b;
    layer6_outputs(4841) <= not a;
    layer6_outputs(4842) <= not b;
    layer6_outputs(4843) <= not (a or b);
    layer6_outputs(4844) <= not b or a;
    layer6_outputs(4845) <= b;
    layer6_outputs(4846) <= not a;
    layer6_outputs(4847) <= not b;
    layer6_outputs(4848) <= a;
    layer6_outputs(4849) <= a or b;
    layer6_outputs(4850) <= not b;
    layer6_outputs(4851) <= not (a xor b);
    layer6_outputs(4852) <= a and not b;
    layer6_outputs(4853) <= a;
    layer6_outputs(4854) <= b;
    layer6_outputs(4855) <= b and not a;
    layer6_outputs(4856) <= a xor b;
    layer6_outputs(4857) <= a xor b;
    layer6_outputs(4858) <= a and b;
    layer6_outputs(4859) <= a and not b;
    layer6_outputs(4860) <= not a;
    layer6_outputs(4861) <= a;
    layer6_outputs(4862) <= a xor b;
    layer6_outputs(4863) <= not a;
    layer6_outputs(4864) <= b and not a;
    layer6_outputs(4865) <= a;
    layer6_outputs(4866) <= b;
    layer6_outputs(4867) <= a and not b;
    layer6_outputs(4868) <= not a;
    layer6_outputs(4869) <= not (a or b);
    layer6_outputs(4870) <= a and b;
    layer6_outputs(4871) <= not b or a;
    layer6_outputs(4872) <= not b;
    layer6_outputs(4873) <= not (a and b);
    layer6_outputs(4874) <= a and not b;
    layer6_outputs(4875) <= a;
    layer6_outputs(4876) <= not a or b;
    layer6_outputs(4877) <= not (a xor b);
    layer6_outputs(4878) <= not a or b;
    layer6_outputs(4879) <= a xor b;
    layer6_outputs(4880) <= a xor b;
    layer6_outputs(4881) <= b;
    layer6_outputs(4882) <= a;
    layer6_outputs(4883) <= a and b;
    layer6_outputs(4884) <= a;
    layer6_outputs(4885) <= not (a or b);
    layer6_outputs(4886) <= b;
    layer6_outputs(4887) <= a and not b;
    layer6_outputs(4888) <= a;
    layer6_outputs(4889) <= not a;
    layer6_outputs(4890) <= a;
    layer6_outputs(4891) <= not a or b;
    layer6_outputs(4892) <= a or b;
    layer6_outputs(4893) <= not (a or b);
    layer6_outputs(4894) <= a;
    layer6_outputs(4895) <= a;
    layer6_outputs(4896) <= not (a xor b);
    layer6_outputs(4897) <= not b or a;
    layer6_outputs(4898) <= not (a and b);
    layer6_outputs(4899) <= not b or a;
    layer6_outputs(4900) <= a and b;
    layer6_outputs(4901) <= not (a and b);
    layer6_outputs(4902) <= not a;
    layer6_outputs(4903) <= b;
    layer6_outputs(4904) <= a and not b;
    layer6_outputs(4905) <= not (a xor b);
    layer6_outputs(4906) <= b;
    layer6_outputs(4907) <= not a;
    layer6_outputs(4908) <= a xor b;
    layer6_outputs(4909) <= a xor b;
    layer6_outputs(4910) <= b;
    layer6_outputs(4911) <= a xor b;
    layer6_outputs(4912) <= a;
    layer6_outputs(4913) <= a xor b;
    layer6_outputs(4914) <= not (a or b);
    layer6_outputs(4915) <= not (a or b);
    layer6_outputs(4916) <= not a;
    layer6_outputs(4917) <= not a or b;
    layer6_outputs(4918) <= not a or b;
    layer6_outputs(4919) <= a xor b;
    layer6_outputs(4920) <= a;
    layer6_outputs(4921) <= b;
    layer6_outputs(4922) <= a xor b;
    layer6_outputs(4923) <= not b or a;
    layer6_outputs(4924) <= a or b;
    layer6_outputs(4925) <= a or b;
    layer6_outputs(4926) <= a xor b;
    layer6_outputs(4927) <= a;
    layer6_outputs(4928) <= a or b;
    layer6_outputs(4929) <= b;
    layer6_outputs(4930) <= a or b;
    layer6_outputs(4931) <= a and not b;
    layer6_outputs(4932) <= not a;
    layer6_outputs(4933) <= b;
    layer6_outputs(4934) <= a;
    layer6_outputs(4935) <= b;
    layer6_outputs(4936) <= a and b;
    layer6_outputs(4937) <= not b;
    layer6_outputs(4938) <= a or b;
    layer6_outputs(4939) <= a;
    layer6_outputs(4940) <= b;
    layer6_outputs(4941) <= b;
    layer6_outputs(4942) <= a;
    layer6_outputs(4943) <= a xor b;
    layer6_outputs(4944) <= b;
    layer6_outputs(4945) <= not (a xor b);
    layer6_outputs(4946) <= b;
    layer6_outputs(4947) <= b;
    layer6_outputs(4948) <= a;
    layer6_outputs(4949) <= not b;
    layer6_outputs(4950) <= a xor b;
    layer6_outputs(4951) <= not (a xor b);
    layer6_outputs(4952) <= not (a xor b);
    layer6_outputs(4953) <= a xor b;
    layer6_outputs(4954) <= a;
    layer6_outputs(4955) <= b;
    layer6_outputs(4956) <= not (a and b);
    layer6_outputs(4957) <= a or b;
    layer6_outputs(4958) <= not b;
    layer6_outputs(4959) <= b;
    layer6_outputs(4960) <= a or b;
    layer6_outputs(4961) <= a and not b;
    layer6_outputs(4962) <= not a;
    layer6_outputs(4963) <= a or b;
    layer6_outputs(4964) <= not (a and b);
    layer6_outputs(4965) <= not (a or b);
    layer6_outputs(4966) <= not (a or b);
    layer6_outputs(4967) <= not a;
    layer6_outputs(4968) <= not a;
    layer6_outputs(4969) <= not b;
    layer6_outputs(4970) <= b;
    layer6_outputs(4971) <= not b;
    layer6_outputs(4972) <= b;
    layer6_outputs(4973) <= a;
    layer6_outputs(4974) <= a xor b;
    layer6_outputs(4975) <= not b;
    layer6_outputs(4976) <= a and not b;
    layer6_outputs(4977) <= a;
    layer6_outputs(4978) <= a xor b;
    layer6_outputs(4979) <= not a;
    layer6_outputs(4980) <= not b;
    layer6_outputs(4981) <= a;
    layer6_outputs(4982) <= not (a xor b);
    layer6_outputs(4983) <= b;
    layer6_outputs(4984) <= a and not b;
    layer6_outputs(4985) <= b and not a;
    layer6_outputs(4986) <= not a;
    layer6_outputs(4987) <= not a;
    layer6_outputs(4988) <= a or b;
    layer6_outputs(4989) <= b;
    layer6_outputs(4990) <= b;
    layer6_outputs(4991) <= not a;
    layer6_outputs(4992) <= not (a or b);
    layer6_outputs(4993) <= a;
    layer6_outputs(4994) <= not a;
    layer6_outputs(4995) <= a;
    layer6_outputs(4996) <= a or b;
    layer6_outputs(4997) <= not a;
    layer6_outputs(4998) <= not (a xor b);
    layer6_outputs(4999) <= not b or a;
    layer6_outputs(5000) <= not b;
    layer6_outputs(5001) <= b;
    layer6_outputs(5002) <= not a or b;
    layer6_outputs(5003) <= b;
    layer6_outputs(5004) <= not (a or b);
    layer6_outputs(5005) <= not a;
    layer6_outputs(5006) <= not a;
    layer6_outputs(5007) <= not b;
    layer6_outputs(5008) <= not a;
    layer6_outputs(5009) <= a;
    layer6_outputs(5010) <= b;
    layer6_outputs(5011) <= b and not a;
    layer6_outputs(5012) <= not a;
    layer6_outputs(5013) <= b;
    layer6_outputs(5014) <= not b;
    layer6_outputs(5015) <= a or b;
    layer6_outputs(5016) <= b;
    layer6_outputs(5017) <= a;
    layer6_outputs(5018) <= not a;
    layer6_outputs(5019) <= not b;
    layer6_outputs(5020) <= not (a xor b);
    layer6_outputs(5021) <= not b;
    layer6_outputs(5022) <= not (a and b);
    layer6_outputs(5023) <= a and not b;
    layer6_outputs(5024) <= a;
    layer6_outputs(5025) <= not b;
    layer6_outputs(5026) <= a;
    layer6_outputs(5027) <= not b or a;
    layer6_outputs(5028) <= a and not b;
    layer6_outputs(5029) <= not (a and b);
    layer6_outputs(5030) <= a xor b;
    layer6_outputs(5031) <= not a;
    layer6_outputs(5032) <= b;
    layer6_outputs(5033) <= not b;
    layer6_outputs(5034) <= b and not a;
    layer6_outputs(5035) <= b and not a;
    layer6_outputs(5036) <= a and b;
    layer6_outputs(5037) <= not (a and b);
    layer6_outputs(5038) <= a or b;
    layer6_outputs(5039) <= not (a and b);
    layer6_outputs(5040) <= not b;
    layer6_outputs(5041) <= a or b;
    layer6_outputs(5042) <= not (a and b);
    layer6_outputs(5043) <= a;
    layer6_outputs(5044) <= not (a or b);
    layer6_outputs(5045) <= a and not b;
    layer6_outputs(5046) <= not b;
    layer6_outputs(5047) <= not (a or b);
    layer6_outputs(5048) <= not b;
    layer6_outputs(5049) <= b;
    layer6_outputs(5050) <= not (a and b);
    layer6_outputs(5051) <= a;
    layer6_outputs(5052) <= not (a xor b);
    layer6_outputs(5053) <= a;
    layer6_outputs(5054) <= b and not a;
    layer6_outputs(5055) <= a and b;
    layer6_outputs(5056) <= a xor b;
    layer6_outputs(5057) <= b;
    layer6_outputs(5058) <= not b;
    layer6_outputs(5059) <= not b;
    layer6_outputs(5060) <= b;
    layer6_outputs(5061) <= not (a and b);
    layer6_outputs(5062) <= b;
    layer6_outputs(5063) <= b;
    layer6_outputs(5064) <= b;
    layer6_outputs(5065) <= a and not b;
    layer6_outputs(5066) <= a and not b;
    layer6_outputs(5067) <= not a or b;
    layer6_outputs(5068) <= not b;
    layer6_outputs(5069) <= a;
    layer6_outputs(5070) <= b;
    layer6_outputs(5071) <= not (a xor b);
    layer6_outputs(5072) <= a;
    layer6_outputs(5073) <= b;
    layer6_outputs(5074) <= a and not b;
    layer6_outputs(5075) <= a;
    layer6_outputs(5076) <= not (a or b);
    layer6_outputs(5077) <= a;
    layer6_outputs(5078) <= a;
    layer6_outputs(5079) <= a;
    layer6_outputs(5080) <= not b or a;
    layer6_outputs(5081) <= a and b;
    layer6_outputs(5082) <= not (a xor b);
    layer6_outputs(5083) <= not b;
    layer6_outputs(5084) <= a and not b;
    layer6_outputs(5085) <= not a;
    layer6_outputs(5086) <= a and b;
    layer6_outputs(5087) <= a;
    layer6_outputs(5088) <= not (a or b);
    layer6_outputs(5089) <= not (a xor b);
    layer6_outputs(5090) <= b and not a;
    layer6_outputs(5091) <= a and not b;
    layer6_outputs(5092) <= not a;
    layer6_outputs(5093) <= a;
    layer6_outputs(5094) <= not (a and b);
    layer6_outputs(5095) <= b;
    layer6_outputs(5096) <= a or b;
    layer6_outputs(5097) <= b and not a;
    layer6_outputs(5098) <= b and not a;
    layer6_outputs(5099) <= b;
    layer6_outputs(5100) <= a;
    layer6_outputs(5101) <= a or b;
    layer6_outputs(5102) <= a xor b;
    layer6_outputs(5103) <= not (a and b);
    layer6_outputs(5104) <= not a or b;
    layer6_outputs(5105) <= not a;
    layer6_outputs(5106) <= b;
    layer6_outputs(5107) <= not a or b;
    layer6_outputs(5108) <= not b;
    layer6_outputs(5109) <= b and not a;
    layer6_outputs(5110) <= not b;
    layer6_outputs(5111) <= not b or a;
    layer6_outputs(5112) <= not a;
    layer6_outputs(5113) <= a or b;
    layer6_outputs(5114) <= not a;
    layer6_outputs(5115) <= not b;
    layer6_outputs(5116) <= not (a or b);
    layer6_outputs(5117) <= not (a xor b);
    layer6_outputs(5118) <= a;
    layer6_outputs(5119) <= a;
    layer6_outputs(5120) <= a and b;
    layer6_outputs(5121) <= not (a or b);
    layer6_outputs(5122) <= b;
    layer6_outputs(5123) <= not b or a;
    layer6_outputs(5124) <= a or b;
    layer6_outputs(5125) <= not a or b;
    layer6_outputs(5126) <= a xor b;
    layer6_outputs(5127) <= b;
    layer6_outputs(5128) <= not (a or b);
    layer6_outputs(5129) <= not a;
    layer6_outputs(5130) <= b and not a;
    layer6_outputs(5131) <= a xor b;
    layer6_outputs(5132) <= a and not b;
    layer6_outputs(5133) <= not a;
    layer6_outputs(5134) <= not a or b;
    layer6_outputs(5135) <= b and not a;
    layer6_outputs(5136) <= not (a xor b);
    layer6_outputs(5137) <= not a;
    layer6_outputs(5138) <= a;
    layer6_outputs(5139) <= a or b;
    layer6_outputs(5140) <= not (a xor b);
    layer6_outputs(5141) <= a and b;
    layer6_outputs(5142) <= a;
    layer6_outputs(5143) <= not (a and b);
    layer6_outputs(5144) <= not (a and b);
    layer6_outputs(5145) <= not b;
    layer6_outputs(5146) <= not b;
    layer6_outputs(5147) <= not b;
    layer6_outputs(5148) <= not (a or b);
    layer6_outputs(5149) <= not a;
    layer6_outputs(5150) <= b and not a;
    layer6_outputs(5151) <= b;
    layer6_outputs(5152) <= not b;
    layer6_outputs(5153) <= not b;
    layer6_outputs(5154) <= not b;
    layer6_outputs(5155) <= a or b;
    layer6_outputs(5156) <= not (a xor b);
    layer6_outputs(5157) <= not a or b;
    layer6_outputs(5158) <= a;
    layer6_outputs(5159) <= not (a xor b);
    layer6_outputs(5160) <= not b or a;
    layer6_outputs(5161) <= not b;
    layer6_outputs(5162) <= not a;
    layer6_outputs(5163) <= not (a or b);
    layer6_outputs(5164) <= a xor b;
    layer6_outputs(5165) <= b;
    layer6_outputs(5166) <= b;
    layer6_outputs(5167) <= b and not a;
    layer6_outputs(5168) <= not a;
    layer6_outputs(5169) <= not b;
    layer6_outputs(5170) <= a xor b;
    layer6_outputs(5171) <= not (a or b);
    layer6_outputs(5172) <= not (a or b);
    layer6_outputs(5173) <= b;
    layer6_outputs(5174) <= a;
    layer6_outputs(5175) <= not a;
    layer6_outputs(5176) <= b and not a;
    layer6_outputs(5177) <= a;
    layer6_outputs(5178) <= not (a xor b);
    layer6_outputs(5179) <= not (a and b);
    layer6_outputs(5180) <= not b;
    layer6_outputs(5181) <= a xor b;
    layer6_outputs(5182) <= not b;
    layer6_outputs(5183) <= b;
    layer6_outputs(5184) <= a xor b;
    layer6_outputs(5185) <= not b;
    layer6_outputs(5186) <= a;
    layer6_outputs(5187) <= b;
    layer6_outputs(5188) <= not a;
    layer6_outputs(5189) <= not b;
    layer6_outputs(5190) <= b;
    layer6_outputs(5191) <= b;
    layer6_outputs(5192) <= not (a or b);
    layer6_outputs(5193) <= a and not b;
    layer6_outputs(5194) <= not (a or b);
    layer6_outputs(5195) <= not a;
    layer6_outputs(5196) <= not b;
    layer6_outputs(5197) <= a and b;
    layer6_outputs(5198) <= not (a or b);
    layer6_outputs(5199) <= b;
    layer6_outputs(5200) <= not b or a;
    layer6_outputs(5201) <= not a;
    layer6_outputs(5202) <= a;
    layer6_outputs(5203) <= not b;
    layer6_outputs(5204) <= not b or a;
    layer6_outputs(5205) <= not (a xor b);
    layer6_outputs(5206) <= a or b;
    layer6_outputs(5207) <= not b;
    layer6_outputs(5208) <= b;
    layer6_outputs(5209) <= a and not b;
    layer6_outputs(5210) <= b and not a;
    layer6_outputs(5211) <= a;
    layer6_outputs(5212) <= not b or a;
    layer6_outputs(5213) <= b;
    layer6_outputs(5214) <= b;
    layer6_outputs(5215) <= not (a xor b);
    layer6_outputs(5216) <= not (a and b);
    layer6_outputs(5217) <= not a;
    layer6_outputs(5218) <= a;
    layer6_outputs(5219) <= a or b;
    layer6_outputs(5220) <= not (a and b);
    layer6_outputs(5221) <= not a or b;
    layer6_outputs(5222) <= not a;
    layer6_outputs(5223) <= a xor b;
    layer6_outputs(5224) <= a;
    layer6_outputs(5225) <= not (a xor b);
    layer6_outputs(5226) <= a or b;
    layer6_outputs(5227) <= a and b;
    layer6_outputs(5228) <= a or b;
    layer6_outputs(5229) <= not (a xor b);
    layer6_outputs(5230) <= not b;
    layer6_outputs(5231) <= not a;
    layer6_outputs(5232) <= not b or a;
    layer6_outputs(5233) <= a and b;
    layer6_outputs(5234) <= not a;
    layer6_outputs(5235) <= not (a or b);
    layer6_outputs(5236) <= not (a and b);
    layer6_outputs(5237) <= a or b;
    layer6_outputs(5238) <= b and not a;
    layer6_outputs(5239) <= b and not a;
    layer6_outputs(5240) <= b;
    layer6_outputs(5241) <= a;
    layer6_outputs(5242) <= not (a and b);
    layer6_outputs(5243) <= not b;
    layer6_outputs(5244) <= a and b;
    layer6_outputs(5245) <= '1';
    layer6_outputs(5246) <= not b;
    layer6_outputs(5247) <= not (a xor b);
    layer6_outputs(5248) <= not (a xor b);
    layer6_outputs(5249) <= not (a or b);
    layer6_outputs(5250) <= not (a or b);
    layer6_outputs(5251) <= not a or b;
    layer6_outputs(5252) <= not a;
    layer6_outputs(5253) <= not (a or b);
    layer6_outputs(5254) <= not a;
    layer6_outputs(5255) <= not b;
    layer6_outputs(5256) <= not (a and b);
    layer6_outputs(5257) <= not a or b;
    layer6_outputs(5258) <= not a or b;
    layer6_outputs(5259) <= a and b;
    layer6_outputs(5260) <= not a;
    layer6_outputs(5261) <= not (a xor b);
    layer6_outputs(5262) <= b;
    layer6_outputs(5263) <= b and not a;
    layer6_outputs(5264) <= not (a and b);
    layer6_outputs(5265) <= a;
    layer6_outputs(5266) <= not (a xor b);
    layer6_outputs(5267) <= a;
    layer6_outputs(5268) <= a xor b;
    layer6_outputs(5269) <= a;
    layer6_outputs(5270) <= a;
    layer6_outputs(5271) <= a;
    layer6_outputs(5272) <= b;
    layer6_outputs(5273) <= a;
    layer6_outputs(5274) <= b;
    layer6_outputs(5275) <= not a;
    layer6_outputs(5276) <= a xor b;
    layer6_outputs(5277) <= not a;
    layer6_outputs(5278) <= not b;
    layer6_outputs(5279) <= a or b;
    layer6_outputs(5280) <= not (a xor b);
    layer6_outputs(5281) <= a xor b;
    layer6_outputs(5282) <= a or b;
    layer6_outputs(5283) <= not a;
    layer6_outputs(5284) <= not b or a;
    layer6_outputs(5285) <= not a;
    layer6_outputs(5286) <= b;
    layer6_outputs(5287) <= not b;
    layer6_outputs(5288) <= not (a xor b);
    layer6_outputs(5289) <= a and b;
    layer6_outputs(5290) <= a and not b;
    layer6_outputs(5291) <= a;
    layer6_outputs(5292) <= b and not a;
    layer6_outputs(5293) <= a;
    layer6_outputs(5294) <= a;
    layer6_outputs(5295) <= b and not a;
    layer6_outputs(5296) <= a and not b;
    layer6_outputs(5297) <= not (a xor b);
    layer6_outputs(5298) <= a xor b;
    layer6_outputs(5299) <= not b;
    layer6_outputs(5300) <= not a or b;
    layer6_outputs(5301) <= b;
    layer6_outputs(5302) <= b;
    layer6_outputs(5303) <= not b;
    layer6_outputs(5304) <= '1';
    layer6_outputs(5305) <= not b;
    layer6_outputs(5306) <= b;
    layer6_outputs(5307) <= not (a xor b);
    layer6_outputs(5308) <= not a;
    layer6_outputs(5309) <= b;
    layer6_outputs(5310) <= b;
    layer6_outputs(5311) <= a and b;
    layer6_outputs(5312) <= not a;
    layer6_outputs(5313) <= b and not a;
    layer6_outputs(5314) <= a;
    layer6_outputs(5315) <= '0';
    layer6_outputs(5316) <= a xor b;
    layer6_outputs(5317) <= b;
    layer6_outputs(5318) <= a;
    layer6_outputs(5319) <= a and b;
    layer6_outputs(5320) <= not (a or b);
    layer6_outputs(5321) <= not b;
    layer6_outputs(5322) <= a and b;
    layer6_outputs(5323) <= not a or b;
    layer6_outputs(5324) <= a xor b;
    layer6_outputs(5325) <= '0';
    layer6_outputs(5326) <= a;
    layer6_outputs(5327) <= not b;
    layer6_outputs(5328) <= not b;
    layer6_outputs(5329) <= b;
    layer6_outputs(5330) <= not (a xor b);
    layer6_outputs(5331) <= b;
    layer6_outputs(5332) <= b;
    layer6_outputs(5333) <= not b;
    layer6_outputs(5334) <= a;
    layer6_outputs(5335) <= b;
    layer6_outputs(5336) <= a and not b;
    layer6_outputs(5337) <= b and not a;
    layer6_outputs(5338) <= not (a or b);
    layer6_outputs(5339) <= not (a xor b);
    layer6_outputs(5340) <= not b;
    layer6_outputs(5341) <= not b;
    layer6_outputs(5342) <= not b;
    layer6_outputs(5343) <= a;
    layer6_outputs(5344) <= a and b;
    layer6_outputs(5345) <= b and not a;
    layer6_outputs(5346) <= not a;
    layer6_outputs(5347) <= not a;
    layer6_outputs(5348) <= a and b;
    layer6_outputs(5349) <= a or b;
    layer6_outputs(5350) <= not a;
    layer6_outputs(5351) <= not a or b;
    layer6_outputs(5352) <= b and not a;
    layer6_outputs(5353) <= b and not a;
    layer6_outputs(5354) <= a;
    layer6_outputs(5355) <= a;
    layer6_outputs(5356) <= a and not b;
    layer6_outputs(5357) <= not (a or b);
    layer6_outputs(5358) <= not b;
    layer6_outputs(5359) <= not (a or b);
    layer6_outputs(5360) <= not b;
    layer6_outputs(5361) <= not a;
    layer6_outputs(5362) <= not (a xor b);
    layer6_outputs(5363) <= a;
    layer6_outputs(5364) <= not b or a;
    layer6_outputs(5365) <= b;
    layer6_outputs(5366) <= b and not a;
    layer6_outputs(5367) <= a;
    layer6_outputs(5368) <= not b;
    layer6_outputs(5369) <= not (a xor b);
    layer6_outputs(5370) <= b;
    layer6_outputs(5371) <= not b;
    layer6_outputs(5372) <= not (a xor b);
    layer6_outputs(5373) <= a and not b;
    layer6_outputs(5374) <= not (a or b);
    layer6_outputs(5375) <= b;
    layer6_outputs(5376) <= not b;
    layer6_outputs(5377) <= not (a and b);
    layer6_outputs(5378) <= a xor b;
    layer6_outputs(5379) <= not a or b;
    layer6_outputs(5380) <= not b or a;
    layer6_outputs(5381) <= not b;
    layer6_outputs(5382) <= a and not b;
    layer6_outputs(5383) <= b;
    layer6_outputs(5384) <= a;
    layer6_outputs(5385) <= a and b;
    layer6_outputs(5386) <= not b;
    layer6_outputs(5387) <= a xor b;
    layer6_outputs(5388) <= not a;
    layer6_outputs(5389) <= not b;
    layer6_outputs(5390) <= a or b;
    layer6_outputs(5391) <= not b or a;
    layer6_outputs(5392) <= a and b;
    layer6_outputs(5393) <= not b;
    layer6_outputs(5394) <= a and not b;
    layer6_outputs(5395) <= not a or b;
    layer6_outputs(5396) <= a xor b;
    layer6_outputs(5397) <= not (a xor b);
    layer6_outputs(5398) <= a and b;
    layer6_outputs(5399) <= not (a xor b);
    layer6_outputs(5400) <= b;
    layer6_outputs(5401) <= b;
    layer6_outputs(5402) <= not (a xor b);
    layer6_outputs(5403) <= not a;
    layer6_outputs(5404) <= b;
    layer6_outputs(5405) <= not b;
    layer6_outputs(5406) <= a xor b;
    layer6_outputs(5407) <= not b;
    layer6_outputs(5408) <= not (a and b);
    layer6_outputs(5409) <= not (a and b);
    layer6_outputs(5410) <= a xor b;
    layer6_outputs(5411) <= a;
    layer6_outputs(5412) <= a xor b;
    layer6_outputs(5413) <= not (a xor b);
    layer6_outputs(5414) <= a xor b;
    layer6_outputs(5415) <= not (a or b);
    layer6_outputs(5416) <= a and not b;
    layer6_outputs(5417) <= not (a and b);
    layer6_outputs(5418) <= a;
    layer6_outputs(5419) <= a and not b;
    layer6_outputs(5420) <= a;
    layer6_outputs(5421) <= not b;
    layer6_outputs(5422) <= not b;
    layer6_outputs(5423) <= not b;
    layer6_outputs(5424) <= not (a xor b);
    layer6_outputs(5425) <= not b;
    layer6_outputs(5426) <= a and b;
    layer6_outputs(5427) <= a and not b;
    layer6_outputs(5428) <= not (a xor b);
    layer6_outputs(5429) <= not (a or b);
    layer6_outputs(5430) <= not (a xor b);
    layer6_outputs(5431) <= not a;
    layer6_outputs(5432) <= not a;
    layer6_outputs(5433) <= not (a or b);
    layer6_outputs(5434) <= a xor b;
    layer6_outputs(5435) <= a and b;
    layer6_outputs(5436) <= a;
    layer6_outputs(5437) <= not a;
    layer6_outputs(5438) <= b;
    layer6_outputs(5439) <= not (a or b);
    layer6_outputs(5440) <= a and not b;
    layer6_outputs(5441) <= not a;
    layer6_outputs(5442) <= not a or b;
    layer6_outputs(5443) <= not b;
    layer6_outputs(5444) <= not b;
    layer6_outputs(5445) <= not b;
    layer6_outputs(5446) <= not b or a;
    layer6_outputs(5447) <= not a;
    layer6_outputs(5448) <= b;
    layer6_outputs(5449) <= not b;
    layer6_outputs(5450) <= not a or b;
    layer6_outputs(5451) <= a and b;
    layer6_outputs(5452) <= b;
    layer6_outputs(5453) <= not (a xor b);
    layer6_outputs(5454) <= a or b;
    layer6_outputs(5455) <= not (a xor b);
    layer6_outputs(5456) <= a;
    layer6_outputs(5457) <= not (a xor b);
    layer6_outputs(5458) <= not b;
    layer6_outputs(5459) <= not b or a;
    layer6_outputs(5460) <= not (a or b);
    layer6_outputs(5461) <= b and not a;
    layer6_outputs(5462) <= a;
    layer6_outputs(5463) <= a;
    layer6_outputs(5464) <= not b or a;
    layer6_outputs(5465) <= b;
    layer6_outputs(5466) <= not (a and b);
    layer6_outputs(5467) <= b and not a;
    layer6_outputs(5468) <= a and b;
    layer6_outputs(5469) <= a or b;
    layer6_outputs(5470) <= a;
    layer6_outputs(5471) <= not (a and b);
    layer6_outputs(5472) <= not (a xor b);
    layer6_outputs(5473) <= a and b;
    layer6_outputs(5474) <= not (a xor b);
    layer6_outputs(5475) <= not a;
    layer6_outputs(5476) <= a or b;
    layer6_outputs(5477) <= not a or b;
    layer6_outputs(5478) <= not a;
    layer6_outputs(5479) <= not a;
    layer6_outputs(5480) <= not b;
    layer6_outputs(5481) <= not b or a;
    layer6_outputs(5482) <= not (a xor b);
    layer6_outputs(5483) <= not a;
    layer6_outputs(5484) <= a or b;
    layer6_outputs(5485) <= not a;
    layer6_outputs(5486) <= a and b;
    layer6_outputs(5487) <= not b or a;
    layer6_outputs(5488) <= b;
    layer6_outputs(5489) <= b and not a;
    layer6_outputs(5490) <= a or b;
    layer6_outputs(5491) <= a;
    layer6_outputs(5492) <= not (a xor b);
    layer6_outputs(5493) <= b and not a;
    layer6_outputs(5494) <= b;
    layer6_outputs(5495) <= a and b;
    layer6_outputs(5496) <= a xor b;
    layer6_outputs(5497) <= not a;
    layer6_outputs(5498) <= not b;
    layer6_outputs(5499) <= a xor b;
    layer6_outputs(5500) <= not (a and b);
    layer6_outputs(5501) <= b;
    layer6_outputs(5502) <= not a;
    layer6_outputs(5503) <= b;
    layer6_outputs(5504) <= not a;
    layer6_outputs(5505) <= a;
    layer6_outputs(5506) <= b;
    layer6_outputs(5507) <= b and not a;
    layer6_outputs(5508) <= b;
    layer6_outputs(5509) <= a and not b;
    layer6_outputs(5510) <= a;
    layer6_outputs(5511) <= b;
    layer6_outputs(5512) <= not a;
    layer6_outputs(5513) <= a xor b;
    layer6_outputs(5514) <= not a or b;
    layer6_outputs(5515) <= not a;
    layer6_outputs(5516) <= not (a and b);
    layer6_outputs(5517) <= not a;
    layer6_outputs(5518) <= a;
    layer6_outputs(5519) <= not a;
    layer6_outputs(5520) <= not a;
    layer6_outputs(5521) <= not (a xor b);
    layer6_outputs(5522) <= b;
    layer6_outputs(5523) <= a and not b;
    layer6_outputs(5524) <= not b;
    layer6_outputs(5525) <= a and b;
    layer6_outputs(5526) <= not b;
    layer6_outputs(5527) <= not (a xor b);
    layer6_outputs(5528) <= a;
    layer6_outputs(5529) <= a;
    layer6_outputs(5530) <= not (a xor b);
    layer6_outputs(5531) <= not (a xor b);
    layer6_outputs(5532) <= not b;
    layer6_outputs(5533) <= not b;
    layer6_outputs(5534) <= not b;
    layer6_outputs(5535) <= not (a or b);
    layer6_outputs(5536) <= not b;
    layer6_outputs(5537) <= not (a xor b);
    layer6_outputs(5538) <= a xor b;
    layer6_outputs(5539) <= not a;
    layer6_outputs(5540) <= not b;
    layer6_outputs(5541) <= a;
    layer6_outputs(5542) <= a or b;
    layer6_outputs(5543) <= a and not b;
    layer6_outputs(5544) <= a;
    layer6_outputs(5545) <= not (a xor b);
    layer6_outputs(5546) <= not (a xor b);
    layer6_outputs(5547) <= not a;
    layer6_outputs(5548) <= not a;
    layer6_outputs(5549) <= not b;
    layer6_outputs(5550) <= not (a xor b);
    layer6_outputs(5551) <= a xor b;
    layer6_outputs(5552) <= not (a xor b);
    layer6_outputs(5553) <= not (a and b);
    layer6_outputs(5554) <= not (a and b);
    layer6_outputs(5555) <= a and b;
    layer6_outputs(5556) <= a;
    layer6_outputs(5557) <= not a;
    layer6_outputs(5558) <= not a;
    layer6_outputs(5559) <= not b or a;
    layer6_outputs(5560) <= b;
    layer6_outputs(5561) <= a xor b;
    layer6_outputs(5562) <= not (a xor b);
    layer6_outputs(5563) <= not a or b;
    layer6_outputs(5564) <= not a;
    layer6_outputs(5565) <= a and b;
    layer6_outputs(5566) <= a;
    layer6_outputs(5567) <= a;
    layer6_outputs(5568) <= not b;
    layer6_outputs(5569) <= a xor b;
    layer6_outputs(5570) <= not a;
    layer6_outputs(5571) <= not b or a;
    layer6_outputs(5572) <= a and b;
    layer6_outputs(5573) <= not a;
    layer6_outputs(5574) <= a;
    layer6_outputs(5575) <= a and b;
    layer6_outputs(5576) <= not b;
    layer6_outputs(5577) <= a and not b;
    layer6_outputs(5578) <= a;
    layer6_outputs(5579) <= b;
    layer6_outputs(5580) <= a;
    layer6_outputs(5581) <= not b or a;
    layer6_outputs(5582) <= a xor b;
    layer6_outputs(5583) <= not (a or b);
    layer6_outputs(5584) <= a or b;
    layer6_outputs(5585) <= not a;
    layer6_outputs(5586) <= not a;
    layer6_outputs(5587) <= b and not a;
    layer6_outputs(5588) <= not a;
    layer6_outputs(5589) <= a and not b;
    layer6_outputs(5590) <= a;
    layer6_outputs(5591) <= not a;
    layer6_outputs(5592) <= not b;
    layer6_outputs(5593) <= not a or b;
    layer6_outputs(5594) <= a xor b;
    layer6_outputs(5595) <= not b;
    layer6_outputs(5596) <= not (a xor b);
    layer6_outputs(5597) <= not b or a;
    layer6_outputs(5598) <= a and b;
    layer6_outputs(5599) <= not a;
    layer6_outputs(5600) <= b and not a;
    layer6_outputs(5601) <= not (a and b);
    layer6_outputs(5602) <= '0';
    layer6_outputs(5603) <= a;
    layer6_outputs(5604) <= not a or b;
    layer6_outputs(5605) <= a xor b;
    layer6_outputs(5606) <= a and not b;
    layer6_outputs(5607) <= b and not a;
    layer6_outputs(5608) <= b and not a;
    layer6_outputs(5609) <= a;
    layer6_outputs(5610) <= not (a xor b);
    layer6_outputs(5611) <= a and not b;
    layer6_outputs(5612) <= a xor b;
    layer6_outputs(5613) <= not (a xor b);
    layer6_outputs(5614) <= b;
    layer6_outputs(5615) <= b;
    layer6_outputs(5616) <= '1';
    layer6_outputs(5617) <= not b or a;
    layer6_outputs(5618) <= not b;
    layer6_outputs(5619) <= a and b;
    layer6_outputs(5620) <= not a or b;
    layer6_outputs(5621) <= a and b;
    layer6_outputs(5622) <= b;
    layer6_outputs(5623) <= a;
    layer6_outputs(5624) <= not a or b;
    layer6_outputs(5625) <= not (a xor b);
    layer6_outputs(5626) <= a xor b;
    layer6_outputs(5627) <= not a;
    layer6_outputs(5628) <= not b or a;
    layer6_outputs(5629) <= b and not a;
    layer6_outputs(5630) <= not (a xor b);
    layer6_outputs(5631) <= not (a or b);
    layer6_outputs(5632) <= not b;
    layer6_outputs(5633) <= a xor b;
    layer6_outputs(5634) <= not b or a;
    layer6_outputs(5635) <= not (a or b);
    layer6_outputs(5636) <= not b or a;
    layer6_outputs(5637) <= not b;
    layer6_outputs(5638) <= not (a xor b);
    layer6_outputs(5639) <= a;
    layer6_outputs(5640) <= not a;
    layer6_outputs(5641) <= not a;
    layer6_outputs(5642) <= a and not b;
    layer6_outputs(5643) <= not a or b;
    layer6_outputs(5644) <= not (a xor b);
    layer6_outputs(5645) <= a;
    layer6_outputs(5646) <= not a;
    layer6_outputs(5647) <= '0';
    layer6_outputs(5648) <= a;
    layer6_outputs(5649) <= not a;
    layer6_outputs(5650) <= a and not b;
    layer6_outputs(5651) <= a xor b;
    layer6_outputs(5652) <= not a or b;
    layer6_outputs(5653) <= not a;
    layer6_outputs(5654) <= not b or a;
    layer6_outputs(5655) <= not (a xor b);
    layer6_outputs(5656) <= a and b;
    layer6_outputs(5657) <= a and b;
    layer6_outputs(5658) <= b and not a;
    layer6_outputs(5659) <= b;
    layer6_outputs(5660) <= not (a and b);
    layer6_outputs(5661) <= a;
    layer6_outputs(5662) <= not b or a;
    layer6_outputs(5663) <= not a;
    layer6_outputs(5664) <= not a;
    layer6_outputs(5665) <= not (a xor b);
    layer6_outputs(5666) <= not b;
    layer6_outputs(5667) <= not (a or b);
    layer6_outputs(5668) <= not b;
    layer6_outputs(5669) <= not b or a;
    layer6_outputs(5670) <= not (a xor b);
    layer6_outputs(5671) <= b;
    layer6_outputs(5672) <= not a;
    layer6_outputs(5673) <= not (a xor b);
    layer6_outputs(5674) <= not a;
    layer6_outputs(5675) <= not (a xor b);
    layer6_outputs(5676) <= not (a and b);
    layer6_outputs(5677) <= not b;
    layer6_outputs(5678) <= a;
    layer6_outputs(5679) <= a;
    layer6_outputs(5680) <= a;
    layer6_outputs(5681) <= not b;
    layer6_outputs(5682) <= not a;
    layer6_outputs(5683) <= b;
    layer6_outputs(5684) <= not a or b;
    layer6_outputs(5685) <= b;
    layer6_outputs(5686) <= not b or a;
    layer6_outputs(5687) <= b;
    layer6_outputs(5688) <= b and not a;
    layer6_outputs(5689) <= b;
    layer6_outputs(5690) <= not a or b;
    layer6_outputs(5691) <= not b;
    layer6_outputs(5692) <= a;
    layer6_outputs(5693) <= b;
    layer6_outputs(5694) <= a;
    layer6_outputs(5695) <= a xor b;
    layer6_outputs(5696) <= not (a or b);
    layer6_outputs(5697) <= not b;
    layer6_outputs(5698) <= not (a xor b);
    layer6_outputs(5699) <= not a;
    layer6_outputs(5700) <= b and not a;
    layer6_outputs(5701) <= not b;
    layer6_outputs(5702) <= not (a or b);
    layer6_outputs(5703) <= not (a xor b);
    layer6_outputs(5704) <= b;
    layer6_outputs(5705) <= not (a and b);
    layer6_outputs(5706) <= b;
    layer6_outputs(5707) <= not a;
    layer6_outputs(5708) <= not (a or b);
    layer6_outputs(5709) <= not a;
    layer6_outputs(5710) <= not (a xor b);
    layer6_outputs(5711) <= b and not a;
    layer6_outputs(5712) <= not (a xor b);
    layer6_outputs(5713) <= not b;
    layer6_outputs(5714) <= not (a or b);
    layer6_outputs(5715) <= not (a xor b);
    layer6_outputs(5716) <= a and not b;
    layer6_outputs(5717) <= not b or a;
    layer6_outputs(5718) <= a;
    layer6_outputs(5719) <= not a;
    layer6_outputs(5720) <= a xor b;
    layer6_outputs(5721) <= not a;
    layer6_outputs(5722) <= not b or a;
    layer6_outputs(5723) <= not b;
    layer6_outputs(5724) <= b and not a;
    layer6_outputs(5725) <= b;
    layer6_outputs(5726) <= a and b;
    layer6_outputs(5727) <= not a;
    layer6_outputs(5728) <= a and b;
    layer6_outputs(5729) <= a;
    layer6_outputs(5730) <= a xor b;
    layer6_outputs(5731) <= a xor b;
    layer6_outputs(5732) <= b;
    layer6_outputs(5733) <= not (a or b);
    layer6_outputs(5734) <= not b or a;
    layer6_outputs(5735) <= a;
    layer6_outputs(5736) <= not (a and b);
    layer6_outputs(5737) <= not (a xor b);
    layer6_outputs(5738) <= a and b;
    layer6_outputs(5739) <= b;
    layer6_outputs(5740) <= b;
    layer6_outputs(5741) <= not b or a;
    layer6_outputs(5742) <= a or b;
    layer6_outputs(5743) <= not a or b;
    layer6_outputs(5744) <= a or b;
    layer6_outputs(5745) <= a;
    layer6_outputs(5746) <= not b;
    layer6_outputs(5747) <= not a or b;
    layer6_outputs(5748) <= not a;
    layer6_outputs(5749) <= b;
    layer6_outputs(5750) <= not b;
    layer6_outputs(5751) <= not (a or b);
    layer6_outputs(5752) <= b and not a;
    layer6_outputs(5753) <= a xor b;
    layer6_outputs(5754) <= not a;
    layer6_outputs(5755) <= not (a xor b);
    layer6_outputs(5756) <= b and not a;
    layer6_outputs(5757) <= not b;
    layer6_outputs(5758) <= b;
    layer6_outputs(5759) <= not (a xor b);
    layer6_outputs(5760) <= a;
    layer6_outputs(5761) <= a or b;
    layer6_outputs(5762) <= not b or a;
    layer6_outputs(5763) <= a;
    layer6_outputs(5764) <= a;
    layer6_outputs(5765) <= b;
    layer6_outputs(5766) <= not (a xor b);
    layer6_outputs(5767) <= not (a and b);
    layer6_outputs(5768) <= b;
    layer6_outputs(5769) <= b and not a;
    layer6_outputs(5770) <= b;
    layer6_outputs(5771) <= not (a or b);
    layer6_outputs(5772) <= a;
    layer6_outputs(5773) <= not a or b;
    layer6_outputs(5774) <= not b;
    layer6_outputs(5775) <= not a;
    layer6_outputs(5776) <= not (a or b);
    layer6_outputs(5777) <= not a or b;
    layer6_outputs(5778) <= not a or b;
    layer6_outputs(5779) <= not (a and b);
    layer6_outputs(5780) <= not (a and b);
    layer6_outputs(5781) <= b and not a;
    layer6_outputs(5782) <= b;
    layer6_outputs(5783) <= not (a xor b);
    layer6_outputs(5784) <= b and not a;
    layer6_outputs(5785) <= a;
    layer6_outputs(5786) <= not a;
    layer6_outputs(5787) <= a xor b;
    layer6_outputs(5788) <= not (a xor b);
    layer6_outputs(5789) <= a or b;
    layer6_outputs(5790) <= a;
    layer6_outputs(5791) <= a and b;
    layer6_outputs(5792) <= not a;
    layer6_outputs(5793) <= not a or b;
    layer6_outputs(5794) <= not (a xor b);
    layer6_outputs(5795) <= a xor b;
    layer6_outputs(5796) <= not a or b;
    layer6_outputs(5797) <= a and not b;
    layer6_outputs(5798) <= not (a xor b);
    layer6_outputs(5799) <= not a;
    layer6_outputs(5800) <= not a;
    layer6_outputs(5801) <= a;
    layer6_outputs(5802) <= not (a or b);
    layer6_outputs(5803) <= a xor b;
    layer6_outputs(5804) <= a;
    layer6_outputs(5805) <= a and b;
    layer6_outputs(5806) <= not a;
    layer6_outputs(5807) <= not (a or b);
    layer6_outputs(5808) <= not a;
    layer6_outputs(5809) <= not a;
    layer6_outputs(5810) <= not a;
    layer6_outputs(5811) <= not (a or b);
    layer6_outputs(5812) <= not a;
    layer6_outputs(5813) <= not (a or b);
    layer6_outputs(5814) <= not a;
    layer6_outputs(5815) <= not b;
    layer6_outputs(5816) <= not (a and b);
    layer6_outputs(5817) <= '0';
    layer6_outputs(5818) <= not b;
    layer6_outputs(5819) <= not a;
    layer6_outputs(5820) <= a and b;
    layer6_outputs(5821) <= b and not a;
    layer6_outputs(5822) <= not (a xor b);
    layer6_outputs(5823) <= a and not b;
    layer6_outputs(5824) <= b;
    layer6_outputs(5825) <= a;
    layer6_outputs(5826) <= a and not b;
    layer6_outputs(5827) <= b;
    layer6_outputs(5828) <= b;
    layer6_outputs(5829) <= a xor b;
    layer6_outputs(5830) <= '1';
    layer6_outputs(5831) <= a and not b;
    layer6_outputs(5832) <= not a;
    layer6_outputs(5833) <= not a;
    layer6_outputs(5834) <= not a or b;
    layer6_outputs(5835) <= b;
    layer6_outputs(5836) <= not b;
    layer6_outputs(5837) <= b;
    layer6_outputs(5838) <= a;
    layer6_outputs(5839) <= not a;
    layer6_outputs(5840) <= a;
    layer6_outputs(5841) <= b;
    layer6_outputs(5842) <= a or b;
    layer6_outputs(5843) <= not b or a;
    layer6_outputs(5844) <= not (a xor b);
    layer6_outputs(5845) <= a and not b;
    layer6_outputs(5846) <= b;
    layer6_outputs(5847) <= a xor b;
    layer6_outputs(5848) <= not a or b;
    layer6_outputs(5849) <= a xor b;
    layer6_outputs(5850) <= not a;
    layer6_outputs(5851) <= b;
    layer6_outputs(5852) <= not a;
    layer6_outputs(5853) <= not b;
    layer6_outputs(5854) <= a and b;
    layer6_outputs(5855) <= b;
    layer6_outputs(5856) <= not b;
    layer6_outputs(5857) <= b;
    layer6_outputs(5858) <= b;
    layer6_outputs(5859) <= not (a and b);
    layer6_outputs(5860) <= not a;
    layer6_outputs(5861) <= not (a xor b);
    layer6_outputs(5862) <= not (a and b);
    layer6_outputs(5863) <= a or b;
    layer6_outputs(5864) <= b;
    layer6_outputs(5865) <= a xor b;
    layer6_outputs(5866) <= a xor b;
    layer6_outputs(5867) <= not (a and b);
    layer6_outputs(5868) <= not (a xor b);
    layer6_outputs(5869) <= not a;
    layer6_outputs(5870) <= not b;
    layer6_outputs(5871) <= b;
    layer6_outputs(5872) <= a;
    layer6_outputs(5873) <= a;
    layer6_outputs(5874) <= not a;
    layer6_outputs(5875) <= a xor b;
    layer6_outputs(5876) <= not (a xor b);
    layer6_outputs(5877) <= not (a and b);
    layer6_outputs(5878) <= b;
    layer6_outputs(5879) <= not b;
    layer6_outputs(5880) <= not b;
    layer6_outputs(5881) <= a xor b;
    layer6_outputs(5882) <= not b;
    layer6_outputs(5883) <= not (a and b);
    layer6_outputs(5884) <= b;
    layer6_outputs(5885) <= not b;
    layer6_outputs(5886) <= not (a xor b);
    layer6_outputs(5887) <= '1';
    layer6_outputs(5888) <= not a;
    layer6_outputs(5889) <= b;
    layer6_outputs(5890) <= a xor b;
    layer6_outputs(5891) <= not a;
    layer6_outputs(5892) <= not a or b;
    layer6_outputs(5893) <= b;
    layer6_outputs(5894) <= not b;
    layer6_outputs(5895) <= not a;
    layer6_outputs(5896) <= b;
    layer6_outputs(5897) <= not (a xor b);
    layer6_outputs(5898) <= b and not a;
    layer6_outputs(5899) <= not (a and b);
    layer6_outputs(5900) <= not a;
    layer6_outputs(5901) <= not (a or b);
    layer6_outputs(5902) <= b and not a;
    layer6_outputs(5903) <= b;
    layer6_outputs(5904) <= not b;
    layer6_outputs(5905) <= not b or a;
    layer6_outputs(5906) <= '0';
    layer6_outputs(5907) <= a and b;
    layer6_outputs(5908) <= not (a xor b);
    layer6_outputs(5909) <= not (a and b);
    layer6_outputs(5910) <= not (a or b);
    layer6_outputs(5911) <= not b;
    layer6_outputs(5912) <= not b or a;
    layer6_outputs(5913) <= not (a xor b);
    layer6_outputs(5914) <= not b or a;
    layer6_outputs(5915) <= b;
    layer6_outputs(5916) <= a and b;
    layer6_outputs(5917) <= b;
    layer6_outputs(5918) <= not b;
    layer6_outputs(5919) <= not a;
    layer6_outputs(5920) <= not a;
    layer6_outputs(5921) <= a xor b;
    layer6_outputs(5922) <= not a;
    layer6_outputs(5923) <= '1';
    layer6_outputs(5924) <= not a;
    layer6_outputs(5925) <= not (a or b);
    layer6_outputs(5926) <= a and not b;
    layer6_outputs(5927) <= not (a and b);
    layer6_outputs(5928) <= not (a xor b);
    layer6_outputs(5929) <= not a;
    layer6_outputs(5930) <= not (a xor b);
    layer6_outputs(5931) <= a;
    layer6_outputs(5932) <= not b;
    layer6_outputs(5933) <= a xor b;
    layer6_outputs(5934) <= not (a and b);
    layer6_outputs(5935) <= a and not b;
    layer6_outputs(5936) <= a xor b;
    layer6_outputs(5937) <= not b;
    layer6_outputs(5938) <= not a;
    layer6_outputs(5939) <= a and b;
    layer6_outputs(5940) <= not (a or b);
    layer6_outputs(5941) <= not a;
    layer6_outputs(5942) <= a or b;
    layer6_outputs(5943) <= not a;
    layer6_outputs(5944) <= b;
    layer6_outputs(5945) <= b and not a;
    layer6_outputs(5946) <= a;
    layer6_outputs(5947) <= a or b;
    layer6_outputs(5948) <= a xor b;
    layer6_outputs(5949) <= not b or a;
    layer6_outputs(5950) <= a and not b;
    layer6_outputs(5951) <= '1';
    layer6_outputs(5952) <= b;
    layer6_outputs(5953) <= not (a or b);
    layer6_outputs(5954) <= b and not a;
    layer6_outputs(5955) <= not a or b;
    layer6_outputs(5956) <= not b;
    layer6_outputs(5957) <= not a;
    layer6_outputs(5958) <= not (a xor b);
    layer6_outputs(5959) <= a and not b;
    layer6_outputs(5960) <= not a or b;
    layer6_outputs(5961) <= '0';
    layer6_outputs(5962) <= not (a xor b);
    layer6_outputs(5963) <= not a;
    layer6_outputs(5964) <= a and not b;
    layer6_outputs(5965) <= not (a or b);
    layer6_outputs(5966) <= not a;
    layer6_outputs(5967) <= not a or b;
    layer6_outputs(5968) <= a and b;
    layer6_outputs(5969) <= not b;
    layer6_outputs(5970) <= a;
    layer6_outputs(5971) <= not (a xor b);
    layer6_outputs(5972) <= b;
    layer6_outputs(5973) <= not b;
    layer6_outputs(5974) <= not a;
    layer6_outputs(5975) <= not (a or b);
    layer6_outputs(5976) <= not b or a;
    layer6_outputs(5977) <= a and b;
    layer6_outputs(5978) <= not b;
    layer6_outputs(5979) <= b;
    layer6_outputs(5980) <= not a;
    layer6_outputs(5981) <= a xor b;
    layer6_outputs(5982) <= not (a xor b);
    layer6_outputs(5983) <= not (a or b);
    layer6_outputs(5984) <= not (a or b);
    layer6_outputs(5985) <= a xor b;
    layer6_outputs(5986) <= b;
    layer6_outputs(5987) <= not a or b;
    layer6_outputs(5988) <= '1';
    layer6_outputs(5989) <= a;
    layer6_outputs(5990) <= a and b;
    layer6_outputs(5991) <= a;
    layer6_outputs(5992) <= a xor b;
    layer6_outputs(5993) <= a or b;
    layer6_outputs(5994) <= not b;
    layer6_outputs(5995) <= a and b;
    layer6_outputs(5996) <= a or b;
    layer6_outputs(5997) <= b;
    layer6_outputs(5998) <= not a;
    layer6_outputs(5999) <= not a;
    layer6_outputs(6000) <= a xor b;
    layer6_outputs(6001) <= a or b;
    layer6_outputs(6002) <= a;
    layer6_outputs(6003) <= not (a and b);
    layer6_outputs(6004) <= a xor b;
    layer6_outputs(6005) <= not a or b;
    layer6_outputs(6006) <= b;
    layer6_outputs(6007) <= not a;
    layer6_outputs(6008) <= b;
    layer6_outputs(6009) <= not b or a;
    layer6_outputs(6010) <= a;
    layer6_outputs(6011) <= not (a and b);
    layer6_outputs(6012) <= not a;
    layer6_outputs(6013) <= a or b;
    layer6_outputs(6014) <= not a;
    layer6_outputs(6015) <= b and not a;
    layer6_outputs(6016) <= b;
    layer6_outputs(6017) <= a;
    layer6_outputs(6018) <= b;
    layer6_outputs(6019) <= not b;
    layer6_outputs(6020) <= not a;
    layer6_outputs(6021) <= a or b;
    layer6_outputs(6022) <= not (a and b);
    layer6_outputs(6023) <= b;
    layer6_outputs(6024) <= a or b;
    layer6_outputs(6025) <= not (a or b);
    layer6_outputs(6026) <= not (a and b);
    layer6_outputs(6027) <= not a;
    layer6_outputs(6028) <= b;
    layer6_outputs(6029) <= b;
    layer6_outputs(6030) <= not (a or b);
    layer6_outputs(6031) <= b;
    layer6_outputs(6032) <= b;
    layer6_outputs(6033) <= a and not b;
    layer6_outputs(6034) <= not b or a;
    layer6_outputs(6035) <= not b;
    layer6_outputs(6036) <= b;
    layer6_outputs(6037) <= not b or a;
    layer6_outputs(6038) <= not (a or b);
    layer6_outputs(6039) <= b and not a;
    layer6_outputs(6040) <= not (a xor b);
    layer6_outputs(6041) <= a or b;
    layer6_outputs(6042) <= not a or b;
    layer6_outputs(6043) <= a xor b;
    layer6_outputs(6044) <= a xor b;
    layer6_outputs(6045) <= b;
    layer6_outputs(6046) <= not b or a;
    layer6_outputs(6047) <= not (a xor b);
    layer6_outputs(6048) <= a xor b;
    layer6_outputs(6049) <= b and not a;
    layer6_outputs(6050) <= a or b;
    layer6_outputs(6051) <= a and not b;
    layer6_outputs(6052) <= not (a xor b);
    layer6_outputs(6053) <= not a or b;
    layer6_outputs(6054) <= not a;
    layer6_outputs(6055) <= b;
    layer6_outputs(6056) <= not (a or b);
    layer6_outputs(6057) <= a;
    layer6_outputs(6058) <= a xor b;
    layer6_outputs(6059) <= a and b;
    layer6_outputs(6060) <= not a;
    layer6_outputs(6061) <= not (a or b);
    layer6_outputs(6062) <= not (a or b);
    layer6_outputs(6063) <= not a;
    layer6_outputs(6064) <= b;
    layer6_outputs(6065) <= a and b;
    layer6_outputs(6066) <= b and not a;
    layer6_outputs(6067) <= not (a or b);
    layer6_outputs(6068) <= not a;
    layer6_outputs(6069) <= b and not a;
    layer6_outputs(6070) <= a;
    layer6_outputs(6071) <= not (a and b);
    layer6_outputs(6072) <= a and b;
    layer6_outputs(6073) <= a xor b;
    layer6_outputs(6074) <= b and not a;
    layer6_outputs(6075) <= not (a xor b);
    layer6_outputs(6076) <= not (a and b);
    layer6_outputs(6077) <= not (a or b);
    layer6_outputs(6078) <= not b;
    layer6_outputs(6079) <= a xor b;
    layer6_outputs(6080) <= not (a xor b);
    layer6_outputs(6081) <= not (a xor b);
    layer6_outputs(6082) <= a xor b;
    layer6_outputs(6083) <= not a;
    layer6_outputs(6084) <= a and b;
    layer6_outputs(6085) <= not b;
    layer6_outputs(6086) <= a;
    layer6_outputs(6087) <= not (a xor b);
    layer6_outputs(6088) <= not b;
    layer6_outputs(6089) <= a xor b;
    layer6_outputs(6090) <= b and not a;
    layer6_outputs(6091) <= not (a or b);
    layer6_outputs(6092) <= a;
    layer6_outputs(6093) <= b;
    layer6_outputs(6094) <= not a;
    layer6_outputs(6095) <= not a;
    layer6_outputs(6096) <= a and b;
    layer6_outputs(6097) <= b;
    layer6_outputs(6098) <= not a;
    layer6_outputs(6099) <= b and not a;
    layer6_outputs(6100) <= not a;
    layer6_outputs(6101) <= a;
    layer6_outputs(6102) <= b and not a;
    layer6_outputs(6103) <= a;
    layer6_outputs(6104) <= a xor b;
    layer6_outputs(6105) <= not b or a;
    layer6_outputs(6106) <= not b or a;
    layer6_outputs(6107) <= b and not a;
    layer6_outputs(6108) <= not b;
    layer6_outputs(6109) <= not a;
    layer6_outputs(6110) <= a;
    layer6_outputs(6111) <= b and not a;
    layer6_outputs(6112) <= not b or a;
    layer6_outputs(6113) <= not (a xor b);
    layer6_outputs(6114) <= not b or a;
    layer6_outputs(6115) <= not b;
    layer6_outputs(6116) <= b;
    layer6_outputs(6117) <= not (a and b);
    layer6_outputs(6118) <= not (a and b);
    layer6_outputs(6119) <= a;
    layer6_outputs(6120) <= b;
    layer6_outputs(6121) <= not (a or b);
    layer6_outputs(6122) <= not b;
    layer6_outputs(6123) <= b and not a;
    layer6_outputs(6124) <= not a or b;
    layer6_outputs(6125) <= not (a xor b);
    layer6_outputs(6126) <= b;
    layer6_outputs(6127) <= not a or b;
    layer6_outputs(6128) <= b;
    layer6_outputs(6129) <= b and not a;
    layer6_outputs(6130) <= b;
    layer6_outputs(6131) <= b;
    layer6_outputs(6132) <= not a;
    layer6_outputs(6133) <= a;
    layer6_outputs(6134) <= a and not b;
    layer6_outputs(6135) <= b and not a;
    layer6_outputs(6136) <= not b;
    layer6_outputs(6137) <= not (a or b);
    layer6_outputs(6138) <= not (a and b);
    layer6_outputs(6139) <= not b;
    layer6_outputs(6140) <= a and b;
    layer6_outputs(6141) <= a xor b;
    layer6_outputs(6142) <= a;
    layer6_outputs(6143) <= a;
    layer6_outputs(6144) <= a or b;
    layer6_outputs(6145) <= not b;
    layer6_outputs(6146) <= a and not b;
    layer6_outputs(6147) <= a and b;
    layer6_outputs(6148) <= not b or a;
    layer6_outputs(6149) <= not (a or b);
    layer6_outputs(6150) <= not b;
    layer6_outputs(6151) <= a and not b;
    layer6_outputs(6152) <= b;
    layer6_outputs(6153) <= a;
    layer6_outputs(6154) <= a and not b;
    layer6_outputs(6155) <= a;
    layer6_outputs(6156) <= not a;
    layer6_outputs(6157) <= not (a xor b);
    layer6_outputs(6158) <= not b or a;
    layer6_outputs(6159) <= not b or a;
    layer6_outputs(6160) <= not (a xor b);
    layer6_outputs(6161) <= not a or b;
    layer6_outputs(6162) <= not a;
    layer6_outputs(6163) <= not (a or b);
    layer6_outputs(6164) <= not (a and b);
    layer6_outputs(6165) <= a;
    layer6_outputs(6166) <= not (a or b);
    layer6_outputs(6167) <= b;
    layer6_outputs(6168) <= a;
    layer6_outputs(6169) <= a and b;
    layer6_outputs(6170) <= a xor b;
    layer6_outputs(6171) <= b;
    layer6_outputs(6172) <= not a;
    layer6_outputs(6173) <= b;
    layer6_outputs(6174) <= not b;
    layer6_outputs(6175) <= b;
    layer6_outputs(6176) <= not b;
    layer6_outputs(6177) <= b and not a;
    layer6_outputs(6178) <= not (a xor b);
    layer6_outputs(6179) <= a xor b;
    layer6_outputs(6180) <= a or b;
    layer6_outputs(6181) <= a xor b;
    layer6_outputs(6182) <= not b or a;
    layer6_outputs(6183) <= not a or b;
    layer6_outputs(6184) <= not (a xor b);
    layer6_outputs(6185) <= a;
    layer6_outputs(6186) <= '1';
    layer6_outputs(6187) <= not a;
    layer6_outputs(6188) <= not a;
    layer6_outputs(6189) <= a;
    layer6_outputs(6190) <= not (a xor b);
    layer6_outputs(6191) <= not a;
    layer6_outputs(6192) <= not (a xor b);
    layer6_outputs(6193) <= b and not a;
    layer6_outputs(6194) <= b;
    layer6_outputs(6195) <= b and not a;
    layer6_outputs(6196) <= not b or a;
    layer6_outputs(6197) <= b and not a;
    layer6_outputs(6198) <= not (a xor b);
    layer6_outputs(6199) <= a and b;
    layer6_outputs(6200) <= not (a or b);
    layer6_outputs(6201) <= not a or b;
    layer6_outputs(6202) <= a and not b;
    layer6_outputs(6203) <= a;
    layer6_outputs(6204) <= not (a or b);
    layer6_outputs(6205) <= a or b;
    layer6_outputs(6206) <= not (a xor b);
    layer6_outputs(6207) <= a and not b;
    layer6_outputs(6208) <= a;
    layer6_outputs(6209) <= not b;
    layer6_outputs(6210) <= b;
    layer6_outputs(6211) <= a xor b;
    layer6_outputs(6212) <= not (a and b);
    layer6_outputs(6213) <= not b;
    layer6_outputs(6214) <= not b or a;
    layer6_outputs(6215) <= not a;
    layer6_outputs(6216) <= b;
    layer6_outputs(6217) <= b;
    layer6_outputs(6218) <= b;
    layer6_outputs(6219) <= not (a or b);
    layer6_outputs(6220) <= a xor b;
    layer6_outputs(6221) <= not (a and b);
    layer6_outputs(6222) <= a;
    layer6_outputs(6223) <= not (a or b);
    layer6_outputs(6224) <= not (a xor b);
    layer6_outputs(6225) <= a and not b;
    layer6_outputs(6226) <= b;
    layer6_outputs(6227) <= not (a xor b);
    layer6_outputs(6228) <= a or b;
    layer6_outputs(6229) <= not a;
    layer6_outputs(6230) <= not b;
    layer6_outputs(6231) <= not a;
    layer6_outputs(6232) <= a;
    layer6_outputs(6233) <= not (a xor b);
    layer6_outputs(6234) <= not b;
    layer6_outputs(6235) <= not b;
    layer6_outputs(6236) <= b and not a;
    layer6_outputs(6237) <= not b;
    layer6_outputs(6238) <= not b or a;
    layer6_outputs(6239) <= '0';
    layer6_outputs(6240) <= not b or a;
    layer6_outputs(6241) <= a and not b;
    layer6_outputs(6242) <= a and not b;
    layer6_outputs(6243) <= not b;
    layer6_outputs(6244) <= a and not b;
    layer6_outputs(6245) <= not a or b;
    layer6_outputs(6246) <= a;
    layer6_outputs(6247) <= not b or a;
    layer6_outputs(6248) <= a and not b;
    layer6_outputs(6249) <= a and b;
    layer6_outputs(6250) <= a or b;
    layer6_outputs(6251) <= not a;
    layer6_outputs(6252) <= not a or b;
    layer6_outputs(6253) <= not b;
    layer6_outputs(6254) <= a;
    layer6_outputs(6255) <= not a or b;
    layer6_outputs(6256) <= not b;
    layer6_outputs(6257) <= not a;
    layer6_outputs(6258) <= a xor b;
    layer6_outputs(6259) <= b and not a;
    layer6_outputs(6260) <= a xor b;
    layer6_outputs(6261) <= not b;
    layer6_outputs(6262) <= not b;
    layer6_outputs(6263) <= not a or b;
    layer6_outputs(6264) <= not (a and b);
    layer6_outputs(6265) <= a;
    layer6_outputs(6266) <= a;
    layer6_outputs(6267) <= not b or a;
    layer6_outputs(6268) <= a and b;
    layer6_outputs(6269) <= not b or a;
    layer6_outputs(6270) <= b;
    layer6_outputs(6271) <= '1';
    layer6_outputs(6272) <= a;
    layer6_outputs(6273) <= a;
    layer6_outputs(6274) <= a xor b;
    layer6_outputs(6275) <= a;
    layer6_outputs(6276) <= a xor b;
    layer6_outputs(6277) <= not a;
    layer6_outputs(6278) <= a;
    layer6_outputs(6279) <= not (a xor b);
    layer6_outputs(6280) <= b and not a;
    layer6_outputs(6281) <= not a;
    layer6_outputs(6282) <= not (a xor b);
    layer6_outputs(6283) <= a xor b;
    layer6_outputs(6284) <= a;
    layer6_outputs(6285) <= b;
    layer6_outputs(6286) <= a xor b;
    layer6_outputs(6287) <= not (a xor b);
    layer6_outputs(6288) <= not b;
    layer6_outputs(6289) <= a xor b;
    layer6_outputs(6290) <= a xor b;
    layer6_outputs(6291) <= a xor b;
    layer6_outputs(6292) <= not a or b;
    layer6_outputs(6293) <= a xor b;
    layer6_outputs(6294) <= not b;
    layer6_outputs(6295) <= not b;
    layer6_outputs(6296) <= a xor b;
    layer6_outputs(6297) <= a xor b;
    layer6_outputs(6298) <= not (a and b);
    layer6_outputs(6299) <= b and not a;
    layer6_outputs(6300) <= not a;
    layer6_outputs(6301) <= a xor b;
    layer6_outputs(6302) <= not a;
    layer6_outputs(6303) <= not (a and b);
    layer6_outputs(6304) <= not (a xor b);
    layer6_outputs(6305) <= not b;
    layer6_outputs(6306) <= b;
    layer6_outputs(6307) <= a;
    layer6_outputs(6308) <= a and not b;
    layer6_outputs(6309) <= not a;
    layer6_outputs(6310) <= not a;
    layer6_outputs(6311) <= b;
    layer6_outputs(6312) <= a;
    layer6_outputs(6313) <= a and b;
    layer6_outputs(6314) <= a;
    layer6_outputs(6315) <= b and not a;
    layer6_outputs(6316) <= not a or b;
    layer6_outputs(6317) <= not (a xor b);
    layer6_outputs(6318) <= a;
    layer6_outputs(6319) <= not a or b;
    layer6_outputs(6320) <= a;
    layer6_outputs(6321) <= not b;
    layer6_outputs(6322) <= b;
    layer6_outputs(6323) <= not b or a;
    layer6_outputs(6324) <= b and not a;
    layer6_outputs(6325) <= not (a xor b);
    layer6_outputs(6326) <= a xor b;
    layer6_outputs(6327) <= not (a xor b);
    layer6_outputs(6328) <= not b;
    layer6_outputs(6329) <= not a;
    layer6_outputs(6330) <= a or b;
    layer6_outputs(6331) <= a and not b;
    layer6_outputs(6332) <= a;
    layer6_outputs(6333) <= b and not a;
    layer6_outputs(6334) <= not b;
    layer6_outputs(6335) <= a and not b;
    layer6_outputs(6336) <= not a;
    layer6_outputs(6337) <= not (a or b);
    layer6_outputs(6338) <= not b or a;
    layer6_outputs(6339) <= a xor b;
    layer6_outputs(6340) <= a;
    layer6_outputs(6341) <= a xor b;
    layer6_outputs(6342) <= not (a xor b);
    layer6_outputs(6343) <= not (a or b);
    layer6_outputs(6344) <= a xor b;
    layer6_outputs(6345) <= not a;
    layer6_outputs(6346) <= a and b;
    layer6_outputs(6347) <= a;
    layer6_outputs(6348) <= not b;
    layer6_outputs(6349) <= not b;
    layer6_outputs(6350) <= b;
    layer6_outputs(6351) <= b;
    layer6_outputs(6352) <= not b;
    layer6_outputs(6353) <= not a;
    layer6_outputs(6354) <= not a or b;
    layer6_outputs(6355) <= not (a xor b);
    layer6_outputs(6356) <= b;
    layer6_outputs(6357) <= not b;
    layer6_outputs(6358) <= a or b;
    layer6_outputs(6359) <= b;
    layer6_outputs(6360) <= a xor b;
    layer6_outputs(6361) <= b and not a;
    layer6_outputs(6362) <= not b;
    layer6_outputs(6363) <= a xor b;
    layer6_outputs(6364) <= not (a and b);
    layer6_outputs(6365) <= not b or a;
    layer6_outputs(6366) <= a and not b;
    layer6_outputs(6367) <= not a;
    layer6_outputs(6368) <= b and not a;
    layer6_outputs(6369) <= b;
    layer6_outputs(6370) <= not a;
    layer6_outputs(6371) <= not b;
    layer6_outputs(6372) <= b;
    layer6_outputs(6373) <= not (a and b);
    layer6_outputs(6374) <= b;
    layer6_outputs(6375) <= b;
    layer6_outputs(6376) <= not a;
    layer6_outputs(6377) <= a;
    layer6_outputs(6378) <= not a;
    layer6_outputs(6379) <= a or b;
    layer6_outputs(6380) <= not b;
    layer6_outputs(6381) <= not b;
    layer6_outputs(6382) <= a;
    layer6_outputs(6383) <= a xor b;
    layer6_outputs(6384) <= not (a xor b);
    layer6_outputs(6385) <= not b;
    layer6_outputs(6386) <= a or b;
    layer6_outputs(6387) <= a and not b;
    layer6_outputs(6388) <= b;
    layer6_outputs(6389) <= a and b;
    layer6_outputs(6390) <= a;
    layer6_outputs(6391) <= not a;
    layer6_outputs(6392) <= not (a or b);
    layer6_outputs(6393) <= a and b;
    layer6_outputs(6394) <= not (a xor b);
    layer6_outputs(6395) <= a;
    layer6_outputs(6396) <= b;
    layer6_outputs(6397) <= not b;
    layer6_outputs(6398) <= '1';
    layer6_outputs(6399) <= b;
    layer6_outputs(6400) <= a or b;
    layer6_outputs(6401) <= not b;
    layer6_outputs(6402) <= not b or a;
    layer6_outputs(6403) <= not (a or b);
    layer6_outputs(6404) <= b;
    layer6_outputs(6405) <= a and b;
    layer6_outputs(6406) <= a xor b;
    layer6_outputs(6407) <= a xor b;
    layer6_outputs(6408) <= a;
    layer6_outputs(6409) <= b;
    layer6_outputs(6410) <= a xor b;
    layer6_outputs(6411) <= not b;
    layer6_outputs(6412) <= not (a xor b);
    layer6_outputs(6413) <= b;
    layer6_outputs(6414) <= not (a and b);
    layer6_outputs(6415) <= not b or a;
    layer6_outputs(6416) <= not a;
    layer6_outputs(6417) <= not b or a;
    layer6_outputs(6418) <= a or b;
    layer6_outputs(6419) <= a and b;
    layer6_outputs(6420) <= not b or a;
    layer6_outputs(6421) <= a and not b;
    layer6_outputs(6422) <= not a or b;
    layer6_outputs(6423) <= a and b;
    layer6_outputs(6424) <= not (a xor b);
    layer6_outputs(6425) <= not a;
    layer6_outputs(6426) <= a xor b;
    layer6_outputs(6427) <= not b;
    layer6_outputs(6428) <= not (a xor b);
    layer6_outputs(6429) <= a;
    layer6_outputs(6430) <= a and not b;
    layer6_outputs(6431) <= a xor b;
    layer6_outputs(6432) <= a and not b;
    layer6_outputs(6433) <= a or b;
    layer6_outputs(6434) <= not (a and b);
    layer6_outputs(6435) <= not a;
    layer6_outputs(6436) <= a or b;
    layer6_outputs(6437) <= a;
    layer6_outputs(6438) <= b and not a;
    layer6_outputs(6439) <= not a;
    layer6_outputs(6440) <= not (a xor b);
    layer6_outputs(6441) <= b;
    layer6_outputs(6442) <= not a;
    layer6_outputs(6443) <= not (a xor b);
    layer6_outputs(6444) <= not b;
    layer6_outputs(6445) <= b;
    layer6_outputs(6446) <= not a or b;
    layer6_outputs(6447) <= not a or b;
    layer6_outputs(6448) <= a and b;
    layer6_outputs(6449) <= not b;
    layer6_outputs(6450) <= a xor b;
    layer6_outputs(6451) <= b;
    layer6_outputs(6452) <= b;
    layer6_outputs(6453) <= b;
    layer6_outputs(6454) <= not a;
    layer6_outputs(6455) <= not b;
    layer6_outputs(6456) <= not (a xor b);
    layer6_outputs(6457) <= b;
    layer6_outputs(6458) <= not a or b;
    layer6_outputs(6459) <= b;
    layer6_outputs(6460) <= a xor b;
    layer6_outputs(6461) <= a;
    layer6_outputs(6462) <= a and b;
    layer6_outputs(6463) <= not a;
    layer6_outputs(6464) <= a and not b;
    layer6_outputs(6465) <= not a;
    layer6_outputs(6466) <= b;
    layer6_outputs(6467) <= a;
    layer6_outputs(6468) <= b and not a;
    layer6_outputs(6469) <= not b or a;
    layer6_outputs(6470) <= not a;
    layer6_outputs(6471) <= a;
    layer6_outputs(6472) <= not b;
    layer6_outputs(6473) <= b;
    layer6_outputs(6474) <= a;
    layer6_outputs(6475) <= '1';
    layer6_outputs(6476) <= not (a xor b);
    layer6_outputs(6477) <= not a;
    layer6_outputs(6478) <= b;
    layer6_outputs(6479) <= a;
    layer6_outputs(6480) <= a xor b;
    layer6_outputs(6481) <= b;
    layer6_outputs(6482) <= not (a or b);
    layer6_outputs(6483) <= a;
    layer6_outputs(6484) <= not b;
    layer6_outputs(6485) <= a;
    layer6_outputs(6486) <= a xor b;
    layer6_outputs(6487) <= not b;
    layer6_outputs(6488) <= not (a or b);
    layer6_outputs(6489) <= a xor b;
    layer6_outputs(6490) <= a and b;
    layer6_outputs(6491) <= a and b;
    layer6_outputs(6492) <= not b;
    layer6_outputs(6493) <= not b;
    layer6_outputs(6494) <= not b;
    layer6_outputs(6495) <= not b;
    layer6_outputs(6496) <= not (a and b);
    layer6_outputs(6497) <= b;
    layer6_outputs(6498) <= a;
    layer6_outputs(6499) <= b;
    layer6_outputs(6500) <= not (a and b);
    layer6_outputs(6501) <= a or b;
    layer6_outputs(6502) <= b;
    layer6_outputs(6503) <= not (a xor b);
    layer6_outputs(6504) <= a;
    layer6_outputs(6505) <= b and not a;
    layer6_outputs(6506) <= not b;
    layer6_outputs(6507) <= b;
    layer6_outputs(6508) <= not a;
    layer6_outputs(6509) <= not a or b;
    layer6_outputs(6510) <= a xor b;
    layer6_outputs(6511) <= a or b;
    layer6_outputs(6512) <= not a or b;
    layer6_outputs(6513) <= not (a xor b);
    layer6_outputs(6514) <= a;
    layer6_outputs(6515) <= not a;
    layer6_outputs(6516) <= not a or b;
    layer6_outputs(6517) <= not a;
    layer6_outputs(6518) <= a;
    layer6_outputs(6519) <= not (a or b);
    layer6_outputs(6520) <= a;
    layer6_outputs(6521) <= not b or a;
    layer6_outputs(6522) <= not (a xor b);
    layer6_outputs(6523) <= not (a xor b);
    layer6_outputs(6524) <= b;
    layer6_outputs(6525) <= a xor b;
    layer6_outputs(6526) <= not a or b;
    layer6_outputs(6527) <= a xor b;
    layer6_outputs(6528) <= not (a and b);
    layer6_outputs(6529) <= not b;
    layer6_outputs(6530) <= a xor b;
    layer6_outputs(6531) <= a;
    layer6_outputs(6532) <= a and not b;
    layer6_outputs(6533) <= a xor b;
    layer6_outputs(6534) <= not (a and b);
    layer6_outputs(6535) <= b;
    layer6_outputs(6536) <= not (a xor b);
    layer6_outputs(6537) <= not (a xor b);
    layer6_outputs(6538) <= a;
    layer6_outputs(6539) <= a xor b;
    layer6_outputs(6540) <= a xor b;
    layer6_outputs(6541) <= not b or a;
    layer6_outputs(6542) <= a or b;
    layer6_outputs(6543) <= not (a or b);
    layer6_outputs(6544) <= b;
    layer6_outputs(6545) <= b and not a;
    layer6_outputs(6546) <= not a;
    layer6_outputs(6547) <= b and not a;
    layer6_outputs(6548) <= a;
    layer6_outputs(6549) <= a;
    layer6_outputs(6550) <= not b;
    layer6_outputs(6551) <= not (a or b);
    layer6_outputs(6552) <= b and not a;
    layer6_outputs(6553) <= not b or a;
    layer6_outputs(6554) <= not (a xor b);
    layer6_outputs(6555) <= a;
    layer6_outputs(6556) <= b and not a;
    layer6_outputs(6557) <= a;
    layer6_outputs(6558) <= not a or b;
    layer6_outputs(6559) <= a xor b;
    layer6_outputs(6560) <= a;
    layer6_outputs(6561) <= not (a and b);
    layer6_outputs(6562) <= a xor b;
    layer6_outputs(6563) <= not b;
    layer6_outputs(6564) <= b;
    layer6_outputs(6565) <= b and not a;
    layer6_outputs(6566) <= not a;
    layer6_outputs(6567) <= not b;
    layer6_outputs(6568) <= a;
    layer6_outputs(6569) <= not a;
    layer6_outputs(6570) <= not a;
    layer6_outputs(6571) <= a and not b;
    layer6_outputs(6572) <= not (a xor b);
    layer6_outputs(6573) <= a xor b;
    layer6_outputs(6574) <= not b;
    layer6_outputs(6575) <= a xor b;
    layer6_outputs(6576) <= not b;
    layer6_outputs(6577) <= not a;
    layer6_outputs(6578) <= not (a or b);
    layer6_outputs(6579) <= a xor b;
    layer6_outputs(6580) <= not b;
    layer6_outputs(6581) <= not b or a;
    layer6_outputs(6582) <= not (a or b);
    layer6_outputs(6583) <= not (a xor b);
    layer6_outputs(6584) <= not a;
    layer6_outputs(6585) <= a and not b;
    layer6_outputs(6586) <= not (a xor b);
    layer6_outputs(6587) <= not (a and b);
    layer6_outputs(6588) <= not b;
    layer6_outputs(6589) <= a;
    layer6_outputs(6590) <= a and not b;
    layer6_outputs(6591) <= not (a and b);
    layer6_outputs(6592) <= b;
    layer6_outputs(6593) <= b;
    layer6_outputs(6594) <= not b;
    layer6_outputs(6595) <= b;
    layer6_outputs(6596) <= not b;
    layer6_outputs(6597) <= not (a xor b);
    layer6_outputs(6598) <= not a;
    layer6_outputs(6599) <= not b;
    layer6_outputs(6600) <= not a;
    layer6_outputs(6601) <= b;
    layer6_outputs(6602) <= not (a xor b);
    layer6_outputs(6603) <= a xor b;
    layer6_outputs(6604) <= not (a and b);
    layer6_outputs(6605) <= a;
    layer6_outputs(6606) <= not a or b;
    layer6_outputs(6607) <= a and not b;
    layer6_outputs(6608) <= not a or b;
    layer6_outputs(6609) <= b;
    layer6_outputs(6610) <= a xor b;
    layer6_outputs(6611) <= b and not a;
    layer6_outputs(6612) <= not (a xor b);
    layer6_outputs(6613) <= not b;
    layer6_outputs(6614) <= not (a xor b);
    layer6_outputs(6615) <= a;
    layer6_outputs(6616) <= a and not b;
    layer6_outputs(6617) <= not a;
    layer6_outputs(6618) <= not a;
    layer6_outputs(6619) <= not a;
    layer6_outputs(6620) <= a or b;
    layer6_outputs(6621) <= not b;
    layer6_outputs(6622) <= not (a or b);
    layer6_outputs(6623) <= a xor b;
    layer6_outputs(6624) <= not b;
    layer6_outputs(6625) <= not a or b;
    layer6_outputs(6626) <= a or b;
    layer6_outputs(6627) <= not (a xor b);
    layer6_outputs(6628) <= not (a and b);
    layer6_outputs(6629) <= b;
    layer6_outputs(6630) <= b;
    layer6_outputs(6631) <= a xor b;
    layer6_outputs(6632) <= not b;
    layer6_outputs(6633) <= not b;
    layer6_outputs(6634) <= a and not b;
    layer6_outputs(6635) <= a;
    layer6_outputs(6636) <= a xor b;
    layer6_outputs(6637) <= a xor b;
    layer6_outputs(6638) <= b and not a;
    layer6_outputs(6639) <= not a;
    layer6_outputs(6640) <= a and b;
    layer6_outputs(6641) <= not a;
    layer6_outputs(6642) <= not (a or b);
    layer6_outputs(6643) <= not b;
    layer6_outputs(6644) <= not a;
    layer6_outputs(6645) <= a;
    layer6_outputs(6646) <= not (a xor b);
    layer6_outputs(6647) <= not b;
    layer6_outputs(6648) <= b;
    layer6_outputs(6649) <= not b;
    layer6_outputs(6650) <= a or b;
    layer6_outputs(6651) <= a and b;
    layer6_outputs(6652) <= not a;
    layer6_outputs(6653) <= a xor b;
    layer6_outputs(6654) <= not b;
    layer6_outputs(6655) <= not b;
    layer6_outputs(6656) <= a xor b;
    layer6_outputs(6657) <= not b or a;
    layer6_outputs(6658) <= not (a xor b);
    layer6_outputs(6659) <= not b;
    layer6_outputs(6660) <= a xor b;
    layer6_outputs(6661) <= not a;
    layer6_outputs(6662) <= b and not a;
    layer6_outputs(6663) <= not b;
    layer6_outputs(6664) <= a xor b;
    layer6_outputs(6665) <= not (a xor b);
    layer6_outputs(6666) <= not (a xor b);
    layer6_outputs(6667) <= b;
    layer6_outputs(6668) <= not b;
    layer6_outputs(6669) <= a xor b;
    layer6_outputs(6670) <= a;
    layer6_outputs(6671) <= a xor b;
    layer6_outputs(6672) <= not b;
    layer6_outputs(6673) <= not (a xor b);
    layer6_outputs(6674) <= '0';
    layer6_outputs(6675) <= not a;
    layer6_outputs(6676) <= not (a or b);
    layer6_outputs(6677) <= b;
    layer6_outputs(6678) <= a or b;
    layer6_outputs(6679) <= not b;
    layer6_outputs(6680) <= not (a xor b);
    layer6_outputs(6681) <= not (a xor b);
    layer6_outputs(6682) <= b;
    layer6_outputs(6683) <= a and not b;
    layer6_outputs(6684) <= not (a xor b);
    layer6_outputs(6685) <= b;
    layer6_outputs(6686) <= '0';
    layer6_outputs(6687) <= a or b;
    layer6_outputs(6688) <= a and b;
    layer6_outputs(6689) <= not b;
    layer6_outputs(6690) <= a;
    layer6_outputs(6691) <= a and not b;
    layer6_outputs(6692) <= a and b;
    layer6_outputs(6693) <= not b;
    layer6_outputs(6694) <= a;
    layer6_outputs(6695) <= a xor b;
    layer6_outputs(6696) <= a xor b;
    layer6_outputs(6697) <= a xor b;
    layer6_outputs(6698) <= not b or a;
    layer6_outputs(6699) <= a xor b;
    layer6_outputs(6700) <= a xor b;
    layer6_outputs(6701) <= not (a xor b);
    layer6_outputs(6702) <= not b or a;
    layer6_outputs(6703) <= b;
    layer6_outputs(6704) <= a xor b;
    layer6_outputs(6705) <= not a;
    layer6_outputs(6706) <= not (a xor b);
    layer6_outputs(6707) <= not a or b;
    layer6_outputs(6708) <= a and b;
    layer6_outputs(6709) <= b;
    layer6_outputs(6710) <= not b;
    layer6_outputs(6711) <= not (a and b);
    layer6_outputs(6712) <= a and not b;
    layer6_outputs(6713) <= not (a or b);
    layer6_outputs(6714) <= a xor b;
    layer6_outputs(6715) <= not b;
    layer6_outputs(6716) <= not (a xor b);
    layer6_outputs(6717) <= a;
    layer6_outputs(6718) <= a or b;
    layer6_outputs(6719) <= not b or a;
    layer6_outputs(6720) <= a;
    layer6_outputs(6721) <= b;
    layer6_outputs(6722) <= not (a or b);
    layer6_outputs(6723) <= not (a or b);
    layer6_outputs(6724) <= not (a and b);
    layer6_outputs(6725) <= a or b;
    layer6_outputs(6726) <= not a or b;
    layer6_outputs(6727) <= not (a xor b);
    layer6_outputs(6728) <= not a;
    layer6_outputs(6729) <= not a;
    layer6_outputs(6730) <= a;
    layer6_outputs(6731) <= b;
    layer6_outputs(6732) <= a;
    layer6_outputs(6733) <= not b;
    layer6_outputs(6734) <= b;
    layer6_outputs(6735) <= not b;
    layer6_outputs(6736) <= not b;
    layer6_outputs(6737) <= not (a xor b);
    layer6_outputs(6738) <= not b;
    layer6_outputs(6739) <= not a;
    layer6_outputs(6740) <= not (a xor b);
    layer6_outputs(6741) <= not (a xor b);
    layer6_outputs(6742) <= not (a xor b);
    layer6_outputs(6743) <= not (a and b);
    layer6_outputs(6744) <= not a;
    layer6_outputs(6745) <= not b;
    layer6_outputs(6746) <= not a or b;
    layer6_outputs(6747) <= not b or a;
    layer6_outputs(6748) <= not a or b;
    layer6_outputs(6749) <= a xor b;
    layer6_outputs(6750) <= not b or a;
    layer6_outputs(6751) <= b;
    layer6_outputs(6752) <= not a;
    layer6_outputs(6753) <= b;
    layer6_outputs(6754) <= not a;
    layer6_outputs(6755) <= not a;
    layer6_outputs(6756) <= b and not a;
    layer6_outputs(6757) <= a and b;
    layer6_outputs(6758) <= b;
    layer6_outputs(6759) <= a;
    layer6_outputs(6760) <= a;
    layer6_outputs(6761) <= not a or b;
    layer6_outputs(6762) <= b;
    layer6_outputs(6763) <= not a;
    layer6_outputs(6764) <= a and not b;
    layer6_outputs(6765) <= not (a or b);
    layer6_outputs(6766) <= not (a or b);
    layer6_outputs(6767) <= a and not b;
    layer6_outputs(6768) <= not b;
    layer6_outputs(6769) <= a xor b;
    layer6_outputs(6770) <= b;
    layer6_outputs(6771) <= a;
    layer6_outputs(6772) <= a or b;
    layer6_outputs(6773) <= a xor b;
    layer6_outputs(6774) <= a or b;
    layer6_outputs(6775) <= not a;
    layer6_outputs(6776) <= a xor b;
    layer6_outputs(6777) <= not (a and b);
    layer6_outputs(6778) <= not b;
    layer6_outputs(6779) <= a or b;
    layer6_outputs(6780) <= not a;
    layer6_outputs(6781) <= b and not a;
    layer6_outputs(6782) <= b;
    layer6_outputs(6783) <= not (a xor b);
    layer6_outputs(6784) <= not b;
    layer6_outputs(6785) <= a;
    layer6_outputs(6786) <= b and not a;
    layer6_outputs(6787) <= a and not b;
    layer6_outputs(6788) <= b and not a;
    layer6_outputs(6789) <= not (a or b);
    layer6_outputs(6790) <= not a or b;
    layer6_outputs(6791) <= a xor b;
    layer6_outputs(6792) <= not (a xor b);
    layer6_outputs(6793) <= a;
    layer6_outputs(6794) <= not (a xor b);
    layer6_outputs(6795) <= not a;
    layer6_outputs(6796) <= a or b;
    layer6_outputs(6797) <= a and not b;
    layer6_outputs(6798) <= not (a xor b);
    layer6_outputs(6799) <= a xor b;
    layer6_outputs(6800) <= not a;
    layer6_outputs(6801) <= a;
    layer6_outputs(6802) <= not (a xor b);
    layer6_outputs(6803) <= a;
    layer6_outputs(6804) <= a xor b;
    layer6_outputs(6805) <= not (a xor b);
    layer6_outputs(6806) <= a or b;
    layer6_outputs(6807) <= not (a or b);
    layer6_outputs(6808) <= a xor b;
    layer6_outputs(6809) <= a xor b;
    layer6_outputs(6810) <= a xor b;
    layer6_outputs(6811) <= b;
    layer6_outputs(6812) <= not a;
    layer6_outputs(6813) <= not (a or b);
    layer6_outputs(6814) <= a or b;
    layer6_outputs(6815) <= b and not a;
    layer6_outputs(6816) <= not (a xor b);
    layer6_outputs(6817) <= not a;
    layer6_outputs(6818) <= not a or b;
    layer6_outputs(6819) <= a;
    layer6_outputs(6820) <= b;
    layer6_outputs(6821) <= not a;
    layer6_outputs(6822) <= b;
    layer6_outputs(6823) <= a;
    layer6_outputs(6824) <= not b or a;
    layer6_outputs(6825) <= not a;
    layer6_outputs(6826) <= not (a xor b);
    layer6_outputs(6827) <= not b;
    layer6_outputs(6828) <= not b;
    layer6_outputs(6829) <= a;
    layer6_outputs(6830) <= a;
    layer6_outputs(6831) <= not b or a;
    layer6_outputs(6832) <= not b;
    layer6_outputs(6833) <= not (a xor b);
    layer6_outputs(6834) <= not (a xor b);
    layer6_outputs(6835) <= b and not a;
    layer6_outputs(6836) <= not a or b;
    layer6_outputs(6837) <= b;
    layer6_outputs(6838) <= not b or a;
    layer6_outputs(6839) <= not a;
    layer6_outputs(6840) <= b and not a;
    layer6_outputs(6841) <= not (a and b);
    layer6_outputs(6842) <= not (a or b);
    layer6_outputs(6843) <= not (a xor b);
    layer6_outputs(6844) <= b;
    layer6_outputs(6845) <= a xor b;
    layer6_outputs(6846) <= a xor b;
    layer6_outputs(6847) <= not (a xor b);
    layer6_outputs(6848) <= a;
    layer6_outputs(6849) <= not a;
    layer6_outputs(6850) <= not (a xor b);
    layer6_outputs(6851) <= not a or b;
    layer6_outputs(6852) <= not (a and b);
    layer6_outputs(6853) <= not a or b;
    layer6_outputs(6854) <= a and b;
    layer6_outputs(6855) <= not (a xor b);
    layer6_outputs(6856) <= b;
    layer6_outputs(6857) <= not (a or b);
    layer6_outputs(6858) <= not a or b;
    layer6_outputs(6859) <= not (a xor b);
    layer6_outputs(6860) <= not a;
    layer6_outputs(6861) <= a xor b;
    layer6_outputs(6862) <= not (a xor b);
    layer6_outputs(6863) <= a and not b;
    layer6_outputs(6864) <= a;
    layer6_outputs(6865) <= b;
    layer6_outputs(6866) <= not a or b;
    layer6_outputs(6867) <= b;
    layer6_outputs(6868) <= b and not a;
    layer6_outputs(6869) <= a;
    layer6_outputs(6870) <= not b or a;
    layer6_outputs(6871) <= not a or b;
    layer6_outputs(6872) <= b and not a;
    layer6_outputs(6873) <= not (a and b);
    layer6_outputs(6874) <= a xor b;
    layer6_outputs(6875) <= a xor b;
    layer6_outputs(6876) <= not b;
    layer6_outputs(6877) <= a or b;
    layer6_outputs(6878) <= b and not a;
    layer6_outputs(6879) <= a or b;
    layer6_outputs(6880) <= b;
    layer6_outputs(6881) <= not b or a;
    layer6_outputs(6882) <= not b or a;
    layer6_outputs(6883) <= b and not a;
    layer6_outputs(6884) <= not b;
    layer6_outputs(6885) <= a xor b;
    layer6_outputs(6886) <= a and b;
    layer6_outputs(6887) <= a and not b;
    layer6_outputs(6888) <= not (a or b);
    layer6_outputs(6889) <= a;
    layer6_outputs(6890) <= a and not b;
    layer6_outputs(6891) <= not b;
    layer6_outputs(6892) <= a;
    layer6_outputs(6893) <= a or b;
    layer6_outputs(6894) <= not a or b;
    layer6_outputs(6895) <= a and not b;
    layer6_outputs(6896) <= a;
    layer6_outputs(6897) <= not (a or b);
    layer6_outputs(6898) <= a;
    layer6_outputs(6899) <= a xor b;
    layer6_outputs(6900) <= a and not b;
    layer6_outputs(6901) <= a and not b;
    layer6_outputs(6902) <= a;
    layer6_outputs(6903) <= a and not b;
    layer6_outputs(6904) <= not a;
    layer6_outputs(6905) <= b;
    layer6_outputs(6906) <= not a;
    layer6_outputs(6907) <= b;
    layer6_outputs(6908) <= b;
    layer6_outputs(6909) <= not (a xor b);
    layer6_outputs(6910) <= not b or a;
    layer6_outputs(6911) <= a and not b;
    layer6_outputs(6912) <= a;
    layer6_outputs(6913) <= not a or b;
    layer6_outputs(6914) <= b and not a;
    layer6_outputs(6915) <= not (a xor b);
    layer6_outputs(6916) <= a and not b;
    layer6_outputs(6917) <= a;
    layer6_outputs(6918) <= not (a xor b);
    layer6_outputs(6919) <= not a;
    layer6_outputs(6920) <= b;
    layer6_outputs(6921) <= not b;
    layer6_outputs(6922) <= not (a and b);
    layer6_outputs(6923) <= not (a xor b);
    layer6_outputs(6924) <= a xor b;
    layer6_outputs(6925) <= not (a xor b);
    layer6_outputs(6926) <= not (a xor b);
    layer6_outputs(6927) <= a xor b;
    layer6_outputs(6928) <= a and not b;
    layer6_outputs(6929) <= not b;
    layer6_outputs(6930) <= a;
    layer6_outputs(6931) <= a or b;
    layer6_outputs(6932) <= not a;
    layer6_outputs(6933) <= a;
    layer6_outputs(6934) <= not b;
    layer6_outputs(6935) <= not a;
    layer6_outputs(6936) <= not b;
    layer6_outputs(6937) <= not a;
    layer6_outputs(6938) <= a;
    layer6_outputs(6939) <= not (a or b);
    layer6_outputs(6940) <= not b;
    layer6_outputs(6941) <= a and not b;
    layer6_outputs(6942) <= a and not b;
    layer6_outputs(6943) <= not b;
    layer6_outputs(6944) <= a and not b;
    layer6_outputs(6945) <= not a;
    layer6_outputs(6946) <= a and not b;
    layer6_outputs(6947) <= not b or a;
    layer6_outputs(6948) <= not (a xor b);
    layer6_outputs(6949) <= b;
    layer6_outputs(6950) <= not (a and b);
    layer6_outputs(6951) <= not (a and b);
    layer6_outputs(6952) <= a;
    layer6_outputs(6953) <= not a;
    layer6_outputs(6954) <= b and not a;
    layer6_outputs(6955) <= a;
    layer6_outputs(6956) <= b;
    layer6_outputs(6957) <= a;
    layer6_outputs(6958) <= not b or a;
    layer6_outputs(6959) <= not a;
    layer6_outputs(6960) <= a;
    layer6_outputs(6961) <= not b or a;
    layer6_outputs(6962) <= a xor b;
    layer6_outputs(6963) <= b and not a;
    layer6_outputs(6964) <= not (a and b);
    layer6_outputs(6965) <= not (a xor b);
    layer6_outputs(6966) <= not (a or b);
    layer6_outputs(6967) <= not (a xor b);
    layer6_outputs(6968) <= a xor b;
    layer6_outputs(6969) <= not b;
    layer6_outputs(6970) <= a or b;
    layer6_outputs(6971) <= not a;
    layer6_outputs(6972) <= b;
    layer6_outputs(6973) <= not a;
    layer6_outputs(6974) <= a;
    layer6_outputs(6975) <= b;
    layer6_outputs(6976) <= b and not a;
    layer6_outputs(6977) <= not b;
    layer6_outputs(6978) <= not b;
    layer6_outputs(6979) <= a;
    layer6_outputs(6980) <= a xor b;
    layer6_outputs(6981) <= not a;
    layer6_outputs(6982) <= b;
    layer6_outputs(6983) <= not (a xor b);
    layer6_outputs(6984) <= not b;
    layer6_outputs(6985) <= a;
    layer6_outputs(6986) <= a;
    layer6_outputs(6987) <= not (a xor b);
    layer6_outputs(6988) <= b;
    layer6_outputs(6989) <= not (a xor b);
    layer6_outputs(6990) <= a xor b;
    layer6_outputs(6991) <= not (a and b);
    layer6_outputs(6992) <= b;
    layer6_outputs(6993) <= b and not a;
    layer6_outputs(6994) <= not b;
    layer6_outputs(6995) <= a;
    layer6_outputs(6996) <= not b;
    layer6_outputs(6997) <= not (a or b);
    layer6_outputs(6998) <= b;
    layer6_outputs(6999) <= not (a xor b);
    layer6_outputs(7000) <= a;
    layer6_outputs(7001) <= b;
    layer6_outputs(7002) <= not a;
    layer6_outputs(7003) <= a xor b;
    layer6_outputs(7004) <= a and not b;
    layer6_outputs(7005) <= not b;
    layer6_outputs(7006) <= a and b;
    layer6_outputs(7007) <= a and b;
    layer6_outputs(7008) <= not (a xor b);
    layer6_outputs(7009) <= not a;
    layer6_outputs(7010) <= b;
    layer6_outputs(7011) <= not (a xor b);
    layer6_outputs(7012) <= a;
    layer6_outputs(7013) <= b;
    layer6_outputs(7014) <= not b;
    layer6_outputs(7015) <= a;
    layer6_outputs(7016) <= b and not a;
    layer6_outputs(7017) <= not (a and b);
    layer6_outputs(7018) <= b;
    layer6_outputs(7019) <= a and not b;
    layer6_outputs(7020) <= not a;
    layer6_outputs(7021) <= not b or a;
    layer6_outputs(7022) <= b and not a;
    layer6_outputs(7023) <= not (a xor b);
    layer6_outputs(7024) <= not b;
    layer6_outputs(7025) <= not b or a;
    layer6_outputs(7026) <= not b;
    layer6_outputs(7027) <= b;
    layer6_outputs(7028) <= not a;
    layer6_outputs(7029) <= a xor b;
    layer6_outputs(7030) <= a;
    layer6_outputs(7031) <= not (a and b);
    layer6_outputs(7032) <= a xor b;
    layer6_outputs(7033) <= not (a xor b);
    layer6_outputs(7034) <= a xor b;
    layer6_outputs(7035) <= not b;
    layer6_outputs(7036) <= not a;
    layer6_outputs(7037) <= not a or b;
    layer6_outputs(7038) <= a;
    layer6_outputs(7039) <= a xor b;
    layer6_outputs(7040) <= not (a or b);
    layer6_outputs(7041) <= a and not b;
    layer6_outputs(7042) <= b;
    layer6_outputs(7043) <= b;
    layer6_outputs(7044) <= not b or a;
    layer6_outputs(7045) <= not b;
    layer6_outputs(7046) <= not a;
    layer6_outputs(7047) <= a xor b;
    layer6_outputs(7048) <= not (a and b);
    layer6_outputs(7049) <= not a;
    layer6_outputs(7050) <= not b;
    layer6_outputs(7051) <= b and not a;
    layer6_outputs(7052) <= not a;
    layer6_outputs(7053) <= not b;
    layer6_outputs(7054) <= not a or b;
    layer6_outputs(7055) <= not (a xor b);
    layer6_outputs(7056) <= a or b;
    layer6_outputs(7057) <= not (a or b);
    layer6_outputs(7058) <= b;
    layer6_outputs(7059) <= b;
    layer6_outputs(7060) <= not b;
    layer6_outputs(7061) <= not a;
    layer6_outputs(7062) <= not b;
    layer6_outputs(7063) <= not (a or b);
    layer6_outputs(7064) <= not a;
    layer6_outputs(7065) <= a xor b;
    layer6_outputs(7066) <= a and not b;
    layer6_outputs(7067) <= a and b;
    layer6_outputs(7068) <= b;
    layer6_outputs(7069) <= not (a xor b);
    layer6_outputs(7070) <= not a;
    layer6_outputs(7071) <= not (a or b);
    layer6_outputs(7072) <= not (a and b);
    layer6_outputs(7073) <= a or b;
    layer6_outputs(7074) <= a xor b;
    layer6_outputs(7075) <= not (a or b);
    layer6_outputs(7076) <= a xor b;
    layer6_outputs(7077) <= a and not b;
    layer6_outputs(7078) <= not (a and b);
    layer6_outputs(7079) <= b;
    layer6_outputs(7080) <= a xor b;
    layer6_outputs(7081) <= b;
    layer6_outputs(7082) <= a or b;
    layer6_outputs(7083) <= not (a xor b);
    layer6_outputs(7084) <= not b;
    layer6_outputs(7085) <= not a;
    layer6_outputs(7086) <= a;
    layer6_outputs(7087) <= not b;
    layer6_outputs(7088) <= b;
    layer6_outputs(7089) <= not b;
    layer6_outputs(7090) <= not (a xor b);
    layer6_outputs(7091) <= b and not a;
    layer6_outputs(7092) <= a xor b;
    layer6_outputs(7093) <= b;
    layer6_outputs(7094) <= not (a or b);
    layer6_outputs(7095) <= not a or b;
    layer6_outputs(7096) <= not a;
    layer6_outputs(7097) <= not a or b;
    layer6_outputs(7098) <= a;
    layer6_outputs(7099) <= not b;
    layer6_outputs(7100) <= a and b;
    layer6_outputs(7101) <= a and not b;
    layer6_outputs(7102) <= b and not a;
    layer6_outputs(7103) <= a and not b;
    layer6_outputs(7104) <= not a;
    layer6_outputs(7105) <= '1';
    layer6_outputs(7106) <= a and b;
    layer6_outputs(7107) <= a and not b;
    layer6_outputs(7108) <= b;
    layer6_outputs(7109) <= not b or a;
    layer6_outputs(7110) <= not a;
    layer6_outputs(7111) <= not b or a;
    layer6_outputs(7112) <= not (a and b);
    layer6_outputs(7113) <= a or b;
    layer6_outputs(7114) <= not b;
    layer6_outputs(7115) <= not b;
    layer6_outputs(7116) <= a;
    layer6_outputs(7117) <= not (a and b);
    layer6_outputs(7118) <= a;
    layer6_outputs(7119) <= not (a or b);
    layer6_outputs(7120) <= a xor b;
    layer6_outputs(7121) <= a xor b;
    layer6_outputs(7122) <= not (a xor b);
    layer6_outputs(7123) <= b and not a;
    layer6_outputs(7124) <= a;
    layer6_outputs(7125) <= not b or a;
    layer6_outputs(7126) <= not a;
    layer6_outputs(7127) <= a xor b;
    layer6_outputs(7128) <= not (a xor b);
    layer6_outputs(7129) <= a and b;
    layer6_outputs(7130) <= not b;
    layer6_outputs(7131) <= b;
    layer6_outputs(7132) <= not a;
    layer6_outputs(7133) <= not (a xor b);
    layer6_outputs(7134) <= not (a and b);
    layer6_outputs(7135) <= not b;
    layer6_outputs(7136) <= not b;
    layer6_outputs(7137) <= a;
    layer6_outputs(7138) <= not (a xor b);
    layer6_outputs(7139) <= b;
    layer6_outputs(7140) <= not a or b;
    layer6_outputs(7141) <= a;
    layer6_outputs(7142) <= b;
    layer6_outputs(7143) <= not (a and b);
    layer6_outputs(7144) <= not (a xor b);
    layer6_outputs(7145) <= b;
    layer6_outputs(7146) <= a and b;
    layer6_outputs(7147) <= a and not b;
    layer6_outputs(7148) <= not b or a;
    layer6_outputs(7149) <= a or b;
    layer6_outputs(7150) <= not (a xor b);
    layer6_outputs(7151) <= not a;
    layer6_outputs(7152) <= b;
    layer6_outputs(7153) <= not (a and b);
    layer6_outputs(7154) <= not (a xor b);
    layer6_outputs(7155) <= not a or b;
    layer6_outputs(7156) <= not b;
    layer6_outputs(7157) <= not a;
    layer6_outputs(7158) <= a or b;
    layer6_outputs(7159) <= not (a xor b);
    layer6_outputs(7160) <= not b;
    layer6_outputs(7161) <= b;
    layer6_outputs(7162) <= not (a xor b);
    layer6_outputs(7163) <= not b;
    layer6_outputs(7164) <= a xor b;
    layer6_outputs(7165) <= not b or a;
    layer6_outputs(7166) <= not b or a;
    layer6_outputs(7167) <= a xor b;
    layer6_outputs(7168) <= a;
    layer6_outputs(7169) <= b;
    layer6_outputs(7170) <= b;
    layer6_outputs(7171) <= a;
    layer6_outputs(7172) <= a xor b;
    layer6_outputs(7173) <= b;
    layer6_outputs(7174) <= a xor b;
    layer6_outputs(7175) <= a or b;
    layer6_outputs(7176) <= a xor b;
    layer6_outputs(7177) <= a;
    layer6_outputs(7178) <= a or b;
    layer6_outputs(7179) <= not a or b;
    layer6_outputs(7180) <= a xor b;
    layer6_outputs(7181) <= not (a and b);
    layer6_outputs(7182) <= a;
    layer6_outputs(7183) <= a xor b;
    layer6_outputs(7184) <= not b or a;
    layer6_outputs(7185) <= not a;
    layer6_outputs(7186) <= b;
    layer6_outputs(7187) <= not b;
    layer6_outputs(7188) <= not b;
    layer6_outputs(7189) <= b;
    layer6_outputs(7190) <= a xor b;
    layer6_outputs(7191) <= a and not b;
    layer6_outputs(7192) <= not (a or b);
    layer6_outputs(7193) <= a;
    layer6_outputs(7194) <= not (a and b);
    layer6_outputs(7195) <= not a or b;
    layer6_outputs(7196) <= not a;
    layer6_outputs(7197) <= b;
    layer6_outputs(7198) <= not b;
    layer6_outputs(7199) <= not a or b;
    layer6_outputs(7200) <= b;
    layer6_outputs(7201) <= b;
    layer6_outputs(7202) <= not a;
    layer6_outputs(7203) <= not b;
    layer6_outputs(7204) <= a and b;
    layer6_outputs(7205) <= not a or b;
    layer6_outputs(7206) <= a and not b;
    layer6_outputs(7207) <= a and b;
    layer6_outputs(7208) <= b and not a;
    layer6_outputs(7209) <= not (a xor b);
    layer6_outputs(7210) <= not a;
    layer6_outputs(7211) <= not b;
    layer6_outputs(7212) <= not (a xor b);
    layer6_outputs(7213) <= not a;
    layer6_outputs(7214) <= a xor b;
    layer6_outputs(7215) <= a;
    layer6_outputs(7216) <= a xor b;
    layer6_outputs(7217) <= not a or b;
    layer6_outputs(7218) <= b;
    layer6_outputs(7219) <= a xor b;
    layer6_outputs(7220) <= not (a xor b);
    layer6_outputs(7221) <= not (a xor b);
    layer6_outputs(7222) <= a xor b;
    layer6_outputs(7223) <= a or b;
    layer6_outputs(7224) <= not (a or b);
    layer6_outputs(7225) <= not (a xor b);
    layer6_outputs(7226) <= not a or b;
    layer6_outputs(7227) <= b;
    layer6_outputs(7228) <= b;
    layer6_outputs(7229) <= not b;
    layer6_outputs(7230) <= a or b;
    layer6_outputs(7231) <= b and not a;
    layer6_outputs(7232) <= not a or b;
    layer6_outputs(7233) <= not a;
    layer6_outputs(7234) <= not (a and b);
    layer6_outputs(7235) <= b;
    layer6_outputs(7236) <= not a;
    layer6_outputs(7237) <= not b;
    layer6_outputs(7238) <= a;
    layer6_outputs(7239) <= not a or b;
    layer6_outputs(7240) <= a;
    layer6_outputs(7241) <= not b;
    layer6_outputs(7242) <= not (a xor b);
    layer6_outputs(7243) <= not a;
    layer6_outputs(7244) <= a;
    layer6_outputs(7245) <= b;
    layer6_outputs(7246) <= not a or b;
    layer6_outputs(7247) <= a xor b;
    layer6_outputs(7248) <= b and not a;
    layer6_outputs(7249) <= a or b;
    layer6_outputs(7250) <= b;
    layer6_outputs(7251) <= not a;
    layer6_outputs(7252) <= a;
    layer6_outputs(7253) <= a;
    layer6_outputs(7254) <= not b;
    layer6_outputs(7255) <= not b or a;
    layer6_outputs(7256) <= b and not a;
    layer6_outputs(7257) <= not (a xor b);
    layer6_outputs(7258) <= not (a xor b);
    layer6_outputs(7259) <= not a;
    layer6_outputs(7260) <= '1';
    layer6_outputs(7261) <= not a or b;
    layer6_outputs(7262) <= not (a and b);
    layer6_outputs(7263) <= a;
    layer6_outputs(7264) <= not b;
    layer6_outputs(7265) <= not b;
    layer6_outputs(7266) <= a;
    layer6_outputs(7267) <= not (a xor b);
    layer6_outputs(7268) <= b;
    layer6_outputs(7269) <= not (a or b);
    layer6_outputs(7270) <= b and not a;
    layer6_outputs(7271) <= b;
    layer6_outputs(7272) <= not b or a;
    layer6_outputs(7273) <= not (a and b);
    layer6_outputs(7274) <= a or b;
    layer6_outputs(7275) <= a;
    layer6_outputs(7276) <= a;
    layer6_outputs(7277) <= a;
    layer6_outputs(7278) <= not b;
    layer6_outputs(7279) <= b;
    layer6_outputs(7280) <= a xor b;
    layer6_outputs(7281) <= not a or b;
    layer6_outputs(7282) <= not (a xor b);
    layer6_outputs(7283) <= not b;
    layer6_outputs(7284) <= a and not b;
    layer6_outputs(7285) <= a;
    layer6_outputs(7286) <= not a;
    layer6_outputs(7287) <= not (a or b);
    layer6_outputs(7288) <= a;
    layer6_outputs(7289) <= b;
    layer6_outputs(7290) <= a or b;
    layer6_outputs(7291) <= not b;
    layer6_outputs(7292) <= b;
    layer6_outputs(7293) <= b;
    layer6_outputs(7294) <= b;
    layer6_outputs(7295) <= not a or b;
    layer6_outputs(7296) <= not a;
    layer6_outputs(7297) <= not a;
    layer6_outputs(7298) <= not (a xor b);
    layer6_outputs(7299) <= a;
    layer6_outputs(7300) <= b and not a;
    layer6_outputs(7301) <= a and not b;
    layer6_outputs(7302) <= b and not a;
    layer6_outputs(7303) <= not a;
    layer6_outputs(7304) <= b;
    layer6_outputs(7305) <= b and not a;
    layer6_outputs(7306) <= not b;
    layer6_outputs(7307) <= b and not a;
    layer6_outputs(7308) <= a;
    layer6_outputs(7309) <= '0';
    layer6_outputs(7310) <= b and not a;
    layer6_outputs(7311) <= b;
    layer6_outputs(7312) <= a and b;
    layer6_outputs(7313) <= not b;
    layer6_outputs(7314) <= a or b;
    layer6_outputs(7315) <= not b;
    layer6_outputs(7316) <= not b;
    layer6_outputs(7317) <= not b;
    layer6_outputs(7318) <= not b;
    layer6_outputs(7319) <= a xor b;
    layer6_outputs(7320) <= a;
    layer6_outputs(7321) <= a or b;
    layer6_outputs(7322) <= b;
    layer6_outputs(7323) <= not b;
    layer6_outputs(7324) <= a xor b;
    layer6_outputs(7325) <= not b or a;
    layer6_outputs(7326) <= a;
    layer6_outputs(7327) <= a;
    layer6_outputs(7328) <= b;
    layer6_outputs(7329) <= not b;
    layer6_outputs(7330) <= a;
    layer6_outputs(7331) <= a xor b;
    layer6_outputs(7332) <= not a;
    layer6_outputs(7333) <= a;
    layer6_outputs(7334) <= not b;
    layer6_outputs(7335) <= not a or b;
    layer6_outputs(7336) <= a and not b;
    layer6_outputs(7337) <= not (a or b);
    layer6_outputs(7338) <= a and not b;
    layer6_outputs(7339) <= b;
    layer6_outputs(7340) <= b;
    layer6_outputs(7341) <= a;
    layer6_outputs(7342) <= not b;
    layer6_outputs(7343) <= not b;
    layer6_outputs(7344) <= not (a xor b);
    layer6_outputs(7345) <= not a;
    layer6_outputs(7346) <= not (a xor b);
    layer6_outputs(7347) <= not b or a;
    layer6_outputs(7348) <= b and not a;
    layer6_outputs(7349) <= not b or a;
    layer6_outputs(7350) <= a;
    layer6_outputs(7351) <= not b or a;
    layer6_outputs(7352) <= not b or a;
    layer6_outputs(7353) <= not (a and b);
    layer6_outputs(7354) <= b;
    layer6_outputs(7355) <= not (a or b);
    layer6_outputs(7356) <= b and not a;
    layer6_outputs(7357) <= b;
    layer6_outputs(7358) <= not (a xor b);
    layer6_outputs(7359) <= a;
    layer6_outputs(7360) <= '1';
    layer6_outputs(7361) <= not b;
    layer6_outputs(7362) <= a or b;
    layer6_outputs(7363) <= a and b;
    layer6_outputs(7364) <= not (a or b);
    layer6_outputs(7365) <= b;
    layer6_outputs(7366) <= not a;
    layer6_outputs(7367) <= not (a xor b);
    layer6_outputs(7368) <= not a or b;
    layer6_outputs(7369) <= a xor b;
    layer6_outputs(7370) <= a and not b;
    layer6_outputs(7371) <= not (a xor b);
    layer6_outputs(7372) <= not (a and b);
    layer6_outputs(7373) <= b and not a;
    layer6_outputs(7374) <= b and not a;
    layer6_outputs(7375) <= not b;
    layer6_outputs(7376) <= not (a or b);
    layer6_outputs(7377) <= a xor b;
    layer6_outputs(7378) <= a;
    layer6_outputs(7379) <= not (a xor b);
    layer6_outputs(7380) <= not a;
    layer6_outputs(7381) <= a and not b;
    layer6_outputs(7382) <= a or b;
    layer6_outputs(7383) <= a;
    layer6_outputs(7384) <= not a;
    layer6_outputs(7385) <= not (a or b);
    layer6_outputs(7386) <= not a;
    layer6_outputs(7387) <= '1';
    layer6_outputs(7388) <= a and not b;
    layer6_outputs(7389) <= not (a xor b);
    layer6_outputs(7390) <= not b;
    layer6_outputs(7391) <= not a;
    layer6_outputs(7392) <= a;
    layer6_outputs(7393) <= b;
    layer6_outputs(7394) <= a;
    layer6_outputs(7395) <= not (a xor b);
    layer6_outputs(7396) <= not a;
    layer6_outputs(7397) <= b and not a;
    layer6_outputs(7398) <= not (a or b);
    layer6_outputs(7399) <= b and not a;
    layer6_outputs(7400) <= not b or a;
    layer6_outputs(7401) <= a;
    layer6_outputs(7402) <= not (a or b);
    layer6_outputs(7403) <= a or b;
    layer6_outputs(7404) <= not a or b;
    layer6_outputs(7405) <= not a;
    layer6_outputs(7406) <= not (a or b);
    layer6_outputs(7407) <= not b or a;
    layer6_outputs(7408) <= not a or b;
    layer6_outputs(7409) <= b;
    layer6_outputs(7410) <= not (a and b);
    layer6_outputs(7411) <= not (a xor b);
    layer6_outputs(7412) <= not a;
    layer6_outputs(7413) <= not (a or b);
    layer6_outputs(7414) <= a xor b;
    layer6_outputs(7415) <= not a or b;
    layer6_outputs(7416) <= b and not a;
    layer6_outputs(7417) <= b and not a;
    layer6_outputs(7418) <= not a or b;
    layer6_outputs(7419) <= not b or a;
    layer6_outputs(7420) <= not (a or b);
    layer6_outputs(7421) <= a xor b;
    layer6_outputs(7422) <= not b;
    layer6_outputs(7423) <= not (a and b);
    layer6_outputs(7424) <= b and not a;
    layer6_outputs(7425) <= not (a or b);
    layer6_outputs(7426) <= not (a xor b);
    layer6_outputs(7427) <= not a;
    layer6_outputs(7428) <= not (a xor b);
    layer6_outputs(7429) <= not a;
    layer6_outputs(7430) <= b;
    layer6_outputs(7431) <= a and not b;
    layer6_outputs(7432) <= not a;
    layer6_outputs(7433) <= not (a or b);
    layer6_outputs(7434) <= not a;
    layer6_outputs(7435) <= not a;
    layer6_outputs(7436) <= not (a xor b);
    layer6_outputs(7437) <= b;
    layer6_outputs(7438) <= not (a or b);
    layer6_outputs(7439) <= a and not b;
    layer6_outputs(7440) <= b;
    layer6_outputs(7441) <= a xor b;
    layer6_outputs(7442) <= b and not a;
    layer6_outputs(7443) <= b;
    layer6_outputs(7444) <= not a;
    layer6_outputs(7445) <= not (a and b);
    layer6_outputs(7446) <= a xor b;
    layer6_outputs(7447) <= not a;
    layer6_outputs(7448) <= not a or b;
    layer6_outputs(7449) <= not b;
    layer6_outputs(7450) <= not (a or b);
    layer6_outputs(7451) <= b;
    layer6_outputs(7452) <= not (a xor b);
    layer6_outputs(7453) <= b;
    layer6_outputs(7454) <= not a;
    layer6_outputs(7455) <= not (a and b);
    layer6_outputs(7456) <= a;
    layer6_outputs(7457) <= a and b;
    layer6_outputs(7458) <= not b;
    layer6_outputs(7459) <= a or b;
    layer6_outputs(7460) <= not (a and b);
    layer6_outputs(7461) <= not a or b;
    layer6_outputs(7462) <= not a or b;
    layer6_outputs(7463) <= b;
    layer6_outputs(7464) <= b;
    layer6_outputs(7465) <= not a;
    layer6_outputs(7466) <= not (a xor b);
    layer6_outputs(7467) <= not (a and b);
    layer6_outputs(7468) <= b;
    layer6_outputs(7469) <= not (a xor b);
    layer6_outputs(7470) <= not (a xor b);
    layer6_outputs(7471) <= not (a or b);
    layer6_outputs(7472) <= not b;
    layer6_outputs(7473) <= b and not a;
    layer6_outputs(7474) <= a and not b;
    layer6_outputs(7475) <= not b;
    layer6_outputs(7476) <= not (a xor b);
    layer6_outputs(7477) <= not a;
    layer6_outputs(7478) <= b;
    layer6_outputs(7479) <= not a;
    layer6_outputs(7480) <= b;
    layer6_outputs(7481) <= not (a or b);
    layer6_outputs(7482) <= b;
    layer6_outputs(7483) <= not a;
    layer6_outputs(7484) <= not a;
    layer6_outputs(7485) <= not (a xor b);
    layer6_outputs(7486) <= b;
    layer6_outputs(7487) <= a;
    layer6_outputs(7488) <= a;
    layer6_outputs(7489) <= b;
    layer6_outputs(7490) <= a or b;
    layer6_outputs(7491) <= not (a or b);
    layer6_outputs(7492) <= not a;
    layer6_outputs(7493) <= not (a xor b);
    layer6_outputs(7494) <= not (a xor b);
    layer6_outputs(7495) <= not a;
    layer6_outputs(7496) <= a xor b;
    layer6_outputs(7497) <= not (a xor b);
    layer6_outputs(7498) <= b and not a;
    layer6_outputs(7499) <= a and not b;
    layer6_outputs(7500) <= a and not b;
    layer6_outputs(7501) <= not a;
    layer6_outputs(7502) <= b;
    layer6_outputs(7503) <= not (a or b);
    layer6_outputs(7504) <= not a;
    layer6_outputs(7505) <= not (a and b);
    layer6_outputs(7506) <= a;
    layer6_outputs(7507) <= not b or a;
    layer6_outputs(7508) <= b;
    layer6_outputs(7509) <= b and not a;
    layer6_outputs(7510) <= not b;
    layer6_outputs(7511) <= a;
    layer6_outputs(7512) <= not a or b;
    layer6_outputs(7513) <= not a;
    layer6_outputs(7514) <= not b;
    layer6_outputs(7515) <= not a;
    layer6_outputs(7516) <= b;
    layer6_outputs(7517) <= not a;
    layer6_outputs(7518) <= not (a xor b);
    layer6_outputs(7519) <= b;
    layer6_outputs(7520) <= b and not a;
    layer6_outputs(7521) <= not b;
    layer6_outputs(7522) <= not b;
    layer6_outputs(7523) <= not a;
    layer6_outputs(7524) <= not (a xor b);
    layer6_outputs(7525) <= not (a xor b);
    layer6_outputs(7526) <= not b;
    layer6_outputs(7527) <= b and not a;
    layer6_outputs(7528) <= not a or b;
    layer6_outputs(7529) <= not b;
    layer6_outputs(7530) <= b;
    layer6_outputs(7531) <= not (a or b);
    layer6_outputs(7532) <= not a;
    layer6_outputs(7533) <= a and not b;
    layer6_outputs(7534) <= b;
    layer6_outputs(7535) <= not a;
    layer6_outputs(7536) <= not (a xor b);
    layer6_outputs(7537) <= not (a xor b);
    layer6_outputs(7538) <= not a;
    layer6_outputs(7539) <= not a;
    layer6_outputs(7540) <= not b;
    layer6_outputs(7541) <= a and b;
    layer6_outputs(7542) <= a and b;
    layer6_outputs(7543) <= not a;
    layer6_outputs(7544) <= not (a and b);
    layer6_outputs(7545) <= a;
    layer6_outputs(7546) <= not b;
    layer6_outputs(7547) <= not (a xor b);
    layer6_outputs(7548) <= not a or b;
    layer6_outputs(7549) <= a xor b;
    layer6_outputs(7550) <= a xor b;
    layer6_outputs(7551) <= a xor b;
    layer6_outputs(7552) <= a or b;
    layer6_outputs(7553) <= b;
    layer6_outputs(7554) <= a;
    layer6_outputs(7555) <= not (a or b);
    layer6_outputs(7556) <= not b;
    layer6_outputs(7557) <= not a;
    layer6_outputs(7558) <= not a;
    layer6_outputs(7559) <= a or b;
    layer6_outputs(7560) <= not (a or b);
    layer6_outputs(7561) <= not a;
    layer6_outputs(7562) <= not (a or b);
    layer6_outputs(7563) <= not (a and b);
    layer6_outputs(7564) <= a xor b;
    layer6_outputs(7565) <= not (a xor b);
    layer6_outputs(7566) <= not a;
    layer6_outputs(7567) <= not b or a;
    layer6_outputs(7568) <= not (a xor b);
    layer6_outputs(7569) <= '0';
    layer6_outputs(7570) <= a and b;
    layer6_outputs(7571) <= not (a xor b);
    layer6_outputs(7572) <= b and not a;
    layer6_outputs(7573) <= a xor b;
    layer6_outputs(7574) <= not b;
    layer6_outputs(7575) <= not (a xor b);
    layer6_outputs(7576) <= not (a or b);
    layer6_outputs(7577) <= not b;
    layer6_outputs(7578) <= not (a xor b);
    layer6_outputs(7579) <= a xor b;
    layer6_outputs(7580) <= b;
    layer6_outputs(7581) <= not b;
    layer6_outputs(7582) <= not (a xor b);
    layer6_outputs(7583) <= b and not a;
    layer6_outputs(7584) <= a;
    layer6_outputs(7585) <= a xor b;
    layer6_outputs(7586) <= a or b;
    layer6_outputs(7587) <= not b;
    layer6_outputs(7588) <= not a;
    layer6_outputs(7589) <= not a;
    layer6_outputs(7590) <= not a or b;
    layer6_outputs(7591) <= a or b;
    layer6_outputs(7592) <= not b;
    layer6_outputs(7593) <= a and not b;
    layer6_outputs(7594) <= a;
    layer6_outputs(7595) <= a xor b;
    layer6_outputs(7596) <= a and not b;
    layer6_outputs(7597) <= not b or a;
    layer6_outputs(7598) <= not a;
    layer6_outputs(7599) <= not b or a;
    layer6_outputs(7600) <= not b;
    layer6_outputs(7601) <= not b or a;
    layer6_outputs(7602) <= a;
    layer6_outputs(7603) <= not b;
    layer6_outputs(7604) <= a xor b;
    layer6_outputs(7605) <= not (a or b);
    layer6_outputs(7606) <= b;
    layer6_outputs(7607) <= not b;
    layer6_outputs(7608) <= a and not b;
    layer6_outputs(7609) <= b and not a;
    layer6_outputs(7610) <= not (a and b);
    layer6_outputs(7611) <= a and b;
    layer6_outputs(7612) <= not (a and b);
    layer6_outputs(7613) <= not a or b;
    layer6_outputs(7614) <= a xor b;
    layer6_outputs(7615) <= not b;
    layer6_outputs(7616) <= not a;
    layer6_outputs(7617) <= b and not a;
    layer6_outputs(7618) <= b;
    layer6_outputs(7619) <= not (a xor b);
    layer6_outputs(7620) <= a;
    layer6_outputs(7621) <= not (a and b);
    layer6_outputs(7622) <= a xor b;
    layer6_outputs(7623) <= b;
    layer6_outputs(7624) <= not b;
    layer6_outputs(7625) <= '0';
    layer6_outputs(7626) <= b;
    layer6_outputs(7627) <= not a;
    layer6_outputs(7628) <= not a;
    layer6_outputs(7629) <= not b;
    layer6_outputs(7630) <= a and b;
    layer6_outputs(7631) <= not a;
    layer6_outputs(7632) <= not b;
    layer6_outputs(7633) <= a xor b;
    layer6_outputs(7634) <= a;
    layer6_outputs(7635) <= not a;
    layer6_outputs(7636) <= a xor b;
    layer6_outputs(7637) <= b;
    layer6_outputs(7638) <= a;
    layer6_outputs(7639) <= not a or b;
    layer6_outputs(7640) <= a and not b;
    layer6_outputs(7641) <= b;
    layer6_outputs(7642) <= not (a xor b);
    layer6_outputs(7643) <= not a or b;
    layer6_outputs(7644) <= a or b;
    layer6_outputs(7645) <= not b or a;
    layer6_outputs(7646) <= not b;
    layer6_outputs(7647) <= a;
    layer6_outputs(7648) <= not a;
    layer6_outputs(7649) <= b;
    layer6_outputs(7650) <= a xor b;
    layer6_outputs(7651) <= not a;
    layer6_outputs(7652) <= not b;
    layer6_outputs(7653) <= not b or a;
    layer6_outputs(7654) <= not (a xor b);
    layer6_outputs(7655) <= '1';
    layer6_outputs(7656) <= b and not a;
    layer6_outputs(7657) <= a and not b;
    layer6_outputs(7658) <= not (a xor b);
    layer6_outputs(7659) <= b;
    layer6_outputs(7660) <= not b;
    layer6_outputs(7661) <= not b or a;
    layer6_outputs(7662) <= not a;
    layer6_outputs(7663) <= b;
    layer6_outputs(7664) <= b;
    layer6_outputs(7665) <= not a;
    layer6_outputs(7666) <= not (a xor b);
    layer6_outputs(7667) <= b and not a;
    layer6_outputs(7668) <= not (a xor b);
    layer6_outputs(7669) <= not b;
    layer6_outputs(7670) <= a or b;
    layer6_outputs(7671) <= not a;
    layer6_outputs(7672) <= not a;
    layer6_outputs(7673) <= not a;
    layer6_outputs(7674) <= a xor b;
    layer6_outputs(7675) <= b;
    layer6_outputs(7676) <= a and b;
    layer6_outputs(7677) <= not b;
    layer6_outputs(7678) <= not (a xor b);
    layer6_outputs(7679) <= not b;
    layer6_outputs(7680) <= b;
    layer6_outputs(7681) <= b;
    layer6_outputs(7682) <= a xor b;
    layer6_outputs(7683) <= a xor b;
    layer6_outputs(7684) <= b;
    layer6_outputs(7685) <= not b;
    layer6_outputs(7686) <= not b;
    layer6_outputs(7687) <= a or b;
    layer6_outputs(7688) <= not a;
    layer6_outputs(7689) <= a;
    layer6_outputs(7690) <= not a;
    layer6_outputs(7691) <= not a;
    layer6_outputs(7692) <= a;
    layer6_outputs(7693) <= a and not b;
    layer6_outputs(7694) <= not a;
    layer6_outputs(7695) <= a;
    layer6_outputs(7696) <= a or b;
    layer6_outputs(7697) <= not (a xor b);
    layer6_outputs(7698) <= not a;
    layer6_outputs(7699) <= not b;
    layer6_outputs(7700) <= b;
    layer6_outputs(7701) <= a xor b;
    layer6_outputs(7702) <= not a;
    layer6_outputs(7703) <= a;
    layer6_outputs(7704) <= not a;
    layer6_outputs(7705) <= a and not b;
    layer6_outputs(7706) <= a xor b;
    layer6_outputs(7707) <= a;
    layer6_outputs(7708) <= b;
    layer6_outputs(7709) <= a xor b;
    layer6_outputs(7710) <= not a or b;
    layer6_outputs(7711) <= a and b;
    layer6_outputs(7712) <= not (a and b);
    layer6_outputs(7713) <= not (a xor b);
    layer6_outputs(7714) <= not a;
    layer6_outputs(7715) <= b and not a;
    layer6_outputs(7716) <= not (a or b);
    layer6_outputs(7717) <= not a;
    layer6_outputs(7718) <= not (a xor b);
    layer6_outputs(7719) <= a xor b;
    layer6_outputs(7720) <= a and not b;
    layer6_outputs(7721) <= not (a or b);
    layer6_outputs(7722) <= a xor b;
    layer6_outputs(7723) <= not (a or b);
    layer6_outputs(7724) <= not b;
    layer6_outputs(7725) <= not (a and b);
    layer6_outputs(7726) <= a;
    layer6_outputs(7727) <= a and not b;
    layer6_outputs(7728) <= not a;
    layer6_outputs(7729) <= b;
    layer6_outputs(7730) <= a;
    layer6_outputs(7731) <= not a or b;
    layer6_outputs(7732) <= not (a and b);
    layer6_outputs(7733) <= b;
    layer6_outputs(7734) <= a xor b;
    layer6_outputs(7735) <= a;
    layer6_outputs(7736) <= not a or b;
    layer6_outputs(7737) <= b;
    layer6_outputs(7738) <= not b;
    layer6_outputs(7739) <= not a;
    layer6_outputs(7740) <= b;
    layer6_outputs(7741) <= not a;
    layer6_outputs(7742) <= not b or a;
    layer6_outputs(7743) <= not b;
    layer6_outputs(7744) <= not b;
    layer6_outputs(7745) <= a xor b;
    layer6_outputs(7746) <= not a;
    layer6_outputs(7747) <= a and b;
    layer6_outputs(7748) <= b and not a;
    layer6_outputs(7749) <= b;
    layer6_outputs(7750) <= not b;
    layer6_outputs(7751) <= a and not b;
    layer6_outputs(7752) <= not b or a;
    layer6_outputs(7753) <= b;
    layer6_outputs(7754) <= not a;
    layer6_outputs(7755) <= a;
    layer6_outputs(7756) <= not a;
    layer6_outputs(7757) <= a xor b;
    layer6_outputs(7758) <= not b;
    layer6_outputs(7759) <= a;
    layer6_outputs(7760) <= '0';
    layer6_outputs(7761) <= a;
    layer6_outputs(7762) <= not b or a;
    layer6_outputs(7763) <= b;
    layer6_outputs(7764) <= not b;
    layer6_outputs(7765) <= not a;
    layer6_outputs(7766) <= not a;
    layer6_outputs(7767) <= not b;
    layer6_outputs(7768) <= not a;
    layer6_outputs(7769) <= not b or a;
    layer6_outputs(7770) <= not a;
    layer6_outputs(7771) <= not a;
    layer6_outputs(7772) <= not (a xor b);
    layer6_outputs(7773) <= not b;
    layer6_outputs(7774) <= '0';
    layer6_outputs(7775) <= a and b;
    layer6_outputs(7776) <= not a;
    layer6_outputs(7777) <= '1';
    layer6_outputs(7778) <= not b;
    layer6_outputs(7779) <= a xor b;
    layer6_outputs(7780) <= b;
    layer6_outputs(7781) <= not b or a;
    layer6_outputs(7782) <= b and not a;
    layer6_outputs(7783) <= a;
    layer6_outputs(7784) <= not a;
    layer6_outputs(7785) <= a and not b;
    layer6_outputs(7786) <= a or b;
    layer6_outputs(7787) <= a xor b;
    layer6_outputs(7788) <= b and not a;
    layer6_outputs(7789) <= not (a or b);
    layer6_outputs(7790) <= a or b;
    layer6_outputs(7791) <= '0';
    layer6_outputs(7792) <= a xor b;
    layer6_outputs(7793) <= not (a and b);
    layer6_outputs(7794) <= not a or b;
    layer6_outputs(7795) <= not a or b;
    layer6_outputs(7796) <= not b;
    layer6_outputs(7797) <= not b;
    layer6_outputs(7798) <= not b or a;
    layer6_outputs(7799) <= not (a xor b);
    layer6_outputs(7800) <= a and not b;
    layer6_outputs(7801) <= not (a xor b);
    layer6_outputs(7802) <= a;
    layer6_outputs(7803) <= not a;
    layer6_outputs(7804) <= a;
    layer6_outputs(7805) <= b;
    layer6_outputs(7806) <= not b or a;
    layer6_outputs(7807) <= not (a or b);
    layer6_outputs(7808) <= b;
    layer6_outputs(7809) <= a;
    layer6_outputs(7810) <= not (a xor b);
    layer6_outputs(7811) <= a;
    layer6_outputs(7812) <= not a;
    layer6_outputs(7813) <= not b or a;
    layer6_outputs(7814) <= not (a or b);
    layer6_outputs(7815) <= not b;
    layer6_outputs(7816) <= not (a and b);
    layer6_outputs(7817) <= not (a or b);
    layer6_outputs(7818) <= not a;
    layer6_outputs(7819) <= b;
    layer6_outputs(7820) <= a;
    layer6_outputs(7821) <= not a;
    layer6_outputs(7822) <= not (a or b);
    layer6_outputs(7823) <= not b;
    layer6_outputs(7824) <= a;
    layer6_outputs(7825) <= not b;
    layer6_outputs(7826) <= not b;
    layer6_outputs(7827) <= b;
    layer6_outputs(7828) <= a xor b;
    layer6_outputs(7829) <= not (a xor b);
    layer6_outputs(7830) <= not a;
    layer6_outputs(7831) <= not b or a;
    layer6_outputs(7832) <= not a;
    layer6_outputs(7833) <= not b;
    layer6_outputs(7834) <= a xor b;
    layer6_outputs(7835) <= not (a xor b);
    layer6_outputs(7836) <= not b or a;
    layer6_outputs(7837) <= b;
    layer6_outputs(7838) <= a and not b;
    layer6_outputs(7839) <= a xor b;
    layer6_outputs(7840) <= a or b;
    layer6_outputs(7841) <= not (a and b);
    layer6_outputs(7842) <= not (a xor b);
    layer6_outputs(7843) <= not b;
    layer6_outputs(7844) <= '1';
    layer6_outputs(7845) <= a;
    layer6_outputs(7846) <= a xor b;
    layer6_outputs(7847) <= not a;
    layer6_outputs(7848) <= '1';
    layer6_outputs(7849) <= a xor b;
    layer6_outputs(7850) <= not a;
    layer6_outputs(7851) <= not a;
    layer6_outputs(7852) <= not (a or b);
    layer6_outputs(7853) <= not b;
    layer6_outputs(7854) <= a xor b;
    layer6_outputs(7855) <= a or b;
    layer6_outputs(7856) <= a or b;
    layer6_outputs(7857) <= not (a xor b);
    layer6_outputs(7858) <= not b or a;
    layer6_outputs(7859) <= a;
    layer6_outputs(7860) <= not b or a;
    layer6_outputs(7861) <= b;
    layer6_outputs(7862) <= b;
    layer6_outputs(7863) <= not a;
    layer6_outputs(7864) <= not a;
    layer6_outputs(7865) <= not (a xor b);
    layer6_outputs(7866) <= not a or b;
    layer6_outputs(7867) <= b and not a;
    layer6_outputs(7868) <= b;
    layer6_outputs(7869) <= a;
    layer6_outputs(7870) <= not b or a;
    layer6_outputs(7871) <= not b;
    layer6_outputs(7872) <= not a;
    layer6_outputs(7873) <= not (a or b);
    layer6_outputs(7874) <= not b;
    layer6_outputs(7875) <= a;
    layer6_outputs(7876) <= b;
    layer6_outputs(7877) <= b and not a;
    layer6_outputs(7878) <= a;
    layer6_outputs(7879) <= b;
    layer6_outputs(7880) <= not a;
    layer6_outputs(7881) <= not (a xor b);
    layer6_outputs(7882) <= not (a or b);
    layer6_outputs(7883) <= b and not a;
    layer6_outputs(7884) <= a;
    layer6_outputs(7885) <= not b;
    layer6_outputs(7886) <= a or b;
    layer6_outputs(7887) <= not a;
    layer6_outputs(7888) <= a xor b;
    layer6_outputs(7889) <= a;
    layer6_outputs(7890) <= a;
    layer6_outputs(7891) <= not (a and b);
    layer6_outputs(7892) <= a;
    layer6_outputs(7893) <= not (a and b);
    layer6_outputs(7894) <= not b;
    layer6_outputs(7895) <= not (a or b);
    layer6_outputs(7896) <= a;
    layer6_outputs(7897) <= a;
    layer6_outputs(7898) <= not a;
    layer6_outputs(7899) <= not b;
    layer6_outputs(7900) <= a;
    layer6_outputs(7901) <= b and not a;
    layer6_outputs(7902) <= a;
    layer6_outputs(7903) <= not a or b;
    layer6_outputs(7904) <= not (a and b);
    layer6_outputs(7905) <= b;
    layer6_outputs(7906) <= not a;
    layer6_outputs(7907) <= not (a and b);
    layer6_outputs(7908) <= a xor b;
    layer6_outputs(7909) <= not (a xor b);
    layer6_outputs(7910) <= a xor b;
    layer6_outputs(7911) <= b and not a;
    layer6_outputs(7912) <= a xor b;
    layer6_outputs(7913) <= not (a xor b);
    layer6_outputs(7914) <= a and b;
    layer6_outputs(7915) <= a and not b;
    layer6_outputs(7916) <= not (a xor b);
    layer6_outputs(7917) <= not a;
    layer6_outputs(7918) <= b and not a;
    layer6_outputs(7919) <= not (a xor b);
    layer6_outputs(7920) <= not (a xor b);
    layer6_outputs(7921) <= not b or a;
    layer6_outputs(7922) <= a xor b;
    layer6_outputs(7923) <= a and not b;
    layer6_outputs(7924) <= not b;
    layer6_outputs(7925) <= not b;
    layer6_outputs(7926) <= b and not a;
    layer6_outputs(7927) <= not (a and b);
    layer6_outputs(7928) <= not b or a;
    layer6_outputs(7929) <= not (a xor b);
    layer6_outputs(7930) <= a and not b;
    layer6_outputs(7931) <= not b;
    layer6_outputs(7932) <= not (a and b);
    layer6_outputs(7933) <= not b;
    layer6_outputs(7934) <= a xor b;
    layer6_outputs(7935) <= a and not b;
    layer6_outputs(7936) <= not (a xor b);
    layer6_outputs(7937) <= a;
    layer6_outputs(7938) <= b and not a;
    layer6_outputs(7939) <= b;
    layer6_outputs(7940) <= not b;
    layer6_outputs(7941) <= a xor b;
    layer6_outputs(7942) <= a;
    layer6_outputs(7943) <= not b or a;
    layer6_outputs(7944) <= a;
    layer6_outputs(7945) <= b;
    layer6_outputs(7946) <= not a;
    layer6_outputs(7947) <= b and not a;
    layer6_outputs(7948) <= not a;
    layer6_outputs(7949) <= a;
    layer6_outputs(7950) <= not b or a;
    layer6_outputs(7951) <= not b or a;
    layer6_outputs(7952) <= a xor b;
    layer6_outputs(7953) <= not a;
    layer6_outputs(7954) <= not a;
    layer6_outputs(7955) <= a xor b;
    layer6_outputs(7956) <= b and not a;
    layer6_outputs(7957) <= a xor b;
    layer6_outputs(7958) <= not (a xor b);
    layer6_outputs(7959) <= '1';
    layer6_outputs(7960) <= b;
    layer6_outputs(7961) <= not (a xor b);
    layer6_outputs(7962) <= a and b;
    layer6_outputs(7963) <= a or b;
    layer6_outputs(7964) <= a and b;
    layer6_outputs(7965) <= b and not a;
    layer6_outputs(7966) <= b;
    layer6_outputs(7967) <= not a;
    layer6_outputs(7968) <= not b;
    layer6_outputs(7969) <= not a;
    layer6_outputs(7970) <= not (a or b);
    layer6_outputs(7971) <= a;
    layer6_outputs(7972) <= a and b;
    layer6_outputs(7973) <= not a or b;
    layer6_outputs(7974) <= not a or b;
    layer6_outputs(7975) <= not (a or b);
    layer6_outputs(7976) <= not (a xor b);
    layer6_outputs(7977) <= not b or a;
    layer6_outputs(7978) <= not b;
    layer6_outputs(7979) <= b and not a;
    layer6_outputs(7980) <= a xor b;
    layer6_outputs(7981) <= not b;
    layer6_outputs(7982) <= not a or b;
    layer6_outputs(7983) <= not b;
    layer6_outputs(7984) <= not b;
    layer6_outputs(7985) <= not b or a;
    layer6_outputs(7986) <= a;
    layer6_outputs(7987) <= not b;
    layer6_outputs(7988) <= a;
    layer6_outputs(7989) <= a;
    layer6_outputs(7990) <= a;
    layer6_outputs(7991) <= not b;
    layer6_outputs(7992) <= not (a or b);
    layer6_outputs(7993) <= b;
    layer6_outputs(7994) <= a;
    layer6_outputs(7995) <= not (a or b);
    layer6_outputs(7996) <= a;
    layer6_outputs(7997) <= not b;
    layer6_outputs(7998) <= a;
    layer6_outputs(7999) <= a;
    layer6_outputs(8000) <= b;
    layer6_outputs(8001) <= not b or a;
    layer6_outputs(8002) <= not b or a;
    layer6_outputs(8003) <= not a;
    layer6_outputs(8004) <= not b or a;
    layer6_outputs(8005) <= not b;
    layer6_outputs(8006) <= not a;
    layer6_outputs(8007) <= b;
    layer6_outputs(8008) <= not b;
    layer6_outputs(8009) <= not b or a;
    layer6_outputs(8010) <= a;
    layer6_outputs(8011) <= not a or b;
    layer6_outputs(8012) <= not (a xor b);
    layer6_outputs(8013) <= a or b;
    layer6_outputs(8014) <= a and not b;
    layer6_outputs(8015) <= a and not b;
    layer6_outputs(8016) <= not (a and b);
    layer6_outputs(8017) <= a xor b;
    layer6_outputs(8018) <= not a;
    layer6_outputs(8019) <= a;
    layer6_outputs(8020) <= a and b;
    layer6_outputs(8021) <= not a or b;
    layer6_outputs(8022) <= not (a or b);
    layer6_outputs(8023) <= a;
    layer6_outputs(8024) <= a;
    layer6_outputs(8025) <= not (a or b);
    layer6_outputs(8026) <= a xor b;
    layer6_outputs(8027) <= a and not b;
    layer6_outputs(8028) <= a;
    layer6_outputs(8029) <= '1';
    layer6_outputs(8030) <= not (a xor b);
    layer6_outputs(8031) <= a and not b;
    layer6_outputs(8032) <= not b;
    layer6_outputs(8033) <= not (a xor b);
    layer6_outputs(8034) <= not (a and b);
    layer6_outputs(8035) <= not a;
    layer6_outputs(8036) <= not b or a;
    layer6_outputs(8037) <= not b or a;
    layer6_outputs(8038) <= not (a xor b);
    layer6_outputs(8039) <= not (a xor b);
    layer6_outputs(8040) <= not a or b;
    layer6_outputs(8041) <= not a;
    layer6_outputs(8042) <= a or b;
    layer6_outputs(8043) <= not b;
    layer6_outputs(8044) <= b;
    layer6_outputs(8045) <= a xor b;
    layer6_outputs(8046) <= not a;
    layer6_outputs(8047) <= not (a and b);
    layer6_outputs(8048) <= a xor b;
    layer6_outputs(8049) <= not b;
    layer6_outputs(8050) <= not (a or b);
    layer6_outputs(8051) <= not (a or b);
    layer6_outputs(8052) <= not (a xor b);
    layer6_outputs(8053) <= a or b;
    layer6_outputs(8054) <= not b;
    layer6_outputs(8055) <= a;
    layer6_outputs(8056) <= a xor b;
    layer6_outputs(8057) <= a;
    layer6_outputs(8058) <= a;
    layer6_outputs(8059) <= not a;
    layer6_outputs(8060) <= a and not b;
    layer6_outputs(8061) <= not b or a;
    layer6_outputs(8062) <= b and not a;
    layer6_outputs(8063) <= '1';
    layer6_outputs(8064) <= b;
    layer6_outputs(8065) <= not a;
    layer6_outputs(8066) <= not b;
    layer6_outputs(8067) <= a and b;
    layer6_outputs(8068) <= b;
    layer6_outputs(8069) <= not a;
    layer6_outputs(8070) <= b;
    layer6_outputs(8071) <= not (a and b);
    layer6_outputs(8072) <= a xor b;
    layer6_outputs(8073) <= not a;
    layer6_outputs(8074) <= a or b;
    layer6_outputs(8075) <= not a;
    layer6_outputs(8076) <= not (a and b);
    layer6_outputs(8077) <= not b or a;
    layer6_outputs(8078) <= a and not b;
    layer6_outputs(8079) <= not b;
    layer6_outputs(8080) <= not a;
    layer6_outputs(8081) <= a xor b;
    layer6_outputs(8082) <= not b or a;
    layer6_outputs(8083) <= a;
    layer6_outputs(8084) <= a and b;
    layer6_outputs(8085) <= not (a and b);
    layer6_outputs(8086) <= b;
    layer6_outputs(8087) <= a xor b;
    layer6_outputs(8088) <= not b;
    layer6_outputs(8089) <= not b or a;
    layer6_outputs(8090) <= b;
    layer6_outputs(8091) <= not (a xor b);
    layer6_outputs(8092) <= not (a xor b);
    layer6_outputs(8093) <= b;
    layer6_outputs(8094) <= not (a xor b);
    layer6_outputs(8095) <= a and not b;
    layer6_outputs(8096) <= b and not a;
    layer6_outputs(8097) <= b;
    layer6_outputs(8098) <= not a;
    layer6_outputs(8099) <= b;
    layer6_outputs(8100) <= a;
    layer6_outputs(8101) <= not a or b;
    layer6_outputs(8102) <= not a or b;
    layer6_outputs(8103) <= not a or b;
    layer6_outputs(8104) <= b;
    layer6_outputs(8105) <= not b or a;
    layer6_outputs(8106) <= not b or a;
    layer6_outputs(8107) <= not (a and b);
    layer6_outputs(8108) <= not (a and b);
    layer6_outputs(8109) <= a and not b;
    layer6_outputs(8110) <= b and not a;
    layer6_outputs(8111) <= a;
    layer6_outputs(8112) <= not b or a;
    layer6_outputs(8113) <= not (a xor b);
    layer6_outputs(8114) <= not a;
    layer6_outputs(8115) <= not b;
    layer6_outputs(8116) <= a;
    layer6_outputs(8117) <= a xor b;
    layer6_outputs(8118) <= not (a xor b);
    layer6_outputs(8119) <= not (a or b);
    layer6_outputs(8120) <= '1';
    layer6_outputs(8121) <= not b;
    layer6_outputs(8122) <= not (a and b);
    layer6_outputs(8123) <= a;
    layer6_outputs(8124) <= a;
    layer6_outputs(8125) <= a xor b;
    layer6_outputs(8126) <= not b;
    layer6_outputs(8127) <= not b;
    layer6_outputs(8128) <= not b;
    layer6_outputs(8129) <= a xor b;
    layer6_outputs(8130) <= a xor b;
    layer6_outputs(8131) <= not (a xor b);
    layer6_outputs(8132) <= not (a and b);
    layer6_outputs(8133) <= a and b;
    layer6_outputs(8134) <= a and not b;
    layer6_outputs(8135) <= b;
    layer6_outputs(8136) <= not b;
    layer6_outputs(8137) <= not (a xor b);
    layer6_outputs(8138) <= b;
    layer6_outputs(8139) <= not b;
    layer6_outputs(8140) <= not a;
    layer6_outputs(8141) <= a or b;
    layer6_outputs(8142) <= a;
    layer6_outputs(8143) <= not (a and b);
    layer6_outputs(8144) <= not a;
    layer6_outputs(8145) <= not (a or b);
    layer6_outputs(8146) <= a;
    layer6_outputs(8147) <= '1';
    layer6_outputs(8148) <= not (a xor b);
    layer6_outputs(8149) <= not b or a;
    layer6_outputs(8150) <= not a;
    layer6_outputs(8151) <= a xor b;
    layer6_outputs(8152) <= b;
    layer6_outputs(8153) <= not b;
    layer6_outputs(8154) <= not b;
    layer6_outputs(8155) <= b;
    layer6_outputs(8156) <= b;
    layer6_outputs(8157) <= not a;
    layer6_outputs(8158) <= not (a xor b);
    layer6_outputs(8159) <= not (a xor b);
    layer6_outputs(8160) <= a and not b;
    layer6_outputs(8161) <= not a;
    layer6_outputs(8162) <= a and not b;
    layer6_outputs(8163) <= not (a xor b);
    layer6_outputs(8164) <= not (a and b);
    layer6_outputs(8165) <= not b;
    layer6_outputs(8166) <= b and not a;
    layer6_outputs(8167) <= not b;
    layer6_outputs(8168) <= not b or a;
    layer6_outputs(8169) <= b;
    layer6_outputs(8170) <= not b or a;
    layer6_outputs(8171) <= not a;
    layer6_outputs(8172) <= a;
    layer6_outputs(8173) <= not b;
    layer6_outputs(8174) <= a xor b;
    layer6_outputs(8175) <= a or b;
    layer6_outputs(8176) <= b and not a;
    layer6_outputs(8177) <= not (a and b);
    layer6_outputs(8178) <= not b or a;
    layer6_outputs(8179) <= not (a xor b);
    layer6_outputs(8180) <= not (a or b);
    layer6_outputs(8181) <= not a;
    layer6_outputs(8182) <= not (a xor b);
    layer6_outputs(8183) <= a;
    layer6_outputs(8184) <= b;
    layer6_outputs(8185) <= not b;
    layer6_outputs(8186) <= b;
    layer6_outputs(8187) <= not b;
    layer6_outputs(8188) <= not a;
    layer6_outputs(8189) <= b and not a;
    layer6_outputs(8190) <= not b;
    layer6_outputs(8191) <= not b;
    layer6_outputs(8192) <= not b;
    layer6_outputs(8193) <= '1';
    layer6_outputs(8194) <= b;
    layer6_outputs(8195) <= a xor b;
    layer6_outputs(8196) <= b and not a;
    layer6_outputs(8197) <= not a;
    layer6_outputs(8198) <= a or b;
    layer6_outputs(8199) <= b;
    layer6_outputs(8200) <= not (a xor b);
    layer6_outputs(8201) <= b;
    layer6_outputs(8202) <= not b;
    layer6_outputs(8203) <= not b;
    layer6_outputs(8204) <= a;
    layer6_outputs(8205) <= a xor b;
    layer6_outputs(8206) <= not a;
    layer6_outputs(8207) <= a;
    layer6_outputs(8208) <= not b;
    layer6_outputs(8209) <= not (a or b);
    layer6_outputs(8210) <= b and not a;
    layer6_outputs(8211) <= not a;
    layer6_outputs(8212) <= not a;
    layer6_outputs(8213) <= a;
    layer6_outputs(8214) <= not (a xor b);
    layer6_outputs(8215) <= b and not a;
    layer6_outputs(8216) <= a or b;
    layer6_outputs(8217) <= not a;
    layer6_outputs(8218) <= not b or a;
    layer6_outputs(8219) <= not (a xor b);
    layer6_outputs(8220) <= a xor b;
    layer6_outputs(8221) <= a and b;
    layer6_outputs(8222) <= a xor b;
    layer6_outputs(8223) <= not (a xor b);
    layer6_outputs(8224) <= not a;
    layer6_outputs(8225) <= not b;
    layer6_outputs(8226) <= a and not b;
    layer6_outputs(8227) <= not b or a;
    layer6_outputs(8228) <= not b or a;
    layer6_outputs(8229) <= not (a xor b);
    layer6_outputs(8230) <= a;
    layer6_outputs(8231) <= not a or b;
    layer6_outputs(8232) <= not b or a;
    layer6_outputs(8233) <= not a or b;
    layer6_outputs(8234) <= a and not b;
    layer6_outputs(8235) <= a and not b;
    layer6_outputs(8236) <= not a;
    layer6_outputs(8237) <= not b;
    layer6_outputs(8238) <= b;
    layer6_outputs(8239) <= not (a and b);
    layer6_outputs(8240) <= b;
    layer6_outputs(8241) <= not (a xor b);
    layer6_outputs(8242) <= a or b;
    layer6_outputs(8243) <= not b or a;
    layer6_outputs(8244) <= b;
    layer6_outputs(8245) <= a;
    layer6_outputs(8246) <= b;
    layer6_outputs(8247) <= not a;
    layer6_outputs(8248) <= not (a and b);
    layer6_outputs(8249) <= a or b;
    layer6_outputs(8250) <= b;
    layer6_outputs(8251) <= b;
    layer6_outputs(8252) <= not a;
    layer6_outputs(8253) <= a or b;
    layer6_outputs(8254) <= a xor b;
    layer6_outputs(8255) <= not b;
    layer6_outputs(8256) <= a xor b;
    layer6_outputs(8257) <= not (a or b);
    layer6_outputs(8258) <= not (a and b);
    layer6_outputs(8259) <= a and b;
    layer6_outputs(8260) <= b;
    layer6_outputs(8261) <= a;
    layer6_outputs(8262) <= a and not b;
    layer6_outputs(8263) <= b;
    layer6_outputs(8264) <= '0';
    layer6_outputs(8265) <= a;
    layer6_outputs(8266) <= a;
    layer6_outputs(8267) <= not (a and b);
    layer6_outputs(8268) <= a;
    layer6_outputs(8269) <= not a or b;
    layer6_outputs(8270) <= not b or a;
    layer6_outputs(8271) <= a or b;
    layer6_outputs(8272) <= b;
    layer6_outputs(8273) <= not (a xor b);
    layer6_outputs(8274) <= not (a xor b);
    layer6_outputs(8275) <= b;
    layer6_outputs(8276) <= not a;
    layer6_outputs(8277) <= not (a xor b);
    layer6_outputs(8278) <= not b;
    layer6_outputs(8279) <= not a or b;
    layer6_outputs(8280) <= b and not a;
    layer6_outputs(8281) <= not a or b;
    layer6_outputs(8282) <= b;
    layer6_outputs(8283) <= not (a and b);
    layer6_outputs(8284) <= a or b;
    layer6_outputs(8285) <= not a or b;
    layer6_outputs(8286) <= not (a or b);
    layer6_outputs(8287) <= a and not b;
    layer6_outputs(8288) <= not (a and b);
    layer6_outputs(8289) <= a;
    layer6_outputs(8290) <= a xor b;
    layer6_outputs(8291) <= not (a xor b);
    layer6_outputs(8292) <= b;
    layer6_outputs(8293) <= b;
    layer6_outputs(8294) <= not a;
    layer6_outputs(8295) <= not b;
    layer6_outputs(8296) <= not b or a;
    layer6_outputs(8297) <= not (a and b);
    layer6_outputs(8298) <= not a;
    layer6_outputs(8299) <= not (a xor b);
    layer6_outputs(8300) <= not b;
    layer6_outputs(8301) <= a and not b;
    layer6_outputs(8302) <= not (a and b);
    layer6_outputs(8303) <= b;
    layer6_outputs(8304) <= not a;
    layer6_outputs(8305) <= a and b;
    layer6_outputs(8306) <= not b;
    layer6_outputs(8307) <= a;
    layer6_outputs(8308) <= a;
    layer6_outputs(8309) <= not b;
    layer6_outputs(8310) <= b and not a;
    layer6_outputs(8311) <= not (a or b);
    layer6_outputs(8312) <= a xor b;
    layer6_outputs(8313) <= a xor b;
    layer6_outputs(8314) <= not a;
    layer6_outputs(8315) <= not (a or b);
    layer6_outputs(8316) <= not a;
    layer6_outputs(8317) <= not b;
    layer6_outputs(8318) <= not b;
    layer6_outputs(8319) <= a;
    layer6_outputs(8320) <= not (a or b);
    layer6_outputs(8321) <= a and b;
    layer6_outputs(8322) <= a or b;
    layer6_outputs(8323) <= not (a and b);
    layer6_outputs(8324) <= not b or a;
    layer6_outputs(8325) <= not (a xor b);
    layer6_outputs(8326) <= a xor b;
    layer6_outputs(8327) <= not (a or b);
    layer6_outputs(8328) <= a or b;
    layer6_outputs(8329) <= '1';
    layer6_outputs(8330) <= not (a xor b);
    layer6_outputs(8331) <= a;
    layer6_outputs(8332) <= a and b;
    layer6_outputs(8333) <= a;
    layer6_outputs(8334) <= a;
    layer6_outputs(8335) <= a;
    layer6_outputs(8336) <= a or b;
    layer6_outputs(8337) <= not a;
    layer6_outputs(8338) <= not b;
    layer6_outputs(8339) <= not b;
    layer6_outputs(8340) <= b;
    layer6_outputs(8341) <= a and b;
    layer6_outputs(8342) <= not a;
    layer6_outputs(8343) <= a or b;
    layer6_outputs(8344) <= not b or a;
    layer6_outputs(8345) <= a;
    layer6_outputs(8346) <= not a or b;
    layer6_outputs(8347) <= not (a xor b);
    layer6_outputs(8348) <= not b or a;
    layer6_outputs(8349) <= '0';
    layer6_outputs(8350) <= not b;
    layer6_outputs(8351) <= a and b;
    layer6_outputs(8352) <= '1';
    layer6_outputs(8353) <= not a;
    layer6_outputs(8354) <= not a;
    layer6_outputs(8355) <= a;
    layer6_outputs(8356) <= a;
    layer6_outputs(8357) <= not b;
    layer6_outputs(8358) <= not (a xor b);
    layer6_outputs(8359) <= not b;
    layer6_outputs(8360) <= not (a xor b);
    layer6_outputs(8361) <= not (a xor b);
    layer6_outputs(8362) <= a and b;
    layer6_outputs(8363) <= '0';
    layer6_outputs(8364) <= b;
    layer6_outputs(8365) <= not (a and b);
    layer6_outputs(8366) <= b and not a;
    layer6_outputs(8367) <= a and b;
    layer6_outputs(8368) <= not a;
    layer6_outputs(8369) <= not a;
    layer6_outputs(8370) <= a xor b;
    layer6_outputs(8371) <= not (a or b);
    layer6_outputs(8372) <= a;
    layer6_outputs(8373) <= not (a or b);
    layer6_outputs(8374) <= a or b;
    layer6_outputs(8375) <= not (a xor b);
    layer6_outputs(8376) <= a;
    layer6_outputs(8377) <= not b;
    layer6_outputs(8378) <= not b;
    layer6_outputs(8379) <= not a;
    layer6_outputs(8380) <= not a;
    layer6_outputs(8381) <= not a;
    layer6_outputs(8382) <= a and not b;
    layer6_outputs(8383) <= a or b;
    layer6_outputs(8384) <= b;
    layer6_outputs(8385) <= b;
    layer6_outputs(8386) <= a;
    layer6_outputs(8387) <= a and b;
    layer6_outputs(8388) <= not b;
    layer6_outputs(8389) <= not b;
    layer6_outputs(8390) <= a;
    layer6_outputs(8391) <= b;
    layer6_outputs(8392) <= not (a xor b);
    layer6_outputs(8393) <= not b;
    layer6_outputs(8394) <= not a or b;
    layer6_outputs(8395) <= not (a and b);
    layer6_outputs(8396) <= a;
    layer6_outputs(8397) <= a;
    layer6_outputs(8398) <= not (a xor b);
    layer6_outputs(8399) <= not b;
    layer6_outputs(8400) <= a;
    layer6_outputs(8401) <= '0';
    layer6_outputs(8402) <= not (a or b);
    layer6_outputs(8403) <= b;
    layer6_outputs(8404) <= not a;
    layer6_outputs(8405) <= not b;
    layer6_outputs(8406) <= a xor b;
    layer6_outputs(8407) <= a xor b;
    layer6_outputs(8408) <= not (a xor b);
    layer6_outputs(8409) <= not b;
    layer6_outputs(8410) <= not a or b;
    layer6_outputs(8411) <= a;
    layer6_outputs(8412) <= b;
    layer6_outputs(8413) <= not (a or b);
    layer6_outputs(8414) <= a;
    layer6_outputs(8415) <= not a;
    layer6_outputs(8416) <= not a or b;
    layer6_outputs(8417) <= '1';
    layer6_outputs(8418) <= a and not b;
    layer6_outputs(8419) <= a or b;
    layer6_outputs(8420) <= a;
    layer6_outputs(8421) <= a;
    layer6_outputs(8422) <= not (a xor b);
    layer6_outputs(8423) <= not a;
    layer6_outputs(8424) <= not b;
    layer6_outputs(8425) <= b;
    layer6_outputs(8426) <= not a or b;
    layer6_outputs(8427) <= not a;
    layer6_outputs(8428) <= not a;
    layer6_outputs(8429) <= a and b;
    layer6_outputs(8430) <= a and not b;
    layer6_outputs(8431) <= a xor b;
    layer6_outputs(8432) <= not b;
    layer6_outputs(8433) <= a and b;
    layer6_outputs(8434) <= not a;
    layer6_outputs(8435) <= a;
    layer6_outputs(8436) <= b and not a;
    layer6_outputs(8437) <= not (a or b);
    layer6_outputs(8438) <= not (a xor b);
    layer6_outputs(8439) <= a;
    layer6_outputs(8440) <= a xor b;
    layer6_outputs(8441) <= b;
    layer6_outputs(8442) <= not b;
    layer6_outputs(8443) <= b;
    layer6_outputs(8444) <= a or b;
    layer6_outputs(8445) <= not b or a;
    layer6_outputs(8446) <= not b;
    layer6_outputs(8447) <= not b;
    layer6_outputs(8448) <= not b or a;
    layer6_outputs(8449) <= a and b;
    layer6_outputs(8450) <= '0';
    layer6_outputs(8451) <= a;
    layer6_outputs(8452) <= not (a or b);
    layer6_outputs(8453) <= not a;
    layer6_outputs(8454) <= not b or a;
    layer6_outputs(8455) <= not a;
    layer6_outputs(8456) <= b;
    layer6_outputs(8457) <= not b or a;
    layer6_outputs(8458) <= not a;
    layer6_outputs(8459) <= not (a or b);
    layer6_outputs(8460) <= not (a xor b);
    layer6_outputs(8461) <= b;
    layer6_outputs(8462) <= a and not b;
    layer6_outputs(8463) <= not (a and b);
    layer6_outputs(8464) <= not (a and b);
    layer6_outputs(8465) <= a;
    layer6_outputs(8466) <= a and b;
    layer6_outputs(8467) <= not b;
    layer6_outputs(8468) <= b;
    layer6_outputs(8469) <= a and b;
    layer6_outputs(8470) <= a xor b;
    layer6_outputs(8471) <= not a;
    layer6_outputs(8472) <= not a;
    layer6_outputs(8473) <= a xor b;
    layer6_outputs(8474) <= b;
    layer6_outputs(8475) <= a;
    layer6_outputs(8476) <= b;
    layer6_outputs(8477) <= not (a or b);
    layer6_outputs(8478) <= not a;
    layer6_outputs(8479) <= a;
    layer6_outputs(8480) <= not b;
    layer6_outputs(8481) <= a;
    layer6_outputs(8482) <= a;
    layer6_outputs(8483) <= not (a or b);
    layer6_outputs(8484) <= not (a or b);
    layer6_outputs(8485) <= a xor b;
    layer6_outputs(8486) <= not (a and b);
    layer6_outputs(8487) <= not b;
    layer6_outputs(8488) <= not b or a;
    layer6_outputs(8489) <= not (a or b);
    layer6_outputs(8490) <= not (a or b);
    layer6_outputs(8491) <= a and not b;
    layer6_outputs(8492) <= not a or b;
    layer6_outputs(8493) <= a xor b;
    layer6_outputs(8494) <= not b;
    layer6_outputs(8495) <= not a;
    layer6_outputs(8496) <= a and not b;
    layer6_outputs(8497) <= a xor b;
    layer6_outputs(8498) <= b;
    layer6_outputs(8499) <= b;
    layer6_outputs(8500) <= b;
    layer6_outputs(8501) <= not (a xor b);
    layer6_outputs(8502) <= not (a or b);
    layer6_outputs(8503) <= a;
    layer6_outputs(8504) <= b;
    layer6_outputs(8505) <= b;
    layer6_outputs(8506) <= not (a xor b);
    layer6_outputs(8507) <= a or b;
    layer6_outputs(8508) <= a xor b;
    layer6_outputs(8509) <= not a or b;
    layer6_outputs(8510) <= not b;
    layer6_outputs(8511) <= not (a xor b);
    layer6_outputs(8512) <= b;
    layer6_outputs(8513) <= not b;
    layer6_outputs(8514) <= not b or a;
    layer6_outputs(8515) <= b and not a;
    layer6_outputs(8516) <= a xor b;
    layer6_outputs(8517) <= not a;
    layer6_outputs(8518) <= not (a xor b);
    layer6_outputs(8519) <= not (a or b);
    layer6_outputs(8520) <= a;
    layer6_outputs(8521) <= not b;
    layer6_outputs(8522) <= a and not b;
    layer6_outputs(8523) <= not (a and b);
    layer6_outputs(8524) <= not b;
    layer6_outputs(8525) <= a xor b;
    layer6_outputs(8526) <= not b;
    layer6_outputs(8527) <= not (a xor b);
    layer6_outputs(8528) <= a xor b;
    layer6_outputs(8529) <= not (a xor b);
    layer6_outputs(8530) <= a;
    layer6_outputs(8531) <= not b;
    layer6_outputs(8532) <= not a or b;
    layer6_outputs(8533) <= not b;
    layer6_outputs(8534) <= not a;
    layer6_outputs(8535) <= not (a xor b);
    layer6_outputs(8536) <= b;
    layer6_outputs(8537) <= b;
    layer6_outputs(8538) <= not (a and b);
    layer6_outputs(8539) <= not a;
    layer6_outputs(8540) <= a and b;
    layer6_outputs(8541) <= a and not b;
    layer6_outputs(8542) <= a;
    layer6_outputs(8543) <= a;
    layer6_outputs(8544) <= a or b;
    layer6_outputs(8545) <= not a;
    layer6_outputs(8546) <= a;
    layer6_outputs(8547) <= a;
    layer6_outputs(8548) <= a and not b;
    layer6_outputs(8549) <= not b;
    layer6_outputs(8550) <= not (a xor b);
    layer6_outputs(8551) <= not a or b;
    layer6_outputs(8552) <= a xor b;
    layer6_outputs(8553) <= not a;
    layer6_outputs(8554) <= a xor b;
    layer6_outputs(8555) <= not b or a;
    layer6_outputs(8556) <= not a;
    layer6_outputs(8557) <= not b or a;
    layer6_outputs(8558) <= b and not a;
    layer6_outputs(8559) <= b;
    layer6_outputs(8560) <= not b;
    layer6_outputs(8561) <= a or b;
    layer6_outputs(8562) <= a and not b;
    layer6_outputs(8563) <= not (a or b);
    layer6_outputs(8564) <= b;
    layer6_outputs(8565) <= not (a or b);
    layer6_outputs(8566) <= a or b;
    layer6_outputs(8567) <= b and not a;
    layer6_outputs(8568) <= not b;
    layer6_outputs(8569) <= a xor b;
    layer6_outputs(8570) <= not (a xor b);
    layer6_outputs(8571) <= not (a xor b);
    layer6_outputs(8572) <= b and not a;
    layer6_outputs(8573) <= a xor b;
    layer6_outputs(8574) <= a or b;
    layer6_outputs(8575) <= b and not a;
    layer6_outputs(8576) <= not (a and b);
    layer6_outputs(8577) <= b and not a;
    layer6_outputs(8578) <= not (a or b);
    layer6_outputs(8579) <= a and b;
    layer6_outputs(8580) <= not a or b;
    layer6_outputs(8581) <= b;
    layer6_outputs(8582) <= not a;
    layer6_outputs(8583) <= not a;
    layer6_outputs(8584) <= not (a xor b);
    layer6_outputs(8585) <= b and not a;
    layer6_outputs(8586) <= not a;
    layer6_outputs(8587) <= not b;
    layer6_outputs(8588) <= b and not a;
    layer6_outputs(8589) <= a;
    layer6_outputs(8590) <= not b;
    layer6_outputs(8591) <= not (a and b);
    layer6_outputs(8592) <= a and not b;
    layer6_outputs(8593) <= not a or b;
    layer6_outputs(8594) <= '1';
    layer6_outputs(8595) <= a;
    layer6_outputs(8596) <= not (a and b);
    layer6_outputs(8597) <= b;
    layer6_outputs(8598) <= a or b;
    layer6_outputs(8599) <= not b;
    layer6_outputs(8600) <= a and not b;
    layer6_outputs(8601) <= not b;
    layer6_outputs(8602) <= b;
    layer6_outputs(8603) <= b and not a;
    layer6_outputs(8604) <= b;
    layer6_outputs(8605) <= not (a xor b);
    layer6_outputs(8606) <= a;
    layer6_outputs(8607) <= a and b;
    layer6_outputs(8608) <= b;
    layer6_outputs(8609) <= b and not a;
    layer6_outputs(8610) <= b and not a;
    layer6_outputs(8611) <= not b;
    layer6_outputs(8612) <= not (a xor b);
    layer6_outputs(8613) <= b and not a;
    layer6_outputs(8614) <= not a;
    layer6_outputs(8615) <= b;
    layer6_outputs(8616) <= not b or a;
    layer6_outputs(8617) <= a;
    layer6_outputs(8618) <= b;
    layer6_outputs(8619) <= not b;
    layer6_outputs(8620) <= a and b;
    layer6_outputs(8621) <= a;
    layer6_outputs(8622) <= a;
    layer6_outputs(8623) <= b;
    layer6_outputs(8624) <= a and not b;
    layer6_outputs(8625) <= not b;
    layer6_outputs(8626) <= a;
    layer6_outputs(8627) <= b;
    layer6_outputs(8628) <= not (a xor b);
    layer6_outputs(8629) <= b;
    layer6_outputs(8630) <= b;
    layer6_outputs(8631) <= not a or b;
    layer6_outputs(8632) <= a;
    layer6_outputs(8633) <= not (a xor b);
    layer6_outputs(8634) <= not a;
    layer6_outputs(8635) <= a and not b;
    layer6_outputs(8636) <= not b;
    layer6_outputs(8637) <= b;
    layer6_outputs(8638) <= a xor b;
    layer6_outputs(8639) <= a and not b;
    layer6_outputs(8640) <= a and not b;
    layer6_outputs(8641) <= b;
    layer6_outputs(8642) <= not (a or b);
    layer6_outputs(8643) <= a or b;
    layer6_outputs(8644) <= a or b;
    layer6_outputs(8645) <= not a;
    layer6_outputs(8646) <= not (a xor b);
    layer6_outputs(8647) <= a or b;
    layer6_outputs(8648) <= not (a xor b);
    layer6_outputs(8649) <= not b;
    layer6_outputs(8650) <= not a;
    layer6_outputs(8651) <= a;
    layer6_outputs(8652) <= a and not b;
    layer6_outputs(8653) <= not a;
    layer6_outputs(8654) <= not a or b;
    layer6_outputs(8655) <= a and b;
    layer6_outputs(8656) <= a xor b;
    layer6_outputs(8657) <= not b;
    layer6_outputs(8658) <= not (a and b);
    layer6_outputs(8659) <= a;
    layer6_outputs(8660) <= not b;
    layer6_outputs(8661) <= not (a and b);
    layer6_outputs(8662) <= b;
    layer6_outputs(8663) <= b;
    layer6_outputs(8664) <= not a;
    layer6_outputs(8665) <= a or b;
    layer6_outputs(8666) <= not (a xor b);
    layer6_outputs(8667) <= a;
    layer6_outputs(8668) <= a xor b;
    layer6_outputs(8669) <= not b or a;
    layer6_outputs(8670) <= not a;
    layer6_outputs(8671) <= a;
    layer6_outputs(8672) <= not (a xor b);
    layer6_outputs(8673) <= not a or b;
    layer6_outputs(8674) <= b and not a;
    layer6_outputs(8675) <= not (a or b);
    layer6_outputs(8676) <= not (a xor b);
    layer6_outputs(8677) <= a and b;
    layer6_outputs(8678) <= a xor b;
    layer6_outputs(8679) <= not a;
    layer6_outputs(8680) <= not b or a;
    layer6_outputs(8681) <= b and not a;
    layer6_outputs(8682) <= a;
    layer6_outputs(8683) <= not b;
    layer6_outputs(8684) <= not (a or b);
    layer6_outputs(8685) <= not (a xor b);
    layer6_outputs(8686) <= a;
    layer6_outputs(8687) <= a;
    layer6_outputs(8688) <= b;
    layer6_outputs(8689) <= not (a and b);
    layer6_outputs(8690) <= not (a xor b);
    layer6_outputs(8691) <= b;
    layer6_outputs(8692) <= not b;
    layer6_outputs(8693) <= b;
    layer6_outputs(8694) <= not a;
    layer6_outputs(8695) <= a;
    layer6_outputs(8696) <= not a;
    layer6_outputs(8697) <= not a;
    layer6_outputs(8698) <= not (a and b);
    layer6_outputs(8699) <= a;
    layer6_outputs(8700) <= not (a and b);
    layer6_outputs(8701) <= a;
    layer6_outputs(8702) <= a xor b;
    layer6_outputs(8703) <= a;
    layer6_outputs(8704) <= a or b;
    layer6_outputs(8705) <= a and b;
    layer6_outputs(8706) <= not (a or b);
    layer6_outputs(8707) <= a xor b;
    layer6_outputs(8708) <= b;
    layer6_outputs(8709) <= not a;
    layer6_outputs(8710) <= a and b;
    layer6_outputs(8711) <= b and not a;
    layer6_outputs(8712) <= b;
    layer6_outputs(8713) <= not b;
    layer6_outputs(8714) <= not (a xor b);
    layer6_outputs(8715) <= a xor b;
    layer6_outputs(8716) <= a;
    layer6_outputs(8717) <= a and b;
    layer6_outputs(8718) <= not a;
    layer6_outputs(8719) <= b;
    layer6_outputs(8720) <= not b;
    layer6_outputs(8721) <= a;
    layer6_outputs(8722) <= b;
    layer6_outputs(8723) <= b;
    layer6_outputs(8724) <= not b;
    layer6_outputs(8725) <= not (a and b);
    layer6_outputs(8726) <= a;
    layer6_outputs(8727) <= not b or a;
    layer6_outputs(8728) <= not (a xor b);
    layer6_outputs(8729) <= not (a xor b);
    layer6_outputs(8730) <= not (a or b);
    layer6_outputs(8731) <= a and b;
    layer6_outputs(8732) <= not b;
    layer6_outputs(8733) <= b;
    layer6_outputs(8734) <= a and b;
    layer6_outputs(8735) <= not (a xor b);
    layer6_outputs(8736) <= not (a xor b);
    layer6_outputs(8737) <= b;
    layer6_outputs(8738) <= not b;
    layer6_outputs(8739) <= a xor b;
    layer6_outputs(8740) <= not (a and b);
    layer6_outputs(8741) <= a xor b;
    layer6_outputs(8742) <= not b or a;
    layer6_outputs(8743) <= b;
    layer6_outputs(8744) <= not a;
    layer6_outputs(8745) <= not (a xor b);
    layer6_outputs(8746) <= not (a and b);
    layer6_outputs(8747) <= not (a xor b);
    layer6_outputs(8748) <= a xor b;
    layer6_outputs(8749) <= a and not b;
    layer6_outputs(8750) <= not (a xor b);
    layer6_outputs(8751) <= b and not a;
    layer6_outputs(8752) <= b;
    layer6_outputs(8753) <= not b;
    layer6_outputs(8754) <= a or b;
    layer6_outputs(8755) <= b;
    layer6_outputs(8756) <= not (a or b);
    layer6_outputs(8757) <= b;
    layer6_outputs(8758) <= a xor b;
    layer6_outputs(8759) <= a and not b;
    layer6_outputs(8760) <= b and not a;
    layer6_outputs(8761) <= not (a and b);
    layer6_outputs(8762) <= a xor b;
    layer6_outputs(8763) <= not a or b;
    layer6_outputs(8764) <= not b;
    layer6_outputs(8765) <= b;
    layer6_outputs(8766) <= not (a xor b);
    layer6_outputs(8767) <= not (a and b);
    layer6_outputs(8768) <= a xor b;
    layer6_outputs(8769) <= not (a and b);
    layer6_outputs(8770) <= not a;
    layer6_outputs(8771) <= a;
    layer6_outputs(8772) <= not (a or b);
    layer6_outputs(8773) <= not a;
    layer6_outputs(8774) <= a or b;
    layer6_outputs(8775) <= a or b;
    layer6_outputs(8776) <= not (a xor b);
    layer6_outputs(8777) <= '0';
    layer6_outputs(8778) <= a xor b;
    layer6_outputs(8779) <= a xor b;
    layer6_outputs(8780) <= not b;
    layer6_outputs(8781) <= not b or a;
    layer6_outputs(8782) <= not a;
    layer6_outputs(8783) <= not b or a;
    layer6_outputs(8784) <= not a;
    layer6_outputs(8785) <= not a;
    layer6_outputs(8786) <= not a;
    layer6_outputs(8787) <= a;
    layer6_outputs(8788) <= a;
    layer6_outputs(8789) <= b and not a;
    layer6_outputs(8790) <= b;
    layer6_outputs(8791) <= not b;
    layer6_outputs(8792) <= b;
    layer6_outputs(8793) <= a;
    layer6_outputs(8794) <= a xor b;
    layer6_outputs(8795) <= a or b;
    layer6_outputs(8796) <= not a or b;
    layer6_outputs(8797) <= not (a or b);
    layer6_outputs(8798) <= not b;
    layer6_outputs(8799) <= not (a xor b);
    layer6_outputs(8800) <= a;
    layer6_outputs(8801) <= not (a xor b);
    layer6_outputs(8802) <= not b;
    layer6_outputs(8803) <= a;
    layer6_outputs(8804) <= not b;
    layer6_outputs(8805) <= a or b;
    layer6_outputs(8806) <= a and not b;
    layer6_outputs(8807) <= not (a xor b);
    layer6_outputs(8808) <= b;
    layer6_outputs(8809) <= a;
    layer6_outputs(8810) <= a and not b;
    layer6_outputs(8811) <= a or b;
    layer6_outputs(8812) <= not a;
    layer6_outputs(8813) <= not a;
    layer6_outputs(8814) <= not b;
    layer6_outputs(8815) <= b;
    layer6_outputs(8816) <= not (a or b);
    layer6_outputs(8817) <= b;
    layer6_outputs(8818) <= b and not a;
    layer6_outputs(8819) <= not b;
    layer6_outputs(8820) <= not b;
    layer6_outputs(8821) <= not b or a;
    layer6_outputs(8822) <= not a;
    layer6_outputs(8823) <= a and b;
    layer6_outputs(8824) <= not a or b;
    layer6_outputs(8825) <= a xor b;
    layer6_outputs(8826) <= not b or a;
    layer6_outputs(8827) <= not b;
    layer6_outputs(8828) <= a and not b;
    layer6_outputs(8829) <= a and b;
    layer6_outputs(8830) <= a xor b;
    layer6_outputs(8831) <= not b;
    layer6_outputs(8832) <= not b;
    layer6_outputs(8833) <= not b or a;
    layer6_outputs(8834) <= a and not b;
    layer6_outputs(8835) <= b;
    layer6_outputs(8836) <= a xor b;
    layer6_outputs(8837) <= not b;
    layer6_outputs(8838) <= a;
    layer6_outputs(8839) <= a and b;
    layer6_outputs(8840) <= not b or a;
    layer6_outputs(8841) <= b and not a;
    layer6_outputs(8842) <= not b or a;
    layer6_outputs(8843) <= not a;
    layer6_outputs(8844) <= a or b;
    layer6_outputs(8845) <= not a;
    layer6_outputs(8846) <= a;
    layer6_outputs(8847) <= not b;
    layer6_outputs(8848) <= b and not a;
    layer6_outputs(8849) <= a or b;
    layer6_outputs(8850) <= not a;
    layer6_outputs(8851) <= not (a xor b);
    layer6_outputs(8852) <= not a;
    layer6_outputs(8853) <= b;
    layer6_outputs(8854) <= b;
    layer6_outputs(8855) <= not b or a;
    layer6_outputs(8856) <= not a;
    layer6_outputs(8857) <= not a;
    layer6_outputs(8858) <= b;
    layer6_outputs(8859) <= b;
    layer6_outputs(8860) <= not (a or b);
    layer6_outputs(8861) <= not (a xor b);
    layer6_outputs(8862) <= not (a xor b);
    layer6_outputs(8863) <= not (a or b);
    layer6_outputs(8864) <= b and not a;
    layer6_outputs(8865) <= b;
    layer6_outputs(8866) <= a;
    layer6_outputs(8867) <= b;
    layer6_outputs(8868) <= not a;
    layer6_outputs(8869) <= a and b;
    layer6_outputs(8870) <= a and b;
    layer6_outputs(8871) <= a and b;
    layer6_outputs(8872) <= not (a and b);
    layer6_outputs(8873) <= a;
    layer6_outputs(8874) <= a;
    layer6_outputs(8875) <= a xor b;
    layer6_outputs(8876) <= a and not b;
    layer6_outputs(8877) <= b and not a;
    layer6_outputs(8878) <= b and not a;
    layer6_outputs(8879) <= a xor b;
    layer6_outputs(8880) <= not a or b;
    layer6_outputs(8881) <= a xor b;
    layer6_outputs(8882) <= a;
    layer6_outputs(8883) <= a and b;
    layer6_outputs(8884) <= a or b;
    layer6_outputs(8885) <= a;
    layer6_outputs(8886) <= not a or b;
    layer6_outputs(8887) <= not b;
    layer6_outputs(8888) <= not b;
    layer6_outputs(8889) <= not a or b;
    layer6_outputs(8890) <= a xor b;
    layer6_outputs(8891) <= not a;
    layer6_outputs(8892) <= not (a or b);
    layer6_outputs(8893) <= not b;
    layer6_outputs(8894) <= a;
    layer6_outputs(8895) <= not a;
    layer6_outputs(8896) <= a;
    layer6_outputs(8897) <= not (a and b);
    layer6_outputs(8898) <= not b or a;
    layer6_outputs(8899) <= a and b;
    layer6_outputs(8900) <= b;
    layer6_outputs(8901) <= not a;
    layer6_outputs(8902) <= not b or a;
    layer6_outputs(8903) <= a;
    layer6_outputs(8904) <= not (a xor b);
    layer6_outputs(8905) <= not b or a;
    layer6_outputs(8906) <= a;
    layer6_outputs(8907) <= not (a xor b);
    layer6_outputs(8908) <= not (a and b);
    layer6_outputs(8909) <= b;
    layer6_outputs(8910) <= b and not a;
    layer6_outputs(8911) <= not (a xor b);
    layer6_outputs(8912) <= a and b;
    layer6_outputs(8913) <= a;
    layer6_outputs(8914) <= a and not b;
    layer6_outputs(8915) <= a and b;
    layer6_outputs(8916) <= a xor b;
    layer6_outputs(8917) <= a or b;
    layer6_outputs(8918) <= a;
    layer6_outputs(8919) <= not b;
    layer6_outputs(8920) <= not a;
    layer6_outputs(8921) <= a and not b;
    layer6_outputs(8922) <= a or b;
    layer6_outputs(8923) <= a and b;
    layer6_outputs(8924) <= not (a xor b);
    layer6_outputs(8925) <= not a;
    layer6_outputs(8926) <= not (a and b);
    layer6_outputs(8927) <= not (a or b);
    layer6_outputs(8928) <= b;
    layer6_outputs(8929) <= not b;
    layer6_outputs(8930) <= a;
    layer6_outputs(8931) <= not a;
    layer6_outputs(8932) <= not (a xor b);
    layer6_outputs(8933) <= not b or a;
    layer6_outputs(8934) <= not (a xor b);
    layer6_outputs(8935) <= not (a and b);
    layer6_outputs(8936) <= not a;
    layer6_outputs(8937) <= a or b;
    layer6_outputs(8938) <= a xor b;
    layer6_outputs(8939) <= b and not a;
    layer6_outputs(8940) <= b;
    layer6_outputs(8941) <= b;
    layer6_outputs(8942) <= a and b;
    layer6_outputs(8943) <= a;
    layer6_outputs(8944) <= not b;
    layer6_outputs(8945) <= not (a xor b);
    layer6_outputs(8946) <= b;
    layer6_outputs(8947) <= b;
    layer6_outputs(8948) <= b;
    layer6_outputs(8949) <= not (a xor b);
    layer6_outputs(8950) <= a and b;
    layer6_outputs(8951) <= not b or a;
    layer6_outputs(8952) <= a xor b;
    layer6_outputs(8953) <= a;
    layer6_outputs(8954) <= not b;
    layer6_outputs(8955) <= not (a and b);
    layer6_outputs(8956) <= not b;
    layer6_outputs(8957) <= not a;
    layer6_outputs(8958) <= b and not a;
    layer6_outputs(8959) <= b and not a;
    layer6_outputs(8960) <= a;
    layer6_outputs(8961) <= not b;
    layer6_outputs(8962) <= not a;
    layer6_outputs(8963) <= not b;
    layer6_outputs(8964) <= a;
    layer6_outputs(8965) <= b;
    layer6_outputs(8966) <= not b;
    layer6_outputs(8967) <= a;
    layer6_outputs(8968) <= not (a xor b);
    layer6_outputs(8969) <= not (a xor b);
    layer6_outputs(8970) <= not (a and b);
    layer6_outputs(8971) <= not (a or b);
    layer6_outputs(8972) <= not b;
    layer6_outputs(8973) <= not (a xor b);
    layer6_outputs(8974) <= a xor b;
    layer6_outputs(8975) <= b and not a;
    layer6_outputs(8976) <= a or b;
    layer6_outputs(8977) <= not (a and b);
    layer6_outputs(8978) <= not a;
    layer6_outputs(8979) <= b;
    layer6_outputs(8980) <= not (a or b);
    layer6_outputs(8981) <= a and b;
    layer6_outputs(8982) <= not a or b;
    layer6_outputs(8983) <= a xor b;
    layer6_outputs(8984) <= b and not a;
    layer6_outputs(8985) <= not (a and b);
    layer6_outputs(8986) <= not (a and b);
    layer6_outputs(8987) <= a and b;
    layer6_outputs(8988) <= not (a and b);
    layer6_outputs(8989) <= b;
    layer6_outputs(8990) <= not (a or b);
    layer6_outputs(8991) <= b;
    layer6_outputs(8992) <= not (a xor b);
    layer6_outputs(8993) <= not (a xor b);
    layer6_outputs(8994) <= not a;
    layer6_outputs(8995) <= not (a or b);
    layer6_outputs(8996) <= a xor b;
    layer6_outputs(8997) <= not (a or b);
    layer6_outputs(8998) <= a xor b;
    layer6_outputs(8999) <= a and not b;
    layer6_outputs(9000) <= a xor b;
    layer6_outputs(9001) <= a;
    layer6_outputs(9002) <= a xor b;
    layer6_outputs(9003) <= not a;
    layer6_outputs(9004) <= not (a or b);
    layer6_outputs(9005) <= not (a or b);
    layer6_outputs(9006) <= b;
    layer6_outputs(9007) <= not (a xor b);
    layer6_outputs(9008) <= not (a or b);
    layer6_outputs(9009) <= not (a or b);
    layer6_outputs(9010) <= not b or a;
    layer6_outputs(9011) <= not a;
    layer6_outputs(9012) <= a and b;
    layer6_outputs(9013) <= not (a and b);
    layer6_outputs(9014) <= a;
    layer6_outputs(9015) <= not (a xor b);
    layer6_outputs(9016) <= a;
    layer6_outputs(9017) <= b;
    layer6_outputs(9018) <= not (a and b);
    layer6_outputs(9019) <= b and not a;
    layer6_outputs(9020) <= not b;
    layer6_outputs(9021) <= b and not a;
    layer6_outputs(9022) <= not a;
    layer6_outputs(9023) <= not b;
    layer6_outputs(9024) <= not b;
    layer6_outputs(9025) <= a or b;
    layer6_outputs(9026) <= not a;
    layer6_outputs(9027) <= not (a xor b);
    layer6_outputs(9028) <= not (a xor b);
    layer6_outputs(9029) <= not b;
    layer6_outputs(9030) <= not (a and b);
    layer6_outputs(9031) <= a;
    layer6_outputs(9032) <= not (a and b);
    layer6_outputs(9033) <= a and not b;
    layer6_outputs(9034) <= not a or b;
    layer6_outputs(9035) <= b;
    layer6_outputs(9036) <= not (a xor b);
    layer6_outputs(9037) <= a;
    layer6_outputs(9038) <= not (a or b);
    layer6_outputs(9039) <= b;
    layer6_outputs(9040) <= not (a and b);
    layer6_outputs(9041) <= not a;
    layer6_outputs(9042) <= a and b;
    layer6_outputs(9043) <= not a;
    layer6_outputs(9044) <= b;
    layer6_outputs(9045) <= a and not b;
    layer6_outputs(9046) <= not a or b;
    layer6_outputs(9047) <= not b or a;
    layer6_outputs(9048) <= not (a xor b);
    layer6_outputs(9049) <= b;
    layer6_outputs(9050) <= a and b;
    layer6_outputs(9051) <= b;
    layer6_outputs(9052) <= b and not a;
    layer6_outputs(9053) <= a;
    layer6_outputs(9054) <= a xor b;
    layer6_outputs(9055) <= not a;
    layer6_outputs(9056) <= a;
    layer6_outputs(9057) <= not (a and b);
    layer6_outputs(9058) <= not (a or b);
    layer6_outputs(9059) <= not (a and b);
    layer6_outputs(9060) <= b;
    layer6_outputs(9061) <= not (a or b);
    layer6_outputs(9062) <= not (a xor b);
    layer6_outputs(9063) <= a and not b;
    layer6_outputs(9064) <= a and not b;
    layer6_outputs(9065) <= not (a or b);
    layer6_outputs(9066) <= a xor b;
    layer6_outputs(9067) <= not (a xor b);
    layer6_outputs(9068) <= not (a or b);
    layer6_outputs(9069) <= not a;
    layer6_outputs(9070) <= not b;
    layer6_outputs(9071) <= not b;
    layer6_outputs(9072) <= b;
    layer6_outputs(9073) <= a xor b;
    layer6_outputs(9074) <= a xor b;
    layer6_outputs(9075) <= not (a or b);
    layer6_outputs(9076) <= a xor b;
    layer6_outputs(9077) <= a xor b;
    layer6_outputs(9078) <= not b;
    layer6_outputs(9079) <= b;
    layer6_outputs(9080) <= not b;
    layer6_outputs(9081) <= not b;
    layer6_outputs(9082) <= not (a xor b);
    layer6_outputs(9083) <= b;
    layer6_outputs(9084) <= a;
    layer6_outputs(9085) <= a and b;
    layer6_outputs(9086) <= not a or b;
    layer6_outputs(9087) <= not a;
    layer6_outputs(9088) <= a;
    layer6_outputs(9089) <= b;
    layer6_outputs(9090) <= not a;
    layer6_outputs(9091) <= not (a and b);
    layer6_outputs(9092) <= a or b;
    layer6_outputs(9093) <= not (a xor b);
    layer6_outputs(9094) <= not b;
    layer6_outputs(9095) <= not b or a;
    layer6_outputs(9096) <= b and not a;
    layer6_outputs(9097) <= not (a xor b);
    layer6_outputs(9098) <= b;
    layer6_outputs(9099) <= a xor b;
    layer6_outputs(9100) <= a xor b;
    layer6_outputs(9101) <= a xor b;
    layer6_outputs(9102) <= not (a xor b);
    layer6_outputs(9103) <= not (a and b);
    layer6_outputs(9104) <= not (a or b);
    layer6_outputs(9105) <= a xor b;
    layer6_outputs(9106) <= a or b;
    layer6_outputs(9107) <= b and not a;
    layer6_outputs(9108) <= a or b;
    layer6_outputs(9109) <= a and not b;
    layer6_outputs(9110) <= not b;
    layer6_outputs(9111) <= b;
    layer6_outputs(9112) <= not a;
    layer6_outputs(9113) <= a and not b;
    layer6_outputs(9114) <= b;
    layer6_outputs(9115) <= a;
    layer6_outputs(9116) <= not a or b;
    layer6_outputs(9117) <= a xor b;
    layer6_outputs(9118) <= a and not b;
    layer6_outputs(9119) <= b;
    layer6_outputs(9120) <= b;
    layer6_outputs(9121) <= not a;
    layer6_outputs(9122) <= not (a or b);
    layer6_outputs(9123) <= a and b;
    layer6_outputs(9124) <= not b or a;
    layer6_outputs(9125) <= b;
    layer6_outputs(9126) <= not (a and b);
    layer6_outputs(9127) <= not a;
    layer6_outputs(9128) <= b;
    layer6_outputs(9129) <= not a;
    layer6_outputs(9130) <= not b;
    layer6_outputs(9131) <= a xor b;
    layer6_outputs(9132) <= not b;
    layer6_outputs(9133) <= not (a xor b);
    layer6_outputs(9134) <= b;
    layer6_outputs(9135) <= not (a xor b);
    layer6_outputs(9136) <= not (a xor b);
    layer6_outputs(9137) <= '1';
    layer6_outputs(9138) <= not (a or b);
    layer6_outputs(9139) <= a;
    layer6_outputs(9140) <= a xor b;
    layer6_outputs(9141) <= a;
    layer6_outputs(9142) <= a;
    layer6_outputs(9143) <= not a or b;
    layer6_outputs(9144) <= a or b;
    layer6_outputs(9145) <= a or b;
    layer6_outputs(9146) <= not a;
    layer6_outputs(9147) <= a;
    layer6_outputs(9148) <= not (a and b);
    layer6_outputs(9149) <= a or b;
    layer6_outputs(9150) <= not b or a;
    layer6_outputs(9151) <= '1';
    layer6_outputs(9152) <= b and not a;
    layer6_outputs(9153) <= not b;
    layer6_outputs(9154) <= b;
    layer6_outputs(9155) <= not (a xor b);
    layer6_outputs(9156) <= not (a xor b);
    layer6_outputs(9157) <= b;
    layer6_outputs(9158) <= a xor b;
    layer6_outputs(9159) <= b;
    layer6_outputs(9160) <= not (a and b);
    layer6_outputs(9161) <= a or b;
    layer6_outputs(9162) <= b and not a;
    layer6_outputs(9163) <= a and b;
    layer6_outputs(9164) <= not (a xor b);
    layer6_outputs(9165) <= a xor b;
    layer6_outputs(9166) <= not (a xor b);
    layer6_outputs(9167) <= a or b;
    layer6_outputs(9168) <= a xor b;
    layer6_outputs(9169) <= b and not a;
    layer6_outputs(9170) <= not b or a;
    layer6_outputs(9171) <= b;
    layer6_outputs(9172) <= b and not a;
    layer6_outputs(9173) <= a;
    layer6_outputs(9174) <= '1';
    layer6_outputs(9175) <= not a or b;
    layer6_outputs(9176) <= a;
    layer6_outputs(9177) <= not a;
    layer6_outputs(9178) <= a;
    layer6_outputs(9179) <= b;
    layer6_outputs(9180) <= a;
    layer6_outputs(9181) <= not a;
    layer6_outputs(9182) <= not a;
    layer6_outputs(9183) <= not (a or b);
    layer6_outputs(9184) <= a xor b;
    layer6_outputs(9185) <= a and b;
    layer6_outputs(9186) <= a xor b;
    layer6_outputs(9187) <= a or b;
    layer6_outputs(9188) <= b;
    layer6_outputs(9189) <= a and not b;
    layer6_outputs(9190) <= not (a or b);
    layer6_outputs(9191) <= not a or b;
    layer6_outputs(9192) <= a;
    layer6_outputs(9193) <= b;
    layer6_outputs(9194) <= a or b;
    layer6_outputs(9195) <= not b;
    layer6_outputs(9196) <= a or b;
    layer6_outputs(9197) <= not a or b;
    layer6_outputs(9198) <= a and not b;
    layer6_outputs(9199) <= a and b;
    layer6_outputs(9200) <= b;
    layer6_outputs(9201) <= not (a and b);
    layer6_outputs(9202) <= a or b;
    layer6_outputs(9203) <= not b or a;
    layer6_outputs(9204) <= not (a or b);
    layer6_outputs(9205) <= not a;
    layer6_outputs(9206) <= not a;
    layer6_outputs(9207) <= not b;
    layer6_outputs(9208) <= b;
    layer6_outputs(9209) <= a xor b;
    layer6_outputs(9210) <= not (a and b);
    layer6_outputs(9211) <= b;
    layer6_outputs(9212) <= a;
    layer6_outputs(9213) <= a and b;
    layer6_outputs(9214) <= a and not b;
    layer6_outputs(9215) <= not a or b;
    layer6_outputs(9216) <= not (a or b);
    layer6_outputs(9217) <= a and not b;
    layer6_outputs(9218) <= not b;
    layer6_outputs(9219) <= not a;
    layer6_outputs(9220) <= a or b;
    layer6_outputs(9221) <= not b or a;
    layer6_outputs(9222) <= a xor b;
    layer6_outputs(9223) <= a and not b;
    layer6_outputs(9224) <= b;
    layer6_outputs(9225) <= a;
    layer6_outputs(9226) <= b;
    layer6_outputs(9227) <= b and not a;
    layer6_outputs(9228) <= not a;
    layer6_outputs(9229) <= not (a or b);
    layer6_outputs(9230) <= a;
    layer6_outputs(9231) <= a;
    layer6_outputs(9232) <= a xor b;
    layer6_outputs(9233) <= not b or a;
    layer6_outputs(9234) <= b;
    layer6_outputs(9235) <= b and not a;
    layer6_outputs(9236) <= b;
    layer6_outputs(9237) <= a;
    layer6_outputs(9238) <= b;
    layer6_outputs(9239) <= a or b;
    layer6_outputs(9240) <= not b or a;
    layer6_outputs(9241) <= not a;
    layer6_outputs(9242) <= a;
    layer6_outputs(9243) <= not (a xor b);
    layer6_outputs(9244) <= a xor b;
    layer6_outputs(9245) <= not a;
    layer6_outputs(9246) <= not (a and b);
    layer6_outputs(9247) <= not (a and b);
    layer6_outputs(9248) <= not b;
    layer6_outputs(9249) <= a and not b;
    layer6_outputs(9250) <= not a;
    layer6_outputs(9251) <= not (a xor b);
    layer6_outputs(9252) <= a xor b;
    layer6_outputs(9253) <= a xor b;
    layer6_outputs(9254) <= a xor b;
    layer6_outputs(9255) <= b;
    layer6_outputs(9256) <= a;
    layer6_outputs(9257) <= not (a or b);
    layer6_outputs(9258) <= not (a or b);
    layer6_outputs(9259) <= not b;
    layer6_outputs(9260) <= a;
    layer6_outputs(9261) <= not a;
    layer6_outputs(9262) <= a or b;
    layer6_outputs(9263) <= not (a and b);
    layer6_outputs(9264) <= '1';
    layer6_outputs(9265) <= not a;
    layer6_outputs(9266) <= b;
    layer6_outputs(9267) <= not a;
    layer6_outputs(9268) <= not a;
    layer6_outputs(9269) <= a and not b;
    layer6_outputs(9270) <= not b;
    layer6_outputs(9271) <= not a;
    layer6_outputs(9272) <= not a;
    layer6_outputs(9273) <= b;
    layer6_outputs(9274) <= a;
    layer6_outputs(9275) <= a and b;
    layer6_outputs(9276) <= not b;
    layer6_outputs(9277) <= a or b;
    layer6_outputs(9278) <= a;
    layer6_outputs(9279) <= a or b;
    layer6_outputs(9280) <= a and not b;
    layer6_outputs(9281) <= not (a xor b);
    layer6_outputs(9282) <= not a;
    layer6_outputs(9283) <= not (a and b);
    layer6_outputs(9284) <= not (a xor b);
    layer6_outputs(9285) <= not b;
    layer6_outputs(9286) <= a;
    layer6_outputs(9287) <= not a;
    layer6_outputs(9288) <= not (a xor b);
    layer6_outputs(9289) <= not b;
    layer6_outputs(9290) <= b;
    layer6_outputs(9291) <= not (a xor b);
    layer6_outputs(9292) <= not b;
    layer6_outputs(9293) <= not (a xor b);
    layer6_outputs(9294) <= a and not b;
    layer6_outputs(9295) <= b;
    layer6_outputs(9296) <= a;
    layer6_outputs(9297) <= a xor b;
    layer6_outputs(9298) <= not b or a;
    layer6_outputs(9299) <= not b;
    layer6_outputs(9300) <= a or b;
    layer6_outputs(9301) <= b and not a;
    layer6_outputs(9302) <= a;
    layer6_outputs(9303) <= not b;
    layer6_outputs(9304) <= a;
    layer6_outputs(9305) <= not b or a;
    layer6_outputs(9306) <= a;
    layer6_outputs(9307) <= a xor b;
    layer6_outputs(9308) <= b;
    layer6_outputs(9309) <= not (a and b);
    layer6_outputs(9310) <= a and not b;
    layer6_outputs(9311) <= not b;
    layer6_outputs(9312) <= a;
    layer6_outputs(9313) <= not b;
    layer6_outputs(9314) <= not b;
    layer6_outputs(9315) <= not b;
    layer6_outputs(9316) <= a;
    layer6_outputs(9317) <= not a or b;
    layer6_outputs(9318) <= a and b;
    layer6_outputs(9319) <= not (a or b);
    layer6_outputs(9320) <= not b;
    layer6_outputs(9321) <= a or b;
    layer6_outputs(9322) <= a;
    layer6_outputs(9323) <= a;
    layer6_outputs(9324) <= a and not b;
    layer6_outputs(9325) <= a;
    layer6_outputs(9326) <= not b;
    layer6_outputs(9327) <= not a;
    layer6_outputs(9328) <= a;
    layer6_outputs(9329) <= a or b;
    layer6_outputs(9330) <= not (a or b);
    layer6_outputs(9331) <= not b;
    layer6_outputs(9332) <= not b;
    layer6_outputs(9333) <= not a or b;
    layer6_outputs(9334) <= a and b;
    layer6_outputs(9335) <= a xor b;
    layer6_outputs(9336) <= not a;
    layer6_outputs(9337) <= not a or b;
    layer6_outputs(9338) <= a and not b;
    layer6_outputs(9339) <= not a;
    layer6_outputs(9340) <= a xor b;
    layer6_outputs(9341) <= not a;
    layer6_outputs(9342) <= not a or b;
    layer6_outputs(9343) <= b;
    layer6_outputs(9344) <= b and not a;
    layer6_outputs(9345) <= b;
    layer6_outputs(9346) <= not (a and b);
    layer6_outputs(9347) <= a;
    layer6_outputs(9348) <= a or b;
    layer6_outputs(9349) <= a or b;
    layer6_outputs(9350) <= not (a and b);
    layer6_outputs(9351) <= a xor b;
    layer6_outputs(9352) <= a;
    layer6_outputs(9353) <= a;
    layer6_outputs(9354) <= a;
    layer6_outputs(9355) <= not b;
    layer6_outputs(9356) <= a xor b;
    layer6_outputs(9357) <= a or b;
    layer6_outputs(9358) <= not (a or b);
    layer6_outputs(9359) <= not (a xor b);
    layer6_outputs(9360) <= b;
    layer6_outputs(9361) <= not b;
    layer6_outputs(9362) <= not a or b;
    layer6_outputs(9363) <= b and not a;
    layer6_outputs(9364) <= a;
    layer6_outputs(9365) <= not a;
    layer6_outputs(9366) <= a;
    layer6_outputs(9367) <= not a;
    layer6_outputs(9368) <= not b;
    layer6_outputs(9369) <= not a or b;
    layer6_outputs(9370) <= a and not b;
    layer6_outputs(9371) <= not (a or b);
    layer6_outputs(9372) <= b;
    layer6_outputs(9373) <= not (a xor b);
    layer6_outputs(9374) <= b and not a;
    layer6_outputs(9375) <= b and not a;
    layer6_outputs(9376) <= a and b;
    layer6_outputs(9377) <= not (a xor b);
    layer6_outputs(9378) <= not (a and b);
    layer6_outputs(9379) <= a xor b;
    layer6_outputs(9380) <= a;
    layer6_outputs(9381) <= not a or b;
    layer6_outputs(9382) <= b;
    layer6_outputs(9383) <= a;
    layer6_outputs(9384) <= not (a and b);
    layer6_outputs(9385) <= not (a xor b);
    layer6_outputs(9386) <= a xor b;
    layer6_outputs(9387) <= b;
    layer6_outputs(9388) <= not (a xor b);
    layer6_outputs(9389) <= not (a and b);
    layer6_outputs(9390) <= not a;
    layer6_outputs(9391) <= a;
    layer6_outputs(9392) <= not a;
    layer6_outputs(9393) <= a or b;
    layer6_outputs(9394) <= a and b;
    layer6_outputs(9395) <= b;
    layer6_outputs(9396) <= b;
    layer6_outputs(9397) <= not (a xor b);
    layer6_outputs(9398) <= not a;
    layer6_outputs(9399) <= not b;
    layer6_outputs(9400) <= b;
    layer6_outputs(9401) <= a;
    layer6_outputs(9402) <= a or b;
    layer6_outputs(9403) <= not (a or b);
    layer6_outputs(9404) <= a;
    layer6_outputs(9405) <= a and not b;
    layer6_outputs(9406) <= a xor b;
    layer6_outputs(9407) <= not b;
    layer6_outputs(9408) <= not a or b;
    layer6_outputs(9409) <= a;
    layer6_outputs(9410) <= '1';
    layer6_outputs(9411) <= not a;
    layer6_outputs(9412) <= a or b;
    layer6_outputs(9413) <= a;
    layer6_outputs(9414) <= not (a xor b);
    layer6_outputs(9415) <= not b or a;
    layer6_outputs(9416) <= a xor b;
    layer6_outputs(9417) <= not (a or b);
    layer6_outputs(9418) <= a;
    layer6_outputs(9419) <= not (a xor b);
    layer6_outputs(9420) <= not b or a;
    layer6_outputs(9421) <= not b;
    layer6_outputs(9422) <= a and b;
    layer6_outputs(9423) <= a xor b;
    layer6_outputs(9424) <= not (a or b);
    layer6_outputs(9425) <= a xor b;
    layer6_outputs(9426) <= not (a xor b);
    layer6_outputs(9427) <= not a or b;
    layer6_outputs(9428) <= not b;
    layer6_outputs(9429) <= b;
    layer6_outputs(9430) <= a and b;
    layer6_outputs(9431) <= a or b;
    layer6_outputs(9432) <= not a;
    layer6_outputs(9433) <= not a;
    layer6_outputs(9434) <= not a;
    layer6_outputs(9435) <= not (a xor b);
    layer6_outputs(9436) <= not a;
    layer6_outputs(9437) <= not a or b;
    layer6_outputs(9438) <= not b;
    layer6_outputs(9439) <= a and not b;
    layer6_outputs(9440) <= b and not a;
    layer6_outputs(9441) <= b and not a;
    layer6_outputs(9442) <= a or b;
    layer6_outputs(9443) <= a and not b;
    layer6_outputs(9444) <= a xor b;
    layer6_outputs(9445) <= a and b;
    layer6_outputs(9446) <= not (a and b);
    layer6_outputs(9447) <= a xor b;
    layer6_outputs(9448) <= not a;
    layer6_outputs(9449) <= a and b;
    layer6_outputs(9450) <= not b;
    layer6_outputs(9451) <= not b;
    layer6_outputs(9452) <= not (a or b);
    layer6_outputs(9453) <= a xor b;
    layer6_outputs(9454) <= a xor b;
    layer6_outputs(9455) <= a and not b;
    layer6_outputs(9456) <= not (a xor b);
    layer6_outputs(9457) <= a and not b;
    layer6_outputs(9458) <= a;
    layer6_outputs(9459) <= not a or b;
    layer6_outputs(9460) <= b;
    layer6_outputs(9461) <= a;
    layer6_outputs(9462) <= a or b;
    layer6_outputs(9463) <= not a;
    layer6_outputs(9464) <= not b;
    layer6_outputs(9465) <= a xor b;
    layer6_outputs(9466) <= a;
    layer6_outputs(9467) <= a xor b;
    layer6_outputs(9468) <= not (a or b);
    layer6_outputs(9469) <= b and not a;
    layer6_outputs(9470) <= a xor b;
    layer6_outputs(9471) <= not b or a;
    layer6_outputs(9472) <= not b;
    layer6_outputs(9473) <= a;
    layer6_outputs(9474) <= b;
    layer6_outputs(9475) <= a;
    layer6_outputs(9476) <= b;
    layer6_outputs(9477) <= not b;
    layer6_outputs(9478) <= a and b;
    layer6_outputs(9479) <= a or b;
    layer6_outputs(9480) <= a or b;
    layer6_outputs(9481) <= a;
    layer6_outputs(9482) <= a xor b;
    layer6_outputs(9483) <= a;
    layer6_outputs(9484) <= not b;
    layer6_outputs(9485) <= not (a xor b);
    layer6_outputs(9486) <= b and not a;
    layer6_outputs(9487) <= not a;
    layer6_outputs(9488) <= not (a and b);
    layer6_outputs(9489) <= a and b;
    layer6_outputs(9490) <= not b or a;
    layer6_outputs(9491) <= not (a xor b);
    layer6_outputs(9492) <= not (a or b);
    layer6_outputs(9493) <= not b;
    layer6_outputs(9494) <= not b;
    layer6_outputs(9495) <= not (a or b);
    layer6_outputs(9496) <= not a or b;
    layer6_outputs(9497) <= not (a and b);
    layer6_outputs(9498) <= b;
    layer6_outputs(9499) <= not a;
    layer6_outputs(9500) <= a;
    layer6_outputs(9501) <= not a;
    layer6_outputs(9502) <= a xor b;
    layer6_outputs(9503) <= not (a and b);
    layer6_outputs(9504) <= a and b;
    layer6_outputs(9505) <= not b;
    layer6_outputs(9506) <= not b;
    layer6_outputs(9507) <= not (a xor b);
    layer6_outputs(9508) <= not b or a;
    layer6_outputs(9509) <= not a or b;
    layer6_outputs(9510) <= not b or a;
    layer6_outputs(9511) <= not b or a;
    layer6_outputs(9512) <= not (a xor b);
    layer6_outputs(9513) <= a xor b;
    layer6_outputs(9514) <= b;
    layer6_outputs(9515) <= not (a or b);
    layer6_outputs(9516) <= a xor b;
    layer6_outputs(9517) <= not (a or b);
    layer6_outputs(9518) <= a;
    layer6_outputs(9519) <= b and not a;
    layer6_outputs(9520) <= b and not a;
    layer6_outputs(9521) <= not (a xor b);
    layer6_outputs(9522) <= a and not b;
    layer6_outputs(9523) <= not (a and b);
    layer6_outputs(9524) <= not (a xor b);
    layer6_outputs(9525) <= b;
    layer6_outputs(9526) <= not a;
    layer6_outputs(9527) <= b;
    layer6_outputs(9528) <= b;
    layer6_outputs(9529) <= not (a or b);
    layer6_outputs(9530) <= not (a or b);
    layer6_outputs(9531) <= a or b;
    layer6_outputs(9532) <= b;
    layer6_outputs(9533) <= not (a xor b);
    layer6_outputs(9534) <= a or b;
    layer6_outputs(9535) <= b;
    layer6_outputs(9536) <= not (a or b);
    layer6_outputs(9537) <= not a;
    layer6_outputs(9538) <= '0';
    layer6_outputs(9539) <= not (a xor b);
    layer6_outputs(9540) <= not b;
    layer6_outputs(9541) <= not b;
    layer6_outputs(9542) <= not a;
    layer6_outputs(9543) <= not (a or b);
    layer6_outputs(9544) <= not a;
    layer6_outputs(9545) <= not a;
    layer6_outputs(9546) <= a and not b;
    layer6_outputs(9547) <= not (a xor b);
    layer6_outputs(9548) <= not b;
    layer6_outputs(9549) <= not b or a;
    layer6_outputs(9550) <= b;
    layer6_outputs(9551) <= not a;
    layer6_outputs(9552) <= a and b;
    layer6_outputs(9553) <= not (a or b);
    layer6_outputs(9554) <= not a;
    layer6_outputs(9555) <= not b;
    layer6_outputs(9556) <= not b;
    layer6_outputs(9557) <= not a;
    layer6_outputs(9558) <= a xor b;
    layer6_outputs(9559) <= '1';
    layer6_outputs(9560) <= b;
    layer6_outputs(9561) <= not (a and b);
    layer6_outputs(9562) <= not a;
    layer6_outputs(9563) <= not (a or b);
    layer6_outputs(9564) <= b and not a;
    layer6_outputs(9565) <= not a;
    layer6_outputs(9566) <= a xor b;
    layer6_outputs(9567) <= not (a or b);
    layer6_outputs(9568) <= b;
    layer6_outputs(9569) <= not a or b;
    layer6_outputs(9570) <= not (a and b);
    layer6_outputs(9571) <= not b;
    layer6_outputs(9572) <= a and not b;
    layer6_outputs(9573) <= a;
    layer6_outputs(9574) <= a xor b;
    layer6_outputs(9575) <= not (a and b);
    layer6_outputs(9576) <= a xor b;
    layer6_outputs(9577) <= not (a xor b);
    layer6_outputs(9578) <= not a;
    layer6_outputs(9579) <= a and b;
    layer6_outputs(9580) <= not (a xor b);
    layer6_outputs(9581) <= not b;
    layer6_outputs(9582) <= b and not a;
    layer6_outputs(9583) <= not (a and b);
    layer6_outputs(9584) <= b;
    layer6_outputs(9585) <= a xor b;
    layer6_outputs(9586) <= a;
    layer6_outputs(9587) <= not a;
    layer6_outputs(9588) <= not b or a;
    layer6_outputs(9589) <= a and not b;
    layer6_outputs(9590) <= b;
    layer6_outputs(9591) <= b;
    layer6_outputs(9592) <= not (a and b);
    layer6_outputs(9593) <= not a or b;
    layer6_outputs(9594) <= a;
    layer6_outputs(9595) <= not b;
    layer6_outputs(9596) <= a xor b;
    layer6_outputs(9597) <= a or b;
    layer6_outputs(9598) <= b and not a;
    layer6_outputs(9599) <= a xor b;
    layer6_outputs(9600) <= a xor b;
    layer6_outputs(9601) <= not (a xor b);
    layer6_outputs(9602) <= not (a or b);
    layer6_outputs(9603) <= not (a xor b);
    layer6_outputs(9604) <= a and not b;
    layer6_outputs(9605) <= a;
    layer6_outputs(9606) <= a and b;
    layer6_outputs(9607) <= b;
    layer6_outputs(9608) <= a;
    layer6_outputs(9609) <= not (a or b);
    layer6_outputs(9610) <= not b;
    layer6_outputs(9611) <= b and not a;
    layer6_outputs(9612) <= b and not a;
    layer6_outputs(9613) <= b and not a;
    layer6_outputs(9614) <= not (a xor b);
    layer6_outputs(9615) <= a;
    layer6_outputs(9616) <= not (a or b);
    layer6_outputs(9617) <= a or b;
    layer6_outputs(9618) <= not a;
    layer6_outputs(9619) <= not a;
    layer6_outputs(9620) <= not (a or b);
    layer6_outputs(9621) <= a and b;
    layer6_outputs(9622) <= not (a xor b);
    layer6_outputs(9623) <= a xor b;
    layer6_outputs(9624) <= a xor b;
    layer6_outputs(9625) <= a or b;
    layer6_outputs(9626) <= a and not b;
    layer6_outputs(9627) <= a;
    layer6_outputs(9628) <= b;
    layer6_outputs(9629) <= a or b;
    layer6_outputs(9630) <= not a;
    layer6_outputs(9631) <= not (a xor b);
    layer6_outputs(9632) <= b;
    layer6_outputs(9633) <= a and b;
    layer6_outputs(9634) <= not (a xor b);
    layer6_outputs(9635) <= not a;
    layer6_outputs(9636) <= a;
    layer6_outputs(9637) <= a;
    layer6_outputs(9638) <= a xor b;
    layer6_outputs(9639) <= a;
    layer6_outputs(9640) <= not (a xor b);
    layer6_outputs(9641) <= not (a xor b);
    layer6_outputs(9642) <= not b or a;
    layer6_outputs(9643) <= not (a or b);
    layer6_outputs(9644) <= a or b;
    layer6_outputs(9645) <= not b or a;
    layer6_outputs(9646) <= not b;
    layer6_outputs(9647) <= b and not a;
    layer6_outputs(9648) <= not b;
    layer6_outputs(9649) <= '0';
    layer6_outputs(9650) <= a and b;
    layer6_outputs(9651) <= not b;
    layer6_outputs(9652) <= a xor b;
    layer6_outputs(9653) <= a and not b;
    layer6_outputs(9654) <= a and b;
    layer6_outputs(9655) <= a and b;
    layer6_outputs(9656) <= not (a or b);
    layer6_outputs(9657) <= not a or b;
    layer6_outputs(9658) <= not (a and b);
    layer6_outputs(9659) <= a xor b;
    layer6_outputs(9660) <= not a or b;
    layer6_outputs(9661) <= b and not a;
    layer6_outputs(9662) <= not (a and b);
    layer6_outputs(9663) <= a xor b;
    layer6_outputs(9664) <= a xor b;
    layer6_outputs(9665) <= b;
    layer6_outputs(9666) <= b;
    layer6_outputs(9667) <= not b;
    layer6_outputs(9668) <= b;
    layer6_outputs(9669) <= not (a or b);
    layer6_outputs(9670) <= a and b;
    layer6_outputs(9671) <= not (a xor b);
    layer6_outputs(9672) <= a and not b;
    layer6_outputs(9673) <= not (a xor b);
    layer6_outputs(9674) <= a xor b;
    layer6_outputs(9675) <= a xor b;
    layer6_outputs(9676) <= not (a and b);
    layer6_outputs(9677) <= not a;
    layer6_outputs(9678) <= a xor b;
    layer6_outputs(9679) <= not a;
    layer6_outputs(9680) <= not a;
    layer6_outputs(9681) <= a;
    layer6_outputs(9682) <= not b;
    layer6_outputs(9683) <= not b;
    layer6_outputs(9684) <= not (a xor b);
    layer6_outputs(9685) <= not (a xor b);
    layer6_outputs(9686) <= b;
    layer6_outputs(9687) <= b;
    layer6_outputs(9688) <= a or b;
    layer6_outputs(9689) <= not a;
    layer6_outputs(9690) <= not b;
    layer6_outputs(9691) <= not (a xor b);
    layer6_outputs(9692) <= b;
    layer6_outputs(9693) <= a xor b;
    layer6_outputs(9694) <= '1';
    layer6_outputs(9695) <= not a;
    layer6_outputs(9696) <= not b;
    layer6_outputs(9697) <= b;
    layer6_outputs(9698) <= a xor b;
    layer6_outputs(9699) <= not a;
    layer6_outputs(9700) <= not a;
    layer6_outputs(9701) <= not a;
    layer6_outputs(9702) <= not a or b;
    layer6_outputs(9703) <= not a;
    layer6_outputs(9704) <= b and not a;
    layer6_outputs(9705) <= not (a xor b);
    layer6_outputs(9706) <= a and not b;
    layer6_outputs(9707) <= b and not a;
    layer6_outputs(9708) <= b;
    layer6_outputs(9709) <= not b;
    layer6_outputs(9710) <= a;
    layer6_outputs(9711) <= not (a or b);
    layer6_outputs(9712) <= not (a xor b);
    layer6_outputs(9713) <= a xor b;
    layer6_outputs(9714) <= not (a and b);
    layer6_outputs(9715) <= not b;
    layer6_outputs(9716) <= a or b;
    layer6_outputs(9717) <= a and b;
    layer6_outputs(9718) <= not b;
    layer6_outputs(9719) <= not b or a;
    layer6_outputs(9720) <= a xor b;
    layer6_outputs(9721) <= not (a xor b);
    layer6_outputs(9722) <= not b;
    layer6_outputs(9723) <= b;
    layer6_outputs(9724) <= not a;
    layer6_outputs(9725) <= not a or b;
    layer6_outputs(9726) <= not (a xor b);
    layer6_outputs(9727) <= a and not b;
    layer6_outputs(9728) <= not a;
    layer6_outputs(9729) <= not (a xor b);
    layer6_outputs(9730) <= not b;
    layer6_outputs(9731) <= b;
    layer6_outputs(9732) <= a;
    layer6_outputs(9733) <= a;
    layer6_outputs(9734) <= not b;
    layer6_outputs(9735) <= b;
    layer6_outputs(9736) <= not (a xor b);
    layer6_outputs(9737) <= not (a or b);
    layer6_outputs(9738) <= a xor b;
    layer6_outputs(9739) <= a and not b;
    layer6_outputs(9740) <= a or b;
    layer6_outputs(9741) <= b;
    layer6_outputs(9742) <= a and b;
    layer6_outputs(9743) <= not (a or b);
    layer6_outputs(9744) <= a xor b;
    layer6_outputs(9745) <= not b;
    layer6_outputs(9746) <= a;
    layer6_outputs(9747) <= b and not a;
    layer6_outputs(9748) <= b;
    layer6_outputs(9749) <= '0';
    layer6_outputs(9750) <= a and not b;
    layer6_outputs(9751) <= not a;
    layer6_outputs(9752) <= a xor b;
    layer6_outputs(9753) <= not (a xor b);
    layer6_outputs(9754) <= a and not b;
    layer6_outputs(9755) <= not a;
    layer6_outputs(9756) <= a or b;
    layer6_outputs(9757) <= not a;
    layer6_outputs(9758) <= not (a xor b);
    layer6_outputs(9759) <= a xor b;
    layer6_outputs(9760) <= a and b;
    layer6_outputs(9761) <= not a;
    layer6_outputs(9762) <= not a;
    layer6_outputs(9763) <= not (a xor b);
    layer6_outputs(9764) <= b;
    layer6_outputs(9765) <= not (a and b);
    layer6_outputs(9766) <= a xor b;
    layer6_outputs(9767) <= not (a xor b);
    layer6_outputs(9768) <= not a;
    layer6_outputs(9769) <= not a or b;
    layer6_outputs(9770) <= a and not b;
    layer6_outputs(9771) <= a or b;
    layer6_outputs(9772) <= b and not a;
    layer6_outputs(9773) <= a xor b;
    layer6_outputs(9774) <= b;
    layer6_outputs(9775) <= not (a and b);
    layer6_outputs(9776) <= not a;
    layer6_outputs(9777) <= a;
    layer6_outputs(9778) <= not b or a;
    layer6_outputs(9779) <= a and not b;
    layer6_outputs(9780) <= a and b;
    layer6_outputs(9781) <= b;
    layer6_outputs(9782) <= b;
    layer6_outputs(9783) <= not b;
    layer6_outputs(9784) <= not (a or b);
    layer6_outputs(9785) <= a or b;
    layer6_outputs(9786) <= not (a xor b);
    layer6_outputs(9787) <= a;
    layer6_outputs(9788) <= a and not b;
    layer6_outputs(9789) <= not b or a;
    layer6_outputs(9790) <= not a;
    layer6_outputs(9791) <= a and not b;
    layer6_outputs(9792) <= a;
    layer6_outputs(9793) <= not b;
    layer6_outputs(9794) <= not a;
    layer6_outputs(9795) <= not a;
    layer6_outputs(9796) <= not (a or b);
    layer6_outputs(9797) <= a;
    layer6_outputs(9798) <= not b;
    layer6_outputs(9799) <= a or b;
    layer6_outputs(9800) <= a and b;
    layer6_outputs(9801) <= not a or b;
    layer6_outputs(9802) <= b;
    layer6_outputs(9803) <= not b;
    layer6_outputs(9804) <= not a;
    layer6_outputs(9805) <= a;
    layer6_outputs(9806) <= a and b;
    layer6_outputs(9807) <= b;
    layer6_outputs(9808) <= not (a and b);
    layer6_outputs(9809) <= not a;
    layer6_outputs(9810) <= not a;
    layer6_outputs(9811) <= not a;
    layer6_outputs(9812) <= not a;
    layer6_outputs(9813) <= not (a xor b);
    layer6_outputs(9814) <= a and b;
    layer6_outputs(9815) <= a and b;
    layer6_outputs(9816) <= not b;
    layer6_outputs(9817) <= not b;
    layer6_outputs(9818) <= not a;
    layer6_outputs(9819) <= a or b;
    layer6_outputs(9820) <= not (a xor b);
    layer6_outputs(9821) <= not a;
    layer6_outputs(9822) <= not (a xor b);
    layer6_outputs(9823) <= a xor b;
    layer6_outputs(9824) <= not (a xor b);
    layer6_outputs(9825) <= a and not b;
    layer6_outputs(9826) <= b;
    layer6_outputs(9827) <= a and b;
    layer6_outputs(9828) <= not (a or b);
    layer6_outputs(9829) <= a xor b;
    layer6_outputs(9830) <= not a;
    layer6_outputs(9831) <= not (a and b);
    layer6_outputs(9832) <= b;
    layer6_outputs(9833) <= a;
    layer6_outputs(9834) <= b;
    layer6_outputs(9835) <= a or b;
    layer6_outputs(9836) <= a;
    layer6_outputs(9837) <= not (a xor b);
    layer6_outputs(9838) <= b;
    layer6_outputs(9839) <= not a;
    layer6_outputs(9840) <= a;
    layer6_outputs(9841) <= a xor b;
    layer6_outputs(9842) <= b;
    layer6_outputs(9843) <= a and b;
    layer6_outputs(9844) <= not a;
    layer6_outputs(9845) <= '1';
    layer6_outputs(9846) <= a xor b;
    layer6_outputs(9847) <= b;
    layer6_outputs(9848) <= not (a xor b);
    layer6_outputs(9849) <= a and b;
    layer6_outputs(9850) <= not b;
    layer6_outputs(9851) <= not a;
    layer6_outputs(9852) <= a and not b;
    layer6_outputs(9853) <= not (a and b);
    layer6_outputs(9854) <= not (a xor b);
    layer6_outputs(9855) <= not (a xor b);
    layer6_outputs(9856) <= a;
    layer6_outputs(9857) <= not b or a;
    layer6_outputs(9858) <= not a or b;
    layer6_outputs(9859) <= b;
    layer6_outputs(9860) <= a;
    layer6_outputs(9861) <= a xor b;
    layer6_outputs(9862) <= b;
    layer6_outputs(9863) <= not (a xor b);
    layer6_outputs(9864) <= a xor b;
    layer6_outputs(9865) <= not a;
    layer6_outputs(9866) <= b;
    layer6_outputs(9867) <= not b;
    layer6_outputs(9868) <= not b;
    layer6_outputs(9869) <= not a;
    layer6_outputs(9870) <= a;
    layer6_outputs(9871) <= not (a and b);
    layer6_outputs(9872) <= not a;
    layer6_outputs(9873) <= not b or a;
    layer6_outputs(9874) <= b;
    layer6_outputs(9875) <= a xor b;
    layer6_outputs(9876) <= not b;
    layer6_outputs(9877) <= not a;
    layer6_outputs(9878) <= not b;
    layer6_outputs(9879) <= a xor b;
    layer6_outputs(9880) <= a xor b;
    layer6_outputs(9881) <= not (a or b);
    layer6_outputs(9882) <= not b;
    layer6_outputs(9883) <= a;
    layer6_outputs(9884) <= not (a and b);
    layer6_outputs(9885) <= not a;
    layer6_outputs(9886) <= not b or a;
    layer6_outputs(9887) <= a or b;
    layer6_outputs(9888) <= b;
    layer6_outputs(9889) <= not (a or b);
    layer6_outputs(9890) <= not (a and b);
    layer6_outputs(9891) <= a or b;
    layer6_outputs(9892) <= a;
    layer6_outputs(9893) <= not a;
    layer6_outputs(9894) <= a and b;
    layer6_outputs(9895) <= b;
    layer6_outputs(9896) <= a xor b;
    layer6_outputs(9897) <= a and not b;
    layer6_outputs(9898) <= a;
    layer6_outputs(9899) <= a;
    layer6_outputs(9900) <= not (a or b);
    layer6_outputs(9901) <= not (a or b);
    layer6_outputs(9902) <= a and not b;
    layer6_outputs(9903) <= a xor b;
    layer6_outputs(9904) <= a and not b;
    layer6_outputs(9905) <= b;
    layer6_outputs(9906) <= '0';
    layer6_outputs(9907) <= not (a xor b);
    layer6_outputs(9908) <= not a;
    layer6_outputs(9909) <= a and b;
    layer6_outputs(9910) <= b;
    layer6_outputs(9911) <= a;
    layer6_outputs(9912) <= not a;
    layer6_outputs(9913) <= a;
    layer6_outputs(9914) <= not a;
    layer6_outputs(9915) <= b;
    layer6_outputs(9916) <= not (a or b);
    layer6_outputs(9917) <= a xor b;
    layer6_outputs(9918) <= not a or b;
    layer6_outputs(9919) <= a xor b;
    layer6_outputs(9920) <= not (a xor b);
    layer6_outputs(9921) <= a;
    layer6_outputs(9922) <= not (a xor b);
    layer6_outputs(9923) <= a or b;
    layer6_outputs(9924) <= not a;
    layer6_outputs(9925) <= not (a xor b);
    layer6_outputs(9926) <= not b;
    layer6_outputs(9927) <= not b;
    layer6_outputs(9928) <= not a;
    layer6_outputs(9929) <= a xor b;
    layer6_outputs(9930) <= not a;
    layer6_outputs(9931) <= not b or a;
    layer6_outputs(9932) <= a and b;
    layer6_outputs(9933) <= not a;
    layer6_outputs(9934) <= a;
    layer6_outputs(9935) <= not (a or b);
    layer6_outputs(9936) <= b and not a;
    layer6_outputs(9937) <= a and not b;
    layer6_outputs(9938) <= not b;
    layer6_outputs(9939) <= not a or b;
    layer6_outputs(9940) <= not b or a;
    layer6_outputs(9941) <= a;
    layer6_outputs(9942) <= b;
    layer6_outputs(9943) <= not (a xor b);
    layer6_outputs(9944) <= not (a xor b);
    layer6_outputs(9945) <= not b or a;
    layer6_outputs(9946) <= a and b;
    layer6_outputs(9947) <= a;
    layer6_outputs(9948) <= b and not a;
    layer6_outputs(9949) <= b and not a;
    layer6_outputs(9950) <= b;
    layer6_outputs(9951) <= not (a xor b);
    layer6_outputs(9952) <= a xor b;
    layer6_outputs(9953) <= b;
    layer6_outputs(9954) <= not (a xor b);
    layer6_outputs(9955) <= a or b;
    layer6_outputs(9956) <= not b;
    layer6_outputs(9957) <= not (a xor b);
    layer6_outputs(9958) <= a and b;
    layer6_outputs(9959) <= not (a xor b);
    layer6_outputs(9960) <= not a;
    layer6_outputs(9961) <= b;
    layer6_outputs(9962) <= b;
    layer6_outputs(9963) <= b;
    layer6_outputs(9964) <= b;
    layer6_outputs(9965) <= not b;
    layer6_outputs(9966) <= not (a xor b);
    layer6_outputs(9967) <= not b or a;
    layer6_outputs(9968) <= a xor b;
    layer6_outputs(9969) <= not b;
    layer6_outputs(9970) <= not a;
    layer6_outputs(9971) <= not a;
    layer6_outputs(9972) <= a;
    layer6_outputs(9973) <= not (a or b);
    layer6_outputs(9974) <= b;
    layer6_outputs(9975) <= b;
    layer6_outputs(9976) <= not b;
    layer6_outputs(9977) <= not a;
    layer6_outputs(9978) <= a and b;
    layer6_outputs(9979) <= a and b;
    layer6_outputs(9980) <= b;
    layer6_outputs(9981) <= not (a xor b);
    layer6_outputs(9982) <= b and not a;
    layer6_outputs(9983) <= a;
    layer6_outputs(9984) <= not a;
    layer6_outputs(9985) <= not a or b;
    layer6_outputs(9986) <= a and not b;
    layer6_outputs(9987) <= a;
    layer6_outputs(9988) <= not b;
    layer6_outputs(9989) <= not a or b;
    layer6_outputs(9990) <= a and b;
    layer6_outputs(9991) <= not a;
    layer6_outputs(9992) <= a and b;
    layer6_outputs(9993) <= b;
    layer6_outputs(9994) <= a xor b;
    layer6_outputs(9995) <= a xor b;
    layer6_outputs(9996) <= not b;
    layer6_outputs(9997) <= not (a or b);
    layer6_outputs(9998) <= not b;
    layer6_outputs(9999) <= b;
    layer6_outputs(10000) <= not (a xor b);
    layer6_outputs(10001) <= b and not a;
    layer6_outputs(10002) <= not (a xor b);
    layer6_outputs(10003) <= not (a xor b);
    layer6_outputs(10004) <= not b;
    layer6_outputs(10005) <= a and not b;
    layer6_outputs(10006) <= a and b;
    layer6_outputs(10007) <= a and not b;
    layer6_outputs(10008) <= not a;
    layer6_outputs(10009) <= b;
    layer6_outputs(10010) <= a and b;
    layer6_outputs(10011) <= not (a xor b);
    layer6_outputs(10012) <= a and not b;
    layer6_outputs(10013) <= not b;
    layer6_outputs(10014) <= b;
    layer6_outputs(10015) <= b and not a;
    layer6_outputs(10016) <= a xor b;
    layer6_outputs(10017) <= not a;
    layer6_outputs(10018) <= a xor b;
    layer6_outputs(10019) <= not a or b;
    layer6_outputs(10020) <= not b or a;
    layer6_outputs(10021) <= not (a or b);
    layer6_outputs(10022) <= a;
    layer6_outputs(10023) <= a;
    layer6_outputs(10024) <= not (a or b);
    layer6_outputs(10025) <= a and b;
    layer6_outputs(10026) <= not (a or b);
    layer6_outputs(10027) <= not b;
    layer6_outputs(10028) <= a xor b;
    layer6_outputs(10029) <= b and not a;
    layer6_outputs(10030) <= b;
    layer6_outputs(10031) <= not (a or b);
    layer6_outputs(10032) <= a;
    layer6_outputs(10033) <= not a;
    layer6_outputs(10034) <= not (a and b);
    layer6_outputs(10035) <= a and not b;
    layer6_outputs(10036) <= a;
    layer6_outputs(10037) <= not (a xor b);
    layer6_outputs(10038) <= not b;
    layer6_outputs(10039) <= not (a xor b);
    layer6_outputs(10040) <= a xor b;
    layer6_outputs(10041) <= a or b;
    layer6_outputs(10042) <= a;
    layer6_outputs(10043) <= a and b;
    layer6_outputs(10044) <= a xor b;
    layer6_outputs(10045) <= not a;
    layer6_outputs(10046) <= '1';
    layer6_outputs(10047) <= not a;
    layer6_outputs(10048) <= not a;
    layer6_outputs(10049) <= not a;
    layer6_outputs(10050) <= not b;
    layer6_outputs(10051) <= a;
    layer6_outputs(10052) <= b and not a;
    layer6_outputs(10053) <= b;
    layer6_outputs(10054) <= not a;
    layer6_outputs(10055) <= not (a and b);
    layer6_outputs(10056) <= not (a and b);
    layer6_outputs(10057) <= a;
    layer6_outputs(10058) <= not b;
    layer6_outputs(10059) <= not (a or b);
    layer6_outputs(10060) <= a xor b;
    layer6_outputs(10061) <= b;
    layer6_outputs(10062) <= b and not a;
    layer6_outputs(10063) <= a xor b;
    layer6_outputs(10064) <= b;
    layer6_outputs(10065) <= not (a xor b);
    layer6_outputs(10066) <= a and not b;
    layer6_outputs(10067) <= not a;
    layer6_outputs(10068) <= b;
    layer6_outputs(10069) <= a;
    layer6_outputs(10070) <= not a;
    layer6_outputs(10071) <= not b or a;
    layer6_outputs(10072) <= not b;
    layer6_outputs(10073) <= b;
    layer6_outputs(10074) <= a xor b;
    layer6_outputs(10075) <= a xor b;
    layer6_outputs(10076) <= not b;
    layer6_outputs(10077) <= not a;
    layer6_outputs(10078) <= not b or a;
    layer6_outputs(10079) <= not a;
    layer6_outputs(10080) <= not b;
    layer6_outputs(10081) <= not a or b;
    layer6_outputs(10082) <= a;
    layer6_outputs(10083) <= not (a xor b);
    layer6_outputs(10084) <= a;
    layer6_outputs(10085) <= not a or b;
    layer6_outputs(10086) <= b;
    layer6_outputs(10087) <= a and b;
    layer6_outputs(10088) <= a and not b;
    layer6_outputs(10089) <= not (a xor b);
    layer6_outputs(10090) <= a xor b;
    layer6_outputs(10091) <= not b or a;
    layer6_outputs(10092) <= a or b;
    layer6_outputs(10093) <= not b;
    layer6_outputs(10094) <= not a;
    layer6_outputs(10095) <= not b or a;
    layer6_outputs(10096) <= a xor b;
    layer6_outputs(10097) <= a xor b;
    layer6_outputs(10098) <= not a or b;
    layer6_outputs(10099) <= a and b;
    layer6_outputs(10100) <= b;
    layer6_outputs(10101) <= not a or b;
    layer6_outputs(10102) <= a and not b;
    layer6_outputs(10103) <= not a or b;
    layer6_outputs(10104) <= not a or b;
    layer6_outputs(10105) <= b;
    layer6_outputs(10106) <= a;
    layer6_outputs(10107) <= not a;
    layer6_outputs(10108) <= a;
    layer6_outputs(10109) <= b;
    layer6_outputs(10110) <= not a or b;
    layer6_outputs(10111) <= a and b;
    layer6_outputs(10112) <= a and not b;
    layer6_outputs(10113) <= b;
    layer6_outputs(10114) <= not (a xor b);
    layer6_outputs(10115) <= a and b;
    layer6_outputs(10116) <= b;
    layer6_outputs(10117) <= not a;
    layer6_outputs(10118) <= a and b;
    layer6_outputs(10119) <= a and not b;
    layer6_outputs(10120) <= a and b;
    layer6_outputs(10121) <= not b;
    layer6_outputs(10122) <= a or b;
    layer6_outputs(10123) <= a xor b;
    layer6_outputs(10124) <= b;
    layer6_outputs(10125) <= not (a xor b);
    layer6_outputs(10126) <= a;
    layer6_outputs(10127) <= b;
    layer6_outputs(10128) <= not a;
    layer6_outputs(10129) <= a;
    layer6_outputs(10130) <= not a or b;
    layer6_outputs(10131) <= not b;
    layer6_outputs(10132) <= a;
    layer6_outputs(10133) <= not a or b;
    layer6_outputs(10134) <= not a;
    layer6_outputs(10135) <= not a;
    layer6_outputs(10136) <= b and not a;
    layer6_outputs(10137) <= not (a xor b);
    layer6_outputs(10138) <= a and b;
    layer6_outputs(10139) <= not b;
    layer6_outputs(10140) <= a;
    layer6_outputs(10141) <= not (a and b);
    layer6_outputs(10142) <= b;
    layer6_outputs(10143) <= not a;
    layer6_outputs(10144) <= a and not b;
    layer6_outputs(10145) <= not (a or b);
    layer6_outputs(10146) <= b and not a;
    layer6_outputs(10147) <= not a;
    layer6_outputs(10148) <= a and not b;
    layer6_outputs(10149) <= not (a xor b);
    layer6_outputs(10150) <= not a;
    layer6_outputs(10151) <= b;
    layer6_outputs(10152) <= not (a xor b);
    layer6_outputs(10153) <= not b;
    layer6_outputs(10154) <= not (a xor b);
    layer6_outputs(10155) <= b;
    layer6_outputs(10156) <= not (a and b);
    layer6_outputs(10157) <= b;
    layer6_outputs(10158) <= not b;
    layer6_outputs(10159) <= not (a xor b);
    layer6_outputs(10160) <= b;
    layer6_outputs(10161) <= a and not b;
    layer6_outputs(10162) <= not b or a;
    layer6_outputs(10163) <= not a;
    layer6_outputs(10164) <= a xor b;
    layer6_outputs(10165) <= b and not a;
    layer6_outputs(10166) <= a xor b;
    layer6_outputs(10167) <= a;
    layer6_outputs(10168) <= not (a xor b);
    layer6_outputs(10169) <= a xor b;
    layer6_outputs(10170) <= not a;
    layer6_outputs(10171) <= a;
    layer6_outputs(10172) <= a;
    layer6_outputs(10173) <= a;
    layer6_outputs(10174) <= not b;
    layer6_outputs(10175) <= b and not a;
    layer6_outputs(10176) <= b and not a;
    layer6_outputs(10177) <= b;
    layer6_outputs(10178) <= not (a xor b);
    layer6_outputs(10179) <= not b;
    layer6_outputs(10180) <= a and b;
    layer6_outputs(10181) <= b and not a;
    layer6_outputs(10182) <= a or b;
    layer6_outputs(10183) <= b;
    layer6_outputs(10184) <= not (a xor b);
    layer6_outputs(10185) <= b;
    layer6_outputs(10186) <= not a;
    layer6_outputs(10187) <= a xor b;
    layer6_outputs(10188) <= a xor b;
    layer6_outputs(10189) <= not a;
    layer6_outputs(10190) <= not (a xor b);
    layer6_outputs(10191) <= not b;
    layer6_outputs(10192) <= not b or a;
    layer6_outputs(10193) <= a xor b;
    layer6_outputs(10194) <= a;
    layer6_outputs(10195) <= b;
    layer6_outputs(10196) <= b;
    layer6_outputs(10197) <= not b;
    layer6_outputs(10198) <= not (a xor b);
    layer6_outputs(10199) <= b and not a;
    layer6_outputs(10200) <= a xor b;
    layer6_outputs(10201) <= not (a and b);
    layer6_outputs(10202) <= b;
    layer6_outputs(10203) <= not b;
    layer6_outputs(10204) <= not a;
    layer6_outputs(10205) <= a;
    layer6_outputs(10206) <= not b;
    layer6_outputs(10207) <= not a;
    layer6_outputs(10208) <= not b or a;
    layer6_outputs(10209) <= b and not a;
    layer6_outputs(10210) <= b and not a;
    layer6_outputs(10211) <= not a or b;
    layer6_outputs(10212) <= not a;
    layer6_outputs(10213) <= b;
    layer6_outputs(10214) <= not (a or b);
    layer6_outputs(10215) <= not (a xor b);
    layer6_outputs(10216) <= a or b;
    layer6_outputs(10217) <= a xor b;
    layer6_outputs(10218) <= not (a xor b);
    layer6_outputs(10219) <= a xor b;
    layer6_outputs(10220) <= not (a xor b);
    layer6_outputs(10221) <= not (a or b);
    layer6_outputs(10222) <= b and not a;
    layer6_outputs(10223) <= a;
    layer6_outputs(10224) <= b;
    layer6_outputs(10225) <= a and b;
    layer6_outputs(10226) <= not (a xor b);
    layer6_outputs(10227) <= not (a or b);
    layer6_outputs(10228) <= not (a or b);
    layer6_outputs(10229) <= not a or b;
    layer6_outputs(10230) <= a and b;
    layer6_outputs(10231) <= b;
    layer6_outputs(10232) <= not b;
    layer6_outputs(10233) <= a and not b;
    layer6_outputs(10234) <= not (a xor b);
    layer6_outputs(10235) <= a and b;
    layer6_outputs(10236) <= not b or a;
    layer6_outputs(10237) <= not b or a;
    layer6_outputs(10238) <= a xor b;
    layer6_outputs(10239) <= not a or b;
    outputs(0) <= b;
    outputs(1) <= a xor b;
    outputs(2) <= a;
    outputs(3) <= not b;
    outputs(4) <= not b;
    outputs(5) <= not b;
    outputs(6) <= b;
    outputs(7) <= not a;
    outputs(8) <= b and not a;
    outputs(9) <= a and not b;
    outputs(10) <= not a;
    outputs(11) <= b;
    outputs(12) <= not (a or b);
    outputs(13) <= not (a or b);
    outputs(14) <= not (a xor b);
    outputs(15) <= a and b;
    outputs(16) <= a xor b;
    outputs(17) <= b;
    outputs(18) <= a;
    outputs(19) <= not (a and b);
    outputs(20) <= a;
    outputs(21) <= a and b;
    outputs(22) <= not (a xor b);
    outputs(23) <= not (a xor b);
    outputs(24) <= a xor b;
    outputs(25) <= not (a xor b);
    outputs(26) <= not a;
    outputs(27) <= a xor b;
    outputs(28) <= not (a xor b);
    outputs(29) <= a xor b;
    outputs(30) <= not a;
    outputs(31) <= b and not a;
    outputs(32) <= b and not a;
    outputs(33) <= not b;
    outputs(34) <= not (a xor b);
    outputs(35) <= b;
    outputs(36) <= a and not b;
    outputs(37) <= a xor b;
    outputs(38) <= not b;
    outputs(39) <= not a;
    outputs(40) <= a and b;
    outputs(41) <= b and not a;
    outputs(42) <= not a;
    outputs(43) <= b;
    outputs(44) <= a;
    outputs(45) <= a or b;
    outputs(46) <= b and not a;
    outputs(47) <= a xor b;
    outputs(48) <= not (a and b);
    outputs(49) <= a and b;
    outputs(50) <= a xor b;
    outputs(51) <= not (a xor b);
    outputs(52) <= a;
    outputs(53) <= not (a xor b);
    outputs(54) <= b;
    outputs(55) <= a or b;
    outputs(56) <= a xor b;
    outputs(57) <= a;
    outputs(58) <= not (a xor b);
    outputs(59) <= not (a xor b);
    outputs(60) <= a;
    outputs(61) <= b;
    outputs(62) <= not a;
    outputs(63) <= not b;
    outputs(64) <= not (a xor b);
    outputs(65) <= not (a xor b);
    outputs(66) <= a;
    outputs(67) <= a;
    outputs(68) <= not a;
    outputs(69) <= not a;
    outputs(70) <= a xor b;
    outputs(71) <= not b;
    outputs(72) <= b;
    outputs(73) <= not a;
    outputs(74) <= not b;
    outputs(75) <= not a;
    outputs(76) <= a or b;
    outputs(77) <= a;
    outputs(78) <= not (a xor b);
    outputs(79) <= b;
    outputs(80) <= a xor b;
    outputs(81) <= a and b;
    outputs(82) <= a;
    outputs(83) <= a;
    outputs(84) <= b;
    outputs(85) <= a;
    outputs(86) <= a;
    outputs(87) <= a and b;
    outputs(88) <= not (a xor b);
    outputs(89) <= not (a xor b);
    outputs(90) <= a or b;
    outputs(91) <= not b;
    outputs(92) <= not b;
    outputs(93) <= a;
    outputs(94) <= a xor b;
    outputs(95) <= not (a and b);
    outputs(96) <= a;
    outputs(97) <= a xor b;
    outputs(98) <= not (a xor b);
    outputs(99) <= not b;
    outputs(100) <= not a;
    outputs(101) <= not b;
    outputs(102) <= a and not b;
    outputs(103) <= not a;
    outputs(104) <= not (a xor b);
    outputs(105) <= a and b;
    outputs(106) <= b;
    outputs(107) <= not b;
    outputs(108) <= b;
    outputs(109) <= not a;
    outputs(110) <= not (a and b);
    outputs(111) <= not b;
    outputs(112) <= not a;
    outputs(113) <= b;
    outputs(114) <= not a;
    outputs(115) <= a;
    outputs(116) <= not (a xor b);
    outputs(117) <= not b;
    outputs(118) <= a;
    outputs(119) <= not a;
    outputs(120) <= not b;
    outputs(121) <= b;
    outputs(122) <= a xor b;
    outputs(123) <= b;
    outputs(124) <= b;
    outputs(125) <= not b;
    outputs(126) <= not (a or b);
    outputs(127) <= not (a xor b);
    outputs(128) <= a xor b;
    outputs(129) <= a and b;
    outputs(130) <= not a;
    outputs(131) <= a;
    outputs(132) <= a;
    outputs(133) <= b;
    outputs(134) <= a or b;
    outputs(135) <= a and b;
    outputs(136) <= a or b;
    outputs(137) <= a and b;
    outputs(138) <= not b;
    outputs(139) <= a and b;
    outputs(140) <= a;
    outputs(141) <= b;
    outputs(142) <= a;
    outputs(143) <= a;
    outputs(144) <= a;
    outputs(145) <= not (a xor b);
    outputs(146) <= not a;
    outputs(147) <= b;
    outputs(148) <= not (a xor b);
    outputs(149) <= not (a xor b);
    outputs(150) <= b;
    outputs(151) <= not b or a;
    outputs(152) <= not a;
    outputs(153) <= a;
    outputs(154) <= b;
    outputs(155) <= not b;
    outputs(156) <= not a;
    outputs(157) <= b;
    outputs(158) <= not (a and b);
    outputs(159) <= not a;
    outputs(160) <= a;
    outputs(161) <= a xor b;
    outputs(162) <= not (a xor b);
    outputs(163) <= b and not a;
    outputs(164) <= not (a xor b);
    outputs(165) <= not a;
    outputs(166) <= not (a and b);
    outputs(167) <= not b or a;
    outputs(168) <= not a;
    outputs(169) <= a and b;
    outputs(170) <= b;
    outputs(171) <= b;
    outputs(172) <= not (a or b);
    outputs(173) <= not (a xor b);
    outputs(174) <= a xor b;
    outputs(175) <= not (a or b);
    outputs(176) <= a xor b;
    outputs(177) <= a xor b;
    outputs(178) <= a xor b;
    outputs(179) <= not (a and b);
    outputs(180) <= not a;
    outputs(181) <= not a;
    outputs(182) <= not (a xor b);
    outputs(183) <= b;
    outputs(184) <= not b;
    outputs(185) <= a xor b;
    outputs(186) <= a xor b;
    outputs(187) <= a xor b;
    outputs(188) <= not a;
    outputs(189) <= not b;
    outputs(190) <= a and not b;
    outputs(191) <= a xor b;
    outputs(192) <= not (a xor b);
    outputs(193) <= a and b;
    outputs(194) <= not (a xor b);
    outputs(195) <= not (a xor b);
    outputs(196) <= not a;
    outputs(197) <= a xor b;
    outputs(198) <= not b;
    outputs(199) <= not a;
    outputs(200) <= a xor b;
    outputs(201) <= not (a xor b);
    outputs(202) <= b;
    outputs(203) <= a xor b;
    outputs(204) <= not a;
    outputs(205) <= a xor b;
    outputs(206) <= a xor b;
    outputs(207) <= a and not b;
    outputs(208) <= a;
    outputs(209) <= not b;
    outputs(210) <= not b;
    outputs(211) <= a;
    outputs(212) <= not b;
    outputs(213) <= b;
    outputs(214) <= a and not b;
    outputs(215) <= a xor b;
    outputs(216) <= not (a xor b);
    outputs(217) <= a;
    outputs(218) <= not b;
    outputs(219) <= not (a xor b);
    outputs(220) <= a xor b;
    outputs(221) <= b;
    outputs(222) <= a;
    outputs(223) <= b;
    outputs(224) <= a;
    outputs(225) <= a and b;
    outputs(226) <= not a;
    outputs(227) <= a xor b;
    outputs(228) <= a xor b;
    outputs(229) <= not (a or b);
    outputs(230) <= b;
    outputs(231) <= a xor b;
    outputs(232) <= a xor b;
    outputs(233) <= not (a or b);
    outputs(234) <= a and not b;
    outputs(235) <= not a;
    outputs(236) <= b;
    outputs(237) <= a;
    outputs(238) <= not (a xor b);
    outputs(239) <= a or b;
    outputs(240) <= not a;
    outputs(241) <= a or b;
    outputs(242) <= not b;
    outputs(243) <= not b;
    outputs(244) <= not b;
    outputs(245) <= b and not a;
    outputs(246) <= a and not b;
    outputs(247) <= a xor b;
    outputs(248) <= not b;
    outputs(249) <= a and not b;
    outputs(250) <= a and not b;
    outputs(251) <= b;
    outputs(252) <= a xor b;
    outputs(253) <= not a;
    outputs(254) <= not a;
    outputs(255) <= b;
    outputs(256) <= b;
    outputs(257) <= a;
    outputs(258) <= not a;
    outputs(259) <= not (a or b);
    outputs(260) <= b;
    outputs(261) <= not a;
    outputs(262) <= not a;
    outputs(263) <= not (a or b);
    outputs(264) <= a and b;
    outputs(265) <= a xor b;
    outputs(266) <= not (a xor b);
    outputs(267) <= not (a or b);
    outputs(268) <= not b or a;
    outputs(269) <= a xor b;
    outputs(270) <= a;
    outputs(271) <= not (a or b);
    outputs(272) <= b and not a;
    outputs(273) <= not a;
    outputs(274) <= not b;
    outputs(275) <= b;
    outputs(276) <= a and not b;
    outputs(277) <= not b;
    outputs(278) <= not a or b;
    outputs(279) <= a xor b;
    outputs(280) <= a and not b;
    outputs(281) <= a;
    outputs(282) <= b;
    outputs(283) <= b;
    outputs(284) <= not a;
    outputs(285) <= b;
    outputs(286) <= a xor b;
    outputs(287) <= not a;
    outputs(288) <= b and not a;
    outputs(289) <= b and not a;
    outputs(290) <= b and not a;
    outputs(291) <= a xor b;
    outputs(292) <= a xor b;
    outputs(293) <= a xor b;
    outputs(294) <= not a or b;
    outputs(295) <= not b;
    outputs(296) <= not a;
    outputs(297) <= a xor b;
    outputs(298) <= a;
    outputs(299) <= not b;
    outputs(300) <= a;
    outputs(301) <= not (a xor b);
    outputs(302) <= b;
    outputs(303) <= not a;
    outputs(304) <= a and b;
    outputs(305) <= b;
    outputs(306) <= not b or a;
    outputs(307) <= not (a xor b);
    outputs(308) <= a xor b;
    outputs(309) <= not (a xor b);
    outputs(310) <= b;
    outputs(311) <= not b;
    outputs(312) <= not a;
    outputs(313) <= not (a xor b);
    outputs(314) <= a xor b;
    outputs(315) <= b;
    outputs(316) <= a and not b;
    outputs(317) <= a xor b;
    outputs(318) <= a;
    outputs(319) <= not b;
    outputs(320) <= a xor b;
    outputs(321) <= b;
    outputs(322) <= a;
    outputs(323) <= not (a xor b);
    outputs(324) <= a xor b;
    outputs(325) <= a xor b;
    outputs(326) <= not a;
    outputs(327) <= a xor b;
    outputs(328) <= not (a xor b);
    outputs(329) <= b;
    outputs(330) <= a;
    outputs(331) <= not (a xor b);
    outputs(332) <= not (a and b);
    outputs(333) <= not (a xor b);
    outputs(334) <= a and not b;
    outputs(335) <= a xor b;
    outputs(336) <= b;
    outputs(337) <= not (a or b);
    outputs(338) <= b and not a;
    outputs(339) <= not b;
    outputs(340) <= not (a xor b);
    outputs(341) <= not (a xor b);
    outputs(342) <= a and b;
    outputs(343) <= not (a or b);
    outputs(344) <= b;
    outputs(345) <= not a;
    outputs(346) <= not (a xor b);
    outputs(347) <= a and not b;
    outputs(348) <= not b;
    outputs(349) <= a;
    outputs(350) <= b and not a;
    outputs(351) <= not b;
    outputs(352) <= b;
    outputs(353) <= a and b;
    outputs(354) <= not (a xor b);
    outputs(355) <= not a;
    outputs(356) <= not (a or b);
    outputs(357) <= not b;
    outputs(358) <= not b;
    outputs(359) <= not b;
    outputs(360) <= a xor b;
    outputs(361) <= not (a xor b);
    outputs(362) <= a and b;
    outputs(363) <= not b;
    outputs(364) <= not (a or b);
    outputs(365) <= a or b;
    outputs(366) <= a and b;
    outputs(367) <= not b;
    outputs(368) <= b;
    outputs(369) <= a xor b;
    outputs(370) <= not (a or b);
    outputs(371) <= b;
    outputs(372) <= not a;
    outputs(373) <= a;
    outputs(374) <= not (a xor b);
    outputs(375) <= not a;
    outputs(376) <= not a;
    outputs(377) <= a;
    outputs(378) <= b;
    outputs(379) <= not (a xor b);
    outputs(380) <= not b;
    outputs(381) <= not a;
    outputs(382) <= not (a and b);
    outputs(383) <= not (a xor b);
    outputs(384) <= a;
    outputs(385) <= b;
    outputs(386) <= a;
    outputs(387) <= a;
    outputs(388) <= a xor b;
    outputs(389) <= a and not b;
    outputs(390) <= not (a and b);
    outputs(391) <= b;
    outputs(392) <= not (a xor b);
    outputs(393) <= not b;
    outputs(394) <= not (a or b);
    outputs(395) <= a;
    outputs(396) <= not b;
    outputs(397) <= a;
    outputs(398) <= a xor b;
    outputs(399) <= not b;
    outputs(400) <= b;
    outputs(401) <= a xor b;
    outputs(402) <= b;
    outputs(403) <= not a;
    outputs(404) <= a and b;
    outputs(405) <= a xor b;
    outputs(406) <= b and not a;
    outputs(407) <= not a or b;
    outputs(408) <= b;
    outputs(409) <= a xor b;
    outputs(410) <= a and not b;
    outputs(411) <= b;
    outputs(412) <= not (a or b);
    outputs(413) <= not a;
    outputs(414) <= a xor b;
    outputs(415) <= not a;
    outputs(416) <= not b;
    outputs(417) <= not (a or b);
    outputs(418) <= a;
    outputs(419) <= not (a or b);
    outputs(420) <= not (a and b);
    outputs(421) <= a or b;
    outputs(422) <= a;
    outputs(423) <= a xor b;
    outputs(424) <= b;
    outputs(425) <= not a;
    outputs(426) <= not (a xor b);
    outputs(427) <= b;
    outputs(428) <= b;
    outputs(429) <= a xor b;
    outputs(430) <= not b;
    outputs(431) <= not a;
    outputs(432) <= b;
    outputs(433) <= not (a xor b);
    outputs(434) <= a xor b;
    outputs(435) <= b;
    outputs(436) <= not (a xor b);
    outputs(437) <= not b;
    outputs(438) <= b;
    outputs(439) <= a xor b;
    outputs(440) <= not a;
    outputs(441) <= b;
    outputs(442) <= b;
    outputs(443) <= a xor b;
    outputs(444) <= a;
    outputs(445) <= not a;
    outputs(446) <= not a;
    outputs(447) <= not b or a;
    outputs(448) <= not a;
    outputs(449) <= a;
    outputs(450) <= not (a xor b);
    outputs(451) <= not (a xor b);
    outputs(452) <= not b;
    outputs(453) <= not b;
    outputs(454) <= not (a xor b);
    outputs(455) <= not (a xor b);
    outputs(456) <= b and not a;
    outputs(457) <= a;
    outputs(458) <= a;
    outputs(459) <= not (a or b);
    outputs(460) <= not (a xor b);
    outputs(461) <= a;
    outputs(462) <= a xor b;
    outputs(463) <= not a;
    outputs(464) <= not b;
    outputs(465) <= a;
    outputs(466) <= b;
    outputs(467) <= a xor b;
    outputs(468) <= b;
    outputs(469) <= not (a or b);
    outputs(470) <= a xor b;
    outputs(471) <= a xor b;
    outputs(472) <= not b;
    outputs(473) <= a xor b;
    outputs(474) <= a xor b;
    outputs(475) <= b;
    outputs(476) <= not a or b;
    outputs(477) <= not (a xor b);
    outputs(478) <= not a;
    outputs(479) <= not (a or b);
    outputs(480) <= b;
    outputs(481) <= a and not b;
    outputs(482) <= not (a xor b);
    outputs(483) <= b;
    outputs(484) <= a xor b;
    outputs(485) <= not b;
    outputs(486) <= b;
    outputs(487) <= a xor b;
    outputs(488) <= b;
    outputs(489) <= not b;
    outputs(490) <= a and b;
    outputs(491) <= b;
    outputs(492) <= a xor b;
    outputs(493) <= a and b;
    outputs(494) <= not b;
    outputs(495) <= not a;
    outputs(496) <= not (a or b);
    outputs(497) <= not (a xor b);
    outputs(498) <= not (a xor b);
    outputs(499) <= a;
    outputs(500) <= b;
    outputs(501) <= a xor b;
    outputs(502) <= not (a xor b);
    outputs(503) <= not b;
    outputs(504) <= a;
    outputs(505) <= not b;
    outputs(506) <= not (a xor b);
    outputs(507) <= not b;
    outputs(508) <= a and b;
    outputs(509) <= a;
    outputs(510) <= not (a xor b);
    outputs(511) <= not a;
    outputs(512) <= not a;
    outputs(513) <= not (a xor b);
    outputs(514) <= not a;
    outputs(515) <= not b or a;
    outputs(516) <= a xor b;
    outputs(517) <= a and not b;
    outputs(518) <= b;
    outputs(519) <= not a;
    outputs(520) <= a xor b;
    outputs(521) <= a and not b;
    outputs(522) <= not (a xor b);
    outputs(523) <= a xor b;
    outputs(524) <= a xor b;
    outputs(525) <= a;
    outputs(526) <= not (a or b);
    outputs(527) <= not b or a;
    outputs(528) <= b;
    outputs(529) <= a and b;
    outputs(530) <= not (a xor b);
    outputs(531) <= not a;
    outputs(532) <= not a;
    outputs(533) <= a xor b;
    outputs(534) <= not b;
    outputs(535) <= b and not a;
    outputs(536) <= a or b;
    outputs(537) <= a;
    outputs(538) <= b and not a;
    outputs(539) <= a xor b;
    outputs(540) <= not a;
    outputs(541) <= a xor b;
    outputs(542) <= a;
    outputs(543) <= not a;
    outputs(544) <= b;
    outputs(545) <= a;
    outputs(546) <= a and not b;
    outputs(547) <= a xor b;
    outputs(548) <= a and b;
    outputs(549) <= not b;
    outputs(550) <= a;
    outputs(551) <= a;
    outputs(552) <= not (a and b);
    outputs(553) <= a and b;
    outputs(554) <= a;
    outputs(555) <= a and b;
    outputs(556) <= b;
    outputs(557) <= a and b;
    outputs(558) <= not b;
    outputs(559) <= b;
    outputs(560) <= b and not a;
    outputs(561) <= a xor b;
    outputs(562) <= a xor b;
    outputs(563) <= a or b;
    outputs(564) <= a xor b;
    outputs(565) <= a xor b;
    outputs(566) <= a and b;
    outputs(567) <= not a or b;
    outputs(568) <= not (a xor b);
    outputs(569) <= b and not a;
    outputs(570) <= not b or a;
    outputs(571) <= a and b;
    outputs(572) <= b;
    outputs(573) <= not b;
    outputs(574) <= not (a or b);
    outputs(575) <= not b;
    outputs(576) <= a xor b;
    outputs(577) <= not b;
    outputs(578) <= a;
    outputs(579) <= a xor b;
    outputs(580) <= not (a or b);
    outputs(581) <= not a or b;
    outputs(582) <= b;
    outputs(583) <= a and not b;
    outputs(584) <= a;
    outputs(585) <= not a;
    outputs(586) <= b and not a;
    outputs(587) <= not b;
    outputs(588) <= not a;
    outputs(589) <= b;
    outputs(590) <= b;
    outputs(591) <= b;
    outputs(592) <= not a;
    outputs(593) <= a;
    outputs(594) <= b;
    outputs(595) <= a xor b;
    outputs(596) <= b and not a;
    outputs(597) <= not a;
    outputs(598) <= a;
    outputs(599) <= not a;
    outputs(600) <= not (a or b);
    outputs(601) <= not b;
    outputs(602) <= b;
    outputs(603) <= not (a xor b);
    outputs(604) <= not (a xor b);
    outputs(605) <= not (a xor b);
    outputs(606) <= a and b;
    outputs(607) <= a;
    outputs(608) <= not b;
    outputs(609) <= not a;
    outputs(610) <= not a;
    outputs(611) <= a;
    outputs(612) <= not (a xor b);
    outputs(613) <= a xor b;
    outputs(614) <= not b;
    outputs(615) <= not (a xor b);
    outputs(616) <= not a;
    outputs(617) <= not (a xor b);
    outputs(618) <= not a;
    outputs(619) <= a;
    outputs(620) <= a;
    outputs(621) <= not a;
    outputs(622) <= b;
    outputs(623) <= not a;
    outputs(624) <= b;
    outputs(625) <= b;
    outputs(626) <= not (a and b);
    outputs(627) <= a;
    outputs(628) <= a xor b;
    outputs(629) <= not b;
    outputs(630) <= not a or b;
    outputs(631) <= a and not b;
    outputs(632) <= not a or b;
    outputs(633) <= not (a xor b);
    outputs(634) <= b;
    outputs(635) <= not (a xor b);
    outputs(636) <= not b;
    outputs(637) <= a and b;
    outputs(638) <= b;
    outputs(639) <= b and not a;
    outputs(640) <= a;
    outputs(641) <= a and not b;
    outputs(642) <= not (a or b);
    outputs(643) <= a;
    outputs(644) <= not (a xor b);
    outputs(645) <= not (a or b);
    outputs(646) <= not b or a;
    outputs(647) <= a;
    outputs(648) <= not (a xor b);
    outputs(649) <= a xor b;
    outputs(650) <= not b;
    outputs(651) <= not (a xor b);
    outputs(652) <= not a;
    outputs(653) <= not b;
    outputs(654) <= a;
    outputs(655) <= b;
    outputs(656) <= not a;
    outputs(657) <= a xor b;
    outputs(658) <= not a;
    outputs(659) <= a xor b;
    outputs(660) <= a xor b;
    outputs(661) <= a xor b;
    outputs(662) <= a xor b;
    outputs(663) <= a;
    outputs(664) <= b;
    outputs(665) <= not b;
    outputs(666) <= a;
    outputs(667) <= a xor b;
    outputs(668) <= '0';
    outputs(669) <= not a;
    outputs(670) <= b;
    outputs(671) <= not b;
    outputs(672) <= not a;
    outputs(673) <= a xor b;
    outputs(674) <= not (a xor b);
    outputs(675) <= a;
    outputs(676) <= not b;
    outputs(677) <= a and b;
    outputs(678) <= a and b;
    outputs(679) <= not a;
    outputs(680) <= a and not b;
    outputs(681) <= not b;
    outputs(682) <= a and not b;
    outputs(683) <= not (a xor b);
    outputs(684) <= a xor b;
    outputs(685) <= not a;
    outputs(686) <= not a;
    outputs(687) <= not a;
    outputs(688) <= not (a xor b);
    outputs(689) <= b;
    outputs(690) <= a and b;
    outputs(691) <= not (a xor b);
    outputs(692) <= not a;
    outputs(693) <= b;
    outputs(694) <= not a;
    outputs(695) <= a and b;
    outputs(696) <= not a or b;
    outputs(697) <= not a;
    outputs(698) <= a;
    outputs(699) <= not a;
    outputs(700) <= not (a xor b);
    outputs(701) <= not a or b;
    outputs(702) <= not (a or b);
    outputs(703) <= not (a xor b);
    outputs(704) <= b and not a;
    outputs(705) <= not (a xor b);
    outputs(706) <= a xor b;
    outputs(707) <= b;
    outputs(708) <= not (a and b);
    outputs(709) <= b;
    outputs(710) <= b;
    outputs(711) <= not (a or b);
    outputs(712) <= a;
    outputs(713) <= not a;
    outputs(714) <= not b or a;
    outputs(715) <= a and b;
    outputs(716) <= not (a and b);
    outputs(717) <= a or b;
    outputs(718) <= a xor b;
    outputs(719) <= a xor b;
    outputs(720) <= not (a or b);
    outputs(721) <= a xor b;
    outputs(722) <= not b or a;
    outputs(723) <= not b or a;
    outputs(724) <= not (a xor b);
    outputs(725) <= a;
    outputs(726) <= not (a or b);
    outputs(727) <= a xor b;
    outputs(728) <= not (a xor b);
    outputs(729) <= b;
    outputs(730) <= not a;
    outputs(731) <= not b or a;
    outputs(732) <= b;
    outputs(733) <= a xor b;
    outputs(734) <= a and not b;
    outputs(735) <= not (a xor b);
    outputs(736) <= not (a and b);
    outputs(737) <= b;
    outputs(738) <= a and b;
    outputs(739) <= not (a or b);
    outputs(740) <= b and not a;
    outputs(741) <= not (a xor b);
    outputs(742) <= a xor b;
    outputs(743) <= b;
    outputs(744) <= not a;
    outputs(745) <= not b;
    outputs(746) <= a;
    outputs(747) <= b;
    outputs(748) <= not (a xor b);
    outputs(749) <= a and b;
    outputs(750) <= not a;
    outputs(751) <= not b or a;
    outputs(752) <= b;
    outputs(753) <= not a;
    outputs(754) <= a xor b;
    outputs(755) <= b;
    outputs(756) <= a and not b;
    outputs(757) <= not (a xor b);
    outputs(758) <= a;
    outputs(759) <= a and not b;
    outputs(760) <= a;
    outputs(761) <= b;
    outputs(762) <= not a;
    outputs(763) <= not (a or b);
    outputs(764) <= a;
    outputs(765) <= not b;
    outputs(766) <= b and not a;
    outputs(767) <= not a;
    outputs(768) <= a;
    outputs(769) <= b;
    outputs(770) <= not b;
    outputs(771) <= not (a xor b);
    outputs(772) <= a xor b;
    outputs(773) <= not b;
    outputs(774) <= a;
    outputs(775) <= not b;
    outputs(776) <= a xor b;
    outputs(777) <= not b;
    outputs(778) <= not b or a;
    outputs(779) <= a;
    outputs(780) <= not b;
    outputs(781) <= not b;
    outputs(782) <= a or b;
    outputs(783) <= not a;
    outputs(784) <= a and b;
    outputs(785) <= not (a xor b);
    outputs(786) <= not (a or b);
    outputs(787) <= a and b;
    outputs(788) <= not (a xor b);
    outputs(789) <= a and not b;
    outputs(790) <= not (a xor b);
    outputs(791) <= not a;
    outputs(792) <= not (a xor b);
    outputs(793) <= a;
    outputs(794) <= a xor b;
    outputs(795) <= a;
    outputs(796) <= b;
    outputs(797) <= b and not a;
    outputs(798) <= not (a xor b);
    outputs(799) <= a or b;
    outputs(800) <= not b;
    outputs(801) <= not a;
    outputs(802) <= not b;
    outputs(803) <= a and b;
    outputs(804) <= b;
    outputs(805) <= not (a xor b);
    outputs(806) <= a xor b;
    outputs(807) <= not a;
    outputs(808) <= b;
    outputs(809) <= not (a xor b);
    outputs(810) <= not b;
    outputs(811) <= not b;
    outputs(812) <= a;
    outputs(813) <= a xor b;
    outputs(814) <= a;
    outputs(815) <= not (a xor b);
    outputs(816) <= not b;
    outputs(817) <= not (a xor b);
    outputs(818) <= a;
    outputs(819) <= not a;
    outputs(820) <= a or b;
    outputs(821) <= not (a xor b);
    outputs(822) <= not (a xor b);
    outputs(823) <= not (a xor b);
    outputs(824) <= not a or b;
    outputs(825) <= not (a or b);
    outputs(826) <= not (a xor b);
    outputs(827) <= not (a or b);
    outputs(828) <= b;
    outputs(829) <= a and not b;
    outputs(830) <= a;
    outputs(831) <= b;
    outputs(832) <= not a;
    outputs(833) <= b;
    outputs(834) <= not b;
    outputs(835) <= a;
    outputs(836) <= a;
    outputs(837) <= b;
    outputs(838) <= a xor b;
    outputs(839) <= not b;
    outputs(840) <= a;
    outputs(841) <= a;
    outputs(842) <= b;
    outputs(843) <= a;
    outputs(844) <= not b;
    outputs(845) <= a;
    outputs(846) <= not a;
    outputs(847) <= not a;
    outputs(848) <= not (a xor b);
    outputs(849) <= not (a or b);
    outputs(850) <= not a;
    outputs(851) <= not b;
    outputs(852) <= not a;
    outputs(853) <= a or b;
    outputs(854) <= not a;
    outputs(855) <= not b;
    outputs(856) <= b;
    outputs(857) <= not b or a;
    outputs(858) <= not a;
    outputs(859) <= b;
    outputs(860) <= a xor b;
    outputs(861) <= not a;
    outputs(862) <= not (a or b);
    outputs(863) <= not a;
    outputs(864) <= b;
    outputs(865) <= a and not b;
    outputs(866) <= a;
    outputs(867) <= not (a or b);
    outputs(868) <= b;
    outputs(869) <= not (a xor b);
    outputs(870) <= b;
    outputs(871) <= not (a and b);
    outputs(872) <= not a;
    outputs(873) <= not (a and b);
    outputs(874) <= a;
    outputs(875) <= not a;
    outputs(876) <= a;
    outputs(877) <= a xor b;
    outputs(878) <= not (a xor b);
    outputs(879) <= not a;
    outputs(880) <= not a;
    outputs(881) <= a;
    outputs(882) <= a;
    outputs(883) <= not (a xor b);
    outputs(884) <= not b;
    outputs(885) <= not a;
    outputs(886) <= a;
    outputs(887) <= a and b;
    outputs(888) <= a;
    outputs(889) <= not b;
    outputs(890) <= b;
    outputs(891) <= not b;
    outputs(892) <= a;
    outputs(893) <= a xor b;
    outputs(894) <= not a;
    outputs(895) <= not (a xor b);
    outputs(896) <= not a;
    outputs(897) <= a or b;
    outputs(898) <= a;
    outputs(899) <= a xor b;
    outputs(900) <= not b;
    outputs(901) <= not (a xor b);
    outputs(902) <= b;
    outputs(903) <= not a or b;
    outputs(904) <= not b;
    outputs(905) <= not (a xor b);
    outputs(906) <= a xor b;
    outputs(907) <= b and not a;
    outputs(908) <= b;
    outputs(909) <= a xor b;
    outputs(910) <= b;
    outputs(911) <= a xor b;
    outputs(912) <= a;
    outputs(913) <= a and not b;
    outputs(914) <= not (a xor b);
    outputs(915) <= a xor b;
    outputs(916) <= a and not b;
    outputs(917) <= a;
    outputs(918) <= b;
    outputs(919) <= a xor b;
    outputs(920) <= a xor b;
    outputs(921) <= not (a xor b);
    outputs(922) <= not b;
    outputs(923) <= a;
    outputs(924) <= a;
    outputs(925) <= b;
    outputs(926) <= not b;
    outputs(927) <= not b or a;
    outputs(928) <= not (a xor b);
    outputs(929) <= b;
    outputs(930) <= not b;
    outputs(931) <= not (a xor b);
    outputs(932) <= a;
    outputs(933) <= a;
    outputs(934) <= not (a xor b);
    outputs(935) <= a;
    outputs(936) <= a xor b;
    outputs(937) <= a and not b;
    outputs(938) <= a;
    outputs(939) <= not a;
    outputs(940) <= not a;
    outputs(941) <= b;
    outputs(942) <= a xor b;
    outputs(943) <= not (a xor b);
    outputs(944) <= a or b;
    outputs(945) <= not a;
    outputs(946) <= a;
    outputs(947) <= not (a or b);
    outputs(948) <= b;
    outputs(949) <= not b;
    outputs(950) <= not b;
    outputs(951) <= not a;
    outputs(952) <= a xor b;
    outputs(953) <= not a;
    outputs(954) <= a and not b;
    outputs(955) <= b;
    outputs(956) <= not b;
    outputs(957) <= not b;
    outputs(958) <= not a or b;
    outputs(959) <= a;
    outputs(960) <= not (a xor b);
    outputs(961) <= not a;
    outputs(962) <= not b or a;
    outputs(963) <= a and not b;
    outputs(964) <= b and not a;
    outputs(965) <= a;
    outputs(966) <= a and b;
    outputs(967) <= b;
    outputs(968) <= not a;
    outputs(969) <= a xor b;
    outputs(970) <= not a;
    outputs(971) <= a;
    outputs(972) <= not a;
    outputs(973) <= a and b;
    outputs(974) <= not a;
    outputs(975) <= b;
    outputs(976) <= a xor b;
    outputs(977) <= not (a xor b);
    outputs(978) <= a xor b;
    outputs(979) <= a and not b;
    outputs(980) <= not a;
    outputs(981) <= not b;
    outputs(982) <= a;
    outputs(983) <= a;
    outputs(984) <= not (a xor b);
    outputs(985) <= not b;
    outputs(986) <= a and not b;
    outputs(987) <= not (a or b);
    outputs(988) <= not b or a;
    outputs(989) <= b and not a;
    outputs(990) <= not b;
    outputs(991) <= not a;
    outputs(992) <= a;
    outputs(993) <= not (a or b);
    outputs(994) <= a and b;
    outputs(995) <= not (a and b);
    outputs(996) <= a and b;
    outputs(997) <= a;
    outputs(998) <= not a;
    outputs(999) <= b;
    outputs(1000) <= a xor b;
    outputs(1001) <= a xor b;
    outputs(1002) <= a and not b;
    outputs(1003) <= a;
    outputs(1004) <= not (a or b);
    outputs(1005) <= not a;
    outputs(1006) <= not b;
    outputs(1007) <= b and not a;
    outputs(1008) <= not b;
    outputs(1009) <= not a;
    outputs(1010) <= a and b;
    outputs(1011) <= a or b;
    outputs(1012) <= a and b;
    outputs(1013) <= not (a xor b);
    outputs(1014) <= a xor b;
    outputs(1015) <= not (a xor b);
    outputs(1016) <= not a;
    outputs(1017) <= b;
    outputs(1018) <= a xor b;
    outputs(1019) <= b;
    outputs(1020) <= a xor b;
    outputs(1021) <= a and not b;
    outputs(1022) <= not b;
    outputs(1023) <= a or b;
    outputs(1024) <= a and not b;
    outputs(1025) <= not b;
    outputs(1026) <= b and not a;
    outputs(1027) <= a and not b;
    outputs(1028) <= b;
    outputs(1029) <= not (a xor b);
    outputs(1030) <= not (a or b);
    outputs(1031) <= a and b;
    outputs(1032) <= not (a or b);
    outputs(1033) <= not (a xor b);
    outputs(1034) <= not (a and b);
    outputs(1035) <= a and b;
    outputs(1036) <= a and not b;
    outputs(1037) <= not (a xor b);
    outputs(1038) <= not (a or b);
    outputs(1039) <= a xor b;
    outputs(1040) <= not a;
    outputs(1041) <= b;
    outputs(1042) <= a or b;
    outputs(1043) <= a and not b;
    outputs(1044) <= not (a xor b);
    outputs(1045) <= a xor b;
    outputs(1046) <= not a;
    outputs(1047) <= a xor b;
    outputs(1048) <= not (a and b);
    outputs(1049) <= a xor b;
    outputs(1050) <= a;
    outputs(1051) <= not (a xor b);
    outputs(1052) <= b and not a;
    outputs(1053) <= b and not a;
    outputs(1054) <= not (a xor b);
    outputs(1055) <= a xor b;
    outputs(1056) <= b;
    outputs(1057) <= a xor b;
    outputs(1058) <= not (a xor b);
    outputs(1059) <= a xor b;
    outputs(1060) <= a xor b;
    outputs(1061) <= a and not b;
    outputs(1062) <= not b;
    outputs(1063) <= a and not b;
    outputs(1064) <= a xor b;
    outputs(1065) <= not a;
    outputs(1066) <= a xor b;
    outputs(1067) <= not a;
    outputs(1068) <= b;
    outputs(1069) <= not (a xor b);
    outputs(1070) <= b;
    outputs(1071) <= not b;
    outputs(1072) <= a xor b;
    outputs(1073) <= not (a xor b);
    outputs(1074) <= not a;
    outputs(1075) <= a xor b;
    outputs(1076) <= a;
    outputs(1077) <= not (a or b);
    outputs(1078) <= not b;
    outputs(1079) <= not b;
    outputs(1080) <= b;
    outputs(1081) <= a;
    outputs(1082) <= not (a xor b);
    outputs(1083) <= a;
    outputs(1084) <= a and not b;
    outputs(1085) <= not (a xor b);
    outputs(1086) <= not (a or b);
    outputs(1087) <= a xor b;
    outputs(1088) <= a xor b;
    outputs(1089) <= a or b;
    outputs(1090) <= a and b;
    outputs(1091) <= b and not a;
    outputs(1092) <= a and b;
    outputs(1093) <= not a or b;
    outputs(1094) <= not (a xor b);
    outputs(1095) <= not (a or b);
    outputs(1096) <= not (a or b);
    outputs(1097) <= b and not a;
    outputs(1098) <= not (a xor b);
    outputs(1099) <= b;
    outputs(1100) <= a;
    outputs(1101) <= not b or a;
    outputs(1102) <= not (a or b);
    outputs(1103) <= not (a or b);
    outputs(1104) <= not (a xor b);
    outputs(1105) <= b and not a;
    outputs(1106) <= a;
    outputs(1107) <= b;
    outputs(1108) <= not a or b;
    outputs(1109) <= not (a or b);
    outputs(1110) <= a xor b;
    outputs(1111) <= a xor b;
    outputs(1112) <= a xor b;
    outputs(1113) <= a and not b;
    outputs(1114) <= b;
    outputs(1115) <= b;
    outputs(1116) <= a xor b;
    outputs(1117) <= a or b;
    outputs(1118) <= b;
    outputs(1119) <= not (a xor b);
    outputs(1120) <= a xor b;
    outputs(1121) <= not b;
    outputs(1122) <= a;
    outputs(1123) <= a xor b;
    outputs(1124) <= a;
    outputs(1125) <= b;
    outputs(1126) <= a xor b;
    outputs(1127) <= not (a xor b);
    outputs(1128) <= not b;
    outputs(1129) <= a xor b;
    outputs(1130) <= a and b;
    outputs(1131) <= a and not b;
    outputs(1132) <= a xor b;
    outputs(1133) <= not b;
    outputs(1134) <= b and not a;
    outputs(1135) <= not (a xor b);
    outputs(1136) <= not (a or b);
    outputs(1137) <= b;
    outputs(1138) <= not (a xor b);
    outputs(1139) <= not a;
    outputs(1140) <= not b or a;
    outputs(1141) <= not (a xor b);
    outputs(1142) <= not a;
    outputs(1143) <= a and not b;
    outputs(1144) <= not (a xor b);
    outputs(1145) <= not (a xor b);
    outputs(1146) <= a xor b;
    outputs(1147) <= not (a xor b);
    outputs(1148) <= a;
    outputs(1149) <= not a;
    outputs(1150) <= not (a xor b);
    outputs(1151) <= not (a or b);
    outputs(1152) <= not b;
    outputs(1153) <= a xor b;
    outputs(1154) <= not a;
    outputs(1155) <= not b;
    outputs(1156) <= a;
    outputs(1157) <= a;
    outputs(1158) <= a or b;
    outputs(1159) <= not (a xor b);
    outputs(1160) <= b and not a;
    outputs(1161) <= a and not b;
    outputs(1162) <= b;
    outputs(1163) <= not a;
    outputs(1164) <= not (a or b);
    outputs(1165) <= a and not b;
    outputs(1166) <= a;
    outputs(1167) <= a xor b;
    outputs(1168) <= not a;
    outputs(1169) <= a;
    outputs(1170) <= a and b;
    outputs(1171) <= a;
    outputs(1172) <= not (a xor b);
    outputs(1173) <= b;
    outputs(1174) <= a xor b;
    outputs(1175) <= not a or b;
    outputs(1176) <= b and not a;
    outputs(1177) <= not (a xor b);
    outputs(1178) <= not b;
    outputs(1179) <= a xor b;
    outputs(1180) <= a;
    outputs(1181) <= b and not a;
    outputs(1182) <= a and not b;
    outputs(1183) <= a xor b;
    outputs(1184) <= a;
    outputs(1185) <= not a;
    outputs(1186) <= b;
    outputs(1187) <= not (a and b);
    outputs(1188) <= b;
    outputs(1189) <= a xor b;
    outputs(1190) <= not (a or b);
    outputs(1191) <= b and not a;
    outputs(1192) <= not (a or b);
    outputs(1193) <= not a;
    outputs(1194) <= not a;
    outputs(1195) <= a and not b;
    outputs(1196) <= a xor b;
    outputs(1197) <= not a;
    outputs(1198) <= a and b;
    outputs(1199) <= not b;
    outputs(1200) <= not (a xor b);
    outputs(1201) <= a and not b;
    outputs(1202) <= a;
    outputs(1203) <= not (a or b);
    outputs(1204) <= a;
    outputs(1205) <= not (a or b);
    outputs(1206) <= not (a or b);
    outputs(1207) <= b;
    outputs(1208) <= a xor b;
    outputs(1209) <= b;
    outputs(1210) <= a xor b;
    outputs(1211) <= not a;
    outputs(1212) <= not (a xor b);
    outputs(1213) <= a and b;
    outputs(1214) <= not b;
    outputs(1215) <= a xor b;
    outputs(1216) <= b;
    outputs(1217) <= b and not a;
    outputs(1218) <= not a;
    outputs(1219) <= not a;
    outputs(1220) <= a and not b;
    outputs(1221) <= b and not a;
    outputs(1222) <= a and not b;
    outputs(1223) <= not b;
    outputs(1224) <= a;
    outputs(1225) <= not (a or b);
    outputs(1226) <= not b;
    outputs(1227) <= not (a or b);
    outputs(1228) <= not a or b;
    outputs(1229) <= a xor b;
    outputs(1230) <= not a;
    outputs(1231) <= a;
    outputs(1232) <= a and b;
    outputs(1233) <= not a;
    outputs(1234) <= not (a xor b);
    outputs(1235) <= a;
    outputs(1236) <= a;
    outputs(1237) <= a xor b;
    outputs(1238) <= not (a xor b);
    outputs(1239) <= a;
    outputs(1240) <= a xor b;
    outputs(1241) <= a;
    outputs(1242) <= b;
    outputs(1243) <= not (a or b);
    outputs(1244) <= b;
    outputs(1245) <= not a;
    outputs(1246) <= a or b;
    outputs(1247) <= a and not b;
    outputs(1248) <= not b;
    outputs(1249) <= a;
    outputs(1250) <= b and not a;
    outputs(1251) <= not (a xor b);
    outputs(1252) <= not a;
    outputs(1253) <= not (a or b);
    outputs(1254) <= a;
    outputs(1255) <= a;
    outputs(1256) <= a xor b;
    outputs(1257) <= not (a xor b);
    outputs(1258) <= b;
    outputs(1259) <= '0';
    outputs(1260) <= b;
    outputs(1261) <= a;
    outputs(1262) <= not b;
    outputs(1263) <= b and not a;
    outputs(1264) <= a xor b;
    outputs(1265) <= a;
    outputs(1266) <= b and not a;
    outputs(1267) <= not (a xor b);
    outputs(1268) <= not (a xor b);
    outputs(1269) <= not (a or b);
    outputs(1270) <= a;
    outputs(1271) <= b and not a;
    outputs(1272) <= a xor b;
    outputs(1273) <= not a;
    outputs(1274) <= a xor b;
    outputs(1275) <= a or b;
    outputs(1276) <= a and b;
    outputs(1277) <= not (a xor b);
    outputs(1278) <= not a;
    outputs(1279) <= not b or a;
    outputs(1280) <= a xor b;
    outputs(1281) <= not (a xor b);
    outputs(1282) <= not b;
    outputs(1283) <= not (a xor b);
    outputs(1284) <= a;
    outputs(1285) <= not (a and b);
    outputs(1286) <= a xor b;
    outputs(1287) <= not b;
    outputs(1288) <= not a;
    outputs(1289) <= a and b;
    outputs(1290) <= not (a xor b);
    outputs(1291) <= a xor b;
    outputs(1292) <= b and not a;
    outputs(1293) <= not b;
    outputs(1294) <= b;
    outputs(1295) <= a xor b;
    outputs(1296) <= not b;
    outputs(1297) <= not (a xor b);
    outputs(1298) <= a and b;
    outputs(1299) <= a and b;
    outputs(1300) <= not (a xor b);
    outputs(1301) <= not b;
    outputs(1302) <= a and b;
    outputs(1303) <= not (a xor b);
    outputs(1304) <= not b;
    outputs(1305) <= not (a xor b);
    outputs(1306) <= b;
    outputs(1307) <= not (a xor b);
    outputs(1308) <= not (a xor b);
    outputs(1309) <= a and not b;
    outputs(1310) <= a xor b;
    outputs(1311) <= b;
    outputs(1312) <= a and b;
    outputs(1313) <= b;
    outputs(1314) <= b;
    outputs(1315) <= a;
    outputs(1316) <= not b;
    outputs(1317) <= a xor b;
    outputs(1318) <= a xor b;
    outputs(1319) <= b;
    outputs(1320) <= not a;
    outputs(1321) <= a xor b;
    outputs(1322) <= b;
    outputs(1323) <= not (a xor b);
    outputs(1324) <= b;
    outputs(1325) <= not a;
    outputs(1326) <= a xor b;
    outputs(1327) <= a xor b;
    outputs(1328) <= not b;
    outputs(1329) <= not (a xor b);
    outputs(1330) <= not (a or b);
    outputs(1331) <= b;
    outputs(1332) <= a xor b;
    outputs(1333) <= a and b;
    outputs(1334) <= a xor b;
    outputs(1335) <= not a;
    outputs(1336) <= a xor b;
    outputs(1337) <= not b;
    outputs(1338) <= b;
    outputs(1339) <= not (a or b);
    outputs(1340) <= not a;
    outputs(1341) <= a and b;
    outputs(1342) <= a;
    outputs(1343) <= not b;
    outputs(1344) <= a;
    outputs(1345) <= b and not a;
    outputs(1346) <= a xor b;
    outputs(1347) <= not (a xor b);
    outputs(1348) <= a xor b;
    outputs(1349) <= b and not a;
    outputs(1350) <= not (a or b);
    outputs(1351) <= not (a xor b);
    outputs(1352) <= not (a xor b);
    outputs(1353) <= b;
    outputs(1354) <= b and not a;
    outputs(1355) <= a xor b;
    outputs(1356) <= not a;
    outputs(1357) <= not (a xor b);
    outputs(1358) <= b and not a;
    outputs(1359) <= not (a xor b);
    outputs(1360) <= not b;
    outputs(1361) <= not (a xor b);
    outputs(1362) <= b and not a;
    outputs(1363) <= a xor b;
    outputs(1364) <= a;
    outputs(1365) <= not a;
    outputs(1366) <= a xor b;
    outputs(1367) <= not (a xor b);
    outputs(1368) <= a;
    outputs(1369) <= not (a xor b);
    outputs(1370) <= not b;
    outputs(1371) <= a;
    outputs(1372) <= not (a xor b);
    outputs(1373) <= not b;
    outputs(1374) <= not b;
    outputs(1375) <= not (a or b);
    outputs(1376) <= b and not a;
    outputs(1377) <= a and b;
    outputs(1378) <= a;
    outputs(1379) <= not a;
    outputs(1380) <= a and not b;
    outputs(1381) <= a and b;
    outputs(1382) <= a xor b;
    outputs(1383) <= not b;
    outputs(1384) <= b and not a;
    outputs(1385) <= not b;
    outputs(1386) <= a and b;
    outputs(1387) <= not (a xor b);
    outputs(1388) <= not (a xor b);
    outputs(1389) <= b;
    outputs(1390) <= not (a xor b);
    outputs(1391) <= a and not b;
    outputs(1392) <= not b;
    outputs(1393) <= b;
    outputs(1394) <= a xor b;
    outputs(1395) <= not (a or b);
    outputs(1396) <= a and not b;
    outputs(1397) <= not b;
    outputs(1398) <= a;
    outputs(1399) <= a;
    outputs(1400) <= b and not a;
    outputs(1401) <= b and not a;
    outputs(1402) <= a or b;
    outputs(1403) <= a and b;
    outputs(1404) <= a;
    outputs(1405) <= a and b;
    outputs(1406) <= not (a and b);
    outputs(1407) <= not (a xor b);
    outputs(1408) <= a and b;
    outputs(1409) <= not b;
    outputs(1410) <= not b;
    outputs(1411) <= b;
    outputs(1412) <= a and not b;
    outputs(1413) <= b;
    outputs(1414) <= b;
    outputs(1415) <= a xor b;
    outputs(1416) <= b;
    outputs(1417) <= a;
    outputs(1418) <= not a;
    outputs(1419) <= not a;
    outputs(1420) <= not (a xor b);
    outputs(1421) <= not (a and b);
    outputs(1422) <= not b;
    outputs(1423) <= a xor b;
    outputs(1424) <= not b;
    outputs(1425) <= b and not a;
    outputs(1426) <= a xor b;
    outputs(1427) <= a xor b;
    outputs(1428) <= not (a xor b);
    outputs(1429) <= not a;
    outputs(1430) <= a;
    outputs(1431) <= a xor b;
    outputs(1432) <= not (a xor b);
    outputs(1433) <= not a;
    outputs(1434) <= a and b;
    outputs(1435) <= not a or b;
    outputs(1436) <= not b;
    outputs(1437) <= not a;
    outputs(1438) <= not (a xor b);
    outputs(1439) <= a;
    outputs(1440) <= b;
    outputs(1441) <= b and not a;
    outputs(1442) <= b;
    outputs(1443) <= a xor b;
    outputs(1444) <= b;
    outputs(1445) <= not (a xor b);
    outputs(1446) <= a and b;
    outputs(1447) <= not b;
    outputs(1448) <= a xor b;
    outputs(1449) <= not b;
    outputs(1450) <= not b;
    outputs(1451) <= b;
    outputs(1452) <= a and not b;
    outputs(1453) <= not b;
    outputs(1454) <= a;
    outputs(1455) <= a and b;
    outputs(1456) <= a and b;
    outputs(1457) <= a xor b;
    outputs(1458) <= a xor b;
    outputs(1459) <= a and not b;
    outputs(1460) <= b and not a;
    outputs(1461) <= not b;
    outputs(1462) <= not b;
    outputs(1463) <= a;
    outputs(1464) <= a xor b;
    outputs(1465) <= a xor b;
    outputs(1466) <= not (a xor b);
    outputs(1467) <= b;
    outputs(1468) <= a;
    outputs(1469) <= a xor b;
    outputs(1470) <= not (a xor b);
    outputs(1471) <= not b;
    outputs(1472) <= not b;
    outputs(1473) <= not (a xor b);
    outputs(1474) <= b;
    outputs(1475) <= b;
    outputs(1476) <= a xor b;
    outputs(1477) <= not (a or b);
    outputs(1478) <= a;
    outputs(1479) <= not b;
    outputs(1480) <= b and not a;
    outputs(1481) <= not b;
    outputs(1482) <= not (a xor b);
    outputs(1483) <= not b;
    outputs(1484) <= not a;
    outputs(1485) <= not (a xor b);
    outputs(1486) <= b and not a;
    outputs(1487) <= a xor b;
    outputs(1488) <= a;
    outputs(1489) <= b;
    outputs(1490) <= not b;
    outputs(1491) <= not (a xor b);
    outputs(1492) <= not a;
    outputs(1493) <= not (a and b);
    outputs(1494) <= not b;
    outputs(1495) <= a;
    outputs(1496) <= a;
    outputs(1497) <= not (a or b);
    outputs(1498) <= a and b;
    outputs(1499) <= not a or b;
    outputs(1500) <= b;
    outputs(1501) <= not a;
    outputs(1502) <= a and not b;
    outputs(1503) <= not b;
    outputs(1504) <= not (a xor b);
    outputs(1505) <= not (a xor b);
    outputs(1506) <= not a;
    outputs(1507) <= not b;
    outputs(1508) <= not a or b;
    outputs(1509) <= not a;
    outputs(1510) <= a xor b;
    outputs(1511) <= a xor b;
    outputs(1512) <= a and b;
    outputs(1513) <= b;
    outputs(1514) <= not (a or b);
    outputs(1515) <= a xor b;
    outputs(1516) <= b and not a;
    outputs(1517) <= not a;
    outputs(1518) <= a and not b;
    outputs(1519) <= not (a xor b);
    outputs(1520) <= b;
    outputs(1521) <= not a;
    outputs(1522) <= not (a xor b);
    outputs(1523) <= a xor b;
    outputs(1524) <= b;
    outputs(1525) <= a;
    outputs(1526) <= a xor b;
    outputs(1527) <= not b;
    outputs(1528) <= not a;
    outputs(1529) <= not b;
    outputs(1530) <= a xor b;
    outputs(1531) <= a;
    outputs(1532) <= not b;
    outputs(1533) <= b and not a;
    outputs(1534) <= not (a xor b);
    outputs(1535) <= not a;
    outputs(1536) <= not b;
    outputs(1537) <= not a;
    outputs(1538) <= a and b;
    outputs(1539) <= a and not b;
    outputs(1540) <= not b;
    outputs(1541) <= not (a xor b);
    outputs(1542) <= a and b;
    outputs(1543) <= a xor b;
    outputs(1544) <= a xor b;
    outputs(1545) <= a and not b;
    outputs(1546) <= b and not a;
    outputs(1547) <= not a;
    outputs(1548) <= a xor b;
    outputs(1549) <= not (a xor b);
    outputs(1550) <= a;
    outputs(1551) <= not a or b;
    outputs(1552) <= a and b;
    outputs(1553) <= not (a xor b);
    outputs(1554) <= a and b;
    outputs(1555) <= not a or b;
    outputs(1556) <= b and not a;
    outputs(1557) <= not a;
    outputs(1558) <= a and not b;
    outputs(1559) <= not a;
    outputs(1560) <= a or b;
    outputs(1561) <= b;
    outputs(1562) <= b and not a;
    outputs(1563) <= a xor b;
    outputs(1564) <= not (a xor b);
    outputs(1565) <= b;
    outputs(1566) <= not b;
    outputs(1567) <= b;
    outputs(1568) <= not b;
    outputs(1569) <= b;
    outputs(1570) <= a and b;
    outputs(1571) <= not (a xor b);
    outputs(1572) <= a xor b;
    outputs(1573) <= not a;
    outputs(1574) <= a;
    outputs(1575) <= a;
    outputs(1576) <= b and not a;
    outputs(1577) <= a xor b;
    outputs(1578) <= b;
    outputs(1579) <= a xor b;
    outputs(1580) <= not (a xor b);
    outputs(1581) <= a xor b;
    outputs(1582) <= a;
    outputs(1583) <= a and b;
    outputs(1584) <= not b;
    outputs(1585) <= a xor b;
    outputs(1586) <= not (a xor b);
    outputs(1587) <= a;
    outputs(1588) <= not a;
    outputs(1589) <= not (a or b);
    outputs(1590) <= a xor b;
    outputs(1591) <= b and not a;
    outputs(1592) <= not (a or b);
    outputs(1593) <= not (a or b);
    outputs(1594) <= b;
    outputs(1595) <= a and b;
    outputs(1596) <= a;
    outputs(1597) <= a xor b;
    outputs(1598) <= a xor b;
    outputs(1599) <= b;
    outputs(1600) <= b and not a;
    outputs(1601) <= not b;
    outputs(1602) <= not (a xor b);
    outputs(1603) <= not (a or b);
    outputs(1604) <= b;
    outputs(1605) <= b;
    outputs(1606) <= not b;
    outputs(1607) <= not (a xor b);
    outputs(1608) <= not (a xor b);
    outputs(1609) <= a;
    outputs(1610) <= not (a xor b);
    outputs(1611) <= b;
    outputs(1612) <= b and not a;
    outputs(1613) <= a xor b;
    outputs(1614) <= not (a xor b);
    outputs(1615) <= a and b;
    outputs(1616) <= not (a xor b);
    outputs(1617) <= a;
    outputs(1618) <= b;
    outputs(1619) <= a and b;
    outputs(1620) <= a and b;
    outputs(1621) <= not (a or b);
    outputs(1622) <= a;
    outputs(1623) <= not a;
    outputs(1624) <= a and not b;
    outputs(1625) <= not (a xor b);
    outputs(1626) <= not (a xor b);
    outputs(1627) <= not a;
    outputs(1628) <= b;
    outputs(1629) <= b;
    outputs(1630) <= a;
    outputs(1631) <= b and not a;
    outputs(1632) <= not (a or b);
    outputs(1633) <= not a;
    outputs(1634) <= a xor b;
    outputs(1635) <= a xor b;
    outputs(1636) <= not b;
    outputs(1637) <= not (a xor b);
    outputs(1638) <= b;
    outputs(1639) <= a xor b;
    outputs(1640) <= not (a xor b);
    outputs(1641) <= not b;
    outputs(1642) <= not a;
    outputs(1643) <= a;
    outputs(1644) <= not (a or b);
    outputs(1645) <= not (a xor b);
    outputs(1646) <= not (a or b);
    outputs(1647) <= a xor b;
    outputs(1648) <= a xor b;
    outputs(1649) <= a and not b;
    outputs(1650) <= not b or a;
    outputs(1651) <= b;
    outputs(1652) <= a xor b;
    outputs(1653) <= not a;
    outputs(1654) <= '0';
    outputs(1655) <= not (a xor b);
    outputs(1656) <= a and b;
    outputs(1657) <= not b;
    outputs(1658) <= b;
    outputs(1659) <= a and not b;
    outputs(1660) <= b and not a;
    outputs(1661) <= not a or b;
    outputs(1662) <= not (a xor b);
    outputs(1663) <= not b;
    outputs(1664) <= not (a or b);
    outputs(1665) <= a xor b;
    outputs(1666) <= not (a xor b);
    outputs(1667) <= a xor b;
    outputs(1668) <= a and not b;
    outputs(1669) <= not a;
    outputs(1670) <= a xor b;
    outputs(1671) <= not (a or b);
    outputs(1672) <= b;
    outputs(1673) <= not (a xor b);
    outputs(1674) <= a;
    outputs(1675) <= not a;
    outputs(1676) <= a xor b;
    outputs(1677) <= b and not a;
    outputs(1678) <= a and b;
    outputs(1679) <= not (a xor b);
    outputs(1680) <= not a;
    outputs(1681) <= a and b;
    outputs(1682) <= not (a xor b);
    outputs(1683) <= not (a or b);
    outputs(1684) <= not (a xor b);
    outputs(1685) <= b;
    outputs(1686) <= a xor b;
    outputs(1687) <= not (a and b);
    outputs(1688) <= a xor b;
    outputs(1689) <= not a;
    outputs(1690) <= not b;
    outputs(1691) <= a xor b;
    outputs(1692) <= b and not a;
    outputs(1693) <= a and not b;
    outputs(1694) <= not a;
    outputs(1695) <= a xor b;
    outputs(1696) <= a xor b;
    outputs(1697) <= a;
    outputs(1698) <= a xor b;
    outputs(1699) <= not a or b;
    outputs(1700) <= b;
    outputs(1701) <= b;
    outputs(1702) <= b;
    outputs(1703) <= a and not b;
    outputs(1704) <= a xor b;
    outputs(1705) <= not b;
    outputs(1706) <= a xor b;
    outputs(1707) <= not b;
    outputs(1708) <= b and not a;
    outputs(1709) <= not b;
    outputs(1710) <= not (a and b);
    outputs(1711) <= not a;
    outputs(1712) <= not (a or b);
    outputs(1713) <= not (a xor b);
    outputs(1714) <= not (a or b);
    outputs(1715) <= a;
    outputs(1716) <= not (a xor b);
    outputs(1717) <= a and not b;
    outputs(1718) <= a and b;
    outputs(1719) <= a;
    outputs(1720) <= not (a xor b);
    outputs(1721) <= not (a or b);
    outputs(1722) <= a and not b;
    outputs(1723) <= a xor b;
    outputs(1724) <= a xor b;
    outputs(1725) <= not b or a;
    outputs(1726) <= not a;
    outputs(1727) <= a;
    outputs(1728) <= b;
    outputs(1729) <= a;
    outputs(1730) <= not (a xor b);
    outputs(1731) <= b;
    outputs(1732) <= not (a xor b);
    outputs(1733) <= not (a or b);
    outputs(1734) <= not (a xor b);
    outputs(1735) <= a;
    outputs(1736) <= a xor b;
    outputs(1737) <= a or b;
    outputs(1738) <= not (a or b);
    outputs(1739) <= not (a or b);
    outputs(1740) <= a xor b;
    outputs(1741) <= not a;
    outputs(1742) <= a xor b;
    outputs(1743) <= not a;
    outputs(1744) <= not (a or b);
    outputs(1745) <= a xor b;
    outputs(1746) <= a and not b;
    outputs(1747) <= a;
    outputs(1748) <= not b;
    outputs(1749) <= a;
    outputs(1750) <= not (a xor b);
    outputs(1751) <= a and not b;
    outputs(1752) <= not a or b;
    outputs(1753) <= a xor b;
    outputs(1754) <= a and b;
    outputs(1755) <= b;
    outputs(1756) <= b and not a;
    outputs(1757) <= b;
    outputs(1758) <= a xor b;
    outputs(1759) <= a xor b;
    outputs(1760) <= a and not b;
    outputs(1761) <= a and b;
    outputs(1762) <= a;
    outputs(1763) <= not a;
    outputs(1764) <= not a;
    outputs(1765) <= a;
    outputs(1766) <= a and b;
    outputs(1767) <= not (a or b);
    outputs(1768) <= b;
    outputs(1769) <= a xor b;
    outputs(1770) <= not a;
    outputs(1771) <= a xor b;
    outputs(1772) <= not (a xor b);
    outputs(1773) <= not (a or b);
    outputs(1774) <= not (a xor b);
    outputs(1775) <= a;
    outputs(1776) <= b and not a;
    outputs(1777) <= a xor b;
    outputs(1778) <= b;
    outputs(1779) <= not (a or b);
    outputs(1780) <= a;
    outputs(1781) <= b;
    outputs(1782) <= not b or a;
    outputs(1783) <= not (a xor b);
    outputs(1784) <= a xor b;
    outputs(1785) <= a;
    outputs(1786) <= a;
    outputs(1787) <= not b;
    outputs(1788) <= not b;
    outputs(1789) <= b and not a;
    outputs(1790) <= a and b;
    outputs(1791) <= a;
    outputs(1792) <= a;
    outputs(1793) <= not (a xor b);
    outputs(1794) <= b;
    outputs(1795) <= not a;
    outputs(1796) <= a;
    outputs(1797) <= a;
    outputs(1798) <= a and b;
    outputs(1799) <= b;
    outputs(1800) <= not b or a;
    outputs(1801) <= a;
    outputs(1802) <= not (a xor b);
    outputs(1803) <= not a or b;
    outputs(1804) <= a xor b;
    outputs(1805) <= a xor b;
    outputs(1806) <= not (a or b);
    outputs(1807) <= a xor b;
    outputs(1808) <= a xor b;
    outputs(1809) <= a and b;
    outputs(1810) <= a;
    outputs(1811) <= not b;
    outputs(1812) <= not a;
    outputs(1813) <= a and b;
    outputs(1814) <= a;
    outputs(1815) <= a xor b;
    outputs(1816) <= a and not b;
    outputs(1817) <= a;
    outputs(1818) <= not b;
    outputs(1819) <= a and b;
    outputs(1820) <= a and b;
    outputs(1821) <= a;
    outputs(1822) <= a and b;
    outputs(1823) <= b and not a;
    outputs(1824) <= not a or b;
    outputs(1825) <= not (a or b);
    outputs(1826) <= not (a and b);
    outputs(1827) <= not a;
    outputs(1828) <= a and not b;
    outputs(1829) <= not (a xor b);
    outputs(1830) <= not a;
    outputs(1831) <= not (a xor b);
    outputs(1832) <= not (a xor b);
    outputs(1833) <= not b;
    outputs(1834) <= not (a xor b);
    outputs(1835) <= not (a xor b);
    outputs(1836) <= not a;
    outputs(1837) <= not a;
    outputs(1838) <= not b;
    outputs(1839) <= not (a xor b);
    outputs(1840) <= b;
    outputs(1841) <= not (a xor b);
    outputs(1842) <= not (a or b);
    outputs(1843) <= a;
    outputs(1844) <= not a;
    outputs(1845) <= a xor b;
    outputs(1846) <= not a;
    outputs(1847) <= not a;
    outputs(1848) <= not b;
    outputs(1849) <= a and b;
    outputs(1850) <= b and not a;
    outputs(1851) <= not (a xor b);
    outputs(1852) <= b and not a;
    outputs(1853) <= not (a or b);
    outputs(1854) <= a;
    outputs(1855) <= a xor b;
    outputs(1856) <= not (a and b);
    outputs(1857) <= not (a xor b);
    outputs(1858) <= not a;
    outputs(1859) <= not b;
    outputs(1860) <= not a;
    outputs(1861) <= not (a xor b);
    outputs(1862) <= b;
    outputs(1863) <= not b;
    outputs(1864) <= not a;
    outputs(1865) <= not b;
    outputs(1866) <= a;
    outputs(1867) <= a and b;
    outputs(1868) <= a and not b;
    outputs(1869) <= b and not a;
    outputs(1870) <= not a;
    outputs(1871) <= not (a xor b);
    outputs(1872) <= a and not b;
    outputs(1873) <= not a;
    outputs(1874) <= b and not a;
    outputs(1875) <= a and not b;
    outputs(1876) <= not (a xor b);
    outputs(1877) <= a xor b;
    outputs(1878) <= not (a xor b);
    outputs(1879) <= a or b;
    outputs(1880) <= a;
    outputs(1881) <= a xor b;
    outputs(1882) <= a xor b;
    outputs(1883) <= not (a xor b);
    outputs(1884) <= a or b;
    outputs(1885) <= a xor b;
    outputs(1886) <= a xor b;
    outputs(1887) <= not (a xor b);
    outputs(1888) <= a or b;
    outputs(1889) <= not a or b;
    outputs(1890) <= not b;
    outputs(1891) <= a;
    outputs(1892) <= a xor b;
    outputs(1893) <= a xor b;
    outputs(1894) <= a;
    outputs(1895) <= a xor b;
    outputs(1896) <= not (a xor b);
    outputs(1897) <= a;
    outputs(1898) <= a and b;
    outputs(1899) <= b and not a;
    outputs(1900) <= a and b;
    outputs(1901) <= not (a or b);
    outputs(1902) <= a and b;
    outputs(1903) <= b;
    outputs(1904) <= not b;
    outputs(1905) <= not (a xor b);
    outputs(1906) <= not (a and b);
    outputs(1907) <= not (a xor b);
    outputs(1908) <= b and not a;
    outputs(1909) <= not a;
    outputs(1910) <= b;
    outputs(1911) <= a;
    outputs(1912) <= b;
    outputs(1913) <= b and not a;
    outputs(1914) <= b;
    outputs(1915) <= a and b;
    outputs(1916) <= not b;
    outputs(1917) <= not a;
    outputs(1918) <= not b;
    outputs(1919) <= a and b;
    outputs(1920) <= a xor b;
    outputs(1921) <= not b;
    outputs(1922) <= a and b;
    outputs(1923) <= not b;
    outputs(1924) <= b;
    outputs(1925) <= a and b;
    outputs(1926) <= a xor b;
    outputs(1927) <= not (a xor b);
    outputs(1928) <= a;
    outputs(1929) <= not (a or b);
    outputs(1930) <= a xor b;
    outputs(1931) <= b and not a;
    outputs(1932) <= a xor b;
    outputs(1933) <= b;
    outputs(1934) <= not a;
    outputs(1935) <= a;
    outputs(1936) <= b;
    outputs(1937) <= b;
    outputs(1938) <= b and not a;
    outputs(1939) <= b;
    outputs(1940) <= b and not a;
    outputs(1941) <= not a;
    outputs(1942) <= a and b;
    outputs(1943) <= b;
    outputs(1944) <= not a;
    outputs(1945) <= a xor b;
    outputs(1946) <= not b;
    outputs(1947) <= a;
    outputs(1948) <= not a;
    outputs(1949) <= a xor b;
    outputs(1950) <= a and b;
    outputs(1951) <= not b;
    outputs(1952) <= not b;
    outputs(1953) <= a xor b;
    outputs(1954) <= a and b;
    outputs(1955) <= not b or a;
    outputs(1956) <= not (a xor b);
    outputs(1957) <= a xor b;
    outputs(1958) <= not (a or b);
    outputs(1959) <= not (a xor b);
    outputs(1960) <= not (a xor b);
    outputs(1961) <= not b;
    outputs(1962) <= not a;
    outputs(1963) <= b;
    outputs(1964) <= not (a xor b);
    outputs(1965) <= a xor b;
    outputs(1966) <= not (a or b);
    outputs(1967) <= not b;
    outputs(1968) <= not a;
    outputs(1969) <= not b;
    outputs(1970) <= b;
    outputs(1971) <= a;
    outputs(1972) <= b;
    outputs(1973) <= a or b;
    outputs(1974) <= not (a or b);
    outputs(1975) <= a;
    outputs(1976) <= b;
    outputs(1977) <= a;
    outputs(1978) <= '1';
    outputs(1979) <= a and not b;
    outputs(1980) <= not (a xor b);
    outputs(1981) <= b;
    outputs(1982) <= not a;
    outputs(1983) <= a xor b;
    outputs(1984) <= b;
    outputs(1985) <= not (a xor b);
    outputs(1986) <= not (a xor b);
    outputs(1987) <= not (a or b);
    outputs(1988) <= a;
    outputs(1989) <= a and not b;
    outputs(1990) <= not b;
    outputs(1991) <= a xor b;
    outputs(1992) <= a or b;
    outputs(1993) <= not a;
    outputs(1994) <= not (a xor b);
    outputs(1995) <= a and b;
    outputs(1996) <= a xor b;
    outputs(1997) <= not (a xor b);
    outputs(1998) <= not a;
    outputs(1999) <= b and not a;
    outputs(2000) <= b;
    outputs(2001) <= a and b;
    outputs(2002) <= a and not b;
    outputs(2003) <= a;
    outputs(2004) <= b;
    outputs(2005) <= a xor b;
    outputs(2006) <= not (a xor b);
    outputs(2007) <= not b;
    outputs(2008) <= b;
    outputs(2009) <= a or b;
    outputs(2010) <= a xor b;
    outputs(2011) <= not (a and b);
    outputs(2012) <= a;
    outputs(2013) <= not b;
    outputs(2014) <= not b;
    outputs(2015) <= b and not a;
    outputs(2016) <= a and b;
    outputs(2017) <= not (a xor b);
    outputs(2018) <= a and b;
    outputs(2019) <= b;
    outputs(2020) <= a xor b;
    outputs(2021) <= not (a xor b);
    outputs(2022) <= b and not a;
    outputs(2023) <= a xor b;
    outputs(2024) <= a xor b;
    outputs(2025) <= not a;
    outputs(2026) <= b;
    outputs(2027) <= a;
    outputs(2028) <= not (a and b);
    outputs(2029) <= not a;
    outputs(2030) <= not a;
    outputs(2031) <= not b;
    outputs(2032) <= b;
    outputs(2033) <= a xor b;
    outputs(2034) <= not (a or b);
    outputs(2035) <= b and not a;
    outputs(2036) <= b;
    outputs(2037) <= not b;
    outputs(2038) <= not (a xor b);
    outputs(2039) <= b and not a;
    outputs(2040) <= b and not a;
    outputs(2041) <= not (a xor b);
    outputs(2042) <= not (a or b);
    outputs(2043) <= a xor b;
    outputs(2044) <= not b;
    outputs(2045) <= not (a xor b);
    outputs(2046) <= not (a or b);
    outputs(2047) <= a xor b;
    outputs(2048) <= a and b;
    outputs(2049) <= not (a xor b);
    outputs(2050) <= a;
    outputs(2051) <= not (a or b);
    outputs(2052) <= not b;
    outputs(2053) <= b;
    outputs(2054) <= not (a xor b);
    outputs(2055) <= a or b;
    outputs(2056) <= a or b;
    outputs(2057) <= b;
    outputs(2058) <= a xor b;
    outputs(2059) <= not (a xor b);
    outputs(2060) <= b;
    outputs(2061) <= not (a xor b);
    outputs(2062) <= not (a xor b);
    outputs(2063) <= not (a xor b);
    outputs(2064) <= not b;
    outputs(2065) <= not (a or b);
    outputs(2066) <= not a;
    outputs(2067) <= a;
    outputs(2068) <= a xor b;
    outputs(2069) <= not a;
    outputs(2070) <= not (a and b);
    outputs(2071) <= b;
    outputs(2072) <= b;
    outputs(2073) <= not b;
    outputs(2074) <= a xor b;
    outputs(2075) <= a;
    outputs(2076) <= not (a xor b);
    outputs(2077) <= not a;
    outputs(2078) <= not (a or b);
    outputs(2079) <= not a;
    outputs(2080) <= not b;
    outputs(2081) <= a and not b;
    outputs(2082) <= not b;
    outputs(2083) <= b;
    outputs(2084) <= not b or a;
    outputs(2085) <= not (a xor b);
    outputs(2086) <= not b;
    outputs(2087) <= a xor b;
    outputs(2088) <= not b or a;
    outputs(2089) <= not a or b;
    outputs(2090) <= a;
    outputs(2091) <= a;
    outputs(2092) <= a and b;
    outputs(2093) <= not (a or b);
    outputs(2094) <= not a or b;
    outputs(2095) <= not a or b;
    outputs(2096) <= a xor b;
    outputs(2097) <= not b;
    outputs(2098) <= not (a xor b);
    outputs(2099) <= a xor b;
    outputs(2100) <= not b or a;
    outputs(2101) <= a;
    outputs(2102) <= not b;
    outputs(2103) <= not (a xor b);
    outputs(2104) <= not a;
    outputs(2105) <= a xor b;
    outputs(2106) <= not a;
    outputs(2107) <= not b;
    outputs(2108) <= a;
    outputs(2109) <= a xor b;
    outputs(2110) <= a xor b;
    outputs(2111) <= a xor b;
    outputs(2112) <= a;
    outputs(2113) <= b;
    outputs(2114) <= not b;
    outputs(2115) <= not a;
    outputs(2116) <= a;
    outputs(2117) <= a and b;
    outputs(2118) <= not (a or b);
    outputs(2119) <= not (a or b);
    outputs(2120) <= a xor b;
    outputs(2121) <= not a;
    outputs(2122) <= b and not a;
    outputs(2123) <= a;
    outputs(2124) <= not (a xor b);
    outputs(2125) <= not a or b;
    outputs(2126) <= not b;
    outputs(2127) <= not a;
    outputs(2128) <= a xor b;
    outputs(2129) <= a;
    outputs(2130) <= b;
    outputs(2131) <= a and b;
    outputs(2132) <= not (a xor b);
    outputs(2133) <= b;
    outputs(2134) <= a or b;
    outputs(2135) <= a and not b;
    outputs(2136) <= a;
    outputs(2137) <= a or b;
    outputs(2138) <= not a;
    outputs(2139) <= b;
    outputs(2140) <= not (a xor b);
    outputs(2141) <= not b;
    outputs(2142) <= not b;
    outputs(2143) <= b and not a;
    outputs(2144) <= a;
    outputs(2145) <= not (a xor b);
    outputs(2146) <= not a;
    outputs(2147) <= a;
    outputs(2148) <= not (a xor b);
    outputs(2149) <= a;
    outputs(2150) <= a;
    outputs(2151) <= not b;
    outputs(2152) <= not a;
    outputs(2153) <= a xor b;
    outputs(2154) <= not a or b;
    outputs(2155) <= not a;
    outputs(2156) <= not (a or b);
    outputs(2157) <= not a;
    outputs(2158) <= not (a xor b);
    outputs(2159) <= a xor b;
    outputs(2160) <= a xor b;
    outputs(2161) <= not (a xor b);
    outputs(2162) <= a;
    outputs(2163) <= not b;
    outputs(2164) <= a xor b;
    outputs(2165) <= a;
    outputs(2166) <= b;
    outputs(2167) <= not b;
    outputs(2168) <= not (a xor b);
    outputs(2169) <= not (a xor b);
    outputs(2170) <= b;
    outputs(2171) <= a xor b;
    outputs(2172) <= not (a xor b);
    outputs(2173) <= not (a and b);
    outputs(2174) <= b;
    outputs(2175) <= not a;
    outputs(2176) <= a xor b;
    outputs(2177) <= a xor b;
    outputs(2178) <= a xor b;
    outputs(2179) <= a xor b;
    outputs(2180) <= not b;
    outputs(2181) <= not (a xor b);
    outputs(2182) <= not (a and b);
    outputs(2183) <= not a;
    outputs(2184) <= not b;
    outputs(2185) <= not a or b;
    outputs(2186) <= a xor b;
    outputs(2187) <= b;
    outputs(2188) <= a xor b;
    outputs(2189) <= not a or b;
    outputs(2190) <= a and not b;
    outputs(2191) <= not b;
    outputs(2192) <= not a;
    outputs(2193) <= a;
    outputs(2194) <= not a or b;
    outputs(2195) <= b;
    outputs(2196) <= a;
    outputs(2197) <= not b;
    outputs(2198) <= not b or a;
    outputs(2199) <= not a or b;
    outputs(2200) <= not (a xor b);
    outputs(2201) <= a xor b;
    outputs(2202) <= not (a xor b);
    outputs(2203) <= b;
    outputs(2204) <= not a;
    outputs(2205) <= not (a xor b);
    outputs(2206) <= not (a xor b);
    outputs(2207) <= not b;
    outputs(2208) <= b;
    outputs(2209) <= b;
    outputs(2210) <= b;
    outputs(2211) <= not (a xor b);
    outputs(2212) <= not b;
    outputs(2213) <= not b;
    outputs(2214) <= a xor b;
    outputs(2215) <= a and not b;
    outputs(2216) <= a xor b;
    outputs(2217) <= a and not b;
    outputs(2218) <= not a;
    outputs(2219) <= a;
    outputs(2220) <= b;
    outputs(2221) <= a xor b;
    outputs(2222) <= not a;
    outputs(2223) <= not (a xor b);
    outputs(2224) <= not (a xor b);
    outputs(2225) <= b;
    outputs(2226) <= not (a xor b);
    outputs(2227) <= not (a xor b);
    outputs(2228) <= not a;
    outputs(2229) <= b;
    outputs(2230) <= not (a xor b);
    outputs(2231) <= a;
    outputs(2232) <= a;
    outputs(2233) <= b;
    outputs(2234) <= not b;
    outputs(2235) <= not a;
    outputs(2236) <= not a;
    outputs(2237) <= b;
    outputs(2238) <= a;
    outputs(2239) <= b;
    outputs(2240) <= a xor b;
    outputs(2241) <= a;
    outputs(2242) <= a xor b;
    outputs(2243) <= b;
    outputs(2244) <= b;
    outputs(2245) <= not a;
    outputs(2246) <= not (a and b);
    outputs(2247) <= not a or b;
    outputs(2248) <= not (a xor b);
    outputs(2249) <= not (a xor b);
    outputs(2250) <= b;
    outputs(2251) <= not a;
    outputs(2252) <= a xor b;
    outputs(2253) <= a xor b;
    outputs(2254) <= a xor b;
    outputs(2255) <= a xor b;
    outputs(2256) <= b and not a;
    outputs(2257) <= not b;
    outputs(2258) <= not b;
    outputs(2259) <= not a;
    outputs(2260) <= not b;
    outputs(2261) <= a;
    outputs(2262) <= not b;
    outputs(2263) <= a xor b;
    outputs(2264) <= not b;
    outputs(2265) <= not b or a;
    outputs(2266) <= not (a xor b);
    outputs(2267) <= not a;
    outputs(2268) <= not a;
    outputs(2269) <= not (a and b);
    outputs(2270) <= a;
    outputs(2271) <= b and not a;
    outputs(2272) <= a xor b;
    outputs(2273) <= a xor b;
    outputs(2274) <= not (a xor b);
    outputs(2275) <= a xor b;
    outputs(2276) <= a xor b;
    outputs(2277) <= not (a xor b);
    outputs(2278) <= a xor b;
    outputs(2279) <= a or b;
    outputs(2280) <= not a;
    outputs(2281) <= a;
    outputs(2282) <= not a;
    outputs(2283) <= not b;
    outputs(2284) <= not a;
    outputs(2285) <= not b or a;
    outputs(2286) <= a xor b;
    outputs(2287) <= not b;
    outputs(2288) <= not a;
    outputs(2289) <= b;
    outputs(2290) <= not a or b;
    outputs(2291) <= not (a xor b);
    outputs(2292) <= a xor b;
    outputs(2293) <= b;
    outputs(2294) <= not b;
    outputs(2295) <= not a;
    outputs(2296) <= a xor b;
    outputs(2297) <= a xor b;
    outputs(2298) <= not b;
    outputs(2299) <= not (a or b);
    outputs(2300) <= a;
    outputs(2301) <= not a;
    outputs(2302) <= b;
    outputs(2303) <= not a;
    outputs(2304) <= a or b;
    outputs(2305) <= not a;
    outputs(2306) <= not b;
    outputs(2307) <= a and b;
    outputs(2308) <= a;
    outputs(2309) <= a and not b;
    outputs(2310) <= not a;
    outputs(2311) <= not b or a;
    outputs(2312) <= a and not b;
    outputs(2313) <= not (a and b);
    outputs(2314) <= a xor b;
    outputs(2315) <= not b;
    outputs(2316) <= not b;
    outputs(2317) <= not (a xor b);
    outputs(2318) <= not b;
    outputs(2319) <= b and not a;
    outputs(2320) <= not (a and b);
    outputs(2321) <= b;
    outputs(2322) <= not b;
    outputs(2323) <= a xor b;
    outputs(2324) <= not b or a;
    outputs(2325) <= a xor b;
    outputs(2326) <= not b;
    outputs(2327) <= b and not a;
    outputs(2328) <= not b;
    outputs(2329) <= a;
    outputs(2330) <= not a or b;
    outputs(2331) <= not a;
    outputs(2332) <= b;
    outputs(2333) <= a and b;
    outputs(2334) <= not b;
    outputs(2335) <= a;
    outputs(2336) <= a;
    outputs(2337) <= a;
    outputs(2338) <= not b or a;
    outputs(2339) <= not (a xor b);
    outputs(2340) <= not (a xor b);
    outputs(2341) <= not b;
    outputs(2342) <= a;
    outputs(2343) <= a;
    outputs(2344) <= a xor b;
    outputs(2345) <= not (a and b);
    outputs(2346) <= b;
    outputs(2347) <= a;
    outputs(2348) <= not a;
    outputs(2349) <= not (a xor b);
    outputs(2350) <= not (a and b);
    outputs(2351) <= a;
    outputs(2352) <= not b;
    outputs(2353) <= not a;
    outputs(2354) <= not a;
    outputs(2355) <= not (a xor b);
    outputs(2356) <= not (a xor b);
    outputs(2357) <= not a;
    outputs(2358) <= not a;
    outputs(2359) <= a xor b;
    outputs(2360) <= a;
    outputs(2361) <= a xor b;
    outputs(2362) <= not (a xor b);
    outputs(2363) <= b;
    outputs(2364) <= a or b;
    outputs(2365) <= not a;
    outputs(2366) <= not b;
    outputs(2367) <= a xor b;
    outputs(2368) <= not (a and b);
    outputs(2369) <= a;
    outputs(2370) <= a xor b;
    outputs(2371) <= not (a and b);
    outputs(2372) <= not b;
    outputs(2373) <= not a or b;
    outputs(2374) <= not (a xor b);
    outputs(2375) <= not (a xor b);
    outputs(2376) <= not b or a;
    outputs(2377) <= not (a or b);
    outputs(2378) <= not a;
    outputs(2379) <= not (a and b);
    outputs(2380) <= not (a xor b);
    outputs(2381) <= not b;
    outputs(2382) <= not a;
    outputs(2383) <= b;
    outputs(2384) <= a;
    outputs(2385) <= not (a xor b);
    outputs(2386) <= a and not b;
    outputs(2387) <= b;
    outputs(2388) <= not b or a;
    outputs(2389) <= a;
    outputs(2390) <= a;
    outputs(2391) <= a;
    outputs(2392) <= not b;
    outputs(2393) <= a xor b;
    outputs(2394) <= not b;
    outputs(2395) <= a or b;
    outputs(2396) <= not (a and b);
    outputs(2397) <= not b;
    outputs(2398) <= not a;
    outputs(2399) <= a;
    outputs(2400) <= a xor b;
    outputs(2401) <= not b;
    outputs(2402) <= not a;
    outputs(2403) <= b;
    outputs(2404) <= b;
    outputs(2405) <= a xor b;
    outputs(2406) <= not a;
    outputs(2407) <= not b or a;
    outputs(2408) <= not b or a;
    outputs(2409) <= not a;
    outputs(2410) <= a and b;
    outputs(2411) <= not b;
    outputs(2412) <= not (a xor b);
    outputs(2413) <= not b;
    outputs(2414) <= b;
    outputs(2415) <= b;
    outputs(2416) <= a or b;
    outputs(2417) <= not (a and b);
    outputs(2418) <= not (a xor b);
    outputs(2419) <= a;
    outputs(2420) <= not (a xor b);
    outputs(2421) <= not (a xor b);
    outputs(2422) <= b and not a;
    outputs(2423) <= not (a xor b);
    outputs(2424) <= b and not a;
    outputs(2425) <= not a;
    outputs(2426) <= a and b;
    outputs(2427) <= a;
    outputs(2428) <= b and not a;
    outputs(2429) <= a;
    outputs(2430) <= not a or b;
    outputs(2431) <= b and not a;
    outputs(2432) <= b;
    outputs(2433) <= not (a xor b);
    outputs(2434) <= a;
    outputs(2435) <= a xor b;
    outputs(2436) <= a xor b;
    outputs(2437) <= not a;
    outputs(2438) <= not b;
    outputs(2439) <= not a or b;
    outputs(2440) <= not b;
    outputs(2441) <= not a;
    outputs(2442) <= a;
    outputs(2443) <= a or b;
    outputs(2444) <= a xor b;
    outputs(2445) <= a;
    outputs(2446) <= a and not b;
    outputs(2447) <= a;
    outputs(2448) <= not a;
    outputs(2449) <= a or b;
    outputs(2450) <= not (a xor b);
    outputs(2451) <= a or b;
    outputs(2452) <= not (a xor b);
    outputs(2453) <= a xor b;
    outputs(2454) <= a;
    outputs(2455) <= not a;
    outputs(2456) <= not b;
    outputs(2457) <= a xor b;
    outputs(2458) <= not b;
    outputs(2459) <= a xor b;
    outputs(2460) <= b and not a;
    outputs(2461) <= a xor b;
    outputs(2462) <= a or b;
    outputs(2463) <= not b or a;
    outputs(2464) <= a;
    outputs(2465) <= not (a xor b);
    outputs(2466) <= not a or b;
    outputs(2467) <= a or b;
    outputs(2468) <= a xor b;
    outputs(2469) <= b;
    outputs(2470) <= not (a xor b);
    outputs(2471) <= a and b;
    outputs(2472) <= not b;
    outputs(2473) <= not b or a;
    outputs(2474) <= not a or b;
    outputs(2475) <= a xor b;
    outputs(2476) <= not b;
    outputs(2477) <= b and not a;
    outputs(2478) <= a and not b;
    outputs(2479) <= not b or a;
    outputs(2480) <= b;
    outputs(2481) <= not b;
    outputs(2482) <= not a;
    outputs(2483) <= not (a xor b);
    outputs(2484) <= a xor b;
    outputs(2485) <= not a or b;
    outputs(2486) <= not a or b;
    outputs(2487) <= not b;
    outputs(2488) <= not (a xor b);
    outputs(2489) <= b;
    outputs(2490) <= not (a xor b);
    outputs(2491) <= a xor b;
    outputs(2492) <= b;
    outputs(2493) <= not (a xor b);
    outputs(2494) <= a;
    outputs(2495) <= not b;
    outputs(2496) <= a and not b;
    outputs(2497) <= not (a xor b);
    outputs(2498) <= b;
    outputs(2499) <= not a;
    outputs(2500) <= not (a and b);
    outputs(2501) <= a or b;
    outputs(2502) <= b;
    outputs(2503) <= a or b;
    outputs(2504) <= not a;
    outputs(2505) <= not a;
    outputs(2506) <= not b;
    outputs(2507) <= b;
    outputs(2508) <= not b;
    outputs(2509) <= not b or a;
    outputs(2510) <= not a;
    outputs(2511) <= not b;
    outputs(2512) <= a and b;
    outputs(2513) <= b and not a;
    outputs(2514) <= a xor b;
    outputs(2515) <= a and not b;
    outputs(2516) <= b;
    outputs(2517) <= a xor b;
    outputs(2518) <= not (a and b);
    outputs(2519) <= not (a xor b);
    outputs(2520) <= not (a xor b);
    outputs(2521) <= not a;
    outputs(2522) <= not b;
    outputs(2523) <= a;
    outputs(2524) <= a;
    outputs(2525) <= not (a xor b);
    outputs(2526) <= not (a xor b);
    outputs(2527) <= a xor b;
    outputs(2528) <= a;
    outputs(2529) <= not (a and b);
    outputs(2530) <= not a;
    outputs(2531) <= not a;
    outputs(2532) <= a;
    outputs(2533) <= not a or b;
    outputs(2534) <= a and b;
    outputs(2535) <= a;
    outputs(2536) <= '1';
    outputs(2537) <= a xor b;
    outputs(2538) <= not b or a;
    outputs(2539) <= a xor b;
    outputs(2540) <= not a or b;
    outputs(2541) <= not (a xor b);
    outputs(2542) <= a;
    outputs(2543) <= a;
    outputs(2544) <= b and not a;
    outputs(2545) <= not (a xor b);
    outputs(2546) <= not b;
    outputs(2547) <= a or b;
    outputs(2548) <= not (a xor b);
    outputs(2549) <= not a;
    outputs(2550) <= not b;
    outputs(2551) <= not b;
    outputs(2552) <= not (a and b);
    outputs(2553) <= a xor b;
    outputs(2554) <= a;
    outputs(2555) <= not (a xor b);
    outputs(2556) <= not a;
    outputs(2557) <= a and not b;
    outputs(2558) <= a xor b;
    outputs(2559) <= b;
    outputs(2560) <= a;
    outputs(2561) <= a xor b;
    outputs(2562) <= not b;
    outputs(2563) <= a xor b;
    outputs(2564) <= a;
    outputs(2565) <= not a;
    outputs(2566) <= a;
    outputs(2567) <= a xor b;
    outputs(2568) <= not b;
    outputs(2569) <= a;
    outputs(2570) <= a xor b;
    outputs(2571) <= b and not a;
    outputs(2572) <= not (a xor b);
    outputs(2573) <= a xor b;
    outputs(2574) <= a;
    outputs(2575) <= b;
    outputs(2576) <= not a;
    outputs(2577) <= b;
    outputs(2578) <= a and b;
    outputs(2579) <= not (a xor b);
    outputs(2580) <= b;
    outputs(2581) <= not b;
    outputs(2582) <= a;
    outputs(2583) <= not b;
    outputs(2584) <= a xor b;
    outputs(2585) <= not b or a;
    outputs(2586) <= a;
    outputs(2587) <= b;
    outputs(2588) <= b and not a;
    outputs(2589) <= not b or a;
    outputs(2590) <= not (a xor b);
    outputs(2591) <= not a;
    outputs(2592) <= not b;
    outputs(2593) <= not b or a;
    outputs(2594) <= a;
    outputs(2595) <= a;
    outputs(2596) <= a xor b;
    outputs(2597) <= b and not a;
    outputs(2598) <= a xor b;
    outputs(2599) <= a xor b;
    outputs(2600) <= a or b;
    outputs(2601) <= not b;
    outputs(2602) <= b;
    outputs(2603) <= not a or b;
    outputs(2604) <= not (a xor b);
    outputs(2605) <= a or b;
    outputs(2606) <= a xor b;
    outputs(2607) <= b;
    outputs(2608) <= a xor b;
    outputs(2609) <= a;
    outputs(2610) <= not (a xor b);
    outputs(2611) <= b;
    outputs(2612) <= b;
    outputs(2613) <= not (a xor b);
    outputs(2614) <= b;
    outputs(2615) <= not (a and b);
    outputs(2616) <= not b;
    outputs(2617) <= a and not b;
    outputs(2618) <= not b;
    outputs(2619) <= not b;
    outputs(2620) <= b;
    outputs(2621) <= not (a or b);
    outputs(2622) <= not (a xor b);
    outputs(2623) <= b;
    outputs(2624) <= not a;
    outputs(2625) <= a xor b;
    outputs(2626) <= a or b;
    outputs(2627) <= not a;
    outputs(2628) <= a;
    outputs(2629) <= not (a or b);
    outputs(2630) <= a;
    outputs(2631) <= not (a and b);
    outputs(2632) <= a xor b;
    outputs(2633) <= not (a and b);
    outputs(2634) <= b;
    outputs(2635) <= a and not b;
    outputs(2636) <= b;
    outputs(2637) <= not a;
    outputs(2638) <= a or b;
    outputs(2639) <= a and b;
    outputs(2640) <= a;
    outputs(2641) <= not (a xor b);
    outputs(2642) <= not b;
    outputs(2643) <= not (a or b);
    outputs(2644) <= a xor b;
    outputs(2645) <= not b;
    outputs(2646) <= a;
    outputs(2647) <= a or b;
    outputs(2648) <= not (a xor b);
    outputs(2649) <= not (a xor b);
    outputs(2650) <= not b or a;
    outputs(2651) <= not a;
    outputs(2652) <= b;
    outputs(2653) <= not b or a;
    outputs(2654) <= not (a xor b);
    outputs(2655) <= a;
    outputs(2656) <= b;
    outputs(2657) <= a;
    outputs(2658) <= a and b;
    outputs(2659) <= not b;
    outputs(2660) <= a;
    outputs(2661) <= a and b;
    outputs(2662) <= not (a and b);
    outputs(2663) <= not (a xor b);
    outputs(2664) <= b;
    outputs(2665) <= not a;
    outputs(2666) <= a;
    outputs(2667) <= a xor b;
    outputs(2668) <= not (a and b);
    outputs(2669) <= not (a xor b);
    outputs(2670) <= a and not b;
    outputs(2671) <= a;
    outputs(2672) <= not b;
    outputs(2673) <= b;
    outputs(2674) <= not (a xor b);
    outputs(2675) <= not (a xor b);
    outputs(2676) <= a;
    outputs(2677) <= a xor b;
    outputs(2678) <= not (a and b);
    outputs(2679) <= a;
    outputs(2680) <= not (a xor b);
    outputs(2681) <= not a;
    outputs(2682) <= not (a and b);
    outputs(2683) <= not b;
    outputs(2684) <= a xor b;
    outputs(2685) <= not a or b;
    outputs(2686) <= not a;
    outputs(2687) <= a or b;
    outputs(2688) <= not b;
    outputs(2689) <= not b;
    outputs(2690) <= a xor b;
    outputs(2691) <= not (a xor b);
    outputs(2692) <= not b;
    outputs(2693) <= a xor b;
    outputs(2694) <= b;
    outputs(2695) <= not (a xor b);
    outputs(2696) <= not (a xor b);
    outputs(2697) <= a xor b;
    outputs(2698) <= a;
    outputs(2699) <= a;
    outputs(2700) <= b;
    outputs(2701) <= not a;
    outputs(2702) <= b and not a;
    outputs(2703) <= not (a xor b);
    outputs(2704) <= not a;
    outputs(2705) <= not b;
    outputs(2706) <= a;
    outputs(2707) <= a;
    outputs(2708) <= not b;
    outputs(2709) <= not b or a;
    outputs(2710) <= a xor b;
    outputs(2711) <= not (a xor b);
    outputs(2712) <= a and b;
    outputs(2713) <= a xor b;
    outputs(2714) <= not (a and b);
    outputs(2715) <= a or b;
    outputs(2716) <= not b;
    outputs(2717) <= a xor b;
    outputs(2718) <= not b or a;
    outputs(2719) <= not (a xor b);
    outputs(2720) <= a;
    outputs(2721) <= b;
    outputs(2722) <= not (a xor b);
    outputs(2723) <= b and not a;
    outputs(2724) <= b;
    outputs(2725) <= a;
    outputs(2726) <= a and not b;
    outputs(2727) <= a;
    outputs(2728) <= b;
    outputs(2729) <= a;
    outputs(2730) <= not a;
    outputs(2731) <= a xor b;
    outputs(2732) <= a xor b;
    outputs(2733) <= b;
    outputs(2734) <= a xor b;
    outputs(2735) <= not a;
    outputs(2736) <= a xor b;
    outputs(2737) <= b;
    outputs(2738) <= b;
    outputs(2739) <= not a;
    outputs(2740) <= a;
    outputs(2741) <= not (a xor b);
    outputs(2742) <= b;
    outputs(2743) <= a;
    outputs(2744) <= a;
    outputs(2745) <= b;
    outputs(2746) <= b;
    outputs(2747) <= a xor b;
    outputs(2748) <= a;
    outputs(2749) <= not (a xor b);
    outputs(2750) <= a or b;
    outputs(2751) <= not (a xor b);
    outputs(2752) <= a xor b;
    outputs(2753) <= a;
    outputs(2754) <= not b;
    outputs(2755) <= not b;
    outputs(2756) <= a;
    outputs(2757) <= b;
    outputs(2758) <= b;
    outputs(2759) <= not (a xor b);
    outputs(2760) <= not a or b;
    outputs(2761) <= b;
    outputs(2762) <= not b;
    outputs(2763) <= b;
    outputs(2764) <= not (a xor b);
    outputs(2765) <= b;
    outputs(2766) <= a or b;
    outputs(2767) <= not (a xor b);
    outputs(2768) <= a xor b;
    outputs(2769) <= b and not a;
    outputs(2770) <= not b;
    outputs(2771) <= not b or a;
    outputs(2772) <= not a;
    outputs(2773) <= a xor b;
    outputs(2774) <= a;
    outputs(2775) <= not b or a;
    outputs(2776) <= a and b;
    outputs(2777) <= not (a and b);
    outputs(2778) <= not (a xor b);
    outputs(2779) <= a;
    outputs(2780) <= b;
    outputs(2781) <= a xor b;
    outputs(2782) <= not b;
    outputs(2783) <= a xor b;
    outputs(2784) <= not a;
    outputs(2785) <= not (a xor b);
    outputs(2786) <= not b or a;
    outputs(2787) <= not (a xor b);
    outputs(2788) <= a xor b;
    outputs(2789) <= a;
    outputs(2790) <= not b;
    outputs(2791) <= a;
    outputs(2792) <= not a;
    outputs(2793) <= a xor b;
    outputs(2794) <= not a;
    outputs(2795) <= b;
    outputs(2796) <= a xor b;
    outputs(2797) <= not a;
    outputs(2798) <= a xor b;
    outputs(2799) <= not (a xor b);
    outputs(2800) <= not (a and b);
    outputs(2801) <= a or b;
    outputs(2802) <= not b;
    outputs(2803) <= not a;
    outputs(2804) <= a xor b;
    outputs(2805) <= b;
    outputs(2806) <= not b;
    outputs(2807) <= a xor b;
    outputs(2808) <= a xor b;
    outputs(2809) <= a and b;
    outputs(2810) <= not a;
    outputs(2811) <= a and b;
    outputs(2812) <= a and b;
    outputs(2813) <= not b;
    outputs(2814) <= a;
    outputs(2815) <= not b;
    outputs(2816) <= a;
    outputs(2817) <= not (a xor b);
    outputs(2818) <= a and b;
    outputs(2819) <= not a or b;
    outputs(2820) <= not b;
    outputs(2821) <= a or b;
    outputs(2822) <= b and not a;
    outputs(2823) <= not (a xor b);
    outputs(2824) <= a;
    outputs(2825) <= not (a xor b);
    outputs(2826) <= a xor b;
    outputs(2827) <= not b;
    outputs(2828) <= not (a xor b);
    outputs(2829) <= not b;
    outputs(2830) <= not a or b;
    outputs(2831) <= a xor b;
    outputs(2832) <= b;
    outputs(2833) <= not b;
    outputs(2834) <= not (a xor b);
    outputs(2835) <= not (a xor b);
    outputs(2836) <= b;
    outputs(2837) <= not a or b;
    outputs(2838) <= a;
    outputs(2839) <= a;
    outputs(2840) <= not a;
    outputs(2841) <= b;
    outputs(2842) <= a xor b;
    outputs(2843) <= not a;
    outputs(2844) <= b;
    outputs(2845) <= a xor b;
    outputs(2846) <= a;
    outputs(2847) <= a and b;
    outputs(2848) <= not (a xor b);
    outputs(2849) <= not (a xor b);
    outputs(2850) <= not (a or b);
    outputs(2851) <= a;
    outputs(2852) <= a xor b;
    outputs(2853) <= a and b;
    outputs(2854) <= b;
    outputs(2855) <= not b;
    outputs(2856) <= not a or b;
    outputs(2857) <= not (a and b);
    outputs(2858) <= not (a and b);
    outputs(2859) <= a xor b;
    outputs(2860) <= not (a xor b);
    outputs(2861) <= not b;
    outputs(2862) <= not b;
    outputs(2863) <= a xor b;
    outputs(2864) <= not b;
    outputs(2865) <= not b;
    outputs(2866) <= not b;
    outputs(2867) <= not (a xor b);
    outputs(2868) <= b;
    outputs(2869) <= a xor b;
    outputs(2870) <= a and not b;
    outputs(2871) <= not b or a;
    outputs(2872) <= not a;
    outputs(2873) <= a;
    outputs(2874) <= a;
    outputs(2875) <= not a;
    outputs(2876) <= not (a and b);
    outputs(2877) <= a or b;
    outputs(2878) <= a xor b;
    outputs(2879) <= not (a and b);
    outputs(2880) <= a xor b;
    outputs(2881) <= not a or b;
    outputs(2882) <= a;
    outputs(2883) <= not b or a;
    outputs(2884) <= not a;
    outputs(2885) <= not b or a;
    outputs(2886) <= not (a xor b);
    outputs(2887) <= a;
    outputs(2888) <= a;
    outputs(2889) <= not b;
    outputs(2890) <= not (a and b);
    outputs(2891) <= a and not b;
    outputs(2892) <= a xor b;
    outputs(2893) <= not (a or b);
    outputs(2894) <= not a or b;
    outputs(2895) <= a xor b;
    outputs(2896) <= a xor b;
    outputs(2897) <= not b;
    outputs(2898) <= a and not b;
    outputs(2899) <= a and not b;
    outputs(2900) <= b;
    outputs(2901) <= a;
    outputs(2902) <= not b;
    outputs(2903) <= not (a xor b);
    outputs(2904) <= a;
    outputs(2905) <= a;
    outputs(2906) <= not b or a;
    outputs(2907) <= not b;
    outputs(2908) <= not a or b;
    outputs(2909) <= b;
    outputs(2910) <= a xor b;
    outputs(2911) <= not (a xor b);
    outputs(2912) <= a xor b;
    outputs(2913) <= a xor b;
    outputs(2914) <= not (a xor b);
    outputs(2915) <= a xor b;
    outputs(2916) <= b and not a;
    outputs(2917) <= not b or a;
    outputs(2918) <= b;
    outputs(2919) <= not a;
    outputs(2920) <= not b or a;
    outputs(2921) <= not (a xor b);
    outputs(2922) <= not a;
    outputs(2923) <= a;
    outputs(2924) <= a;
    outputs(2925) <= a xor b;
    outputs(2926) <= a;
    outputs(2927) <= a xor b;
    outputs(2928) <= a xor b;
    outputs(2929) <= a;
    outputs(2930) <= a xor b;
    outputs(2931) <= not (a and b);
    outputs(2932) <= a and not b;
    outputs(2933) <= not b;
    outputs(2934) <= a xor b;
    outputs(2935) <= not (a xor b);
    outputs(2936) <= a or b;
    outputs(2937) <= a or b;
    outputs(2938) <= not (a xor b);
    outputs(2939) <= a;
    outputs(2940) <= a and b;
    outputs(2941) <= not b or a;
    outputs(2942) <= a xor b;
    outputs(2943) <= not b;
    outputs(2944) <= not a;
    outputs(2945) <= b and not a;
    outputs(2946) <= a or b;
    outputs(2947) <= b and not a;
    outputs(2948) <= a xor b;
    outputs(2949) <= not a or b;
    outputs(2950) <= not b;
    outputs(2951) <= not b or a;
    outputs(2952) <= a xor b;
    outputs(2953) <= not (a and b);
    outputs(2954) <= not (a xor b);
    outputs(2955) <= a or b;
    outputs(2956) <= not b;
    outputs(2957) <= a xor b;
    outputs(2958) <= b;
    outputs(2959) <= a xor b;
    outputs(2960) <= a xor b;
    outputs(2961) <= b;
    outputs(2962) <= b;
    outputs(2963) <= not b;
    outputs(2964) <= not (a or b);
    outputs(2965) <= a xor b;
    outputs(2966) <= a xor b;
    outputs(2967) <= not a or b;
    outputs(2968) <= not a;
    outputs(2969) <= a;
    outputs(2970) <= not b;
    outputs(2971) <= not (a xor b);
    outputs(2972) <= not (a xor b);
    outputs(2973) <= not (a xor b);
    outputs(2974) <= b;
    outputs(2975) <= a;
    outputs(2976) <= not (a xor b);
    outputs(2977) <= b;
    outputs(2978) <= not (a or b);
    outputs(2979) <= a;
    outputs(2980) <= not b or a;
    outputs(2981) <= not a;
    outputs(2982) <= not b;
    outputs(2983) <= b;
    outputs(2984) <= not b or a;
    outputs(2985) <= a and not b;
    outputs(2986) <= a;
    outputs(2987) <= not (a xor b);
    outputs(2988) <= a xor b;
    outputs(2989) <= a;
    outputs(2990) <= not a;
    outputs(2991) <= b;
    outputs(2992) <= a xor b;
    outputs(2993) <= a xor b;
    outputs(2994) <= not b;
    outputs(2995) <= not (a xor b);
    outputs(2996) <= not (a xor b);
    outputs(2997) <= not (a xor b);
    outputs(2998) <= a xor b;
    outputs(2999) <= not (a or b);
    outputs(3000) <= not a;
    outputs(3001) <= a xor b;
    outputs(3002) <= not b;
    outputs(3003) <= not (a xor b);
    outputs(3004) <= a xor b;
    outputs(3005) <= not (a xor b);
    outputs(3006) <= not b;
    outputs(3007) <= not (a or b);
    outputs(3008) <= not a;
    outputs(3009) <= not a;
    outputs(3010) <= b;
    outputs(3011) <= not b or a;
    outputs(3012) <= not a;
    outputs(3013) <= a xor b;
    outputs(3014) <= a xor b;
    outputs(3015) <= not b or a;
    outputs(3016) <= b and not a;
    outputs(3017) <= not (a or b);
    outputs(3018) <= not (a xor b);
    outputs(3019) <= not b;
    outputs(3020) <= b and not a;
    outputs(3021) <= b;
    outputs(3022) <= not (a or b);
    outputs(3023) <= not b;
    outputs(3024) <= a;
    outputs(3025) <= not b or a;
    outputs(3026) <= not (a xor b);
    outputs(3027) <= not (a xor b);
    outputs(3028) <= a and b;
    outputs(3029) <= not (a xor b);
    outputs(3030) <= b;
    outputs(3031) <= b;
    outputs(3032) <= a;
    outputs(3033) <= not a;
    outputs(3034) <= not a;
    outputs(3035) <= not (a xor b);
    outputs(3036) <= not b;
    outputs(3037) <= b;
    outputs(3038) <= a xor b;
    outputs(3039) <= not b;
    outputs(3040) <= b;
    outputs(3041) <= not (a xor b);
    outputs(3042) <= not a;
    outputs(3043) <= not (a xor b);
    outputs(3044) <= a xor b;
    outputs(3045) <= not (a or b);
    outputs(3046) <= not (a xor b);
    outputs(3047) <= not b;
    outputs(3048) <= not a or b;
    outputs(3049) <= not (a xor b);
    outputs(3050) <= not a;
    outputs(3051) <= b;
    outputs(3052) <= not (a xor b);
    outputs(3053) <= not b;
    outputs(3054) <= a;
    outputs(3055) <= b;
    outputs(3056) <= a or b;
    outputs(3057) <= a xor b;
    outputs(3058) <= not (a xor b);
    outputs(3059) <= not b;
    outputs(3060) <= not a or b;
    outputs(3061) <= not a;
    outputs(3062) <= not a;
    outputs(3063) <= a xor b;
    outputs(3064) <= b;
    outputs(3065) <= a;
    outputs(3066) <= not a;
    outputs(3067) <= a;
    outputs(3068) <= not (a and b);
    outputs(3069) <= b;
    outputs(3070) <= not a;
    outputs(3071) <= not a;
    outputs(3072) <= a;
    outputs(3073) <= not a;
    outputs(3074) <= not (a xor b);
    outputs(3075) <= a xor b;
    outputs(3076) <= a;
    outputs(3077) <= not a;
    outputs(3078) <= not (a and b);
    outputs(3079) <= a or b;
    outputs(3080) <= a and not b;
    outputs(3081) <= not b;
    outputs(3082) <= not b;
    outputs(3083) <= not b or a;
    outputs(3084) <= a;
    outputs(3085) <= a;
    outputs(3086) <= a or b;
    outputs(3087) <= not b;
    outputs(3088) <= a and not b;
    outputs(3089) <= a and b;
    outputs(3090) <= not b or a;
    outputs(3091) <= not (a xor b);
    outputs(3092) <= b;
    outputs(3093) <= not (a xor b);
    outputs(3094) <= b;
    outputs(3095) <= not (a xor b);
    outputs(3096) <= not (a xor b);
    outputs(3097) <= b and not a;
    outputs(3098) <= a and not b;
    outputs(3099) <= not b;
    outputs(3100) <= not (a xor b);
    outputs(3101) <= a and not b;
    outputs(3102) <= not b;
    outputs(3103) <= not (a xor b);
    outputs(3104) <= not (a xor b);
    outputs(3105) <= not (a xor b);
    outputs(3106) <= not b;
    outputs(3107) <= not a;
    outputs(3108) <= a;
    outputs(3109) <= a xor b;
    outputs(3110) <= a;
    outputs(3111) <= a xor b;
    outputs(3112) <= not b;
    outputs(3113) <= not (a or b);
    outputs(3114) <= a and not b;
    outputs(3115) <= not a;
    outputs(3116) <= not b;
    outputs(3117) <= not (a or b);
    outputs(3118) <= not b;
    outputs(3119) <= not b;
    outputs(3120) <= not b;
    outputs(3121) <= not (a xor b);
    outputs(3122) <= b;
    outputs(3123) <= a xor b;
    outputs(3124) <= not b or a;
    outputs(3125) <= b;
    outputs(3126) <= a and not b;
    outputs(3127) <= a xor b;
    outputs(3128) <= b and not a;
    outputs(3129) <= a or b;
    outputs(3130) <= b;
    outputs(3131) <= b and not a;
    outputs(3132) <= not (a xor b);
    outputs(3133) <= b;
    outputs(3134) <= b;
    outputs(3135) <= not b;
    outputs(3136) <= not a;
    outputs(3137) <= not (a and b);
    outputs(3138) <= b;
    outputs(3139) <= a xor b;
    outputs(3140) <= a xor b;
    outputs(3141) <= a xor b;
    outputs(3142) <= not b;
    outputs(3143) <= a xor b;
    outputs(3144) <= a xor b;
    outputs(3145) <= a xor b;
    outputs(3146) <= b and not a;
    outputs(3147) <= not (a or b);
    outputs(3148) <= not a or b;
    outputs(3149) <= a xor b;
    outputs(3150) <= not a;
    outputs(3151) <= not a;
    outputs(3152) <= not a or b;
    outputs(3153) <= a;
    outputs(3154) <= a and not b;
    outputs(3155) <= a xor b;
    outputs(3156) <= a;
    outputs(3157) <= not a;
    outputs(3158) <= b;
    outputs(3159) <= not a;
    outputs(3160) <= b;
    outputs(3161) <= not (a xor b);
    outputs(3162) <= b and not a;
    outputs(3163) <= b;
    outputs(3164) <= not (a and b);
    outputs(3165) <= a or b;
    outputs(3166) <= not (a and b);
    outputs(3167) <= not (a xor b);
    outputs(3168) <= b;
    outputs(3169) <= a;
    outputs(3170) <= not (a xor b);
    outputs(3171) <= a;
    outputs(3172) <= a xor b;
    outputs(3173) <= not a or b;
    outputs(3174) <= not (a xor b);
    outputs(3175) <= a;
    outputs(3176) <= a and not b;
    outputs(3177) <= a and not b;
    outputs(3178) <= not a or b;
    outputs(3179) <= not a;
    outputs(3180) <= a;
    outputs(3181) <= not b or a;
    outputs(3182) <= a xor b;
    outputs(3183) <= a;
    outputs(3184) <= a xor b;
    outputs(3185) <= not (a xor b);
    outputs(3186) <= not (a and b);
    outputs(3187) <= not a;
    outputs(3188) <= a xor b;
    outputs(3189) <= not (a xor b);
    outputs(3190) <= a xor b;
    outputs(3191) <= not b;
    outputs(3192) <= not a;
    outputs(3193) <= a xor b;
    outputs(3194) <= a and b;
    outputs(3195) <= not b;
    outputs(3196) <= a or b;
    outputs(3197) <= not b;
    outputs(3198) <= a xor b;
    outputs(3199) <= not a;
    outputs(3200) <= a and not b;
    outputs(3201) <= not b or a;
    outputs(3202) <= a xor b;
    outputs(3203) <= not (a xor b);
    outputs(3204) <= a and not b;
    outputs(3205) <= not b;
    outputs(3206) <= a and b;
    outputs(3207) <= a or b;
    outputs(3208) <= a;
    outputs(3209) <= a xor b;
    outputs(3210) <= b;
    outputs(3211) <= not a;
    outputs(3212) <= a;
    outputs(3213) <= a and not b;
    outputs(3214) <= a;
    outputs(3215) <= b;
    outputs(3216) <= a and not b;
    outputs(3217) <= a and b;
    outputs(3218) <= not (a xor b);
    outputs(3219) <= not (a xor b);
    outputs(3220) <= not (a and b);
    outputs(3221) <= not b;
    outputs(3222) <= not (a xor b);
    outputs(3223) <= not (a xor b);
    outputs(3224) <= not a;
    outputs(3225) <= not (a xor b);
    outputs(3226) <= not a;
    outputs(3227) <= b;
    outputs(3228) <= b;
    outputs(3229) <= not b or a;
    outputs(3230) <= a and b;
    outputs(3231) <= a and not b;
    outputs(3232) <= not a;
    outputs(3233) <= a;
    outputs(3234) <= b;
    outputs(3235) <= a xor b;
    outputs(3236) <= a xor b;
    outputs(3237) <= not (a xor b);
    outputs(3238) <= b;
    outputs(3239) <= not (a xor b);
    outputs(3240) <= not b;
    outputs(3241) <= not (a or b);
    outputs(3242) <= b;
    outputs(3243) <= not b or a;
    outputs(3244) <= not b;
    outputs(3245) <= not a;
    outputs(3246) <= a;
    outputs(3247) <= a xor b;
    outputs(3248) <= not (a xor b);
    outputs(3249) <= not b;
    outputs(3250) <= not (a xor b);
    outputs(3251) <= b and not a;
    outputs(3252) <= a;
    outputs(3253) <= b;
    outputs(3254) <= a xor b;
    outputs(3255) <= a;
    outputs(3256) <= a and b;
    outputs(3257) <= not a or b;
    outputs(3258) <= b;
    outputs(3259) <= b and not a;
    outputs(3260) <= not (a and b);
    outputs(3261) <= b;
    outputs(3262) <= a xor b;
    outputs(3263) <= b and not a;
    outputs(3264) <= a and not b;
    outputs(3265) <= not (a xor b);
    outputs(3266) <= not (a xor b);
    outputs(3267) <= b;
    outputs(3268) <= not a or b;
    outputs(3269) <= a;
    outputs(3270) <= a;
    outputs(3271) <= not a;
    outputs(3272) <= not b;
    outputs(3273) <= a or b;
    outputs(3274) <= a and b;
    outputs(3275) <= b;
    outputs(3276) <= not (a xor b);
    outputs(3277) <= not a or b;
    outputs(3278) <= a;
    outputs(3279) <= a and b;
    outputs(3280) <= not (a and b);
    outputs(3281) <= b and not a;
    outputs(3282) <= not b;
    outputs(3283) <= b;
    outputs(3284) <= a;
    outputs(3285) <= b;
    outputs(3286) <= b;
    outputs(3287) <= not (a xor b);
    outputs(3288) <= not (a xor b);
    outputs(3289) <= a or b;
    outputs(3290) <= not (a or b);
    outputs(3291) <= not (a and b);
    outputs(3292) <= b;
    outputs(3293) <= a and b;
    outputs(3294) <= not a or b;
    outputs(3295) <= a;
    outputs(3296) <= a and not b;
    outputs(3297) <= b;
    outputs(3298) <= not (a and b);
    outputs(3299) <= not b;
    outputs(3300) <= a or b;
    outputs(3301) <= not b;
    outputs(3302) <= not b;
    outputs(3303) <= not b;
    outputs(3304) <= b;
    outputs(3305) <= b;
    outputs(3306) <= a xor b;
    outputs(3307) <= a or b;
    outputs(3308) <= not b;
    outputs(3309) <= b;
    outputs(3310) <= a;
    outputs(3311) <= a;
    outputs(3312) <= a xor b;
    outputs(3313) <= not a or b;
    outputs(3314) <= a xor b;
    outputs(3315) <= b;
    outputs(3316) <= a;
    outputs(3317) <= not (a or b);
    outputs(3318) <= b;
    outputs(3319) <= a;
    outputs(3320) <= a and b;
    outputs(3321) <= not (a xor b);
    outputs(3322) <= a and not b;
    outputs(3323) <= not (a xor b);
    outputs(3324) <= not a or b;
    outputs(3325) <= not a or b;
    outputs(3326) <= a;
    outputs(3327) <= a;
    outputs(3328) <= a and b;
    outputs(3329) <= not a;
    outputs(3330) <= b;
    outputs(3331) <= a;
    outputs(3332) <= not a;
    outputs(3333) <= a xor b;
    outputs(3334) <= a;
    outputs(3335) <= a and not b;
    outputs(3336) <= a;
    outputs(3337) <= not (a xor b);
    outputs(3338) <= a xor b;
    outputs(3339) <= a xor b;
    outputs(3340) <= a and not b;
    outputs(3341) <= a xor b;
    outputs(3342) <= a and b;
    outputs(3343) <= not (a xor b);
    outputs(3344) <= not (a and b);
    outputs(3345) <= a and b;
    outputs(3346) <= not (a or b);
    outputs(3347) <= not (a xor b);
    outputs(3348) <= not b;
    outputs(3349) <= not a;
    outputs(3350) <= not (a xor b);
    outputs(3351) <= a;
    outputs(3352) <= b;
    outputs(3353) <= not (a xor b);
    outputs(3354) <= not b or a;
    outputs(3355) <= not (a and b);
    outputs(3356) <= b and not a;
    outputs(3357) <= b;
    outputs(3358) <= a;
    outputs(3359) <= a;
    outputs(3360) <= a and b;
    outputs(3361) <= not b or a;
    outputs(3362) <= a;
    outputs(3363) <= b and not a;
    outputs(3364) <= not a or b;
    outputs(3365) <= a xor b;
    outputs(3366) <= not a;
    outputs(3367) <= not (a xor b);
    outputs(3368) <= a and not b;
    outputs(3369) <= a;
    outputs(3370) <= not b;
    outputs(3371) <= not (a xor b);
    outputs(3372) <= not a;
    outputs(3373) <= not a;
    outputs(3374) <= a xor b;
    outputs(3375) <= not a;
    outputs(3376) <= not b;
    outputs(3377) <= a xor b;
    outputs(3378) <= b;
    outputs(3379) <= not b;
    outputs(3380) <= a and not b;
    outputs(3381) <= b;
    outputs(3382) <= not (a xor b);
    outputs(3383) <= a and b;
    outputs(3384) <= not (a xor b);
    outputs(3385) <= not a or b;
    outputs(3386) <= a xor b;
    outputs(3387) <= not a;
    outputs(3388) <= b;
    outputs(3389) <= a xor b;
    outputs(3390) <= a;
    outputs(3391) <= not a or b;
    outputs(3392) <= a xor b;
    outputs(3393) <= not (a xor b);
    outputs(3394) <= a xor b;
    outputs(3395) <= b and not a;
    outputs(3396) <= a or b;
    outputs(3397) <= not (a xor b);
    outputs(3398) <= not (a xor b);
    outputs(3399) <= a xor b;
    outputs(3400) <= a and not b;
    outputs(3401) <= a;
    outputs(3402) <= b;
    outputs(3403) <= not b;
    outputs(3404) <= not b;
    outputs(3405) <= b;
    outputs(3406) <= not (a xor b);
    outputs(3407) <= b;
    outputs(3408) <= not (a or b);
    outputs(3409) <= b;
    outputs(3410) <= a xor b;
    outputs(3411) <= not a;
    outputs(3412) <= a;
    outputs(3413) <= a;
    outputs(3414) <= not a;
    outputs(3415) <= a xor b;
    outputs(3416) <= not a or b;
    outputs(3417) <= not a;
    outputs(3418) <= not (a and b);
    outputs(3419) <= a and not b;
    outputs(3420) <= a xor b;
    outputs(3421) <= b;
    outputs(3422) <= not (a xor b);
    outputs(3423) <= a xor b;
    outputs(3424) <= b;
    outputs(3425) <= not a;
    outputs(3426) <= b;
    outputs(3427) <= a xor b;
    outputs(3428) <= a and b;
    outputs(3429) <= b;
    outputs(3430) <= not b;
    outputs(3431) <= a and b;
    outputs(3432) <= b;
    outputs(3433) <= not (a xor b);
    outputs(3434) <= not a;
    outputs(3435) <= not a;
    outputs(3436) <= not b;
    outputs(3437) <= not b;
    outputs(3438) <= a;
    outputs(3439) <= a xor b;
    outputs(3440) <= not (a xor b);
    outputs(3441) <= a;
    outputs(3442) <= b;
    outputs(3443) <= not a or b;
    outputs(3444) <= b and not a;
    outputs(3445) <= not b;
    outputs(3446) <= a;
    outputs(3447) <= a xor b;
    outputs(3448) <= not b;
    outputs(3449) <= not (a xor b);
    outputs(3450) <= not a;
    outputs(3451) <= not (a xor b);
    outputs(3452) <= not b;
    outputs(3453) <= a;
    outputs(3454) <= not (a xor b);
    outputs(3455) <= not a;
    outputs(3456) <= not b;
    outputs(3457) <= not a;
    outputs(3458) <= not (a xor b);
    outputs(3459) <= not a;
    outputs(3460) <= not (a and b);
    outputs(3461) <= a and b;
    outputs(3462) <= a;
    outputs(3463) <= b;
    outputs(3464) <= not b or a;
    outputs(3465) <= not (a or b);
    outputs(3466) <= b;
    outputs(3467) <= a and not b;
    outputs(3468) <= not b;
    outputs(3469) <= not (a xor b);
    outputs(3470) <= b;
    outputs(3471) <= a xor b;
    outputs(3472) <= b;
    outputs(3473) <= a;
    outputs(3474) <= not b;
    outputs(3475) <= not b;
    outputs(3476) <= not (a xor b);
    outputs(3477) <= b;
    outputs(3478) <= a and b;
    outputs(3479) <= not (a xor b);
    outputs(3480) <= a and not b;
    outputs(3481) <= not (a or b);
    outputs(3482) <= not (a xor b);
    outputs(3483) <= not b;
    outputs(3484) <= a;
    outputs(3485) <= a xor b;
    outputs(3486) <= a xor b;
    outputs(3487) <= not (a xor b);
    outputs(3488) <= b and not a;
    outputs(3489) <= not a;
    outputs(3490) <= not b;
    outputs(3491) <= a;
    outputs(3492) <= b;
    outputs(3493) <= not a;
    outputs(3494) <= b;
    outputs(3495) <= not b or a;
    outputs(3496) <= not (a and b);
    outputs(3497) <= a and b;
    outputs(3498) <= not a or b;
    outputs(3499) <= a xor b;
    outputs(3500) <= a xor b;
    outputs(3501) <= a;
    outputs(3502) <= a xor b;
    outputs(3503) <= not (a xor b);
    outputs(3504) <= not b;
    outputs(3505) <= not b;
    outputs(3506) <= not (a xor b);
    outputs(3507) <= not (a xor b);
    outputs(3508) <= not a or b;
    outputs(3509) <= b;
    outputs(3510) <= not a;
    outputs(3511) <= not b or a;
    outputs(3512) <= a xor b;
    outputs(3513) <= not a;
    outputs(3514) <= not a or b;
    outputs(3515) <= a;
    outputs(3516) <= a xor b;
    outputs(3517) <= not b or a;
    outputs(3518) <= not (a xor b);
    outputs(3519) <= not a;
    outputs(3520) <= not b;
    outputs(3521) <= not a;
    outputs(3522) <= not b or a;
    outputs(3523) <= not a;
    outputs(3524) <= not (a xor b);
    outputs(3525) <= a;
    outputs(3526) <= a xor b;
    outputs(3527) <= not a;
    outputs(3528) <= not b;
    outputs(3529) <= not b;
    outputs(3530) <= a;
    outputs(3531) <= not (a xor b);
    outputs(3532) <= not a;
    outputs(3533) <= a;
    outputs(3534) <= a xor b;
    outputs(3535) <= not a or b;
    outputs(3536) <= b and not a;
    outputs(3537) <= a;
    outputs(3538) <= not b;
    outputs(3539) <= not (a xor b);
    outputs(3540) <= not a;
    outputs(3541) <= not (a xor b);
    outputs(3542) <= not b;
    outputs(3543) <= a xor b;
    outputs(3544) <= a and b;
    outputs(3545) <= b and not a;
    outputs(3546) <= b;
    outputs(3547) <= not a;
    outputs(3548) <= not b or a;
    outputs(3549) <= not a;
    outputs(3550) <= not (a xor b);
    outputs(3551) <= not (a xor b);
    outputs(3552) <= a xor b;
    outputs(3553) <= a;
    outputs(3554) <= a;
    outputs(3555) <= a and not b;
    outputs(3556) <= not b;
    outputs(3557) <= a;
    outputs(3558) <= not a;
    outputs(3559) <= not a;
    outputs(3560) <= not b;
    outputs(3561) <= a;
    outputs(3562) <= not b;
    outputs(3563) <= not b;
    outputs(3564) <= a;
    outputs(3565) <= not b;
    outputs(3566) <= not a or b;
    outputs(3567) <= not b;
    outputs(3568) <= b and not a;
    outputs(3569) <= b;
    outputs(3570) <= not a;
    outputs(3571) <= b;
    outputs(3572) <= not (a and b);
    outputs(3573) <= a;
    outputs(3574) <= not (a xor b);
    outputs(3575) <= not a or b;
    outputs(3576) <= a xor b;
    outputs(3577) <= a;
    outputs(3578) <= not b;
    outputs(3579) <= not (a or b);
    outputs(3580) <= a;
    outputs(3581) <= a or b;
    outputs(3582) <= a xor b;
    outputs(3583) <= not (a xor b);
    outputs(3584) <= not (a or b);
    outputs(3585) <= not b;
    outputs(3586) <= a xor b;
    outputs(3587) <= b;
    outputs(3588) <= not (a xor b);
    outputs(3589) <= not a;
    outputs(3590) <= a;
    outputs(3591) <= a xor b;
    outputs(3592) <= a and b;
    outputs(3593) <= a xor b;
    outputs(3594) <= b and not a;
    outputs(3595) <= not a or b;
    outputs(3596) <= b and not a;
    outputs(3597) <= not b;
    outputs(3598) <= b;
    outputs(3599) <= a and not b;
    outputs(3600) <= not a;
    outputs(3601) <= not a or b;
    outputs(3602) <= not a;
    outputs(3603) <= not a;
    outputs(3604) <= not a;
    outputs(3605) <= b;
    outputs(3606) <= not b;
    outputs(3607) <= not a;
    outputs(3608) <= not (a xor b);
    outputs(3609) <= not a;
    outputs(3610) <= not b;
    outputs(3611) <= not a;
    outputs(3612) <= a xor b;
    outputs(3613) <= not b;
    outputs(3614) <= not b;
    outputs(3615) <= b;
    outputs(3616) <= a xor b;
    outputs(3617) <= not (a or b);
    outputs(3618) <= a;
    outputs(3619) <= b and not a;
    outputs(3620) <= a;
    outputs(3621) <= not a;
    outputs(3622) <= not a;
    outputs(3623) <= not b;
    outputs(3624) <= a;
    outputs(3625) <= not (a xor b);
    outputs(3626) <= not b;
    outputs(3627) <= a xor b;
    outputs(3628) <= not (a xor b);
    outputs(3629) <= not b;
    outputs(3630) <= not (a and b);
    outputs(3631) <= not b or a;
    outputs(3632) <= b and not a;
    outputs(3633) <= not a or b;
    outputs(3634) <= not a;
    outputs(3635) <= not b;
    outputs(3636) <= not (a xor b);
    outputs(3637) <= b;
    outputs(3638) <= b;
    outputs(3639) <= a or b;
    outputs(3640) <= b;
    outputs(3641) <= a xor b;
    outputs(3642) <= not a;
    outputs(3643) <= a;
    outputs(3644) <= a xor b;
    outputs(3645) <= not b or a;
    outputs(3646) <= not (a xor b);
    outputs(3647) <= not b or a;
    outputs(3648) <= not b;
    outputs(3649) <= b;
    outputs(3650) <= b;
    outputs(3651) <= not b;
    outputs(3652) <= not (a or b);
    outputs(3653) <= not b;
    outputs(3654) <= not (a and b);
    outputs(3655) <= a;
    outputs(3656) <= not a;
    outputs(3657) <= a;
    outputs(3658) <= not a;
    outputs(3659) <= a;
    outputs(3660) <= b;
    outputs(3661) <= a or b;
    outputs(3662) <= not b;
    outputs(3663) <= a xor b;
    outputs(3664) <= a and not b;
    outputs(3665) <= not b;
    outputs(3666) <= a xor b;
    outputs(3667) <= b;
    outputs(3668) <= not (a xor b);
    outputs(3669) <= a or b;
    outputs(3670) <= not b;
    outputs(3671) <= not b;
    outputs(3672) <= b;
    outputs(3673) <= a and not b;
    outputs(3674) <= a or b;
    outputs(3675) <= a xor b;
    outputs(3676) <= a and not b;
    outputs(3677) <= b;
    outputs(3678) <= not b;
    outputs(3679) <= not a;
    outputs(3680) <= a xor b;
    outputs(3681) <= not b;
    outputs(3682) <= a xor b;
    outputs(3683) <= b;
    outputs(3684) <= b and not a;
    outputs(3685) <= not b or a;
    outputs(3686) <= not a;
    outputs(3687) <= not b;
    outputs(3688) <= not b;
    outputs(3689) <= b;
    outputs(3690) <= a;
    outputs(3691) <= not (a xor b);
    outputs(3692) <= a and b;
    outputs(3693) <= a and b;
    outputs(3694) <= not (a or b);
    outputs(3695) <= b;
    outputs(3696) <= not a;
    outputs(3697) <= not a;
    outputs(3698) <= not a;
    outputs(3699) <= not b;
    outputs(3700) <= b;
    outputs(3701) <= not b;
    outputs(3702) <= b;
    outputs(3703) <= a xor b;
    outputs(3704) <= a or b;
    outputs(3705) <= not (a xor b);
    outputs(3706) <= a and b;
    outputs(3707) <= b;
    outputs(3708) <= a and not b;
    outputs(3709) <= a xor b;
    outputs(3710) <= not a;
    outputs(3711) <= not a;
    outputs(3712) <= not a;
    outputs(3713) <= a and not b;
    outputs(3714) <= a xor b;
    outputs(3715) <= not a;
    outputs(3716) <= a xor b;
    outputs(3717) <= not b;
    outputs(3718) <= a;
    outputs(3719) <= a and not b;
    outputs(3720) <= b and not a;
    outputs(3721) <= not a;
    outputs(3722) <= a xor b;
    outputs(3723) <= not (a xor b);
    outputs(3724) <= b;
    outputs(3725) <= a;
    outputs(3726) <= not (a xor b);
    outputs(3727) <= not (a and b);
    outputs(3728) <= a and not b;
    outputs(3729) <= not a;
    outputs(3730) <= not a;
    outputs(3731) <= not a;
    outputs(3732) <= b;
    outputs(3733) <= a and not b;
    outputs(3734) <= not a;
    outputs(3735) <= not a or b;
    outputs(3736) <= a and not b;
    outputs(3737) <= not a or b;
    outputs(3738) <= not a;
    outputs(3739) <= not (a xor b);
    outputs(3740) <= not (a xor b);
    outputs(3741) <= a xor b;
    outputs(3742) <= b;
    outputs(3743) <= a and b;
    outputs(3744) <= a;
    outputs(3745) <= not b;
    outputs(3746) <= not b;
    outputs(3747) <= a xor b;
    outputs(3748) <= b;
    outputs(3749) <= not a;
    outputs(3750) <= a xor b;
    outputs(3751) <= not a;
    outputs(3752) <= not (a xor b);
    outputs(3753) <= not b or a;
    outputs(3754) <= not a or b;
    outputs(3755) <= b and not a;
    outputs(3756) <= b;
    outputs(3757) <= a;
    outputs(3758) <= not (a xor b);
    outputs(3759) <= not b;
    outputs(3760) <= not a;
    outputs(3761) <= a;
    outputs(3762) <= not a;
    outputs(3763) <= a and not b;
    outputs(3764) <= b;
    outputs(3765) <= not b;
    outputs(3766) <= a xor b;
    outputs(3767) <= not b;
    outputs(3768) <= b and not a;
    outputs(3769) <= b;
    outputs(3770) <= a and not b;
    outputs(3771) <= not (a xor b);
    outputs(3772) <= not a;
    outputs(3773) <= not b or a;
    outputs(3774) <= b;
    outputs(3775) <= a xor b;
    outputs(3776) <= b and not a;
    outputs(3777) <= not b;
    outputs(3778) <= a xor b;
    outputs(3779) <= not (a or b);
    outputs(3780) <= not b;
    outputs(3781) <= not (a xor b);
    outputs(3782) <= not (a xor b);
    outputs(3783) <= not a;
    outputs(3784) <= b and not a;
    outputs(3785) <= not (a xor b);
    outputs(3786) <= a and not b;
    outputs(3787) <= a and b;
    outputs(3788) <= not b;
    outputs(3789) <= a xor b;
    outputs(3790) <= not (a and b);
    outputs(3791) <= not b or a;
    outputs(3792) <= not (a xor b);
    outputs(3793) <= not a;
    outputs(3794) <= a xor b;
    outputs(3795) <= not (a xor b);
    outputs(3796) <= not a;
    outputs(3797) <= not (a xor b);
    outputs(3798) <= not (a xor b);
    outputs(3799) <= not b;
    outputs(3800) <= not a;
    outputs(3801) <= not b;
    outputs(3802) <= not (a or b);
    outputs(3803) <= a xor b;
    outputs(3804) <= not (a xor b);
    outputs(3805) <= a xor b;
    outputs(3806) <= a;
    outputs(3807) <= b;
    outputs(3808) <= a xor b;
    outputs(3809) <= not (a or b);
    outputs(3810) <= not b;
    outputs(3811) <= not b or a;
    outputs(3812) <= a xor b;
    outputs(3813) <= not b or a;
    outputs(3814) <= a;
    outputs(3815) <= b;
    outputs(3816) <= not (a xor b);
    outputs(3817) <= a and b;
    outputs(3818) <= b;
    outputs(3819) <= not a;
    outputs(3820) <= not (a xor b);
    outputs(3821) <= not b;
    outputs(3822) <= a xor b;
    outputs(3823) <= a xor b;
    outputs(3824) <= a xor b;
    outputs(3825) <= not (a xor b);
    outputs(3826) <= not b;
    outputs(3827) <= a and b;
    outputs(3828) <= not a;
    outputs(3829) <= not b;
    outputs(3830) <= not a;
    outputs(3831) <= not b;
    outputs(3832) <= a;
    outputs(3833) <= not (a xor b);
    outputs(3834) <= a;
    outputs(3835) <= a and b;
    outputs(3836) <= b;
    outputs(3837) <= not (a and b);
    outputs(3838) <= not (a xor b);
    outputs(3839) <= not a;
    outputs(3840) <= a and b;
    outputs(3841) <= a;
    outputs(3842) <= not (a or b);
    outputs(3843) <= not b;
    outputs(3844) <= b;
    outputs(3845) <= b and not a;
    outputs(3846) <= b and not a;
    outputs(3847) <= not a;
    outputs(3848) <= not (a or b);
    outputs(3849) <= a;
    outputs(3850) <= a xor b;
    outputs(3851) <= a and b;
    outputs(3852) <= not (a and b);
    outputs(3853) <= b;
    outputs(3854) <= a;
    outputs(3855) <= not a;
    outputs(3856) <= not (a or b);
    outputs(3857) <= not (a and b);
    outputs(3858) <= b;
    outputs(3859) <= not a;
    outputs(3860) <= not (a and b);
    outputs(3861) <= not a;
    outputs(3862) <= not a;
    outputs(3863) <= a xor b;
    outputs(3864) <= not b;
    outputs(3865) <= not (a xor b);
    outputs(3866) <= b and not a;
    outputs(3867) <= a and not b;
    outputs(3868) <= a;
    outputs(3869) <= not (a and b);
    outputs(3870) <= not (a xor b);
    outputs(3871) <= a;
    outputs(3872) <= a;
    outputs(3873) <= not (a xor b);
    outputs(3874) <= not (a xor b);
    outputs(3875) <= not (a and b);
    outputs(3876) <= not b;
    outputs(3877) <= b;
    outputs(3878) <= not a;
    outputs(3879) <= not (a or b);
    outputs(3880) <= not (a xor b);
    outputs(3881) <= a xor b;
    outputs(3882) <= b and not a;
    outputs(3883) <= a;
    outputs(3884) <= a xor b;
    outputs(3885) <= not b;
    outputs(3886) <= not b;
    outputs(3887) <= a xor b;
    outputs(3888) <= not (a or b);
    outputs(3889) <= b and not a;
    outputs(3890) <= a xor b;
    outputs(3891) <= a;
    outputs(3892) <= not b;
    outputs(3893) <= not (a or b);
    outputs(3894) <= a and not b;
    outputs(3895) <= b;
    outputs(3896) <= a or b;
    outputs(3897) <= a;
    outputs(3898) <= not b;
    outputs(3899) <= b;
    outputs(3900) <= not (a xor b);
    outputs(3901) <= not a;
    outputs(3902) <= b;
    outputs(3903) <= not a;
    outputs(3904) <= b;
    outputs(3905) <= not (a or b);
    outputs(3906) <= not b or a;
    outputs(3907) <= not (a xor b);
    outputs(3908) <= a or b;
    outputs(3909) <= not b;
    outputs(3910) <= b and not a;
    outputs(3911) <= b;
    outputs(3912) <= a;
    outputs(3913) <= b and not a;
    outputs(3914) <= not (a xor b);
    outputs(3915) <= not (a xor b);
    outputs(3916) <= not (a or b);
    outputs(3917) <= a xor b;
    outputs(3918) <= not (a xor b);
    outputs(3919) <= not (a xor b);
    outputs(3920) <= a or b;
    outputs(3921) <= not (a or b);
    outputs(3922) <= not (a xor b);
    outputs(3923) <= not (a xor b);
    outputs(3924) <= a xor b;
    outputs(3925) <= not (a xor b);
    outputs(3926) <= a and not b;
    outputs(3927) <= not b or a;
    outputs(3928) <= a xor b;
    outputs(3929) <= not (a xor b);
    outputs(3930) <= a;
    outputs(3931) <= not b;
    outputs(3932) <= b;
    outputs(3933) <= a and not b;
    outputs(3934) <= not a;
    outputs(3935) <= not b or a;
    outputs(3936) <= a;
    outputs(3937) <= a and not b;
    outputs(3938) <= not b;
    outputs(3939) <= b;
    outputs(3940) <= not (a or b);
    outputs(3941) <= b;
    outputs(3942) <= not (a xor b);
    outputs(3943) <= b;
    outputs(3944) <= not b;
    outputs(3945) <= a and b;
    outputs(3946) <= not a;
    outputs(3947) <= a;
    outputs(3948) <= b;
    outputs(3949) <= not a;
    outputs(3950) <= not b;
    outputs(3951) <= not (a or b);
    outputs(3952) <= not a;
    outputs(3953) <= not a;
    outputs(3954) <= b;
    outputs(3955) <= not (a xor b);
    outputs(3956) <= b and not a;
    outputs(3957) <= b;
    outputs(3958) <= a xor b;
    outputs(3959) <= a xor b;
    outputs(3960) <= not (a xor b);
    outputs(3961) <= not b;
    outputs(3962) <= a;
    outputs(3963) <= a and b;
    outputs(3964) <= a;
    outputs(3965) <= not (a and b);
    outputs(3966) <= not (a xor b);
    outputs(3967) <= not (a xor b);
    outputs(3968) <= not a;
    outputs(3969) <= a xor b;
    outputs(3970) <= a xor b;
    outputs(3971) <= a xor b;
    outputs(3972) <= a xor b;
    outputs(3973) <= a;
    outputs(3974) <= a and not b;
    outputs(3975) <= a or b;
    outputs(3976) <= a and b;
    outputs(3977) <= not (a xor b);
    outputs(3978) <= not a;
    outputs(3979) <= not (a xor b);
    outputs(3980) <= not (a or b);
    outputs(3981) <= not b;
    outputs(3982) <= not a;
    outputs(3983) <= a and b;
    outputs(3984) <= not a or b;
    outputs(3985) <= not (a xor b);
    outputs(3986) <= a;
    outputs(3987) <= not b or a;
    outputs(3988) <= a xor b;
    outputs(3989) <= not (a and b);
    outputs(3990) <= not b;
    outputs(3991) <= not a;
    outputs(3992) <= b;
    outputs(3993) <= not (a xor b);
    outputs(3994) <= not b;
    outputs(3995) <= not (a or b);
    outputs(3996) <= not b;
    outputs(3997) <= b and not a;
    outputs(3998) <= b;
    outputs(3999) <= a xor b;
    outputs(4000) <= a and not b;
    outputs(4001) <= a xor b;
    outputs(4002) <= a;
    outputs(4003) <= b;
    outputs(4004) <= a xor b;
    outputs(4005) <= a and not b;
    outputs(4006) <= not (a xor b);
    outputs(4007) <= not (a or b);
    outputs(4008) <= b;
    outputs(4009) <= a xor b;
    outputs(4010) <= not b or a;
    outputs(4011) <= not (a xor b);
    outputs(4012) <= not a;
    outputs(4013) <= a;
    outputs(4014) <= not (a or b);
    outputs(4015) <= not (a xor b);
    outputs(4016) <= not a or b;
    outputs(4017) <= not (a or b);
    outputs(4018) <= not (a or b);
    outputs(4019) <= not (a xor b);
    outputs(4020) <= a xor b;
    outputs(4021) <= a xor b;
    outputs(4022) <= not a;
    outputs(4023) <= a xor b;
    outputs(4024) <= not (a or b);
    outputs(4025) <= a or b;
    outputs(4026) <= a xor b;
    outputs(4027) <= not b;
    outputs(4028) <= not b;
    outputs(4029) <= a or b;
    outputs(4030) <= not b;
    outputs(4031) <= a;
    outputs(4032) <= a and not b;
    outputs(4033) <= not (a and b);
    outputs(4034) <= a or b;
    outputs(4035) <= b and not a;
    outputs(4036) <= a;
    outputs(4037) <= not b;
    outputs(4038) <= b;
    outputs(4039) <= a;
    outputs(4040) <= b;
    outputs(4041) <= not (a xor b);
    outputs(4042) <= not a;
    outputs(4043) <= not b;
    outputs(4044) <= not (a or b);
    outputs(4045) <= b and not a;
    outputs(4046) <= a xor b;
    outputs(4047) <= a and b;
    outputs(4048) <= b;
    outputs(4049) <= not (a xor b);
    outputs(4050) <= not a;
    outputs(4051) <= not (a or b);
    outputs(4052) <= a and b;
    outputs(4053) <= not a;
    outputs(4054) <= a;
    outputs(4055) <= not (a xor b);
    outputs(4056) <= not a;
    outputs(4057) <= b;
    outputs(4058) <= not a;
    outputs(4059) <= a xor b;
    outputs(4060) <= not (a xor b);
    outputs(4061) <= not a or b;
    outputs(4062) <= b;
    outputs(4063) <= not a;
    outputs(4064) <= not (a xor b);
    outputs(4065) <= b;
    outputs(4066) <= a xor b;
    outputs(4067) <= a;
    outputs(4068) <= not a;
    outputs(4069) <= b;
    outputs(4070) <= a xor b;
    outputs(4071) <= a;
    outputs(4072) <= b;
    outputs(4073) <= not a;
    outputs(4074) <= a and not b;
    outputs(4075) <= a;
    outputs(4076) <= not (a xor b);
    outputs(4077) <= not b;
    outputs(4078) <= a and b;
    outputs(4079) <= a or b;
    outputs(4080) <= not b;
    outputs(4081) <= b;
    outputs(4082) <= a xor b;
    outputs(4083) <= not b;
    outputs(4084) <= not b or a;
    outputs(4085) <= b;
    outputs(4086) <= not b;
    outputs(4087) <= b;
    outputs(4088) <= a;
    outputs(4089) <= a xor b;
    outputs(4090) <= not a or b;
    outputs(4091) <= not a;
    outputs(4092) <= not b;
    outputs(4093) <= b and not a;
    outputs(4094) <= not a;
    outputs(4095) <= a and b;
    outputs(4096) <= a and b;
    outputs(4097) <= not (a and b);
    outputs(4098) <= a and b;
    outputs(4099) <= a xor b;
    outputs(4100) <= a and not b;
    outputs(4101) <= not (a or b);
    outputs(4102) <= a xor b;
    outputs(4103) <= b;
    outputs(4104) <= not b or a;
    outputs(4105) <= not b;
    outputs(4106) <= not (a xor b);
    outputs(4107) <= not (a xor b);
    outputs(4108) <= a;
    outputs(4109) <= a and b;
    outputs(4110) <= not a;
    outputs(4111) <= not b;
    outputs(4112) <= not (a xor b);
    outputs(4113) <= a;
    outputs(4114) <= not b;
    outputs(4115) <= not a;
    outputs(4116) <= a and not b;
    outputs(4117) <= a xor b;
    outputs(4118) <= not a;
    outputs(4119) <= not a;
    outputs(4120) <= not a;
    outputs(4121) <= a and not b;
    outputs(4122) <= not a or b;
    outputs(4123) <= a xor b;
    outputs(4124) <= a xor b;
    outputs(4125) <= not (a xor b);
    outputs(4126) <= not (a xor b);
    outputs(4127) <= a and b;
    outputs(4128) <= not (a xor b);
    outputs(4129) <= not a;
    outputs(4130) <= not b;
    outputs(4131) <= a and not b;
    outputs(4132) <= a;
    outputs(4133) <= a;
    outputs(4134) <= not (a xor b);
    outputs(4135) <= not (a xor b);
    outputs(4136) <= not b;
    outputs(4137) <= not (a or b);
    outputs(4138) <= a or b;
    outputs(4139) <= not (a xor b);
    outputs(4140) <= not (a xor b);
    outputs(4141) <= b;
    outputs(4142) <= a;
    outputs(4143) <= a;
    outputs(4144) <= not (a xor b);
    outputs(4145) <= not b;
    outputs(4146) <= b;
    outputs(4147) <= not a;
    outputs(4148) <= a;
    outputs(4149) <= not a;
    outputs(4150) <= a;
    outputs(4151) <= not (a or b);
    outputs(4152) <= not (a or b);
    outputs(4153) <= a xor b;
    outputs(4154) <= a;
    outputs(4155) <= a;
    outputs(4156) <= not (a xor b);
    outputs(4157) <= not b;
    outputs(4158) <= not b or a;
    outputs(4159) <= a xor b;
    outputs(4160) <= not a;
    outputs(4161) <= not b;
    outputs(4162) <= a;
    outputs(4163) <= a and not b;
    outputs(4164) <= a and not b;
    outputs(4165) <= a;
    outputs(4166) <= not b;
    outputs(4167) <= a and not b;
    outputs(4168) <= not (a xor b);
    outputs(4169) <= a xor b;
    outputs(4170) <= a;
    outputs(4171) <= b;
    outputs(4172) <= a and not b;
    outputs(4173) <= b;
    outputs(4174) <= a xor b;
    outputs(4175) <= not a;
    outputs(4176) <= a;
    outputs(4177) <= b;
    outputs(4178) <= not b;
    outputs(4179) <= b and not a;
    outputs(4180) <= not b;
    outputs(4181) <= a;
    outputs(4182) <= a xor b;
    outputs(4183) <= b;
    outputs(4184) <= b;
    outputs(4185) <= not (a xor b);
    outputs(4186) <= a xor b;
    outputs(4187) <= not a;
    outputs(4188) <= not a;
    outputs(4189) <= b;
    outputs(4190) <= not b;
    outputs(4191) <= a;
    outputs(4192) <= not b;
    outputs(4193) <= b;
    outputs(4194) <= b;
    outputs(4195) <= not (a xor b);
    outputs(4196) <= a xor b;
    outputs(4197) <= a and not b;
    outputs(4198) <= a xor b;
    outputs(4199) <= not a;
    outputs(4200) <= a xor b;
    outputs(4201) <= not (a xor b);
    outputs(4202) <= a xor b;
    outputs(4203) <= a and b;
    outputs(4204) <= not (a xor b);
    outputs(4205) <= not a;
    outputs(4206) <= not b;
    outputs(4207) <= b;
    outputs(4208) <= not a;
    outputs(4209) <= b;
    outputs(4210) <= not a;
    outputs(4211) <= not (a xor b);
    outputs(4212) <= a xor b;
    outputs(4213) <= a or b;
    outputs(4214) <= not b;
    outputs(4215) <= a xor b;
    outputs(4216) <= a and b;
    outputs(4217) <= a;
    outputs(4218) <= a;
    outputs(4219) <= not (a xor b);
    outputs(4220) <= b and not a;
    outputs(4221) <= not a;
    outputs(4222) <= not b;
    outputs(4223) <= not (a xor b);
    outputs(4224) <= not a;
    outputs(4225) <= not a;
    outputs(4226) <= not b;
    outputs(4227) <= a xor b;
    outputs(4228) <= a and b;
    outputs(4229) <= a;
    outputs(4230) <= not a;
    outputs(4231) <= a and b;
    outputs(4232) <= not (a xor b);
    outputs(4233) <= b;
    outputs(4234) <= not (a xor b);
    outputs(4235) <= a xor b;
    outputs(4236) <= a;
    outputs(4237) <= not b;
    outputs(4238) <= not a;
    outputs(4239) <= a;
    outputs(4240) <= not a;
    outputs(4241) <= not a;
    outputs(4242) <= not a;
    outputs(4243) <= a;
    outputs(4244) <= a xor b;
    outputs(4245) <= b and not a;
    outputs(4246) <= b and not a;
    outputs(4247) <= not b;
    outputs(4248) <= b;
    outputs(4249) <= a;
    outputs(4250) <= a xor b;
    outputs(4251) <= not a;
    outputs(4252) <= not a;
    outputs(4253) <= not a;
    outputs(4254) <= a or b;
    outputs(4255) <= a xor b;
    outputs(4256) <= not a;
    outputs(4257) <= not (a xor b);
    outputs(4258) <= not a;
    outputs(4259) <= a xor b;
    outputs(4260) <= not (a xor b);
    outputs(4261) <= b and not a;
    outputs(4262) <= a and not b;
    outputs(4263) <= a;
    outputs(4264) <= not b;
    outputs(4265) <= a xor b;
    outputs(4266) <= not a;
    outputs(4267) <= not b;
    outputs(4268) <= a xor b;
    outputs(4269) <= not b;
    outputs(4270) <= not (a and b);
    outputs(4271) <= not b or a;
    outputs(4272) <= b;
    outputs(4273) <= not b;
    outputs(4274) <= a xor b;
    outputs(4275) <= a xor b;
    outputs(4276) <= a and not b;
    outputs(4277) <= b;
    outputs(4278) <= b;
    outputs(4279) <= b;
    outputs(4280) <= not (a xor b);
    outputs(4281) <= a;
    outputs(4282) <= not (a or b);
    outputs(4283) <= a xor b;
    outputs(4284) <= a xor b;
    outputs(4285) <= a xor b;
    outputs(4286) <= b;
    outputs(4287) <= not b;
    outputs(4288) <= not b;
    outputs(4289) <= a;
    outputs(4290) <= not b;
    outputs(4291) <= not a;
    outputs(4292) <= b;
    outputs(4293) <= not b;
    outputs(4294) <= a or b;
    outputs(4295) <= a;
    outputs(4296) <= b;
    outputs(4297) <= a and not b;
    outputs(4298) <= not a;
    outputs(4299) <= b;
    outputs(4300) <= not a;
    outputs(4301) <= a;
    outputs(4302) <= not b;
    outputs(4303) <= not (a xor b);
    outputs(4304) <= a;
    outputs(4305) <= not b;
    outputs(4306) <= b;
    outputs(4307) <= not (a or b);
    outputs(4308) <= a xor b;
    outputs(4309) <= not b;
    outputs(4310) <= a;
    outputs(4311) <= not (a xor b);
    outputs(4312) <= not b;
    outputs(4313) <= not b;
    outputs(4314) <= a and not b;
    outputs(4315) <= not b;
    outputs(4316) <= a;
    outputs(4317) <= not b or a;
    outputs(4318) <= not (a xor b);
    outputs(4319) <= a xor b;
    outputs(4320) <= not (a xor b);
    outputs(4321) <= b;
    outputs(4322) <= not (a xor b);
    outputs(4323) <= not (a or b);
    outputs(4324) <= a xor b;
    outputs(4325) <= not (a or b);
    outputs(4326) <= a;
    outputs(4327) <= a or b;
    outputs(4328) <= a or b;
    outputs(4329) <= a xor b;
    outputs(4330) <= a xor b;
    outputs(4331) <= not (a xor b);
    outputs(4332) <= not b;
    outputs(4333) <= a;
    outputs(4334) <= a xor b;
    outputs(4335) <= not (a xor b);
    outputs(4336) <= not (a xor b);
    outputs(4337) <= b and not a;
    outputs(4338) <= a and not b;
    outputs(4339) <= not (a and b);
    outputs(4340) <= not b;
    outputs(4341) <= not a;
    outputs(4342) <= a or b;
    outputs(4343) <= not b;
    outputs(4344) <= not b;
    outputs(4345) <= not b;
    outputs(4346) <= not b;
    outputs(4347) <= a xor b;
    outputs(4348) <= not b;
    outputs(4349) <= b and not a;
    outputs(4350) <= a and not b;
    outputs(4351) <= a;
    outputs(4352) <= a xor b;
    outputs(4353) <= b;
    outputs(4354) <= not (a xor b);
    outputs(4355) <= not (a xor b);
    outputs(4356) <= a xor b;
    outputs(4357) <= a;
    outputs(4358) <= b;
    outputs(4359) <= a xor b;
    outputs(4360) <= not (a xor b);
    outputs(4361) <= not (a or b);
    outputs(4362) <= b and not a;
    outputs(4363) <= not b;
    outputs(4364) <= a;
    outputs(4365) <= a xor b;
    outputs(4366) <= not (a xor b);
    outputs(4367) <= not b;
    outputs(4368) <= not b;
    outputs(4369) <= a xor b;
    outputs(4370) <= not a;
    outputs(4371) <= not a;
    outputs(4372) <= not (a xor b);
    outputs(4373) <= not b;
    outputs(4374) <= not a;
    outputs(4375) <= a or b;
    outputs(4376) <= not b;
    outputs(4377) <= not b;
    outputs(4378) <= not (a xor b);
    outputs(4379) <= b and not a;
    outputs(4380) <= a;
    outputs(4381) <= a xor b;
    outputs(4382) <= a xor b;
    outputs(4383) <= not a;
    outputs(4384) <= not (a xor b);
    outputs(4385) <= not b;
    outputs(4386) <= not b;
    outputs(4387) <= not a or b;
    outputs(4388) <= not (a and b);
    outputs(4389) <= b;
    outputs(4390) <= a;
    outputs(4391) <= not (a xor b);
    outputs(4392) <= not b;
    outputs(4393) <= not a or b;
    outputs(4394) <= a xor b;
    outputs(4395) <= a;
    outputs(4396) <= a xor b;
    outputs(4397) <= not (a xor b);
    outputs(4398) <= not b;
    outputs(4399) <= b;
    outputs(4400) <= b;
    outputs(4401) <= a and not b;
    outputs(4402) <= not b or a;
    outputs(4403) <= a and b;
    outputs(4404) <= not (a xor b);
    outputs(4405) <= not (a or b);
    outputs(4406) <= not (a or b);
    outputs(4407) <= b;
    outputs(4408) <= not a;
    outputs(4409) <= not a;
    outputs(4410) <= a xor b;
    outputs(4411) <= not b;
    outputs(4412) <= a xor b;
    outputs(4413) <= a xor b;
    outputs(4414) <= not b;
    outputs(4415) <= a and b;
    outputs(4416) <= a;
    outputs(4417) <= not b;
    outputs(4418) <= b;
    outputs(4419) <= a xor b;
    outputs(4420) <= not b;
    outputs(4421) <= not a or b;
    outputs(4422) <= not b;
    outputs(4423) <= a;
    outputs(4424) <= not (a xor b);
    outputs(4425) <= not (a or b);
    outputs(4426) <= a;
    outputs(4427) <= not a;
    outputs(4428) <= not b;
    outputs(4429) <= a;
    outputs(4430) <= b;
    outputs(4431) <= not (a xor b);
    outputs(4432) <= b;
    outputs(4433) <= a and not b;
    outputs(4434) <= not b;
    outputs(4435) <= a and b;
    outputs(4436) <= b;
    outputs(4437) <= not a;
    outputs(4438) <= a xor b;
    outputs(4439) <= a xor b;
    outputs(4440) <= b;
    outputs(4441) <= not (a xor b);
    outputs(4442) <= not a;
    outputs(4443) <= b;
    outputs(4444) <= b and not a;
    outputs(4445) <= not (a xor b);
    outputs(4446) <= a and not b;
    outputs(4447) <= a xor b;
    outputs(4448) <= not a;
    outputs(4449) <= b;
    outputs(4450) <= b and not a;
    outputs(4451) <= not b;
    outputs(4452) <= not b;
    outputs(4453) <= not a;
    outputs(4454) <= a xor b;
    outputs(4455) <= not a;
    outputs(4456) <= not b;
    outputs(4457) <= a xor b;
    outputs(4458) <= not (a xor b);
    outputs(4459) <= not a;
    outputs(4460) <= b;
    outputs(4461) <= a and b;
    outputs(4462) <= b and not a;
    outputs(4463) <= not b;
    outputs(4464) <= a xor b;
    outputs(4465) <= a xor b;
    outputs(4466) <= a and not b;
    outputs(4467) <= not b;
    outputs(4468) <= not b;
    outputs(4469) <= a xor b;
    outputs(4470) <= a xor b;
    outputs(4471) <= not (a xor b);
    outputs(4472) <= a;
    outputs(4473) <= not (a or b);
    outputs(4474) <= not b or a;
    outputs(4475) <= b;
    outputs(4476) <= not b;
    outputs(4477) <= a;
    outputs(4478) <= b;
    outputs(4479) <= not a or b;
    outputs(4480) <= not b;
    outputs(4481) <= not a;
    outputs(4482) <= not (a xor b);
    outputs(4483) <= b and not a;
    outputs(4484) <= b;
    outputs(4485) <= not (a xor b);
    outputs(4486) <= b;
    outputs(4487) <= not b;
    outputs(4488) <= b and not a;
    outputs(4489) <= not (a xor b);
    outputs(4490) <= not (a xor b);
    outputs(4491) <= not (a xor b);
    outputs(4492) <= a;
    outputs(4493) <= not (a xor b);
    outputs(4494) <= a xor b;
    outputs(4495) <= a and b;
    outputs(4496) <= not b;
    outputs(4497) <= b;
    outputs(4498) <= not b or a;
    outputs(4499) <= not (a xor b);
    outputs(4500) <= a and not b;
    outputs(4501) <= not a;
    outputs(4502) <= not (a and b);
    outputs(4503) <= not b or a;
    outputs(4504) <= b and not a;
    outputs(4505) <= not b;
    outputs(4506) <= a and b;
    outputs(4507) <= a;
    outputs(4508) <= b and not a;
    outputs(4509) <= not a;
    outputs(4510) <= b;
    outputs(4511) <= not (a xor b);
    outputs(4512) <= not b;
    outputs(4513) <= a and not b;
    outputs(4514) <= not a;
    outputs(4515) <= not (a xor b);
    outputs(4516) <= not (a or b);
    outputs(4517) <= a;
    outputs(4518) <= not a;
    outputs(4519) <= not (a xor b);
    outputs(4520) <= b and not a;
    outputs(4521) <= b;
    outputs(4522) <= a;
    outputs(4523) <= b and not a;
    outputs(4524) <= not b;
    outputs(4525) <= a xor b;
    outputs(4526) <= b;
    outputs(4527) <= not b;
    outputs(4528) <= a or b;
    outputs(4529) <= a xor b;
    outputs(4530) <= not (a and b);
    outputs(4531) <= not (a xor b);
    outputs(4532) <= a xor b;
    outputs(4533) <= b;
    outputs(4534) <= b;
    outputs(4535) <= a xor b;
    outputs(4536) <= a xor b;
    outputs(4537) <= a;
    outputs(4538) <= not b;
    outputs(4539) <= b;
    outputs(4540) <= not a;
    outputs(4541) <= b and not a;
    outputs(4542) <= a;
    outputs(4543) <= not (a xor b);
    outputs(4544) <= a xor b;
    outputs(4545) <= a;
    outputs(4546) <= not b;
    outputs(4547) <= not (a xor b);
    outputs(4548) <= a and not b;
    outputs(4549) <= a;
    outputs(4550) <= b;
    outputs(4551) <= b;
    outputs(4552) <= b and not a;
    outputs(4553) <= not (a xor b);
    outputs(4554) <= not (a xor b);
    outputs(4555) <= not (a xor b);
    outputs(4556) <= not a;
    outputs(4557) <= b;
    outputs(4558) <= a;
    outputs(4559) <= b and not a;
    outputs(4560) <= not a;
    outputs(4561) <= not (a xor b);
    outputs(4562) <= a;
    outputs(4563) <= a;
    outputs(4564) <= a;
    outputs(4565) <= a and b;
    outputs(4566) <= not b;
    outputs(4567) <= not b;
    outputs(4568) <= b;
    outputs(4569) <= not a or b;
    outputs(4570) <= not a;
    outputs(4571) <= not a;
    outputs(4572) <= b and not a;
    outputs(4573) <= not b;
    outputs(4574) <= a or b;
    outputs(4575) <= b and not a;
    outputs(4576) <= not a;
    outputs(4577) <= b;
    outputs(4578) <= not a;
    outputs(4579) <= b and not a;
    outputs(4580) <= not b;
    outputs(4581) <= a;
    outputs(4582) <= not (a xor b);
    outputs(4583) <= a;
    outputs(4584) <= not (a xor b);
    outputs(4585) <= a and b;
    outputs(4586) <= not (a xor b);
    outputs(4587) <= not a or b;
    outputs(4588) <= a;
    outputs(4589) <= a;
    outputs(4590) <= not b;
    outputs(4591) <= b and not a;
    outputs(4592) <= not b;
    outputs(4593) <= a;
    outputs(4594) <= a;
    outputs(4595) <= a xor b;
    outputs(4596) <= not b;
    outputs(4597) <= not (a or b);
    outputs(4598) <= a;
    outputs(4599) <= not (a xor b);
    outputs(4600) <= a and b;
    outputs(4601) <= not a;
    outputs(4602) <= not (a xor b);
    outputs(4603) <= not b;
    outputs(4604) <= not (a xor b);
    outputs(4605) <= not a;
    outputs(4606) <= a;
    outputs(4607) <= a xor b;
    outputs(4608) <= not (a and b);
    outputs(4609) <= not b or a;
    outputs(4610) <= a;
    outputs(4611) <= not (a xor b);
    outputs(4612) <= a and b;
    outputs(4613) <= a xor b;
    outputs(4614) <= a xor b;
    outputs(4615) <= b and not a;
    outputs(4616) <= not b;
    outputs(4617) <= a or b;
    outputs(4618) <= not a;
    outputs(4619) <= b;
    outputs(4620) <= a;
    outputs(4621) <= a;
    outputs(4622) <= a xor b;
    outputs(4623) <= not (a xor b);
    outputs(4624) <= b;
    outputs(4625) <= not (a xor b);
    outputs(4626) <= b and not a;
    outputs(4627) <= b and not a;
    outputs(4628) <= not b;
    outputs(4629) <= a;
    outputs(4630) <= a xor b;
    outputs(4631) <= not b or a;
    outputs(4632) <= not (a and b);
    outputs(4633) <= a and b;
    outputs(4634) <= b and not a;
    outputs(4635) <= not b;
    outputs(4636) <= not a;
    outputs(4637) <= b;
    outputs(4638) <= not b;
    outputs(4639) <= not a;
    outputs(4640) <= not a;
    outputs(4641) <= a and b;
    outputs(4642) <= not b or a;
    outputs(4643) <= not a;
    outputs(4644) <= a;
    outputs(4645) <= not (a xor b);
    outputs(4646) <= not (a and b);
    outputs(4647) <= not b;
    outputs(4648) <= not b;
    outputs(4649) <= a;
    outputs(4650) <= a xor b;
    outputs(4651) <= not (a or b);
    outputs(4652) <= b;
    outputs(4653) <= a;
    outputs(4654) <= not (a xor b);
    outputs(4655) <= b and not a;
    outputs(4656) <= a and not b;
    outputs(4657) <= not (a and b);
    outputs(4658) <= not a;
    outputs(4659) <= not b;
    outputs(4660) <= b;
    outputs(4661) <= not (a and b);
    outputs(4662) <= a xor b;
    outputs(4663) <= a xor b;
    outputs(4664) <= not a;
    outputs(4665) <= not b or a;
    outputs(4666) <= a xor b;
    outputs(4667) <= a;
    outputs(4668) <= b;
    outputs(4669) <= not (a xor b);
    outputs(4670) <= a and b;
    outputs(4671) <= a xor b;
    outputs(4672) <= a or b;
    outputs(4673) <= a;
    outputs(4674) <= a;
    outputs(4675) <= a xor b;
    outputs(4676) <= a or b;
    outputs(4677) <= a;
    outputs(4678) <= a xor b;
    outputs(4679) <= not b;
    outputs(4680) <= not b or a;
    outputs(4681) <= b;
    outputs(4682) <= not a or b;
    outputs(4683) <= a;
    outputs(4684) <= not (a xor b);
    outputs(4685) <= a and b;
    outputs(4686) <= not (a xor b);
    outputs(4687) <= not b;
    outputs(4688) <= b;
    outputs(4689) <= not a;
    outputs(4690) <= not (a and b);
    outputs(4691) <= not (a or b);
    outputs(4692) <= not b;
    outputs(4693) <= b;
    outputs(4694) <= not a or b;
    outputs(4695) <= not (a xor b);
    outputs(4696) <= not (a xor b);
    outputs(4697) <= a;
    outputs(4698) <= not b or a;
    outputs(4699) <= a xor b;
    outputs(4700) <= not (a or b);
    outputs(4701) <= not a or b;
    outputs(4702) <= not b;
    outputs(4703) <= a and not b;
    outputs(4704) <= not b;
    outputs(4705) <= b;
    outputs(4706) <= a;
    outputs(4707) <= b and not a;
    outputs(4708) <= a or b;
    outputs(4709) <= not b;
    outputs(4710) <= a xor b;
    outputs(4711) <= not (a or b);
    outputs(4712) <= b;
    outputs(4713) <= a xor b;
    outputs(4714) <= not a or b;
    outputs(4715) <= not (a xor b);
    outputs(4716) <= b;
    outputs(4717) <= not b;
    outputs(4718) <= b;
    outputs(4719) <= a;
    outputs(4720) <= a;
    outputs(4721) <= not a;
    outputs(4722) <= b;
    outputs(4723) <= not a;
    outputs(4724) <= b;
    outputs(4725) <= a and b;
    outputs(4726) <= a;
    outputs(4727) <= not (a xor b);
    outputs(4728) <= not a;
    outputs(4729) <= a and not b;
    outputs(4730) <= a and b;
    outputs(4731) <= not (a xor b);
    outputs(4732) <= b;
    outputs(4733) <= not a or b;
    outputs(4734) <= not b;
    outputs(4735) <= a;
    outputs(4736) <= not (a xor b);
    outputs(4737) <= not a;
    outputs(4738) <= not a;
    outputs(4739) <= b and not a;
    outputs(4740) <= not (a xor b);
    outputs(4741) <= a and b;
    outputs(4742) <= not a;
    outputs(4743) <= not a;
    outputs(4744) <= b;
    outputs(4745) <= a and not b;
    outputs(4746) <= not b;
    outputs(4747) <= not a;
    outputs(4748) <= not b;
    outputs(4749) <= not b;
    outputs(4750) <= not a or b;
    outputs(4751) <= a;
    outputs(4752) <= not a;
    outputs(4753) <= not (a and b);
    outputs(4754) <= a and not b;
    outputs(4755) <= a and not b;
    outputs(4756) <= b;
    outputs(4757) <= a and not b;
    outputs(4758) <= not (a and b);
    outputs(4759) <= b;
    outputs(4760) <= not (a xor b);
    outputs(4761) <= not (a xor b);
    outputs(4762) <= b;
    outputs(4763) <= not a;
    outputs(4764) <= a;
    outputs(4765) <= not a;
    outputs(4766) <= a and b;
    outputs(4767) <= not (a or b);
    outputs(4768) <= b;
    outputs(4769) <= not a;
    outputs(4770) <= a and b;
    outputs(4771) <= a xor b;
    outputs(4772) <= a and b;
    outputs(4773) <= a and b;
    outputs(4774) <= a and not b;
    outputs(4775) <= a;
    outputs(4776) <= a;
    outputs(4777) <= a xor b;
    outputs(4778) <= not b;
    outputs(4779) <= b;
    outputs(4780) <= a;
    outputs(4781) <= a and b;
    outputs(4782) <= a and b;
    outputs(4783) <= b;
    outputs(4784) <= not (a or b);
    outputs(4785) <= not b;
    outputs(4786) <= not (a xor b);
    outputs(4787) <= not a;
    outputs(4788) <= a and b;
    outputs(4789) <= b and not a;
    outputs(4790) <= a;
    outputs(4791) <= a xor b;
    outputs(4792) <= a;
    outputs(4793) <= not a;
    outputs(4794) <= b;
    outputs(4795) <= not b;
    outputs(4796) <= a xor b;
    outputs(4797) <= b and not a;
    outputs(4798) <= a xor b;
    outputs(4799) <= not (a xor b);
    outputs(4800) <= not (a xor b);
    outputs(4801) <= a;
    outputs(4802) <= not (a xor b);
    outputs(4803) <= b;
    outputs(4804) <= a and not b;
    outputs(4805) <= not (a xor b);
    outputs(4806) <= a xor b;
    outputs(4807) <= not b;
    outputs(4808) <= a xor b;
    outputs(4809) <= a;
    outputs(4810) <= a xor b;
    outputs(4811) <= a;
    outputs(4812) <= b;
    outputs(4813) <= a or b;
    outputs(4814) <= a and not b;
    outputs(4815) <= a;
    outputs(4816) <= b;
    outputs(4817) <= b and not a;
    outputs(4818) <= a xor b;
    outputs(4819) <= b;
    outputs(4820) <= not a;
    outputs(4821) <= not b;
    outputs(4822) <= not (a xor b);
    outputs(4823) <= b;
    outputs(4824) <= a xor b;
    outputs(4825) <= not a;
    outputs(4826) <= a and b;
    outputs(4827) <= a xor b;
    outputs(4828) <= not (a xor b);
    outputs(4829) <= not a;
    outputs(4830) <= b;
    outputs(4831) <= not (a xor b);
    outputs(4832) <= not b;
    outputs(4833) <= a;
    outputs(4834) <= not a;
    outputs(4835) <= not b;
    outputs(4836) <= b;
    outputs(4837) <= not a;
    outputs(4838) <= b;
    outputs(4839) <= b;
    outputs(4840) <= a xor b;
    outputs(4841) <= a xor b;
    outputs(4842) <= not (a xor b);
    outputs(4843) <= not b;
    outputs(4844) <= b;
    outputs(4845) <= not (a xor b);
    outputs(4846) <= a and b;
    outputs(4847) <= b and not a;
    outputs(4848) <= not (a xor b);
    outputs(4849) <= a;
    outputs(4850) <= b;
    outputs(4851) <= b;
    outputs(4852) <= not (a xor b);
    outputs(4853) <= b;
    outputs(4854) <= not b;
    outputs(4855) <= not (a xor b);
    outputs(4856) <= not (a xor b);
    outputs(4857) <= not b or a;
    outputs(4858) <= not (a xor b);
    outputs(4859) <= a xor b;
    outputs(4860) <= not (a xor b);
    outputs(4861) <= a;
    outputs(4862) <= b and not a;
    outputs(4863) <= a and not b;
    outputs(4864) <= not a;
    outputs(4865) <= b and not a;
    outputs(4866) <= a xor b;
    outputs(4867) <= b and not a;
    outputs(4868) <= b;
    outputs(4869) <= not a;
    outputs(4870) <= a and not b;
    outputs(4871) <= not b;
    outputs(4872) <= not (a xor b);
    outputs(4873) <= b and not a;
    outputs(4874) <= not (a xor b);
    outputs(4875) <= not b;
    outputs(4876) <= a xor b;
    outputs(4877) <= not (a and b);
    outputs(4878) <= a;
    outputs(4879) <= not (a xor b);
    outputs(4880) <= not b;
    outputs(4881) <= b and not a;
    outputs(4882) <= b;
    outputs(4883) <= not (a xor b);
    outputs(4884) <= not b;
    outputs(4885) <= not b;
    outputs(4886) <= not (a xor b);
    outputs(4887) <= a;
    outputs(4888) <= b and not a;
    outputs(4889) <= not (a xor b);
    outputs(4890) <= a and b;
    outputs(4891) <= not a or b;
    outputs(4892) <= b and not a;
    outputs(4893) <= not a;
    outputs(4894) <= a xor b;
    outputs(4895) <= not (a xor b);
    outputs(4896) <= a;
    outputs(4897) <= a and not b;
    outputs(4898) <= not (a or b);
    outputs(4899) <= not a;
    outputs(4900) <= not (a or b);
    outputs(4901) <= b;
    outputs(4902) <= not a;
    outputs(4903) <= a or b;
    outputs(4904) <= not a;
    outputs(4905) <= not (a xor b);
    outputs(4906) <= not b;
    outputs(4907) <= b;
    outputs(4908) <= a and not b;
    outputs(4909) <= a;
    outputs(4910) <= a xor b;
    outputs(4911) <= not a;
    outputs(4912) <= a or b;
    outputs(4913) <= b and not a;
    outputs(4914) <= not (a xor b);
    outputs(4915) <= not (a and b);
    outputs(4916) <= a or b;
    outputs(4917) <= not (a or b);
    outputs(4918) <= a xor b;
    outputs(4919) <= not a or b;
    outputs(4920) <= not (a xor b);
    outputs(4921) <= not (a xor b);
    outputs(4922) <= not (a xor b);
    outputs(4923) <= not a;
    outputs(4924) <= not (a xor b);
    outputs(4925) <= not a;
    outputs(4926) <= not a;
    outputs(4927) <= not b;
    outputs(4928) <= a and not b;
    outputs(4929) <= a;
    outputs(4930) <= not a;
    outputs(4931) <= not (a xor b);
    outputs(4932) <= a and not b;
    outputs(4933) <= not b;
    outputs(4934) <= not a;
    outputs(4935) <= not b;
    outputs(4936) <= not b;
    outputs(4937) <= a xor b;
    outputs(4938) <= not a;
    outputs(4939) <= b;
    outputs(4940) <= not (a or b);
    outputs(4941) <= not a;
    outputs(4942) <= a;
    outputs(4943) <= not (a or b);
    outputs(4944) <= a and not b;
    outputs(4945) <= b;
    outputs(4946) <= b;
    outputs(4947) <= not (a xor b);
    outputs(4948) <= not a;
    outputs(4949) <= not a;
    outputs(4950) <= a and not b;
    outputs(4951) <= a;
    outputs(4952) <= a and b;
    outputs(4953) <= not a;
    outputs(4954) <= a xor b;
    outputs(4955) <= b and not a;
    outputs(4956) <= a and b;
    outputs(4957) <= a;
    outputs(4958) <= a xor b;
    outputs(4959) <= not b;
    outputs(4960) <= b and not a;
    outputs(4961) <= not (a xor b);
    outputs(4962) <= a and not b;
    outputs(4963) <= a xor b;
    outputs(4964) <= b and not a;
    outputs(4965) <= a;
    outputs(4966) <= not a;
    outputs(4967) <= a xor b;
    outputs(4968) <= not (a xor b);
    outputs(4969) <= not b;
    outputs(4970) <= a and not b;
    outputs(4971) <= not b;
    outputs(4972) <= b and not a;
    outputs(4973) <= not (a or b);
    outputs(4974) <= a xor b;
    outputs(4975) <= b and not a;
    outputs(4976) <= b and not a;
    outputs(4977) <= not a;
    outputs(4978) <= a;
    outputs(4979) <= b;
    outputs(4980) <= not a;
    outputs(4981) <= b;
    outputs(4982) <= not (a xor b);
    outputs(4983) <= not a;
    outputs(4984) <= a xor b;
    outputs(4985) <= b;
    outputs(4986) <= not (a xor b);
    outputs(4987) <= b and not a;
    outputs(4988) <= not (a xor b);
    outputs(4989) <= b;
    outputs(4990) <= not a;
    outputs(4991) <= a;
    outputs(4992) <= a xor b;
    outputs(4993) <= b;
    outputs(4994) <= a xor b;
    outputs(4995) <= b;
    outputs(4996) <= a xor b;
    outputs(4997) <= not a;
    outputs(4998) <= a xor b;
    outputs(4999) <= a;
    outputs(5000) <= a;
    outputs(5001) <= a xor b;
    outputs(5002) <= a and b;
    outputs(5003) <= not (a xor b);
    outputs(5004) <= not a;
    outputs(5005) <= not (a xor b);
    outputs(5006) <= a and not b;
    outputs(5007) <= not (a xor b);
    outputs(5008) <= a or b;
    outputs(5009) <= not b;
    outputs(5010) <= not a;
    outputs(5011) <= b;
    outputs(5012) <= not a;
    outputs(5013) <= b;
    outputs(5014) <= b;
    outputs(5015) <= b and not a;
    outputs(5016) <= a xor b;
    outputs(5017) <= a and not b;
    outputs(5018) <= not b or a;
    outputs(5019) <= not a;
    outputs(5020) <= b;
    outputs(5021) <= a or b;
    outputs(5022) <= not (a xor b);
    outputs(5023) <= a xor b;
    outputs(5024) <= a;
    outputs(5025) <= a xor b;
    outputs(5026) <= not (a xor b);
    outputs(5027) <= a xor b;
    outputs(5028) <= b;
    outputs(5029) <= not b;
    outputs(5030) <= not b;
    outputs(5031) <= not (a xor b);
    outputs(5032) <= b and not a;
    outputs(5033) <= not (a or b);
    outputs(5034) <= b;
    outputs(5035) <= b and not a;
    outputs(5036) <= a xor b;
    outputs(5037) <= a xor b;
    outputs(5038) <= not a;
    outputs(5039) <= b;
    outputs(5040) <= a;
    outputs(5041) <= a and not b;
    outputs(5042) <= not a;
    outputs(5043) <= a xor b;
    outputs(5044) <= not b or a;
    outputs(5045) <= b;
    outputs(5046) <= a xor b;
    outputs(5047) <= not (a or b);
    outputs(5048) <= b;
    outputs(5049) <= not a;
    outputs(5050) <= not a;
    outputs(5051) <= a and not b;
    outputs(5052) <= not (a xor b);
    outputs(5053) <= a;
    outputs(5054) <= b;
    outputs(5055) <= not a;
    outputs(5056) <= a xor b;
    outputs(5057) <= a xor b;
    outputs(5058) <= b and not a;
    outputs(5059) <= a and b;
    outputs(5060) <= not a;
    outputs(5061) <= a xor b;
    outputs(5062) <= not (a or b);
    outputs(5063) <= b and not a;
    outputs(5064) <= not (a xor b);
    outputs(5065) <= not (a xor b);
    outputs(5066) <= not b or a;
    outputs(5067) <= a xor b;
    outputs(5068) <= b;
    outputs(5069) <= not (a xor b);
    outputs(5070) <= a or b;
    outputs(5071) <= a xor b;
    outputs(5072) <= a xor b;
    outputs(5073) <= b;
    outputs(5074) <= not a;
    outputs(5075) <= a xor b;
    outputs(5076) <= not (a xor b);
    outputs(5077) <= not b;
    outputs(5078) <= b;
    outputs(5079) <= not (a xor b);
    outputs(5080) <= not (a xor b);
    outputs(5081) <= a;
    outputs(5082) <= a and b;
    outputs(5083) <= a;
    outputs(5084) <= not a;
    outputs(5085) <= not (a xor b);
    outputs(5086) <= a;
    outputs(5087) <= a;
    outputs(5088) <= not b or a;
    outputs(5089) <= not b;
    outputs(5090) <= b and not a;
    outputs(5091) <= not (a or b);
    outputs(5092) <= a;
    outputs(5093) <= not b;
    outputs(5094) <= a or b;
    outputs(5095) <= not b;
    outputs(5096) <= a xor b;
    outputs(5097) <= not b;
    outputs(5098) <= a xor b;
    outputs(5099) <= b;
    outputs(5100) <= a and not b;
    outputs(5101) <= a xor b;
    outputs(5102) <= a and not b;
    outputs(5103) <= not (a xor b);
    outputs(5104) <= a;
    outputs(5105) <= not (a xor b);
    outputs(5106) <= not b or a;
    outputs(5107) <= not (a xor b);
    outputs(5108) <= b and not a;
    outputs(5109) <= a and not b;
    outputs(5110) <= a and not b;
    outputs(5111) <= a xor b;
    outputs(5112) <= a xor b;
    outputs(5113) <= not (a xor b);
    outputs(5114) <= a and b;
    outputs(5115) <= a xor b;
    outputs(5116) <= not b;
    outputs(5117) <= a;
    outputs(5118) <= a xor b;
    outputs(5119) <= not (a or b);
    outputs(5120) <= not a;
    outputs(5121) <= a;
    outputs(5122) <= b;
    outputs(5123) <= not b;
    outputs(5124) <= not b;
    outputs(5125) <= b;
    outputs(5126) <= a;
    outputs(5127) <= a;
    outputs(5128) <= not (a xor b);
    outputs(5129) <= not b;
    outputs(5130) <= a xor b;
    outputs(5131) <= a and b;
    outputs(5132) <= not (a xor b);
    outputs(5133) <= not (a xor b);
    outputs(5134) <= a;
    outputs(5135) <= not a or b;
    outputs(5136) <= not a;
    outputs(5137) <= not a;
    outputs(5138) <= a;
    outputs(5139) <= not b;
    outputs(5140) <= not (a xor b);
    outputs(5141) <= a;
    outputs(5142) <= a xor b;
    outputs(5143) <= a xor b;
    outputs(5144) <= a xor b;
    outputs(5145) <= not b;
    outputs(5146) <= not (a xor b);
    outputs(5147) <= a xor b;
    outputs(5148) <= not a;
    outputs(5149) <= a or b;
    outputs(5150) <= not a;
    outputs(5151) <= not b;
    outputs(5152) <= not b or a;
    outputs(5153) <= a xor b;
    outputs(5154) <= not a;
    outputs(5155) <= not (a and b);
    outputs(5156) <= a xor b;
    outputs(5157) <= a xor b;
    outputs(5158) <= not b;
    outputs(5159) <= a;
    outputs(5160) <= not a;
    outputs(5161) <= not a;
    outputs(5162) <= a;
    outputs(5163) <= a;
    outputs(5164) <= not (a and b);
    outputs(5165) <= not a;
    outputs(5166) <= not (a xor b);
    outputs(5167) <= b;
    outputs(5168) <= not (a xor b);
    outputs(5169) <= not b;
    outputs(5170) <= not a;
    outputs(5171) <= not (a or b);
    outputs(5172) <= a;
    outputs(5173) <= a and not b;
    outputs(5174) <= a xor b;
    outputs(5175) <= b;
    outputs(5176) <= not (a or b);
    outputs(5177) <= b;
    outputs(5178) <= a;
    outputs(5179) <= a xor b;
    outputs(5180) <= not (a and b);
    outputs(5181) <= a and b;
    outputs(5182) <= a xor b;
    outputs(5183) <= a and not b;
    outputs(5184) <= not a or b;
    outputs(5185) <= b;
    outputs(5186) <= not (a xor b);
    outputs(5187) <= not (a or b);
    outputs(5188) <= a xor b;
    outputs(5189) <= a;
    outputs(5190) <= a;
    outputs(5191) <= a xor b;
    outputs(5192) <= a or b;
    outputs(5193) <= not a;
    outputs(5194) <= a;
    outputs(5195) <= not b or a;
    outputs(5196) <= a and not b;
    outputs(5197) <= a xor b;
    outputs(5198) <= b;
    outputs(5199) <= a;
    outputs(5200) <= a;
    outputs(5201) <= a xor b;
    outputs(5202) <= not (a xor b);
    outputs(5203) <= a or b;
    outputs(5204) <= a and not b;
    outputs(5205) <= b;
    outputs(5206) <= not (a xor b);
    outputs(5207) <= not b;
    outputs(5208) <= a xor b;
    outputs(5209) <= b;
    outputs(5210) <= not a;
    outputs(5211) <= a xor b;
    outputs(5212) <= b;
    outputs(5213) <= not (a xor b);
    outputs(5214) <= not a;
    outputs(5215) <= not b;
    outputs(5216) <= not (a xor b);
    outputs(5217) <= a and b;
    outputs(5218) <= not (a xor b);
    outputs(5219) <= a xor b;
    outputs(5220) <= a and b;
    outputs(5221) <= not a or b;
    outputs(5222) <= not b;
    outputs(5223) <= a;
    outputs(5224) <= a;
    outputs(5225) <= a;
    outputs(5226) <= b;
    outputs(5227) <= a;
    outputs(5228) <= not b;
    outputs(5229) <= a xor b;
    outputs(5230) <= a and not b;
    outputs(5231) <= b;
    outputs(5232) <= b;
    outputs(5233) <= a and b;
    outputs(5234) <= b;
    outputs(5235) <= a or b;
    outputs(5236) <= not b;
    outputs(5237) <= a;
    outputs(5238) <= not a;
    outputs(5239) <= b and not a;
    outputs(5240) <= not (a xor b);
    outputs(5241) <= not (a xor b);
    outputs(5242) <= a;
    outputs(5243) <= a and not b;
    outputs(5244) <= not b or a;
    outputs(5245) <= not (a xor b);
    outputs(5246) <= not b;
    outputs(5247) <= not (a xor b);
    outputs(5248) <= not a;
    outputs(5249) <= not (a xor b);
    outputs(5250) <= a xor b;
    outputs(5251) <= not (a xor b);
    outputs(5252) <= a;
    outputs(5253) <= not b or a;
    outputs(5254) <= b;
    outputs(5255) <= not (a and b);
    outputs(5256) <= not (a xor b);
    outputs(5257) <= not b;
    outputs(5258) <= not a;
    outputs(5259) <= not a or b;
    outputs(5260) <= not b;
    outputs(5261) <= not (a xor b);
    outputs(5262) <= b;
    outputs(5263) <= not a or b;
    outputs(5264) <= not a;
    outputs(5265) <= not (a xor b);
    outputs(5266) <= not (a xor b);
    outputs(5267) <= not a;
    outputs(5268) <= a xor b;
    outputs(5269) <= b;
    outputs(5270) <= a xor b;
    outputs(5271) <= not b;
    outputs(5272) <= a;
    outputs(5273) <= a xor b;
    outputs(5274) <= a xor b;
    outputs(5275) <= a;
    outputs(5276) <= not (a xor b);
    outputs(5277) <= not a;
    outputs(5278) <= not b;
    outputs(5279) <= not b or a;
    outputs(5280) <= b;
    outputs(5281) <= not b or a;
    outputs(5282) <= not a;
    outputs(5283) <= a and not b;
    outputs(5284) <= a xor b;
    outputs(5285) <= not a or b;
    outputs(5286) <= not b;
    outputs(5287) <= not (a xor b);
    outputs(5288) <= a and not b;
    outputs(5289) <= b and not a;
    outputs(5290) <= a and b;
    outputs(5291) <= not a;
    outputs(5292) <= not b;
    outputs(5293) <= not b or a;
    outputs(5294) <= b;
    outputs(5295) <= b;
    outputs(5296) <= not (a xor b);
    outputs(5297) <= not b;
    outputs(5298) <= not a;
    outputs(5299) <= a;
    outputs(5300) <= not (a or b);
    outputs(5301) <= not (a xor b);
    outputs(5302) <= a;
    outputs(5303) <= not (a xor b);
    outputs(5304) <= a xor b;
    outputs(5305) <= a xor b;
    outputs(5306) <= a xor b;
    outputs(5307) <= a;
    outputs(5308) <= a and b;
    outputs(5309) <= not (a xor b);
    outputs(5310) <= not b;
    outputs(5311) <= not (a xor b);
    outputs(5312) <= not b;
    outputs(5313) <= not a;
    outputs(5314) <= not (a xor b);
    outputs(5315) <= not a;
    outputs(5316) <= a xor b;
    outputs(5317) <= a xor b;
    outputs(5318) <= not a;
    outputs(5319) <= a xor b;
    outputs(5320) <= not (a xor b);
    outputs(5321) <= a xor b;
    outputs(5322) <= not (a xor b);
    outputs(5323) <= not (a xor b);
    outputs(5324) <= a or b;
    outputs(5325) <= not a;
    outputs(5326) <= not a;
    outputs(5327) <= b;
    outputs(5328) <= a and b;
    outputs(5329) <= a and not b;
    outputs(5330) <= not (a xor b);
    outputs(5331) <= a xor b;
    outputs(5332) <= not (a xor b);
    outputs(5333) <= a xor b;
    outputs(5334) <= b;
    outputs(5335) <= b and not a;
    outputs(5336) <= a;
    outputs(5337) <= not a;
    outputs(5338) <= a xor b;
    outputs(5339) <= a xor b;
    outputs(5340) <= b;
    outputs(5341) <= not a;
    outputs(5342) <= not (a xor b);
    outputs(5343) <= b;
    outputs(5344) <= a and not b;
    outputs(5345) <= not a;
    outputs(5346) <= a;
    outputs(5347) <= not (a xor b);
    outputs(5348) <= a;
    outputs(5349) <= a;
    outputs(5350) <= not b;
    outputs(5351) <= not (a xor b);
    outputs(5352) <= not a;
    outputs(5353) <= a xor b;
    outputs(5354) <= a;
    outputs(5355) <= not a;
    outputs(5356) <= not (a and b);
    outputs(5357) <= b;
    outputs(5358) <= not b;
    outputs(5359) <= a xor b;
    outputs(5360) <= a and not b;
    outputs(5361) <= a xor b;
    outputs(5362) <= a and not b;
    outputs(5363) <= b;
    outputs(5364) <= b;
    outputs(5365) <= not a;
    outputs(5366) <= b;
    outputs(5367) <= not a or b;
    outputs(5368) <= not b or a;
    outputs(5369) <= a and b;
    outputs(5370) <= a and b;
    outputs(5371) <= not (a xor b);
    outputs(5372) <= not (a or b);
    outputs(5373) <= a xor b;
    outputs(5374) <= not b;
    outputs(5375) <= not a;
    outputs(5376) <= b;
    outputs(5377) <= not b or a;
    outputs(5378) <= not b;
    outputs(5379) <= a;
    outputs(5380) <= not (a xor b);
    outputs(5381) <= not b;
    outputs(5382) <= a;
    outputs(5383) <= a xor b;
    outputs(5384) <= not (a or b);
    outputs(5385) <= a xor b;
    outputs(5386) <= a;
    outputs(5387) <= b;
    outputs(5388) <= a xor b;
    outputs(5389) <= not (a xor b);
    outputs(5390) <= b;
    outputs(5391) <= not a;
    outputs(5392) <= b and not a;
    outputs(5393) <= a;
    outputs(5394) <= a;
    outputs(5395) <= a xor b;
    outputs(5396) <= not a;
    outputs(5397) <= b;
    outputs(5398) <= a;
    outputs(5399) <= not a;
    outputs(5400) <= a xor b;
    outputs(5401) <= b;
    outputs(5402) <= a and not b;
    outputs(5403) <= a xor b;
    outputs(5404) <= a xor b;
    outputs(5405) <= a xor b;
    outputs(5406) <= a xor b;
    outputs(5407) <= not a;
    outputs(5408) <= not b;
    outputs(5409) <= not b;
    outputs(5410) <= a xor b;
    outputs(5411) <= not (a xor b);
    outputs(5412) <= not a;
    outputs(5413) <= a xor b;
    outputs(5414) <= not a;
    outputs(5415) <= a;
    outputs(5416) <= not b;
    outputs(5417) <= a xor b;
    outputs(5418) <= b;
    outputs(5419) <= a xor b;
    outputs(5420) <= a xor b;
    outputs(5421) <= a;
    outputs(5422) <= not (a xor b);
    outputs(5423) <= not (a xor b);
    outputs(5424) <= not b;
    outputs(5425) <= not (a xor b);
    outputs(5426) <= not a;
    outputs(5427) <= not (a or b);
    outputs(5428) <= a and b;
    outputs(5429) <= not (a xor b);
    outputs(5430) <= a;
    outputs(5431) <= a and not b;
    outputs(5432) <= a xor b;
    outputs(5433) <= not (a xor b);
    outputs(5434) <= a xor b;
    outputs(5435) <= a or b;
    outputs(5436) <= b and not a;
    outputs(5437) <= a xor b;
    outputs(5438) <= b;
    outputs(5439) <= not (a xor b);
    outputs(5440) <= not b;
    outputs(5441) <= a;
    outputs(5442) <= b;
    outputs(5443) <= not a;
    outputs(5444) <= not b;
    outputs(5445) <= not a;
    outputs(5446) <= b;
    outputs(5447) <= a or b;
    outputs(5448) <= not a or b;
    outputs(5449) <= a;
    outputs(5450) <= a xor b;
    outputs(5451) <= b and not a;
    outputs(5452) <= a xor b;
    outputs(5453) <= b;
    outputs(5454) <= not a or b;
    outputs(5455) <= a xor b;
    outputs(5456) <= not b;
    outputs(5457) <= not (a and b);
    outputs(5458) <= not b or a;
    outputs(5459) <= a xor b;
    outputs(5460) <= a xor b;
    outputs(5461) <= a;
    outputs(5462) <= not (a xor b);
    outputs(5463) <= a and not b;
    outputs(5464) <= not b;
    outputs(5465) <= not b;
    outputs(5466) <= not a;
    outputs(5467) <= not (a xor b);
    outputs(5468) <= a xor b;
    outputs(5469) <= a;
    outputs(5470) <= a;
    outputs(5471) <= a;
    outputs(5472) <= not b;
    outputs(5473) <= not a;
    outputs(5474) <= not a;
    outputs(5475) <= not a;
    outputs(5476) <= not a;
    outputs(5477) <= not (a and b);
    outputs(5478) <= a xor b;
    outputs(5479) <= not a;
    outputs(5480) <= not b or a;
    outputs(5481) <= a;
    outputs(5482) <= a or b;
    outputs(5483) <= b;
    outputs(5484) <= a xor b;
    outputs(5485) <= a xor b;
    outputs(5486) <= not (a xor b);
    outputs(5487) <= b and not a;
    outputs(5488) <= not a;
    outputs(5489) <= not a or b;
    outputs(5490) <= a xor b;
    outputs(5491) <= not a;
    outputs(5492) <= a and not b;
    outputs(5493) <= not a;
    outputs(5494) <= b;
    outputs(5495) <= a;
    outputs(5496) <= not a;
    outputs(5497) <= not (a xor b);
    outputs(5498) <= a xor b;
    outputs(5499) <= not b;
    outputs(5500) <= not a or b;
    outputs(5501) <= a;
    outputs(5502) <= a xor b;
    outputs(5503) <= not (a xor b);
    outputs(5504) <= not a;
    outputs(5505) <= not a or b;
    outputs(5506) <= not b;
    outputs(5507) <= a xor b;
    outputs(5508) <= not a;
    outputs(5509) <= not (a xor b);
    outputs(5510) <= not a;
    outputs(5511) <= not a;
    outputs(5512) <= a xor b;
    outputs(5513) <= not (a xor b);
    outputs(5514) <= not (a xor b);
    outputs(5515) <= a;
    outputs(5516) <= not (a xor b);
    outputs(5517) <= b;
    outputs(5518) <= not (a xor b);
    outputs(5519) <= a;
    outputs(5520) <= a xor b;
    outputs(5521) <= b and not a;
    outputs(5522) <= a and b;
    outputs(5523) <= not a;
    outputs(5524) <= not (a xor b);
    outputs(5525) <= a xor b;
    outputs(5526) <= not a;
    outputs(5527) <= not (a xor b);
    outputs(5528) <= not a or b;
    outputs(5529) <= a xor b;
    outputs(5530) <= not b;
    outputs(5531) <= a xor b;
    outputs(5532) <= a;
    outputs(5533) <= a or b;
    outputs(5534) <= b;
    outputs(5535) <= b;
    outputs(5536) <= b;
    outputs(5537) <= not b;
    outputs(5538) <= not b;
    outputs(5539) <= a;
    outputs(5540) <= not a;
    outputs(5541) <= not (a xor b);
    outputs(5542) <= a xor b;
    outputs(5543) <= b and not a;
    outputs(5544) <= not b;
    outputs(5545) <= a xor b;
    outputs(5546) <= not (a xor b);
    outputs(5547) <= a xor b;
    outputs(5548) <= not b;
    outputs(5549) <= b;
    outputs(5550) <= not (a xor b);
    outputs(5551) <= not (a xor b);
    outputs(5552) <= a;
    outputs(5553) <= a xor b;
    outputs(5554) <= not (a xor b);
    outputs(5555) <= not a;
    outputs(5556) <= not b;
    outputs(5557) <= not (a xor b);
    outputs(5558) <= a or b;
    outputs(5559) <= a xor b;
    outputs(5560) <= b;
    outputs(5561) <= a;
    outputs(5562) <= not a;
    outputs(5563) <= a;
    outputs(5564) <= a xor b;
    outputs(5565) <= not b or a;
    outputs(5566) <= a and b;
    outputs(5567) <= a xor b;
    outputs(5568) <= not a;
    outputs(5569) <= b;
    outputs(5570) <= a;
    outputs(5571) <= not b;
    outputs(5572) <= not (a and b);
    outputs(5573) <= a xor b;
    outputs(5574) <= b;
    outputs(5575) <= a and b;
    outputs(5576) <= not a;
    outputs(5577) <= not b;
    outputs(5578) <= a xor b;
    outputs(5579) <= not (a or b);
    outputs(5580) <= not a;
    outputs(5581) <= not (a xor b);
    outputs(5582) <= a;
    outputs(5583) <= not a;
    outputs(5584) <= a;
    outputs(5585) <= b;
    outputs(5586) <= a xor b;
    outputs(5587) <= not a;
    outputs(5588) <= not (a xor b);
    outputs(5589) <= not (a xor b);
    outputs(5590) <= not (a xor b);
    outputs(5591) <= not (a xor b);
    outputs(5592) <= a;
    outputs(5593) <= b and not a;
    outputs(5594) <= not (a xor b);
    outputs(5595) <= a;
    outputs(5596) <= not b;
    outputs(5597) <= b;
    outputs(5598) <= not (a xor b);
    outputs(5599) <= not a;
    outputs(5600) <= not (a and b);
    outputs(5601) <= not b;
    outputs(5602) <= a;
    outputs(5603) <= b;
    outputs(5604) <= b;
    outputs(5605) <= not a;
    outputs(5606) <= not a;
    outputs(5607) <= a;
    outputs(5608) <= a;
    outputs(5609) <= not b;
    outputs(5610) <= not (a xor b);
    outputs(5611) <= not (a xor b);
    outputs(5612) <= a xor b;
    outputs(5613) <= not (a xor b);
    outputs(5614) <= a xor b;
    outputs(5615) <= not b;
    outputs(5616) <= a;
    outputs(5617) <= a;
    outputs(5618) <= not (a xor b);
    outputs(5619) <= not b;
    outputs(5620) <= a xor b;
    outputs(5621) <= not b or a;
    outputs(5622) <= b;
    outputs(5623) <= b and not a;
    outputs(5624) <= b and not a;
    outputs(5625) <= b;
    outputs(5626) <= b;
    outputs(5627) <= b;
    outputs(5628) <= not b;
    outputs(5629) <= a xor b;
    outputs(5630) <= not a;
    outputs(5631) <= not (a xor b);
    outputs(5632) <= not (a or b);
    outputs(5633) <= a or b;
    outputs(5634) <= not b;
    outputs(5635) <= not b;
    outputs(5636) <= b;
    outputs(5637) <= a xor b;
    outputs(5638) <= a and b;
    outputs(5639) <= a xor b;
    outputs(5640) <= a or b;
    outputs(5641) <= not a;
    outputs(5642) <= not (a xor b);
    outputs(5643) <= not b;
    outputs(5644) <= b;
    outputs(5645) <= not b;
    outputs(5646) <= a xor b;
    outputs(5647) <= not a;
    outputs(5648) <= not (a xor b);
    outputs(5649) <= not a or b;
    outputs(5650) <= a xor b;
    outputs(5651) <= not (a xor b);
    outputs(5652) <= b;
    outputs(5653) <= not (a xor b);
    outputs(5654) <= b and not a;
    outputs(5655) <= a xor b;
    outputs(5656) <= not b;
    outputs(5657) <= not (a xor b);
    outputs(5658) <= a or b;
    outputs(5659) <= not a;
    outputs(5660) <= a xor b;
    outputs(5661) <= a xor b;
    outputs(5662) <= not (a xor b);
    outputs(5663) <= not b;
    outputs(5664) <= b;
    outputs(5665) <= not b or a;
    outputs(5666) <= not b;
    outputs(5667) <= a and b;
    outputs(5668) <= b;
    outputs(5669) <= not b;
    outputs(5670) <= b and not a;
    outputs(5671) <= b;
    outputs(5672) <= not a;
    outputs(5673) <= a xor b;
    outputs(5674) <= a xor b;
    outputs(5675) <= a;
    outputs(5676) <= a or b;
    outputs(5677) <= not b;
    outputs(5678) <= a xor b;
    outputs(5679) <= not b;
    outputs(5680) <= a xor b;
    outputs(5681) <= a xor b;
    outputs(5682) <= b;
    outputs(5683) <= not a or b;
    outputs(5684) <= b;
    outputs(5685) <= not b;
    outputs(5686) <= a xor b;
    outputs(5687) <= a;
    outputs(5688) <= a;
    outputs(5689) <= not a or b;
    outputs(5690) <= a or b;
    outputs(5691) <= not a;
    outputs(5692) <= a;
    outputs(5693) <= a;
    outputs(5694) <= not b;
    outputs(5695) <= not (a or b);
    outputs(5696) <= b;
    outputs(5697) <= not a or b;
    outputs(5698) <= not (a xor b);
    outputs(5699) <= a xor b;
    outputs(5700) <= not b;
    outputs(5701) <= not (a xor b);
    outputs(5702) <= a xor b;
    outputs(5703) <= not b;
    outputs(5704) <= b;
    outputs(5705) <= not a;
    outputs(5706) <= not (a and b);
    outputs(5707) <= not a;
    outputs(5708) <= not a;
    outputs(5709) <= a;
    outputs(5710) <= not (a and b);
    outputs(5711) <= a;
    outputs(5712) <= a xor b;
    outputs(5713) <= b;
    outputs(5714) <= not (a xor b);
    outputs(5715) <= not (a xor b);
    outputs(5716) <= a or b;
    outputs(5717) <= not (a xor b);
    outputs(5718) <= not b;
    outputs(5719) <= not a;
    outputs(5720) <= b;
    outputs(5721) <= a and not b;
    outputs(5722) <= not (a and b);
    outputs(5723) <= b;
    outputs(5724) <= not b;
    outputs(5725) <= not b;
    outputs(5726) <= a xor b;
    outputs(5727) <= a and b;
    outputs(5728) <= not b;
    outputs(5729) <= a and b;
    outputs(5730) <= not (a xor b);
    outputs(5731) <= a xor b;
    outputs(5732) <= a xor b;
    outputs(5733) <= not b;
    outputs(5734) <= b and not a;
    outputs(5735) <= b;
    outputs(5736) <= a xor b;
    outputs(5737) <= not b;
    outputs(5738) <= not (a or b);
    outputs(5739) <= a and b;
    outputs(5740) <= not a;
    outputs(5741) <= a xor b;
    outputs(5742) <= not b or a;
    outputs(5743) <= not a;
    outputs(5744) <= not b;
    outputs(5745) <= a;
    outputs(5746) <= b;
    outputs(5747) <= not b or a;
    outputs(5748) <= a and b;
    outputs(5749) <= a;
    outputs(5750) <= not b;
    outputs(5751) <= not a;
    outputs(5752) <= not (a xor b);
    outputs(5753) <= not a;
    outputs(5754) <= b;
    outputs(5755) <= a and b;
    outputs(5756) <= not a;
    outputs(5757) <= a xor b;
    outputs(5758) <= not a;
    outputs(5759) <= not (a and b);
    outputs(5760) <= b;
    outputs(5761) <= not (a xor b);
    outputs(5762) <= a xor b;
    outputs(5763) <= a xor b;
    outputs(5764) <= not (a xor b);
    outputs(5765) <= b;
    outputs(5766) <= not (a xor b);
    outputs(5767) <= a;
    outputs(5768) <= not a or b;
    outputs(5769) <= not (a xor b);
    outputs(5770) <= not a;
    outputs(5771) <= a or b;
    outputs(5772) <= not a or b;
    outputs(5773) <= b;
    outputs(5774) <= not (a or b);
    outputs(5775) <= not (a xor b);
    outputs(5776) <= b;
    outputs(5777) <= a;
    outputs(5778) <= a xor b;
    outputs(5779) <= b;
    outputs(5780) <= not (a xor b);
    outputs(5781) <= not (a xor b);
    outputs(5782) <= a xor b;
    outputs(5783) <= not (a or b);
    outputs(5784) <= not a or b;
    outputs(5785) <= a xor b;
    outputs(5786) <= b;
    outputs(5787) <= a;
    outputs(5788) <= a and not b;
    outputs(5789) <= not (a xor b);
    outputs(5790) <= a xor b;
    outputs(5791) <= a xor b;
    outputs(5792) <= not a;
    outputs(5793) <= not a;
    outputs(5794) <= not (a xor b);
    outputs(5795) <= a and not b;
    outputs(5796) <= a xor b;
    outputs(5797) <= not (a xor b);
    outputs(5798) <= not b;
    outputs(5799) <= a or b;
    outputs(5800) <= a;
    outputs(5801) <= a and not b;
    outputs(5802) <= a xor b;
    outputs(5803) <= not a;
    outputs(5804) <= b;
    outputs(5805) <= b;
    outputs(5806) <= a xor b;
    outputs(5807) <= a xor b;
    outputs(5808) <= a xor b;
    outputs(5809) <= b;
    outputs(5810) <= not a or b;
    outputs(5811) <= not a;
    outputs(5812) <= not b;
    outputs(5813) <= a xor b;
    outputs(5814) <= not (a xor b);
    outputs(5815) <= b;
    outputs(5816) <= a xor b;
    outputs(5817) <= a;
    outputs(5818) <= not (a xor b);
    outputs(5819) <= a;
    outputs(5820) <= not a;
    outputs(5821) <= b;
    outputs(5822) <= not a or b;
    outputs(5823) <= a and b;
    outputs(5824) <= not (a and b);
    outputs(5825) <= not b;
    outputs(5826) <= a and b;
    outputs(5827) <= a and b;
    outputs(5828) <= b;
    outputs(5829) <= not b;
    outputs(5830) <= a xor b;
    outputs(5831) <= not (a xor b);
    outputs(5832) <= a;
    outputs(5833) <= not b;
    outputs(5834) <= not (a xor b);
    outputs(5835) <= a xor b;
    outputs(5836) <= not b or a;
    outputs(5837) <= a or b;
    outputs(5838) <= not (a xor b);
    outputs(5839) <= not a;
    outputs(5840) <= not (a xor b);
    outputs(5841) <= not b;
    outputs(5842) <= not (a or b);
    outputs(5843) <= not (a and b);
    outputs(5844) <= a xor b;
    outputs(5845) <= not (a xor b);
    outputs(5846) <= not a;
    outputs(5847) <= not b;
    outputs(5848) <= not (a xor b);
    outputs(5849) <= a and b;
    outputs(5850) <= not b;
    outputs(5851) <= a xor b;
    outputs(5852) <= a xor b;
    outputs(5853) <= not (a xor b);
    outputs(5854) <= not (a xor b);
    outputs(5855) <= a and not b;
    outputs(5856) <= b;
    outputs(5857) <= a;
    outputs(5858) <= b;
    outputs(5859) <= a or b;
    outputs(5860) <= not a;
    outputs(5861) <= a and not b;
    outputs(5862) <= not (a xor b);
    outputs(5863) <= a;
    outputs(5864) <= a and b;
    outputs(5865) <= not b;
    outputs(5866) <= not b;
    outputs(5867) <= not (a xor b);
    outputs(5868) <= not b;
    outputs(5869) <= not (a xor b);
    outputs(5870) <= not (a xor b);
    outputs(5871) <= not a;
    outputs(5872) <= not a or b;
    outputs(5873) <= a xor b;
    outputs(5874) <= not b;
    outputs(5875) <= a xor b;
    outputs(5876) <= not (a and b);
    outputs(5877) <= b;
    outputs(5878) <= not b;
    outputs(5879) <= not a;
    outputs(5880) <= not (a xor b);
    outputs(5881) <= not b or a;
    outputs(5882) <= a;
    outputs(5883) <= not (a xor b);
    outputs(5884) <= a and b;
    outputs(5885) <= not b;
    outputs(5886) <= a and not b;
    outputs(5887) <= not (a or b);
    outputs(5888) <= not (a xor b);
    outputs(5889) <= not (a xor b);
    outputs(5890) <= not a;
    outputs(5891) <= a and b;
    outputs(5892) <= not b;
    outputs(5893) <= not a;
    outputs(5894) <= not b;
    outputs(5895) <= a and not b;
    outputs(5896) <= b;
    outputs(5897) <= not b;
    outputs(5898) <= a;
    outputs(5899) <= not b or a;
    outputs(5900) <= a xor b;
    outputs(5901) <= b;
    outputs(5902) <= a xor b;
    outputs(5903) <= not b or a;
    outputs(5904) <= not a or b;
    outputs(5905) <= a xor b;
    outputs(5906) <= a xor b;
    outputs(5907) <= a;
    outputs(5908) <= a xor b;
    outputs(5909) <= a and not b;
    outputs(5910) <= a xor b;
    outputs(5911) <= not b;
    outputs(5912) <= a xor b;
    outputs(5913) <= a xor b;
    outputs(5914) <= a and not b;
    outputs(5915) <= a xor b;
    outputs(5916) <= a;
    outputs(5917) <= not a;
    outputs(5918) <= a;
    outputs(5919) <= a;
    outputs(5920) <= a;
    outputs(5921) <= a xor b;
    outputs(5922) <= not a;
    outputs(5923) <= b;
    outputs(5924) <= not (a or b);
    outputs(5925) <= a xor b;
    outputs(5926) <= b;
    outputs(5927) <= b;
    outputs(5928) <= a;
    outputs(5929) <= a xor b;
    outputs(5930) <= not a;
    outputs(5931) <= not (a and b);
    outputs(5932) <= a xor b;
    outputs(5933) <= b;
    outputs(5934) <= b;
    outputs(5935) <= b;
    outputs(5936) <= not b or a;
    outputs(5937) <= b;
    outputs(5938) <= not a or b;
    outputs(5939) <= not (a and b);
    outputs(5940) <= a xor b;
    outputs(5941) <= a xor b;
    outputs(5942) <= not (a xor b);
    outputs(5943) <= not b;
    outputs(5944) <= b;
    outputs(5945) <= a;
    outputs(5946) <= a;
    outputs(5947) <= not a;
    outputs(5948) <= b and not a;
    outputs(5949) <= a and b;
    outputs(5950) <= b and not a;
    outputs(5951) <= not a or b;
    outputs(5952) <= not b or a;
    outputs(5953) <= not (a xor b);
    outputs(5954) <= b;
    outputs(5955) <= not (a xor b);
    outputs(5956) <= a xor b;
    outputs(5957) <= b;
    outputs(5958) <= not a;
    outputs(5959) <= not (a xor b);
    outputs(5960) <= a xor b;
    outputs(5961) <= not a;
    outputs(5962) <= a xor b;
    outputs(5963) <= not a;
    outputs(5964) <= a;
    outputs(5965) <= b;
    outputs(5966) <= not (a and b);
    outputs(5967) <= b;
    outputs(5968) <= a and not b;
    outputs(5969) <= not (a and b);
    outputs(5970) <= not b;
    outputs(5971) <= b;
    outputs(5972) <= a or b;
    outputs(5973) <= a xor b;
    outputs(5974) <= a and not b;
    outputs(5975) <= a xor b;
    outputs(5976) <= not (a xor b);
    outputs(5977) <= not b or a;
    outputs(5978) <= not a;
    outputs(5979) <= b;
    outputs(5980) <= not a;
    outputs(5981) <= not (a xor b);
    outputs(5982) <= a xor b;
    outputs(5983) <= b;
    outputs(5984) <= not b;
    outputs(5985) <= b;
    outputs(5986) <= not b or a;
    outputs(5987) <= not b or a;
    outputs(5988) <= not a;
    outputs(5989) <= not (a or b);
    outputs(5990) <= not b;
    outputs(5991) <= a xor b;
    outputs(5992) <= not a;
    outputs(5993) <= b;
    outputs(5994) <= not b;
    outputs(5995) <= a;
    outputs(5996) <= a xor b;
    outputs(5997) <= not a;
    outputs(5998) <= a;
    outputs(5999) <= not a or b;
    outputs(6000) <= b;
    outputs(6001) <= not (a and b);
    outputs(6002) <= a;
    outputs(6003) <= not b;
    outputs(6004) <= b and not a;
    outputs(6005) <= a;
    outputs(6006) <= not a;
    outputs(6007) <= a xor b;
    outputs(6008) <= not (a xor b);
    outputs(6009) <= not a;
    outputs(6010) <= not (a xor b);
    outputs(6011) <= not a;
    outputs(6012) <= a and b;
    outputs(6013) <= a;
    outputs(6014) <= not b or a;
    outputs(6015) <= not b or a;
    outputs(6016) <= not (a and b);
    outputs(6017) <= a and not b;
    outputs(6018) <= a xor b;
    outputs(6019) <= not (a or b);
    outputs(6020) <= not a;
    outputs(6021) <= not (a xor b);
    outputs(6022) <= a xor b;
    outputs(6023) <= a and b;
    outputs(6024) <= not (a xor b);
    outputs(6025) <= a xor b;
    outputs(6026) <= b;
    outputs(6027) <= b;
    outputs(6028) <= not a;
    outputs(6029) <= not a;
    outputs(6030) <= not (a xor b);
    outputs(6031) <= a xor b;
    outputs(6032) <= not b;
    outputs(6033) <= a;
    outputs(6034) <= not b;
    outputs(6035) <= not (a or b);
    outputs(6036) <= a xor b;
    outputs(6037) <= not b;
    outputs(6038) <= not a;
    outputs(6039) <= a;
    outputs(6040) <= a;
    outputs(6041) <= b and not a;
    outputs(6042) <= b and not a;
    outputs(6043) <= b;
    outputs(6044) <= a xor b;
    outputs(6045) <= not a;
    outputs(6046) <= b and not a;
    outputs(6047) <= b;
    outputs(6048) <= not (a and b);
    outputs(6049) <= not b or a;
    outputs(6050) <= a xor b;
    outputs(6051) <= not (a xor b);
    outputs(6052) <= a or b;
    outputs(6053) <= not a;
    outputs(6054) <= not (a xor b);
    outputs(6055) <= not a;
    outputs(6056) <= not a or b;
    outputs(6057) <= a;
    outputs(6058) <= not a or b;
    outputs(6059) <= not (a or b);
    outputs(6060) <= a;
    outputs(6061) <= b;
    outputs(6062) <= not (a or b);
    outputs(6063) <= not b;
    outputs(6064) <= not a;
    outputs(6065) <= not (a xor b);
    outputs(6066) <= not a;
    outputs(6067) <= not b;
    outputs(6068) <= not a;
    outputs(6069) <= a and b;
    outputs(6070) <= not a;
    outputs(6071) <= a;
    outputs(6072) <= not b or a;
    outputs(6073) <= not (a and b);
    outputs(6074) <= a xor b;
    outputs(6075) <= a xor b;
    outputs(6076) <= b;
    outputs(6077) <= not a;
    outputs(6078) <= b;
    outputs(6079) <= not a;
    outputs(6080) <= a;
    outputs(6081) <= not a or b;
    outputs(6082) <= not (a xor b);
    outputs(6083) <= a xor b;
    outputs(6084) <= b;
    outputs(6085) <= a or b;
    outputs(6086) <= b and not a;
    outputs(6087) <= not b;
    outputs(6088) <= a xor b;
    outputs(6089) <= b;
    outputs(6090) <= not (a xor b);
    outputs(6091) <= a xor b;
    outputs(6092) <= a and b;
    outputs(6093) <= not (a or b);
    outputs(6094) <= a;
    outputs(6095) <= not a;
    outputs(6096) <= not (a xor b);
    outputs(6097) <= not b;
    outputs(6098) <= a xor b;
    outputs(6099) <= a;
    outputs(6100) <= b;
    outputs(6101) <= b;
    outputs(6102) <= a;
    outputs(6103) <= a;
    outputs(6104) <= a xor b;
    outputs(6105) <= b;
    outputs(6106) <= not a;
    outputs(6107) <= not (a xor b);
    outputs(6108) <= not (a xor b);
    outputs(6109) <= a xor b;
    outputs(6110) <= b;
    outputs(6111) <= not (a xor b);
    outputs(6112) <= not b;
    outputs(6113) <= not (a xor b);
    outputs(6114) <= a;
    outputs(6115) <= a xor b;
    outputs(6116) <= a xor b;
    outputs(6117) <= not (a xor b);
    outputs(6118) <= b and not a;
    outputs(6119) <= a;
    outputs(6120) <= not (a xor b);
    outputs(6121) <= not b or a;
    outputs(6122) <= b;
    outputs(6123) <= a xor b;
    outputs(6124) <= not a or b;
    outputs(6125) <= not b;
    outputs(6126) <= a;
    outputs(6127) <= a xor b;
    outputs(6128) <= b;
    outputs(6129) <= not a;
    outputs(6130) <= a or b;
    outputs(6131) <= not b;
    outputs(6132) <= a xor b;
    outputs(6133) <= not (a xor b);
    outputs(6134) <= not a;
    outputs(6135) <= not b;
    outputs(6136) <= a;
    outputs(6137) <= a xor b;
    outputs(6138) <= b and not a;
    outputs(6139) <= b;
    outputs(6140) <= a and b;
    outputs(6141) <= not (a xor b);
    outputs(6142) <= a;
    outputs(6143) <= not (a xor b);
    outputs(6144) <= not a;
    outputs(6145) <= a;
    outputs(6146) <= not a;
    outputs(6147) <= a xor b;
    outputs(6148) <= a;
    outputs(6149) <= not b;
    outputs(6150) <= not a or b;
    outputs(6151) <= not a;
    outputs(6152) <= not (a or b);
    outputs(6153) <= a or b;
    outputs(6154) <= b;
    outputs(6155) <= not b;
    outputs(6156) <= b;
    outputs(6157) <= b;
    outputs(6158) <= not a or b;
    outputs(6159) <= not b;
    outputs(6160) <= a xor b;
    outputs(6161) <= not a;
    outputs(6162) <= not a;
    outputs(6163) <= b;
    outputs(6164) <= not b;
    outputs(6165) <= a;
    outputs(6166) <= a;
    outputs(6167) <= not a or b;
    outputs(6168) <= a xor b;
    outputs(6169) <= not a;
    outputs(6170) <= a xor b;
    outputs(6171) <= b;
    outputs(6172) <= a;
    outputs(6173) <= not a;
    outputs(6174) <= not (a xor b);
    outputs(6175) <= not b;
    outputs(6176) <= not (a xor b);
    outputs(6177) <= a xor b;
    outputs(6178) <= a;
    outputs(6179) <= not a;
    outputs(6180) <= not (a or b);
    outputs(6181) <= not a;
    outputs(6182) <= a and b;
    outputs(6183) <= not (a and b);
    outputs(6184) <= a and not b;
    outputs(6185) <= not a;
    outputs(6186) <= a;
    outputs(6187) <= b;
    outputs(6188) <= not (a and b);
    outputs(6189) <= b;
    outputs(6190) <= a;
    outputs(6191) <= not a;
    outputs(6192) <= not b;
    outputs(6193) <= not b;
    outputs(6194) <= b and not a;
    outputs(6195) <= a;
    outputs(6196) <= a and b;
    outputs(6197) <= b;
    outputs(6198) <= a;
    outputs(6199) <= not b;
    outputs(6200) <= a and not b;
    outputs(6201) <= not a;
    outputs(6202) <= not a;
    outputs(6203) <= not a or b;
    outputs(6204) <= a and b;
    outputs(6205) <= a xor b;
    outputs(6206) <= b;
    outputs(6207) <= not b;
    outputs(6208) <= a;
    outputs(6209) <= not (a xor b);
    outputs(6210) <= b and not a;
    outputs(6211) <= not a;
    outputs(6212) <= b;
    outputs(6213) <= not b;
    outputs(6214) <= not (a or b);
    outputs(6215) <= b;
    outputs(6216) <= not a;
    outputs(6217) <= not (a or b);
    outputs(6218) <= not (a and b);
    outputs(6219) <= not (a or b);
    outputs(6220) <= a xor b;
    outputs(6221) <= a xor b;
    outputs(6222) <= a xor b;
    outputs(6223) <= not (a or b);
    outputs(6224) <= a;
    outputs(6225) <= not b;
    outputs(6226) <= a xor b;
    outputs(6227) <= not a;
    outputs(6228) <= not a or b;
    outputs(6229) <= a xor b;
    outputs(6230) <= not b;
    outputs(6231) <= not a;
    outputs(6232) <= b;
    outputs(6233) <= a xor b;
    outputs(6234) <= not (a xor b);
    outputs(6235) <= not (a xor b);
    outputs(6236) <= not (a xor b);
    outputs(6237) <= a;
    outputs(6238) <= not a or b;
    outputs(6239) <= not b;
    outputs(6240) <= not (a xor b);
    outputs(6241) <= not (a or b);
    outputs(6242) <= a and not b;
    outputs(6243) <= b;
    outputs(6244) <= a xor b;
    outputs(6245) <= b;
    outputs(6246) <= not (a or b);
    outputs(6247) <= not a;
    outputs(6248) <= not b;
    outputs(6249) <= not a;
    outputs(6250) <= a;
    outputs(6251) <= a and b;
    outputs(6252) <= not a;
    outputs(6253) <= not b;
    outputs(6254) <= a and b;
    outputs(6255) <= b and not a;
    outputs(6256) <= not b;
    outputs(6257) <= a;
    outputs(6258) <= b;
    outputs(6259) <= not (a xor b);
    outputs(6260) <= b;
    outputs(6261) <= not a;
    outputs(6262) <= not (a or b);
    outputs(6263) <= not (a xor b);
    outputs(6264) <= not b;
    outputs(6265) <= not (a xor b);
    outputs(6266) <= not b;
    outputs(6267) <= not a;
    outputs(6268) <= not a;
    outputs(6269) <= not b;
    outputs(6270) <= not a or b;
    outputs(6271) <= a;
    outputs(6272) <= a and not b;
    outputs(6273) <= not (a or b);
    outputs(6274) <= a;
    outputs(6275) <= a and b;
    outputs(6276) <= b;
    outputs(6277) <= b;
    outputs(6278) <= a;
    outputs(6279) <= not (a xor b);
    outputs(6280) <= not (a xor b);
    outputs(6281) <= a and not b;
    outputs(6282) <= a xor b;
    outputs(6283) <= not b;
    outputs(6284) <= b;
    outputs(6285) <= not a;
    outputs(6286) <= not b;
    outputs(6287) <= a and not b;
    outputs(6288) <= a and b;
    outputs(6289) <= not b;
    outputs(6290) <= not (a xor b);
    outputs(6291) <= not b;
    outputs(6292) <= a and b;
    outputs(6293) <= a;
    outputs(6294) <= not (a xor b);
    outputs(6295) <= a and not b;
    outputs(6296) <= b and not a;
    outputs(6297) <= a xor b;
    outputs(6298) <= not a;
    outputs(6299) <= not (a xor b);
    outputs(6300) <= b;
    outputs(6301) <= not b or a;
    outputs(6302) <= not a or b;
    outputs(6303) <= not b;
    outputs(6304) <= not (a xor b);
    outputs(6305) <= not a;
    outputs(6306) <= not b;
    outputs(6307) <= not a;
    outputs(6308) <= b;
    outputs(6309) <= not (a xor b);
    outputs(6310) <= not a;
    outputs(6311) <= b;
    outputs(6312) <= not a;
    outputs(6313) <= not (a and b);
    outputs(6314) <= not a;
    outputs(6315) <= a;
    outputs(6316) <= not b or a;
    outputs(6317) <= not (a and b);
    outputs(6318) <= not b;
    outputs(6319) <= a or b;
    outputs(6320) <= a;
    outputs(6321) <= a;
    outputs(6322) <= a xor b;
    outputs(6323) <= a xor b;
    outputs(6324) <= not (a xor b);
    outputs(6325) <= b;
    outputs(6326) <= not b;
    outputs(6327) <= a;
    outputs(6328) <= a xor b;
    outputs(6329) <= not a;
    outputs(6330) <= b;
    outputs(6331) <= not a;
    outputs(6332) <= not (a and b);
    outputs(6333) <= not (a xor b);
    outputs(6334) <= a xor b;
    outputs(6335) <= a;
    outputs(6336) <= not b or a;
    outputs(6337) <= not b;
    outputs(6338) <= a;
    outputs(6339) <= not a;
    outputs(6340) <= not a;
    outputs(6341) <= not a;
    outputs(6342) <= not (a or b);
    outputs(6343) <= b and not a;
    outputs(6344) <= a and not b;
    outputs(6345) <= not a;
    outputs(6346) <= b;
    outputs(6347) <= not b;
    outputs(6348) <= not b;
    outputs(6349) <= a and not b;
    outputs(6350) <= not b;
    outputs(6351) <= not a;
    outputs(6352) <= b;
    outputs(6353) <= not (a or b);
    outputs(6354) <= not (a xor b);
    outputs(6355) <= not b;
    outputs(6356) <= not a;
    outputs(6357) <= not (a and b);
    outputs(6358) <= not b;
    outputs(6359) <= a and b;
    outputs(6360) <= a and b;
    outputs(6361) <= a;
    outputs(6362) <= a and b;
    outputs(6363) <= not b or a;
    outputs(6364) <= not (a or b);
    outputs(6365) <= b;
    outputs(6366) <= a and b;
    outputs(6367) <= a;
    outputs(6368) <= a xor b;
    outputs(6369) <= a or b;
    outputs(6370) <= not (a or b);
    outputs(6371) <= b;
    outputs(6372) <= a xor b;
    outputs(6373) <= not b;
    outputs(6374) <= a xor b;
    outputs(6375) <= not b;
    outputs(6376) <= not a;
    outputs(6377) <= a and b;
    outputs(6378) <= not (a and b);
    outputs(6379) <= a and not b;
    outputs(6380) <= not b;
    outputs(6381) <= b;
    outputs(6382) <= b;
    outputs(6383) <= a xor b;
    outputs(6384) <= b;
    outputs(6385) <= not (a or b);
    outputs(6386) <= a and not b;
    outputs(6387) <= not b;
    outputs(6388) <= not (a xor b);
    outputs(6389) <= not a;
    outputs(6390) <= not b;
    outputs(6391) <= a;
    outputs(6392) <= b;
    outputs(6393) <= a xor b;
    outputs(6394) <= b and not a;
    outputs(6395) <= a xor b;
    outputs(6396) <= not b;
    outputs(6397) <= a and b;
    outputs(6398) <= not (a and b);
    outputs(6399) <= not a;
    outputs(6400) <= not (a xor b);
    outputs(6401) <= a and b;
    outputs(6402) <= a;
    outputs(6403) <= a;
    outputs(6404) <= not a;
    outputs(6405) <= not (a or b);
    outputs(6406) <= a xor b;
    outputs(6407) <= b and not a;
    outputs(6408) <= a xor b;
    outputs(6409) <= not (a xor b);
    outputs(6410) <= b;
    outputs(6411) <= a;
    outputs(6412) <= a or b;
    outputs(6413) <= not (a xor b);
    outputs(6414) <= a and b;
    outputs(6415) <= a xor b;
    outputs(6416) <= a xor b;
    outputs(6417) <= not (a or b);
    outputs(6418) <= a;
    outputs(6419) <= b and not a;
    outputs(6420) <= not a;
    outputs(6421) <= not b;
    outputs(6422) <= a xor b;
    outputs(6423) <= a xor b;
    outputs(6424) <= not b or a;
    outputs(6425) <= a xor b;
    outputs(6426) <= a and not b;
    outputs(6427) <= a and b;
    outputs(6428) <= not b;
    outputs(6429) <= a;
    outputs(6430) <= not (a or b);
    outputs(6431) <= a or b;
    outputs(6432) <= not b;
    outputs(6433) <= a and not b;
    outputs(6434) <= not b;
    outputs(6435) <= a xor b;
    outputs(6436) <= a;
    outputs(6437) <= a xor b;
    outputs(6438) <= not b;
    outputs(6439) <= not (a or b);
    outputs(6440) <= a;
    outputs(6441) <= b;
    outputs(6442) <= a;
    outputs(6443) <= a xor b;
    outputs(6444) <= b and not a;
    outputs(6445) <= a and b;
    outputs(6446) <= a;
    outputs(6447) <= not b;
    outputs(6448) <= not (a xor b);
    outputs(6449) <= a;
    outputs(6450) <= a;
    outputs(6451) <= not a;
    outputs(6452) <= b;
    outputs(6453) <= not (a xor b);
    outputs(6454) <= b;
    outputs(6455) <= b and not a;
    outputs(6456) <= not (a or b);
    outputs(6457) <= not (a and b);
    outputs(6458) <= not (a or b);
    outputs(6459) <= not a;
    outputs(6460) <= not b;
    outputs(6461) <= a xor b;
    outputs(6462) <= not (a xor b);
    outputs(6463) <= a;
    outputs(6464) <= not b;
    outputs(6465) <= b;
    outputs(6466) <= not b;
    outputs(6467) <= not b or a;
    outputs(6468) <= not b;
    outputs(6469) <= a;
    outputs(6470) <= a;
    outputs(6471) <= b and not a;
    outputs(6472) <= not (a or b);
    outputs(6473) <= a and b;
    outputs(6474) <= a;
    outputs(6475) <= b;
    outputs(6476) <= b;
    outputs(6477) <= not a or b;
    outputs(6478) <= not (a xor b);
    outputs(6479) <= a xor b;
    outputs(6480) <= a;
    outputs(6481) <= b and not a;
    outputs(6482) <= a xor b;
    outputs(6483) <= a xor b;
    outputs(6484) <= not a or b;
    outputs(6485) <= a and not b;
    outputs(6486) <= a and not b;
    outputs(6487) <= not (a xor b);
    outputs(6488) <= not b;
    outputs(6489) <= b;
    outputs(6490) <= a;
    outputs(6491) <= not b;
    outputs(6492) <= b;
    outputs(6493) <= a and b;
    outputs(6494) <= not b;
    outputs(6495) <= not b;
    outputs(6496) <= a;
    outputs(6497) <= not (a and b);
    outputs(6498) <= a xor b;
    outputs(6499) <= b;
    outputs(6500) <= a;
    outputs(6501) <= not b;
    outputs(6502) <= a;
    outputs(6503) <= a and not b;
    outputs(6504) <= b and not a;
    outputs(6505) <= a;
    outputs(6506) <= a or b;
    outputs(6507) <= not a;
    outputs(6508) <= not b;
    outputs(6509) <= not a;
    outputs(6510) <= not a;
    outputs(6511) <= b;
    outputs(6512) <= b;
    outputs(6513) <= b;
    outputs(6514) <= a xor b;
    outputs(6515) <= a;
    outputs(6516) <= not a;
    outputs(6517) <= b;
    outputs(6518) <= not (a xor b);
    outputs(6519) <= not b;
    outputs(6520) <= a and not b;
    outputs(6521) <= a xor b;
    outputs(6522) <= not (a or b);
    outputs(6523) <= not a;
    outputs(6524) <= not (a xor b);
    outputs(6525) <= not a;
    outputs(6526) <= not (a xor b);
    outputs(6527) <= a or b;
    outputs(6528) <= a xor b;
    outputs(6529) <= a and not b;
    outputs(6530) <= not a or b;
    outputs(6531) <= not b;
    outputs(6532) <= not (a xor b);
    outputs(6533) <= b;
    outputs(6534) <= a xor b;
    outputs(6535) <= not (a xor b);
    outputs(6536) <= not a;
    outputs(6537) <= b;
    outputs(6538) <= b;
    outputs(6539) <= b;
    outputs(6540) <= a xor b;
    outputs(6541) <= a xor b;
    outputs(6542) <= not (a xor b);
    outputs(6543) <= b;
    outputs(6544) <= not a;
    outputs(6545) <= not (a xor b);
    outputs(6546) <= b;
    outputs(6547) <= b and not a;
    outputs(6548) <= a and not b;
    outputs(6549) <= a xor b;
    outputs(6550) <= not b;
    outputs(6551) <= not a;
    outputs(6552) <= a xor b;
    outputs(6553) <= b;
    outputs(6554) <= not a;
    outputs(6555) <= not (a xor b);
    outputs(6556) <= b and not a;
    outputs(6557) <= a and not b;
    outputs(6558) <= a and b;
    outputs(6559) <= not a;
    outputs(6560) <= not (a xor b);
    outputs(6561) <= not (a xor b);
    outputs(6562) <= not b;
    outputs(6563) <= not (a or b);
    outputs(6564) <= b;
    outputs(6565) <= not a;
    outputs(6566) <= not (a or b);
    outputs(6567) <= not (a xor b);
    outputs(6568) <= not a;
    outputs(6569) <= a and b;
    outputs(6570) <= a xor b;
    outputs(6571) <= a;
    outputs(6572) <= a;
    outputs(6573) <= a xor b;
    outputs(6574) <= not b;
    outputs(6575) <= a xor b;
    outputs(6576) <= not a;
    outputs(6577) <= not b;
    outputs(6578) <= not b or a;
    outputs(6579) <= not (a xor b);
    outputs(6580) <= not b;
    outputs(6581) <= not a;
    outputs(6582) <= not a;
    outputs(6583) <= a xor b;
    outputs(6584) <= a;
    outputs(6585) <= not a;
    outputs(6586) <= a;
    outputs(6587) <= not (a xor b);
    outputs(6588) <= b and not a;
    outputs(6589) <= a and b;
    outputs(6590) <= b;
    outputs(6591) <= b;
    outputs(6592) <= not a;
    outputs(6593) <= b;
    outputs(6594) <= b;
    outputs(6595) <= b;
    outputs(6596) <= not b;
    outputs(6597) <= b;
    outputs(6598) <= a xor b;
    outputs(6599) <= b and not a;
    outputs(6600) <= not a;
    outputs(6601) <= not b;
    outputs(6602) <= a and not b;
    outputs(6603) <= b;
    outputs(6604) <= a and not b;
    outputs(6605) <= a;
    outputs(6606) <= b;
    outputs(6607) <= not a;
    outputs(6608) <= not b;
    outputs(6609) <= a xor b;
    outputs(6610) <= not b;
    outputs(6611) <= not (a xor b);
    outputs(6612) <= b;
    outputs(6613) <= b and not a;
    outputs(6614) <= not b or a;
    outputs(6615) <= a xor b;
    outputs(6616) <= not (a xor b);
    outputs(6617) <= a and not b;
    outputs(6618) <= not b;
    outputs(6619) <= b;
    outputs(6620) <= not (a xor b);
    outputs(6621) <= b;
    outputs(6622) <= a xor b;
    outputs(6623) <= not (a xor b);
    outputs(6624) <= b;
    outputs(6625) <= a;
    outputs(6626) <= not a;
    outputs(6627) <= not (a xor b);
    outputs(6628) <= b;
    outputs(6629) <= a xor b;
    outputs(6630) <= not (a xor b);
    outputs(6631) <= not b;
    outputs(6632) <= a xor b;
    outputs(6633) <= not b or a;
    outputs(6634) <= not (a and b);
    outputs(6635) <= not a;
    outputs(6636) <= not (a xor b);
    outputs(6637) <= not b or a;
    outputs(6638) <= b;
    outputs(6639) <= not b;
    outputs(6640) <= not (a xor b);
    outputs(6641) <= not (a and b);
    outputs(6642) <= not a;
    outputs(6643) <= b;
    outputs(6644) <= not a;
    outputs(6645) <= a;
    outputs(6646) <= b;
    outputs(6647) <= b;
    outputs(6648) <= b and not a;
    outputs(6649) <= a and b;
    outputs(6650) <= b and not a;
    outputs(6651) <= b;
    outputs(6652) <= b;
    outputs(6653) <= b and not a;
    outputs(6654) <= not (a or b);
    outputs(6655) <= a;
    outputs(6656) <= not (a xor b);
    outputs(6657) <= not (a xor b);
    outputs(6658) <= not b;
    outputs(6659) <= b;
    outputs(6660) <= a and not b;
    outputs(6661) <= not (a xor b);
    outputs(6662) <= b;
    outputs(6663) <= not (a or b);
    outputs(6664) <= not (a xor b);
    outputs(6665) <= not (a xor b);
    outputs(6666) <= b;
    outputs(6667) <= not (a or b);
    outputs(6668) <= a;
    outputs(6669) <= not (a xor b);
    outputs(6670) <= not a;
    outputs(6671) <= not a or b;
    outputs(6672) <= a;
    outputs(6673) <= a and b;
    outputs(6674) <= a and b;
    outputs(6675) <= not b or a;
    outputs(6676) <= not (a and b);
    outputs(6677) <= not a;
    outputs(6678) <= a;
    outputs(6679) <= not b or a;
    outputs(6680) <= not (a xor b);
    outputs(6681) <= a xor b;
    outputs(6682) <= not b;
    outputs(6683) <= b;
    outputs(6684) <= a and not b;
    outputs(6685) <= not a;
    outputs(6686) <= a xor b;
    outputs(6687) <= a;
    outputs(6688) <= not a;
    outputs(6689) <= b;
    outputs(6690) <= a;
    outputs(6691) <= a xor b;
    outputs(6692) <= a;
    outputs(6693) <= a xor b;
    outputs(6694) <= a and not b;
    outputs(6695) <= not (a or b);
    outputs(6696) <= a;
    outputs(6697) <= not b;
    outputs(6698) <= b;
    outputs(6699) <= a;
    outputs(6700) <= not b;
    outputs(6701) <= not (a xor b);
    outputs(6702) <= not a;
    outputs(6703) <= a and b;
    outputs(6704) <= a and b;
    outputs(6705) <= a xor b;
    outputs(6706) <= not (a xor b);
    outputs(6707) <= b;
    outputs(6708) <= not a;
    outputs(6709) <= not b;
    outputs(6710) <= not a;
    outputs(6711) <= not (a xor b);
    outputs(6712) <= b;
    outputs(6713) <= not a;
    outputs(6714) <= a;
    outputs(6715) <= b;
    outputs(6716) <= not (a xor b);
    outputs(6717) <= not b;
    outputs(6718) <= not a;
    outputs(6719) <= not a;
    outputs(6720) <= a and not b;
    outputs(6721) <= a;
    outputs(6722) <= a;
    outputs(6723) <= not (a or b);
    outputs(6724) <= b;
    outputs(6725) <= not b;
    outputs(6726) <= a;
    outputs(6727) <= not a;
    outputs(6728) <= a xor b;
    outputs(6729) <= a xor b;
    outputs(6730) <= not a;
    outputs(6731) <= b;
    outputs(6732) <= not a;
    outputs(6733) <= not b or a;
    outputs(6734) <= b;
    outputs(6735) <= a;
    outputs(6736) <= a xor b;
    outputs(6737) <= not (a or b);
    outputs(6738) <= not (a xor b);
    outputs(6739) <= a and b;
    outputs(6740) <= b;
    outputs(6741) <= a;
    outputs(6742) <= not b;
    outputs(6743) <= a;
    outputs(6744) <= not (a or b);
    outputs(6745) <= b;
    outputs(6746) <= not (a or b);
    outputs(6747) <= a;
    outputs(6748) <= not b;
    outputs(6749) <= not a;
    outputs(6750) <= b;
    outputs(6751) <= b and not a;
    outputs(6752) <= a;
    outputs(6753) <= not a;
    outputs(6754) <= not (a xor b);
    outputs(6755) <= not a;
    outputs(6756) <= not (a or b);
    outputs(6757) <= a and not b;
    outputs(6758) <= a;
    outputs(6759) <= a or b;
    outputs(6760) <= not a;
    outputs(6761) <= a xor b;
    outputs(6762) <= a and b;
    outputs(6763) <= a and not b;
    outputs(6764) <= not (a xor b);
    outputs(6765) <= not (a xor b);
    outputs(6766) <= a xor b;
    outputs(6767) <= a xor b;
    outputs(6768) <= not b;
    outputs(6769) <= b;
    outputs(6770) <= a xor b;
    outputs(6771) <= not a;
    outputs(6772) <= a;
    outputs(6773) <= not (a or b);
    outputs(6774) <= a xor b;
    outputs(6775) <= not (a xor b);
    outputs(6776) <= not a;
    outputs(6777) <= b and not a;
    outputs(6778) <= a;
    outputs(6779) <= not (a xor b);
    outputs(6780) <= a;
    outputs(6781) <= not a;
    outputs(6782) <= not b;
    outputs(6783) <= not b or a;
    outputs(6784) <= not (a xor b);
    outputs(6785) <= a xor b;
    outputs(6786) <= not b;
    outputs(6787) <= not (a xor b);
    outputs(6788) <= not b;
    outputs(6789) <= not a;
    outputs(6790) <= a;
    outputs(6791) <= not a;
    outputs(6792) <= a and not b;
    outputs(6793) <= not b;
    outputs(6794) <= not a;
    outputs(6795) <= b;
    outputs(6796) <= b and not a;
    outputs(6797) <= not (a xor b);
    outputs(6798) <= not a;
    outputs(6799) <= not (a or b);
    outputs(6800) <= a;
    outputs(6801) <= not (a xor b);
    outputs(6802) <= not (a and b);
    outputs(6803) <= a and not b;
    outputs(6804) <= not a;
    outputs(6805) <= b and not a;
    outputs(6806) <= not a;
    outputs(6807) <= not a;
    outputs(6808) <= not (a xor b);
    outputs(6809) <= not (a xor b);
    outputs(6810) <= b;
    outputs(6811) <= a;
    outputs(6812) <= a and b;
    outputs(6813) <= not b;
    outputs(6814) <= not a;
    outputs(6815) <= not a;
    outputs(6816) <= a and b;
    outputs(6817) <= a or b;
    outputs(6818) <= a and b;
    outputs(6819) <= not (a xor b);
    outputs(6820) <= not b;
    outputs(6821) <= not (a or b);
    outputs(6822) <= not b;
    outputs(6823) <= a xor b;
    outputs(6824) <= a or b;
    outputs(6825) <= b;
    outputs(6826) <= not (a xor b);
    outputs(6827) <= not b;
    outputs(6828) <= not (a xor b);
    outputs(6829) <= not b;
    outputs(6830) <= not (a xor b);
    outputs(6831) <= a xor b;
    outputs(6832) <= a or b;
    outputs(6833) <= b and not a;
    outputs(6834) <= b and not a;
    outputs(6835) <= b and not a;
    outputs(6836) <= a and not b;
    outputs(6837) <= not (a and b);
    outputs(6838) <= b;
    outputs(6839) <= a;
    outputs(6840) <= a;
    outputs(6841) <= b;
    outputs(6842) <= a xor b;
    outputs(6843) <= a;
    outputs(6844) <= not a;
    outputs(6845) <= a xor b;
    outputs(6846) <= a xor b;
    outputs(6847) <= not b;
    outputs(6848) <= a or b;
    outputs(6849) <= a and b;
    outputs(6850) <= not (a or b);
    outputs(6851) <= a xor b;
    outputs(6852) <= not (a xor b);
    outputs(6853) <= not b;
    outputs(6854) <= a xor b;
    outputs(6855) <= b and not a;
    outputs(6856) <= not (a xor b);
    outputs(6857) <= b;
    outputs(6858) <= not b or a;
    outputs(6859) <= not a;
    outputs(6860) <= a and b;
    outputs(6861) <= b;
    outputs(6862) <= b;
    outputs(6863) <= not (a or b);
    outputs(6864) <= not a;
    outputs(6865) <= a;
    outputs(6866) <= not (a or b);
    outputs(6867) <= not a;
    outputs(6868) <= a xor b;
    outputs(6869) <= not a;
    outputs(6870) <= a xor b;
    outputs(6871) <= not a;
    outputs(6872) <= a;
    outputs(6873) <= a and not b;
    outputs(6874) <= a xor b;
    outputs(6875) <= not (a or b);
    outputs(6876) <= a and b;
    outputs(6877) <= not a;
    outputs(6878) <= not (a or b);
    outputs(6879) <= b;
    outputs(6880) <= a and b;
    outputs(6881) <= a and not b;
    outputs(6882) <= b;
    outputs(6883) <= not a;
    outputs(6884) <= not (a xor b);
    outputs(6885) <= not b;
    outputs(6886) <= not a or b;
    outputs(6887) <= b;
    outputs(6888) <= a xor b;
    outputs(6889) <= a and not b;
    outputs(6890) <= a and not b;
    outputs(6891) <= b;
    outputs(6892) <= not b;
    outputs(6893) <= b;
    outputs(6894) <= not (a xor b);
    outputs(6895) <= not a;
    outputs(6896) <= not (a xor b);
    outputs(6897) <= b;
    outputs(6898) <= a;
    outputs(6899) <= a;
    outputs(6900) <= not b or a;
    outputs(6901) <= a xor b;
    outputs(6902) <= not a;
    outputs(6903) <= a;
    outputs(6904) <= b and not a;
    outputs(6905) <= a xor b;
    outputs(6906) <= b;
    outputs(6907) <= a and b;
    outputs(6908) <= not b;
    outputs(6909) <= not a;
    outputs(6910) <= not (a or b);
    outputs(6911) <= b;
    outputs(6912) <= not a;
    outputs(6913) <= not b;
    outputs(6914) <= a and not b;
    outputs(6915) <= not a;
    outputs(6916) <= a and b;
    outputs(6917) <= not b;
    outputs(6918) <= not (a xor b);
    outputs(6919) <= not b;
    outputs(6920) <= a xor b;
    outputs(6921) <= a;
    outputs(6922) <= b;
    outputs(6923) <= a;
    outputs(6924) <= a and b;
    outputs(6925) <= a and not b;
    outputs(6926) <= a;
    outputs(6927) <= b;
    outputs(6928) <= a and b;
    outputs(6929) <= a;
    outputs(6930) <= not a or b;
    outputs(6931) <= not a;
    outputs(6932) <= not b;
    outputs(6933) <= not a;
    outputs(6934) <= not b or a;
    outputs(6935) <= not a;
    outputs(6936) <= a xor b;
    outputs(6937) <= a and not b;
    outputs(6938) <= not b;
    outputs(6939) <= b and not a;
    outputs(6940) <= not (a xor b);
    outputs(6941) <= not a;
    outputs(6942) <= not (a or b);
    outputs(6943) <= a xor b;
    outputs(6944) <= not a;
    outputs(6945) <= not a;
    outputs(6946) <= not (a xor b);
    outputs(6947) <= not (a or b);
    outputs(6948) <= not (a or b);
    outputs(6949) <= a xor b;
    outputs(6950) <= a and b;
    outputs(6951) <= not b;
    outputs(6952) <= a xor b;
    outputs(6953) <= a;
    outputs(6954) <= b;
    outputs(6955) <= a xor b;
    outputs(6956) <= not (a xor b);
    outputs(6957) <= not a;
    outputs(6958) <= b;
    outputs(6959) <= b;
    outputs(6960) <= b;
    outputs(6961) <= b;
    outputs(6962) <= not (a xor b);
    outputs(6963) <= a xor b;
    outputs(6964) <= a;
    outputs(6965) <= not (a or b);
    outputs(6966) <= not (a xor b);
    outputs(6967) <= b and not a;
    outputs(6968) <= a and b;
    outputs(6969) <= a and b;
    outputs(6970) <= not (a xor b);
    outputs(6971) <= not b;
    outputs(6972) <= not a;
    outputs(6973) <= not (a xor b);
    outputs(6974) <= a xor b;
    outputs(6975) <= b;
    outputs(6976) <= a and not b;
    outputs(6977) <= not (a xor b);
    outputs(6978) <= not (a xor b);
    outputs(6979) <= a;
    outputs(6980) <= b;
    outputs(6981) <= a and not b;
    outputs(6982) <= a;
    outputs(6983) <= a;
    outputs(6984) <= not b;
    outputs(6985) <= a and b;
    outputs(6986) <= not b;
    outputs(6987) <= not a;
    outputs(6988) <= b;
    outputs(6989) <= a or b;
    outputs(6990) <= not b;
    outputs(6991) <= not a;
    outputs(6992) <= a xor b;
    outputs(6993) <= b and not a;
    outputs(6994) <= a;
    outputs(6995) <= not (a xor b);
    outputs(6996) <= not a;
    outputs(6997) <= not b;
    outputs(6998) <= a xor b;
    outputs(6999) <= not (a xor b);
    outputs(7000) <= b;
    outputs(7001) <= not (a and b);
    outputs(7002) <= not (a xor b);
    outputs(7003) <= b;
    outputs(7004) <= not a;
    outputs(7005) <= a or b;
    outputs(7006) <= not (a or b);
    outputs(7007) <= not (a and b);
    outputs(7008) <= a;
    outputs(7009) <= not a;
    outputs(7010) <= not (a xor b);
    outputs(7011) <= a and not b;
    outputs(7012) <= not a;
    outputs(7013) <= not b;
    outputs(7014) <= not (a xor b);
    outputs(7015) <= a;
    outputs(7016) <= a;
    outputs(7017) <= b;
    outputs(7018) <= not a;
    outputs(7019) <= b;
    outputs(7020) <= b;
    outputs(7021) <= a xor b;
    outputs(7022) <= not (a xor b);
    outputs(7023) <= a;
    outputs(7024) <= a;
    outputs(7025) <= a;
    outputs(7026) <= b;
    outputs(7027) <= b;
    outputs(7028) <= a xor b;
    outputs(7029) <= a;
    outputs(7030) <= b and not a;
    outputs(7031) <= a xor b;
    outputs(7032) <= b and not a;
    outputs(7033) <= a xor b;
    outputs(7034) <= b;
    outputs(7035) <= not (a or b);
    outputs(7036) <= not (a xor b);
    outputs(7037) <= b;
    outputs(7038) <= a;
    outputs(7039) <= a;
    outputs(7040) <= b;
    outputs(7041) <= a;
    outputs(7042) <= not a;
    outputs(7043) <= a xor b;
    outputs(7044) <= a;
    outputs(7045) <= not (a or b);
    outputs(7046) <= not a;
    outputs(7047) <= a and not b;
    outputs(7048) <= b;
    outputs(7049) <= a xor b;
    outputs(7050) <= b and not a;
    outputs(7051) <= not b;
    outputs(7052) <= a;
    outputs(7053) <= not a;
    outputs(7054) <= not a;
    outputs(7055) <= a and b;
    outputs(7056) <= a;
    outputs(7057) <= a xor b;
    outputs(7058) <= a xor b;
    outputs(7059) <= not (a or b);
    outputs(7060) <= not a;
    outputs(7061) <= not b or a;
    outputs(7062) <= not (a xor b);
    outputs(7063) <= not a;
    outputs(7064) <= a xor b;
    outputs(7065) <= a or b;
    outputs(7066) <= a;
    outputs(7067) <= a;
    outputs(7068) <= a xor b;
    outputs(7069) <= b;
    outputs(7070) <= not (a or b);
    outputs(7071) <= not (a or b);
    outputs(7072) <= a xor b;
    outputs(7073) <= a xor b;
    outputs(7074) <= not b;
    outputs(7075) <= a and b;
    outputs(7076) <= b;
    outputs(7077) <= b;
    outputs(7078) <= not (a and b);
    outputs(7079) <= not (a xor b);
    outputs(7080) <= not (a xor b);
    outputs(7081) <= not (a xor b);
    outputs(7082) <= not a or b;
    outputs(7083) <= b;
    outputs(7084) <= b and not a;
    outputs(7085) <= b and not a;
    outputs(7086) <= not a or b;
    outputs(7087) <= not (a xor b);
    outputs(7088) <= not a;
    outputs(7089) <= not b;
    outputs(7090) <= b;
    outputs(7091) <= not (a or b);
    outputs(7092) <= b;
    outputs(7093) <= a;
    outputs(7094) <= a;
    outputs(7095) <= a xor b;
    outputs(7096) <= not (a and b);
    outputs(7097) <= not (a xor b);
    outputs(7098) <= b and not a;
    outputs(7099) <= b and not a;
    outputs(7100) <= a;
    outputs(7101) <= not b;
    outputs(7102) <= not (a xor b);
    outputs(7103) <= a;
    outputs(7104) <= a;
    outputs(7105) <= not b;
    outputs(7106) <= not (a xor b);
    outputs(7107) <= b;
    outputs(7108) <= a and not b;
    outputs(7109) <= not b;
    outputs(7110) <= a;
    outputs(7111) <= b;
    outputs(7112) <= a xor b;
    outputs(7113) <= b;
    outputs(7114) <= a or b;
    outputs(7115) <= a;
    outputs(7116) <= not (a xor b);
    outputs(7117) <= a xor b;
    outputs(7118) <= b and not a;
    outputs(7119) <= a and not b;
    outputs(7120) <= a xor b;
    outputs(7121) <= a;
    outputs(7122) <= not b;
    outputs(7123) <= a and not b;
    outputs(7124) <= b;
    outputs(7125) <= a and b;
    outputs(7126) <= b;
    outputs(7127) <= not (a or b);
    outputs(7128) <= a and b;
    outputs(7129) <= not (a xor b);
    outputs(7130) <= a xor b;
    outputs(7131) <= not (a or b);
    outputs(7132) <= not b;
    outputs(7133) <= not (a xor b);
    outputs(7134) <= a;
    outputs(7135) <= b;
    outputs(7136) <= not a;
    outputs(7137) <= not (a or b);
    outputs(7138) <= a and b;
    outputs(7139) <= a and b;
    outputs(7140) <= b and not a;
    outputs(7141) <= a xor b;
    outputs(7142) <= a xor b;
    outputs(7143) <= a and b;
    outputs(7144) <= a;
    outputs(7145) <= not (a xor b);
    outputs(7146) <= a;
    outputs(7147) <= not b;
    outputs(7148) <= not a;
    outputs(7149) <= not (a xor b);
    outputs(7150) <= not b;
    outputs(7151) <= a;
    outputs(7152) <= a;
    outputs(7153) <= b;
    outputs(7154) <= b and not a;
    outputs(7155) <= a;
    outputs(7156) <= not b or a;
    outputs(7157) <= not (a or b);
    outputs(7158) <= a xor b;
    outputs(7159) <= b;
    outputs(7160) <= not (a xor b);
    outputs(7161) <= not a;
    outputs(7162) <= not a;
    outputs(7163) <= b;
    outputs(7164) <= not (a xor b);
    outputs(7165) <= b and not a;
    outputs(7166) <= not (a or b);
    outputs(7167) <= not a;
    outputs(7168) <= a xor b;
    outputs(7169) <= a xor b;
    outputs(7170) <= b;
    outputs(7171) <= b and not a;
    outputs(7172) <= not b;
    outputs(7173) <= not b;
    outputs(7174) <= not b;
    outputs(7175) <= not b;
    outputs(7176) <= a xor b;
    outputs(7177) <= a xor b;
    outputs(7178) <= not a;
    outputs(7179) <= not (a xor b);
    outputs(7180) <= a or b;
    outputs(7181) <= a and b;
    outputs(7182) <= not b or a;
    outputs(7183) <= a and b;
    outputs(7184) <= not a;
    outputs(7185) <= a xor b;
    outputs(7186) <= not (a or b);
    outputs(7187) <= not (a or b);
    outputs(7188) <= not (a xor b);
    outputs(7189) <= not b;
    outputs(7190) <= b and not a;
    outputs(7191) <= b;
    outputs(7192) <= a;
    outputs(7193) <= a xor b;
    outputs(7194) <= not b or a;
    outputs(7195) <= a;
    outputs(7196) <= not a;
    outputs(7197) <= a xor b;
    outputs(7198) <= a xor b;
    outputs(7199) <= not a;
    outputs(7200) <= b;
    outputs(7201) <= not a or b;
    outputs(7202) <= b;
    outputs(7203) <= a xor b;
    outputs(7204) <= b;
    outputs(7205) <= b;
    outputs(7206) <= a;
    outputs(7207) <= b and not a;
    outputs(7208) <= not b or a;
    outputs(7209) <= not b;
    outputs(7210) <= b;
    outputs(7211) <= not a;
    outputs(7212) <= a xor b;
    outputs(7213) <= not (a xor b);
    outputs(7214) <= b;
    outputs(7215) <= a and not b;
    outputs(7216) <= not a;
    outputs(7217) <= not a;
    outputs(7218) <= not a;
    outputs(7219) <= b;
    outputs(7220) <= a xor b;
    outputs(7221) <= not b;
    outputs(7222) <= a and b;
    outputs(7223) <= not a;
    outputs(7224) <= not b;
    outputs(7225) <= a and not b;
    outputs(7226) <= not a;
    outputs(7227) <= not b;
    outputs(7228) <= a;
    outputs(7229) <= not a;
    outputs(7230) <= not a or b;
    outputs(7231) <= a or b;
    outputs(7232) <= not (a xor b);
    outputs(7233) <= a or b;
    outputs(7234) <= not (a or b);
    outputs(7235) <= not (a xor b);
    outputs(7236) <= not (a xor b);
    outputs(7237) <= not a;
    outputs(7238) <= not b;
    outputs(7239) <= b;
    outputs(7240) <= a;
    outputs(7241) <= not a or b;
    outputs(7242) <= not (a xor b);
    outputs(7243) <= not (a xor b);
    outputs(7244) <= not a;
    outputs(7245) <= not a;
    outputs(7246) <= not b;
    outputs(7247) <= not b;
    outputs(7248) <= b and not a;
    outputs(7249) <= a xor b;
    outputs(7250) <= a xor b;
    outputs(7251) <= a;
    outputs(7252) <= a;
    outputs(7253) <= not (a and b);
    outputs(7254) <= a;
    outputs(7255) <= not b;
    outputs(7256) <= a xor b;
    outputs(7257) <= b;
    outputs(7258) <= b and not a;
    outputs(7259) <= a and b;
    outputs(7260) <= not b;
    outputs(7261) <= not (a xor b);
    outputs(7262) <= a and not b;
    outputs(7263) <= b and not a;
    outputs(7264) <= a xor b;
    outputs(7265) <= a and not b;
    outputs(7266) <= not a;
    outputs(7267) <= not a;
    outputs(7268) <= not a;
    outputs(7269) <= b and not a;
    outputs(7270) <= not b;
    outputs(7271) <= a;
    outputs(7272) <= a;
    outputs(7273) <= b;
    outputs(7274) <= b;
    outputs(7275) <= a;
    outputs(7276) <= not b;
    outputs(7277) <= not (a xor b);
    outputs(7278) <= a and b;
    outputs(7279) <= not b;
    outputs(7280) <= not b;
    outputs(7281) <= a xor b;
    outputs(7282) <= not (a xor b);
    outputs(7283) <= b;
    outputs(7284) <= a;
    outputs(7285) <= b and not a;
    outputs(7286) <= b;
    outputs(7287) <= a;
    outputs(7288) <= b and not a;
    outputs(7289) <= not (a or b);
    outputs(7290) <= b;
    outputs(7291) <= a;
    outputs(7292) <= not b;
    outputs(7293) <= b;
    outputs(7294) <= not (a or b);
    outputs(7295) <= not (a xor b);
    outputs(7296) <= a xor b;
    outputs(7297) <= b;
    outputs(7298) <= b;
    outputs(7299) <= b;
    outputs(7300) <= not a or b;
    outputs(7301) <= a and not b;
    outputs(7302) <= b;
    outputs(7303) <= a and b;
    outputs(7304) <= b and not a;
    outputs(7305) <= b;
    outputs(7306) <= not b;
    outputs(7307) <= not (a and b);
    outputs(7308) <= not b;
    outputs(7309) <= a and not b;
    outputs(7310) <= not a;
    outputs(7311) <= b;
    outputs(7312) <= a;
    outputs(7313) <= not b;
    outputs(7314) <= a;
    outputs(7315) <= not b;
    outputs(7316) <= not (a xor b);
    outputs(7317) <= b;
    outputs(7318) <= not (a or b);
    outputs(7319) <= not a;
    outputs(7320) <= a and b;
    outputs(7321) <= a xor b;
    outputs(7322) <= not a;
    outputs(7323) <= a xor b;
    outputs(7324) <= not b;
    outputs(7325) <= a;
    outputs(7326) <= b and not a;
    outputs(7327) <= a xor b;
    outputs(7328) <= not a;
    outputs(7329) <= a;
    outputs(7330) <= a xor b;
    outputs(7331) <= not b;
    outputs(7332) <= not (a xor b);
    outputs(7333) <= a or b;
    outputs(7334) <= not b;
    outputs(7335) <= not b;
    outputs(7336) <= a;
    outputs(7337) <= not a;
    outputs(7338) <= a xor b;
    outputs(7339) <= not (a xor b);
    outputs(7340) <= a xor b;
    outputs(7341) <= not (a xor b);
    outputs(7342) <= not (a xor b);
    outputs(7343) <= not (a xor b);
    outputs(7344) <= not b;
    outputs(7345) <= a;
    outputs(7346) <= not a;
    outputs(7347) <= b;
    outputs(7348) <= not b;
    outputs(7349) <= not (a xor b);
    outputs(7350) <= a and not b;
    outputs(7351) <= not a;
    outputs(7352) <= not (a and b);
    outputs(7353) <= not a;
    outputs(7354) <= not a;
    outputs(7355) <= a;
    outputs(7356) <= not a;
    outputs(7357) <= a and b;
    outputs(7358) <= not (a xor b);
    outputs(7359) <= not b;
    outputs(7360) <= b and not a;
    outputs(7361) <= a xor b;
    outputs(7362) <= b;
    outputs(7363) <= not b;
    outputs(7364) <= a and not b;
    outputs(7365) <= a xor b;
    outputs(7366) <= not (a xor b);
    outputs(7367) <= a and b;
    outputs(7368) <= a xor b;
    outputs(7369) <= not a or b;
    outputs(7370) <= not (a xor b);
    outputs(7371) <= not a;
    outputs(7372) <= not a or b;
    outputs(7373) <= not (a xor b);
    outputs(7374) <= b;
    outputs(7375) <= a and not b;
    outputs(7376) <= not b;
    outputs(7377) <= a and not b;
    outputs(7378) <= a;
    outputs(7379) <= not (a xor b);
    outputs(7380) <= a;
    outputs(7381) <= a or b;
    outputs(7382) <= a xor b;
    outputs(7383) <= not a;
    outputs(7384) <= not b;
    outputs(7385) <= a xor b;
    outputs(7386) <= not b;
    outputs(7387) <= a xor b;
    outputs(7388) <= a xor b;
    outputs(7389) <= not b or a;
    outputs(7390) <= b;
    outputs(7391) <= a xor b;
    outputs(7392) <= a xor b;
    outputs(7393) <= not a;
    outputs(7394) <= a xor b;
    outputs(7395) <= a and b;
    outputs(7396) <= not (a or b);
    outputs(7397) <= b and not a;
    outputs(7398) <= b;
    outputs(7399) <= not b;
    outputs(7400) <= a;
    outputs(7401) <= not (a xor b);
    outputs(7402) <= a and b;
    outputs(7403) <= not a or b;
    outputs(7404) <= not (a xor b);
    outputs(7405) <= b and not a;
    outputs(7406) <= b;
    outputs(7407) <= not (a xor b);
    outputs(7408) <= a;
    outputs(7409) <= not (a xor b);
    outputs(7410) <= b;
    outputs(7411) <= not b;
    outputs(7412) <= not b;
    outputs(7413) <= a xor b;
    outputs(7414) <= not a;
    outputs(7415) <= a;
    outputs(7416) <= a xor b;
    outputs(7417) <= b;
    outputs(7418) <= a;
    outputs(7419) <= not a or b;
    outputs(7420) <= not (a or b);
    outputs(7421) <= not (a xor b);
    outputs(7422) <= a;
    outputs(7423) <= not (a xor b);
    outputs(7424) <= not a;
    outputs(7425) <= not (a or b);
    outputs(7426) <= a xor b;
    outputs(7427) <= a xor b;
    outputs(7428) <= a;
    outputs(7429) <= not (a or b);
    outputs(7430) <= not a;
    outputs(7431) <= b;
    outputs(7432) <= not a;
    outputs(7433) <= not (a xor b);
    outputs(7434) <= not (a xor b);
    outputs(7435) <= a xor b;
    outputs(7436) <= a xor b;
    outputs(7437) <= not b;
    outputs(7438) <= b;
    outputs(7439) <= a and not b;
    outputs(7440) <= not a;
    outputs(7441) <= not (a or b);
    outputs(7442) <= b and not a;
    outputs(7443) <= a xor b;
    outputs(7444) <= a;
    outputs(7445) <= not (a xor b);
    outputs(7446) <= not (a or b);
    outputs(7447) <= a or b;
    outputs(7448) <= a;
    outputs(7449) <= b;
    outputs(7450) <= b and not a;
    outputs(7451) <= a xor b;
    outputs(7452) <= a or b;
    outputs(7453) <= not (a xor b);
    outputs(7454) <= not (a or b);
    outputs(7455) <= not (a or b);
    outputs(7456) <= a and not b;
    outputs(7457) <= a;
    outputs(7458) <= not a;
    outputs(7459) <= a xor b;
    outputs(7460) <= not (a or b);
    outputs(7461) <= not (a or b);
    outputs(7462) <= not (a xor b);
    outputs(7463) <= b;
    outputs(7464) <= a and not b;
    outputs(7465) <= not b;
    outputs(7466) <= not a;
    outputs(7467) <= not (a xor b);
    outputs(7468) <= not b;
    outputs(7469) <= not b;
    outputs(7470) <= a xor b;
    outputs(7471) <= not b;
    outputs(7472) <= not a;
    outputs(7473) <= not b;
    outputs(7474) <= not (a xor b);
    outputs(7475) <= not b;
    outputs(7476) <= not (a and b);
    outputs(7477) <= not (a or b);
    outputs(7478) <= not a;
    outputs(7479) <= not b;
    outputs(7480) <= a xor b;
    outputs(7481) <= not (a xor b);
    outputs(7482) <= a;
    outputs(7483) <= not a;
    outputs(7484) <= b and not a;
    outputs(7485) <= not a;
    outputs(7486) <= not (a or b);
    outputs(7487) <= not (a xor b);
    outputs(7488) <= b and not a;
    outputs(7489) <= not b;
    outputs(7490) <= not a;
    outputs(7491) <= a xor b;
    outputs(7492) <= a xor b;
    outputs(7493) <= a and b;
    outputs(7494) <= not (a xor b);
    outputs(7495) <= a xor b;
    outputs(7496) <= b;
    outputs(7497) <= not a;
    outputs(7498) <= not b;
    outputs(7499) <= not (a xor b);
    outputs(7500) <= not a;
    outputs(7501) <= a;
    outputs(7502) <= not b;
    outputs(7503) <= a and b;
    outputs(7504) <= b;
    outputs(7505) <= not (a xor b);
    outputs(7506) <= not (a or b);
    outputs(7507) <= not b;
    outputs(7508) <= a;
    outputs(7509) <= a and not b;
    outputs(7510) <= a and not b;
    outputs(7511) <= a;
    outputs(7512) <= not a;
    outputs(7513) <= a xor b;
    outputs(7514) <= b and not a;
    outputs(7515) <= a;
    outputs(7516) <= not b or a;
    outputs(7517) <= a xor b;
    outputs(7518) <= b;
    outputs(7519) <= b;
    outputs(7520) <= not a;
    outputs(7521) <= not b;
    outputs(7522) <= not a or b;
    outputs(7523) <= not (a xor b);
    outputs(7524) <= not b;
    outputs(7525) <= b;
    outputs(7526) <= not a;
    outputs(7527) <= not (a or b);
    outputs(7528) <= not b;
    outputs(7529) <= a xor b;
    outputs(7530) <= not b;
    outputs(7531) <= b;
    outputs(7532) <= not (a or b);
    outputs(7533) <= b and not a;
    outputs(7534) <= a and not b;
    outputs(7535) <= not b;
    outputs(7536) <= a and not b;
    outputs(7537) <= not (a xor b);
    outputs(7538) <= not a;
    outputs(7539) <= a;
    outputs(7540) <= not a;
    outputs(7541) <= b and not a;
    outputs(7542) <= b and not a;
    outputs(7543) <= a;
    outputs(7544) <= not (a xor b);
    outputs(7545) <= not (a xor b);
    outputs(7546) <= not b;
    outputs(7547) <= b;
    outputs(7548) <= b and not a;
    outputs(7549) <= a and not b;
    outputs(7550) <= a;
    outputs(7551) <= not a;
    outputs(7552) <= not b;
    outputs(7553) <= a and b;
    outputs(7554) <= a;
    outputs(7555) <= a;
    outputs(7556) <= not a or b;
    outputs(7557) <= a xor b;
    outputs(7558) <= a and not b;
    outputs(7559) <= not (a or b);
    outputs(7560) <= b;
    outputs(7561) <= not b;
    outputs(7562) <= not (a xor b);
    outputs(7563) <= not b;
    outputs(7564) <= a and not b;
    outputs(7565) <= a xor b;
    outputs(7566) <= a and not b;
    outputs(7567) <= not a;
    outputs(7568) <= not (a xor b);
    outputs(7569) <= a;
    outputs(7570) <= not (a xor b);
    outputs(7571) <= not (a xor b);
    outputs(7572) <= a xor b;
    outputs(7573) <= not b;
    outputs(7574) <= a xor b;
    outputs(7575) <= not a;
    outputs(7576) <= not b;
    outputs(7577) <= not a;
    outputs(7578) <= not (a xor b);
    outputs(7579) <= not (a xor b);
    outputs(7580) <= a and not b;
    outputs(7581) <= a and not b;
    outputs(7582) <= a or b;
    outputs(7583) <= not (a or b);
    outputs(7584) <= not (a xor b);
    outputs(7585) <= b;
    outputs(7586) <= not (a xor b);
    outputs(7587) <= not a;
    outputs(7588) <= not b;
    outputs(7589) <= not a;
    outputs(7590) <= not (a xor b);
    outputs(7591) <= not (a or b);
    outputs(7592) <= not b;
    outputs(7593) <= not (a xor b);
    outputs(7594) <= a xor b;
    outputs(7595) <= not (a or b);
    outputs(7596) <= a and not b;
    outputs(7597) <= not (a or b);
    outputs(7598) <= a and b;
    outputs(7599) <= not a;
    outputs(7600) <= not (a xor b);
    outputs(7601) <= not (a or b);
    outputs(7602) <= not b;
    outputs(7603) <= not (a xor b);
    outputs(7604) <= a xor b;
    outputs(7605) <= not a;
    outputs(7606) <= not (a xor b);
    outputs(7607) <= not (a xor b);
    outputs(7608) <= not (a or b);
    outputs(7609) <= a and b;
    outputs(7610) <= not a or b;
    outputs(7611) <= b;
    outputs(7612) <= a xor b;
    outputs(7613) <= not (a xor b);
    outputs(7614) <= not (a xor b);
    outputs(7615) <= a and not b;
    outputs(7616) <= a;
    outputs(7617) <= a;
    outputs(7618) <= a;
    outputs(7619) <= b;
    outputs(7620) <= not (a xor b);
    outputs(7621) <= not b;
    outputs(7622) <= not (a xor b);
    outputs(7623) <= a xor b;
    outputs(7624) <= b;
    outputs(7625) <= a;
    outputs(7626) <= not a;
    outputs(7627) <= a and b;
    outputs(7628) <= not (a xor b);
    outputs(7629) <= b;
    outputs(7630) <= not a;
    outputs(7631) <= a and not b;
    outputs(7632) <= b;
    outputs(7633) <= not (a xor b);
    outputs(7634) <= not (a and b);
    outputs(7635) <= a and b;
    outputs(7636) <= a and b;
    outputs(7637) <= not a;
    outputs(7638) <= b;
    outputs(7639) <= a and b;
    outputs(7640) <= not a;
    outputs(7641) <= not b;
    outputs(7642) <= not (a xor b);
    outputs(7643) <= not (a xor b);
    outputs(7644) <= a xor b;
    outputs(7645) <= b and not a;
    outputs(7646) <= a xor b;
    outputs(7647) <= a xor b;
    outputs(7648) <= a and not b;
    outputs(7649) <= not a;
    outputs(7650) <= b;
    outputs(7651) <= a xor b;
    outputs(7652) <= not a;
    outputs(7653) <= not (a and b);
    outputs(7654) <= not a;
    outputs(7655) <= a and not b;
    outputs(7656) <= not (a xor b);
    outputs(7657) <= b;
    outputs(7658) <= a;
    outputs(7659) <= b and not a;
    outputs(7660) <= a xor b;
    outputs(7661) <= b and not a;
    outputs(7662) <= b and not a;
    outputs(7663) <= a xor b;
    outputs(7664) <= a;
    outputs(7665) <= b;
    outputs(7666) <= a;
    outputs(7667) <= b;
    outputs(7668) <= not b;
    outputs(7669) <= a;
    outputs(7670) <= not a;
    outputs(7671) <= not (a xor b);
    outputs(7672) <= not a;
    outputs(7673) <= not (a or b);
    outputs(7674) <= not a;
    outputs(7675) <= a;
    outputs(7676) <= not b;
    outputs(7677) <= not b;
    outputs(7678) <= a xor b;
    outputs(7679) <= b and not a;
    outputs(7680) <= not b;
    outputs(7681) <= not b;
    outputs(7682) <= not a;
    outputs(7683) <= a xor b;
    outputs(7684) <= a;
    outputs(7685) <= not (a xor b);
    outputs(7686) <= a xor b;
    outputs(7687) <= b and not a;
    outputs(7688) <= not b or a;
    outputs(7689) <= not a or b;
    outputs(7690) <= b and not a;
    outputs(7691) <= a;
    outputs(7692) <= a and b;
    outputs(7693) <= a and not b;
    outputs(7694) <= b;
    outputs(7695) <= not a;
    outputs(7696) <= a;
    outputs(7697) <= b and not a;
    outputs(7698) <= a xor b;
    outputs(7699) <= not b;
    outputs(7700) <= a;
    outputs(7701) <= not a;
    outputs(7702) <= not b;
    outputs(7703) <= not b or a;
    outputs(7704) <= a xor b;
    outputs(7705) <= a;
    outputs(7706) <= a and b;
    outputs(7707) <= not a;
    outputs(7708) <= not (a xor b);
    outputs(7709) <= not (a xor b);
    outputs(7710) <= not a;
    outputs(7711) <= b;
    outputs(7712) <= not (a or b);
    outputs(7713) <= not b;
    outputs(7714) <= not b;
    outputs(7715) <= a xor b;
    outputs(7716) <= not b;
    outputs(7717) <= b;
    outputs(7718) <= b;
    outputs(7719) <= b;
    outputs(7720) <= a;
    outputs(7721) <= not (a or b);
    outputs(7722) <= a;
    outputs(7723) <= not (a and b);
    outputs(7724) <= not (a xor b);
    outputs(7725) <= a xor b;
    outputs(7726) <= not b;
    outputs(7727) <= a and b;
    outputs(7728) <= b;
    outputs(7729) <= not (a xor b);
    outputs(7730) <= a;
    outputs(7731) <= not a or b;
    outputs(7732) <= a;
    outputs(7733) <= a;
    outputs(7734) <= a;
    outputs(7735) <= a and b;
    outputs(7736) <= a and not b;
    outputs(7737) <= not (a and b);
    outputs(7738) <= not (a xor b);
    outputs(7739) <= not a;
    outputs(7740) <= b;
    outputs(7741) <= a xor b;
    outputs(7742) <= a xor b;
    outputs(7743) <= not b;
    outputs(7744) <= a and not b;
    outputs(7745) <= not b;
    outputs(7746) <= b and not a;
    outputs(7747) <= b;
    outputs(7748) <= a and b;
    outputs(7749) <= not (a or b);
    outputs(7750) <= b;
    outputs(7751) <= b;
    outputs(7752) <= a xor b;
    outputs(7753) <= not (a xor b);
    outputs(7754) <= not a;
    outputs(7755) <= a;
    outputs(7756) <= not b;
    outputs(7757) <= not b;
    outputs(7758) <= a xor b;
    outputs(7759) <= a and not b;
    outputs(7760) <= not (a or b);
    outputs(7761) <= a or b;
    outputs(7762) <= not (a xor b);
    outputs(7763) <= not (a or b);
    outputs(7764) <= not b;
    outputs(7765) <= not a or b;
    outputs(7766) <= a;
    outputs(7767) <= b;
    outputs(7768) <= a xor b;
    outputs(7769) <= not a;
    outputs(7770) <= not b or a;
    outputs(7771) <= not (a and b);
    outputs(7772) <= not b;
    outputs(7773) <= b;
    outputs(7774) <= a and b;
    outputs(7775) <= not (a xor b);
    outputs(7776) <= a and not b;
    outputs(7777) <= b;
    outputs(7778) <= b;
    outputs(7779) <= not a;
    outputs(7780) <= a;
    outputs(7781) <= not (a xor b);
    outputs(7782) <= not (a or b);
    outputs(7783) <= b and not a;
    outputs(7784) <= a;
    outputs(7785) <= not (a xor b);
    outputs(7786) <= not (a xor b);
    outputs(7787) <= not (a xor b);
    outputs(7788) <= not (a or b);
    outputs(7789) <= not a;
    outputs(7790) <= a;
    outputs(7791) <= a xor b;
    outputs(7792) <= b;
    outputs(7793) <= not a;
    outputs(7794) <= a;
    outputs(7795) <= a xor b;
    outputs(7796) <= not a;
    outputs(7797) <= not b;
    outputs(7798) <= not b;
    outputs(7799) <= a;
    outputs(7800) <= a or b;
    outputs(7801) <= a xor b;
    outputs(7802) <= a;
    outputs(7803) <= not b;
    outputs(7804) <= not (a xor b);
    outputs(7805) <= a xor b;
    outputs(7806) <= a;
    outputs(7807) <= a xor b;
    outputs(7808) <= not a;
    outputs(7809) <= b;
    outputs(7810) <= a;
    outputs(7811) <= a;
    outputs(7812) <= a xor b;
    outputs(7813) <= not (a xor b);
    outputs(7814) <= not b;
    outputs(7815) <= not (a or b);
    outputs(7816) <= b and not a;
    outputs(7817) <= a xor b;
    outputs(7818) <= b;
    outputs(7819) <= not (a xor b);
    outputs(7820) <= b;
    outputs(7821) <= a xor b;
    outputs(7822) <= b and not a;
    outputs(7823) <= a and b;
    outputs(7824) <= not a or b;
    outputs(7825) <= not (a xor b);
    outputs(7826) <= a and not b;
    outputs(7827) <= a xor b;
    outputs(7828) <= not (a xor b);
    outputs(7829) <= not (a or b);
    outputs(7830) <= not a;
    outputs(7831) <= a;
    outputs(7832) <= not (a xor b);
    outputs(7833) <= a or b;
    outputs(7834) <= not (a xor b);
    outputs(7835) <= a and b;
    outputs(7836) <= b;
    outputs(7837) <= a xor b;
    outputs(7838) <= a xor b;
    outputs(7839) <= not a;
    outputs(7840) <= not b;
    outputs(7841) <= not b;
    outputs(7842) <= a and b;
    outputs(7843) <= a xor b;
    outputs(7844) <= not (a or b);
    outputs(7845) <= not (a or b);
    outputs(7846) <= b and not a;
    outputs(7847) <= not (a xor b);
    outputs(7848) <= a xor b;
    outputs(7849) <= a and b;
    outputs(7850) <= not a;
    outputs(7851) <= not a;
    outputs(7852) <= a xor b;
    outputs(7853) <= a xor b;
    outputs(7854) <= not b;
    outputs(7855) <= b;
    outputs(7856) <= not b;
    outputs(7857) <= not (a or b);
    outputs(7858) <= not b;
    outputs(7859) <= not (a and b);
    outputs(7860) <= a xor b;
    outputs(7861) <= not (a xor b);
    outputs(7862) <= not (a and b);
    outputs(7863) <= not b;
    outputs(7864) <= not (a xor b);
    outputs(7865) <= not a or b;
    outputs(7866) <= not (a xor b);
    outputs(7867) <= not (a xor b);
    outputs(7868) <= a;
    outputs(7869) <= not b;
    outputs(7870) <= a;
    outputs(7871) <= not b;
    outputs(7872) <= a and b;
    outputs(7873) <= b;
    outputs(7874) <= b and not a;
    outputs(7875) <= a;
    outputs(7876) <= a and b;
    outputs(7877) <= a or b;
    outputs(7878) <= a;
    outputs(7879) <= not (a or b);
    outputs(7880) <= not b;
    outputs(7881) <= not (a xor b);
    outputs(7882) <= not (a xor b);
    outputs(7883) <= not b or a;
    outputs(7884) <= not a;
    outputs(7885) <= b and not a;
    outputs(7886) <= not (a or b);
    outputs(7887) <= a xor b;
    outputs(7888) <= a;
    outputs(7889) <= a xor b;
    outputs(7890) <= a;
    outputs(7891) <= b;
    outputs(7892) <= a xor b;
    outputs(7893) <= a xor b;
    outputs(7894) <= not (a xor b);
    outputs(7895) <= a and not b;
    outputs(7896) <= a or b;
    outputs(7897) <= a xor b;
    outputs(7898) <= not b;
    outputs(7899) <= a xor b;
    outputs(7900) <= not b or a;
    outputs(7901) <= not b;
    outputs(7902) <= a xor b;
    outputs(7903) <= a;
    outputs(7904) <= b and not a;
    outputs(7905) <= not (a or b);
    outputs(7906) <= not (a xor b);
    outputs(7907) <= b and not a;
    outputs(7908) <= b and not a;
    outputs(7909) <= a and b;
    outputs(7910) <= a xor b;
    outputs(7911) <= not (a and b);
    outputs(7912) <= b and not a;
    outputs(7913) <= a;
    outputs(7914) <= not (a xor b);
    outputs(7915) <= a xor b;
    outputs(7916) <= a;
    outputs(7917) <= a;
    outputs(7918) <= not a;
    outputs(7919) <= b;
    outputs(7920) <= not (a xor b);
    outputs(7921) <= b;
    outputs(7922) <= not b;
    outputs(7923) <= a;
    outputs(7924) <= b;
    outputs(7925) <= not b;
    outputs(7926) <= a;
    outputs(7927) <= a xor b;
    outputs(7928) <= not (a xor b);
    outputs(7929) <= not (a and b);
    outputs(7930) <= a;
    outputs(7931) <= not (a and b);
    outputs(7932) <= a xor b;
    outputs(7933) <= a;
    outputs(7934) <= a and not b;
    outputs(7935) <= not a;
    outputs(7936) <= a xor b;
    outputs(7937) <= not a;
    outputs(7938) <= b;
    outputs(7939) <= a and b;
    outputs(7940) <= a and not b;
    outputs(7941) <= not (a xor b);
    outputs(7942) <= not (a xor b);
    outputs(7943) <= not (a xor b);
    outputs(7944) <= a;
    outputs(7945) <= not (a xor b);
    outputs(7946) <= not b;
    outputs(7947) <= not (a xor b);
    outputs(7948) <= not a;
    outputs(7949) <= not a;
    outputs(7950) <= b;
    outputs(7951) <= not a;
    outputs(7952) <= not (a xor b);
    outputs(7953) <= a and not b;
    outputs(7954) <= not b;
    outputs(7955) <= not (a or b);
    outputs(7956) <= not a or b;
    outputs(7957) <= a;
    outputs(7958) <= not a;
    outputs(7959) <= not a;
    outputs(7960) <= a xor b;
    outputs(7961) <= a;
    outputs(7962) <= a;
    outputs(7963) <= a;
    outputs(7964) <= a xor b;
    outputs(7965) <= not b;
    outputs(7966) <= not a;
    outputs(7967) <= a xor b;
    outputs(7968) <= a xor b;
    outputs(7969) <= b;
    outputs(7970) <= a xor b;
    outputs(7971) <= a and b;
    outputs(7972) <= not (a xor b);
    outputs(7973) <= not a;
    outputs(7974) <= b;
    outputs(7975) <= b;
    outputs(7976) <= not b;
    outputs(7977) <= not b;
    outputs(7978) <= b;
    outputs(7979) <= a;
    outputs(7980) <= not (a xor b);
    outputs(7981) <= a;
    outputs(7982) <= not (a xor b);
    outputs(7983) <= a and b;
    outputs(7984) <= not a or b;
    outputs(7985) <= a xor b;
    outputs(7986) <= a xor b;
    outputs(7987) <= not a;
    outputs(7988) <= not (a xor b);
    outputs(7989) <= not (a xor b);
    outputs(7990) <= b and not a;
    outputs(7991) <= a and b;
    outputs(7992) <= not a;
    outputs(7993) <= not a;
    outputs(7994) <= not (a and b);
    outputs(7995) <= b and not a;
    outputs(7996) <= a;
    outputs(7997) <= not a;
    outputs(7998) <= a;
    outputs(7999) <= not (a or b);
    outputs(8000) <= b;
    outputs(8001) <= not (a or b);
    outputs(8002) <= b;
    outputs(8003) <= b and not a;
    outputs(8004) <= not (a xor b);
    outputs(8005) <= a;
    outputs(8006) <= a and b;
    outputs(8007) <= b and not a;
    outputs(8008) <= b;
    outputs(8009) <= b and not a;
    outputs(8010) <= not a;
    outputs(8011) <= a;
    outputs(8012) <= not (a xor b);
    outputs(8013) <= not (a xor b);
    outputs(8014) <= not (a xor b);
    outputs(8015) <= not b;
    outputs(8016) <= a;
    outputs(8017) <= not (a xor b);
    outputs(8018) <= a xor b;
    outputs(8019) <= not a;
    outputs(8020) <= a;
    outputs(8021) <= not b;
    outputs(8022) <= a and b;
    outputs(8023) <= b and not a;
    outputs(8024) <= a xor b;
    outputs(8025) <= b;
    outputs(8026) <= a xor b;
    outputs(8027) <= not a;
    outputs(8028) <= b;
    outputs(8029) <= b;
    outputs(8030) <= a;
    outputs(8031) <= not (a or b);
    outputs(8032) <= not a or b;
    outputs(8033) <= a and not b;
    outputs(8034) <= b;
    outputs(8035) <= a xor b;
    outputs(8036) <= not (a xor b);
    outputs(8037) <= a;
    outputs(8038) <= a;
    outputs(8039) <= a;
    outputs(8040) <= not a;
    outputs(8041) <= a and not b;
    outputs(8042) <= a and b;
    outputs(8043) <= b and not a;
    outputs(8044) <= a;
    outputs(8045) <= not b;
    outputs(8046) <= b and not a;
    outputs(8047) <= not (a xor b);
    outputs(8048) <= not a;
    outputs(8049) <= b;
    outputs(8050) <= not a;
    outputs(8051) <= b and not a;
    outputs(8052) <= not b;
    outputs(8053) <= a xor b;
    outputs(8054) <= b;
    outputs(8055) <= b;
    outputs(8056) <= not b or a;
    outputs(8057) <= a;
    outputs(8058) <= not b;
    outputs(8059) <= a xor b;
    outputs(8060) <= b and not a;
    outputs(8061) <= a;
    outputs(8062) <= not a;
    outputs(8063) <= a and b;
    outputs(8064) <= a;
    outputs(8065) <= not (a xor b);
    outputs(8066) <= a xor b;
    outputs(8067) <= not (a xor b);
    outputs(8068) <= not (a or b);
    outputs(8069) <= a;
    outputs(8070) <= b;
    outputs(8071) <= b;
    outputs(8072) <= b and not a;
    outputs(8073) <= a;
    outputs(8074) <= not (a xor b);
    outputs(8075) <= a;
    outputs(8076) <= not b;
    outputs(8077) <= a xor b;
    outputs(8078) <= a xor b;
    outputs(8079) <= a;
    outputs(8080) <= not b;
    outputs(8081) <= not a;
    outputs(8082) <= not b;
    outputs(8083) <= a xor b;
    outputs(8084) <= not b or a;
    outputs(8085) <= not (a or b);
    outputs(8086) <= a xor b;
    outputs(8087) <= not a;
    outputs(8088) <= a xor b;
    outputs(8089) <= not (a xor b);
    outputs(8090) <= not (a or b);
    outputs(8091) <= not a or b;
    outputs(8092) <= not (a xor b);
    outputs(8093) <= not (a or b);
    outputs(8094) <= a xor b;
    outputs(8095) <= not (a or b);
    outputs(8096) <= not (a or b);
    outputs(8097) <= not a or b;
    outputs(8098) <= a xor b;
    outputs(8099) <= not (a xor b);
    outputs(8100) <= not (a xor b);
    outputs(8101) <= b;
    outputs(8102) <= not (a and b);
    outputs(8103) <= not (a xor b);
    outputs(8104) <= a xor b;
    outputs(8105) <= a and b;
    outputs(8106) <= not (a xor b);
    outputs(8107) <= not a;
    outputs(8108) <= not b;
    outputs(8109) <= b and not a;
    outputs(8110) <= not a;
    outputs(8111) <= a xor b;
    outputs(8112) <= not (a xor b);
    outputs(8113) <= b and not a;
    outputs(8114) <= not b or a;
    outputs(8115) <= not b;
    outputs(8116) <= a or b;
    outputs(8117) <= not b;
    outputs(8118) <= not (a xor b);
    outputs(8119) <= a and not b;
    outputs(8120) <= not (a xor b);
    outputs(8121) <= b;
    outputs(8122) <= not (a xor b);
    outputs(8123) <= not a;
    outputs(8124) <= b;
    outputs(8125) <= not a;
    outputs(8126) <= not a;
    outputs(8127) <= not (a or b);
    outputs(8128) <= b and not a;
    outputs(8129) <= a;
    outputs(8130) <= a;
    outputs(8131) <= not b;
    outputs(8132) <= a;
    outputs(8133) <= a;
    outputs(8134) <= a xor b;
    outputs(8135) <= a xor b;
    outputs(8136) <= a xor b;
    outputs(8137) <= a or b;
    outputs(8138) <= b;
    outputs(8139) <= not a;
    outputs(8140) <= a xor b;
    outputs(8141) <= b;
    outputs(8142) <= not b;
    outputs(8143) <= a and b;
    outputs(8144) <= a xor b;
    outputs(8145) <= a;
    outputs(8146) <= not (a xor b);
    outputs(8147) <= not (a or b);
    outputs(8148) <= a xor b;
    outputs(8149) <= a xor b;
    outputs(8150) <= a;
    outputs(8151) <= not (a xor b);
    outputs(8152) <= b;
    outputs(8153) <= not (a or b);
    outputs(8154) <= a;
    outputs(8155) <= not (a xor b);
    outputs(8156) <= not b or a;
    outputs(8157) <= a xor b;
    outputs(8158) <= not (a xor b);
    outputs(8159) <= not (a xor b);
    outputs(8160) <= b;
    outputs(8161) <= not b;
    outputs(8162) <= a xor b;
    outputs(8163) <= a;
    outputs(8164) <= a and b;
    outputs(8165) <= b;
    outputs(8166) <= not (a xor b);
    outputs(8167) <= not b;
    outputs(8168) <= not b;
    outputs(8169) <= a;
    outputs(8170) <= b;
    outputs(8171) <= a and b;
    outputs(8172) <= a xor b;
    outputs(8173) <= not b;
    outputs(8174) <= not a or b;
    outputs(8175) <= a and not b;
    outputs(8176) <= a xor b;
    outputs(8177) <= not a;
    outputs(8178) <= not b;
    outputs(8179) <= b;
    outputs(8180) <= a and b;
    outputs(8181) <= b and not a;
    outputs(8182) <= not a;
    outputs(8183) <= a;
    outputs(8184) <= not a;
    outputs(8185) <= a xor b;
    outputs(8186) <= a and b;
    outputs(8187) <= not (a xor b);
    outputs(8188) <= a xor b;
    outputs(8189) <= not (a xor b);
    outputs(8190) <= not (a or b);
    outputs(8191) <= not b;
    outputs(8192) <= not (a xor b);
    outputs(8193) <= not (a xor b);
    outputs(8194) <= not (a xor b);
    outputs(8195) <= not b;
    outputs(8196) <= a and b;
    outputs(8197) <= not (a xor b);
    outputs(8198) <= not (a xor b);
    outputs(8199) <= b;
    outputs(8200) <= a or b;
    outputs(8201) <= not b or a;
    outputs(8202) <= not a;
    outputs(8203) <= b;
    outputs(8204) <= not a or b;
    outputs(8205) <= not a or b;
    outputs(8206) <= b;
    outputs(8207) <= not (a xor b);
    outputs(8208) <= not b or a;
    outputs(8209) <= a xor b;
    outputs(8210) <= a;
    outputs(8211) <= a;
    outputs(8212) <= a xor b;
    outputs(8213) <= not (a xor b);
    outputs(8214) <= a xor b;
    outputs(8215) <= not a;
    outputs(8216) <= b;
    outputs(8217) <= not (a xor b);
    outputs(8218) <= a;
    outputs(8219) <= a xor b;
    outputs(8220) <= b and not a;
    outputs(8221) <= a xor b;
    outputs(8222) <= a;
    outputs(8223) <= not a or b;
    outputs(8224) <= not a;
    outputs(8225) <= b;
    outputs(8226) <= not (a xor b);
    outputs(8227) <= a xor b;
    outputs(8228) <= b;
    outputs(8229) <= a xor b;
    outputs(8230) <= not (a xor b);
    outputs(8231) <= b;
    outputs(8232) <= a or b;
    outputs(8233) <= b;
    outputs(8234) <= not (a and b);
    outputs(8235) <= b;
    outputs(8236) <= a or b;
    outputs(8237) <= b and not a;
    outputs(8238) <= not (a and b);
    outputs(8239) <= not (a xor b);
    outputs(8240) <= a;
    outputs(8241) <= not b;
    outputs(8242) <= not a;
    outputs(8243) <= a xor b;
    outputs(8244) <= not (a xor b);
    outputs(8245) <= not (a xor b);
    outputs(8246) <= not b or a;
    outputs(8247) <= b;
    outputs(8248) <= not a;
    outputs(8249) <= b;
    outputs(8250) <= not a or b;
    outputs(8251) <= a;
    outputs(8252) <= a;
    outputs(8253) <= a or b;
    outputs(8254) <= a xor b;
    outputs(8255) <= not (a xor b);
    outputs(8256) <= b;
    outputs(8257) <= not b or a;
    outputs(8258) <= not b or a;
    outputs(8259) <= not (a xor b);
    outputs(8260) <= b;
    outputs(8261) <= a or b;
    outputs(8262) <= a and b;
    outputs(8263) <= a or b;
    outputs(8264) <= b;
    outputs(8265) <= b;
    outputs(8266) <= not (a xor b);
    outputs(8267) <= a;
    outputs(8268) <= not b;
    outputs(8269) <= not b;
    outputs(8270) <= b and not a;
    outputs(8271) <= not (a and b);
    outputs(8272) <= not b;
    outputs(8273) <= b;
    outputs(8274) <= not b;
    outputs(8275) <= not (a or b);
    outputs(8276) <= a;
    outputs(8277) <= a or b;
    outputs(8278) <= a xor b;
    outputs(8279) <= not (a xor b);
    outputs(8280) <= not (a xor b);
    outputs(8281) <= b;
    outputs(8282) <= not (a xor b);
    outputs(8283) <= not a or b;
    outputs(8284) <= not a;
    outputs(8285) <= not a or b;
    outputs(8286) <= not b;
    outputs(8287) <= b;
    outputs(8288) <= b;
    outputs(8289) <= a and not b;
    outputs(8290) <= a;
    outputs(8291) <= not b or a;
    outputs(8292) <= not (a xor b);
    outputs(8293) <= a xor b;
    outputs(8294) <= a;
    outputs(8295) <= not (a xor b);
    outputs(8296) <= a or b;
    outputs(8297) <= not (a xor b);
    outputs(8298) <= a xor b;
    outputs(8299) <= a;
    outputs(8300) <= not (a xor b);
    outputs(8301) <= not b;
    outputs(8302) <= a or b;
    outputs(8303) <= not (a and b);
    outputs(8304) <= not (a xor b);
    outputs(8305) <= a;
    outputs(8306) <= a xor b;
    outputs(8307) <= not b or a;
    outputs(8308) <= not a;
    outputs(8309) <= a;
    outputs(8310) <= a;
    outputs(8311) <= not (a xor b);
    outputs(8312) <= not b;
    outputs(8313) <= not a;
    outputs(8314) <= a;
    outputs(8315) <= a xor b;
    outputs(8316) <= not (a xor b);
    outputs(8317) <= not a;
    outputs(8318) <= not a;
    outputs(8319) <= a xor b;
    outputs(8320) <= b;
    outputs(8321) <= not (a and b);
    outputs(8322) <= not a;
    outputs(8323) <= a;
    outputs(8324) <= a xor b;
    outputs(8325) <= not a;
    outputs(8326) <= a xor b;
    outputs(8327) <= a and not b;
    outputs(8328) <= b and not a;
    outputs(8329) <= not b;
    outputs(8330) <= not a;
    outputs(8331) <= a xor b;
    outputs(8332) <= not (a xor b);
    outputs(8333) <= not (a xor b);
    outputs(8334) <= a xor b;
    outputs(8335) <= not a;
    outputs(8336) <= not (a xor b);
    outputs(8337) <= not (a xor b);
    outputs(8338) <= a;
    outputs(8339) <= a;
    outputs(8340) <= not a;
    outputs(8341) <= not a;
    outputs(8342) <= a;
    outputs(8343) <= a and b;
    outputs(8344) <= not a;
    outputs(8345) <= b;
    outputs(8346) <= not (a xor b);
    outputs(8347) <= a and not b;
    outputs(8348) <= not (a xor b);
    outputs(8349) <= not (a xor b);
    outputs(8350) <= a or b;
    outputs(8351) <= a;
    outputs(8352) <= a;
    outputs(8353) <= b and not a;
    outputs(8354) <= b and not a;
    outputs(8355) <= a and b;
    outputs(8356) <= not a;
    outputs(8357) <= not a;
    outputs(8358) <= a xor b;
    outputs(8359) <= b;
    outputs(8360) <= not (a xor b);
    outputs(8361) <= not b;
    outputs(8362) <= a and b;
    outputs(8363) <= not b or a;
    outputs(8364) <= not (a xor b);
    outputs(8365) <= a xor b;
    outputs(8366) <= a and b;
    outputs(8367) <= a and not b;
    outputs(8368) <= not (a xor b);
    outputs(8369) <= not b;
    outputs(8370) <= not (a xor b);
    outputs(8371) <= not a;
    outputs(8372) <= a;
    outputs(8373) <= a;
    outputs(8374) <= not (a xor b);
    outputs(8375) <= a;
    outputs(8376) <= a;
    outputs(8377) <= not (a or b);
    outputs(8378) <= a xor b;
    outputs(8379) <= not a;
    outputs(8380) <= not (a or b);
    outputs(8381) <= not (a xor b);
    outputs(8382) <= not (a xor b);
    outputs(8383) <= not b or a;
    outputs(8384) <= not a or b;
    outputs(8385) <= b;
    outputs(8386) <= not a;
    outputs(8387) <= not a;
    outputs(8388) <= not b or a;
    outputs(8389) <= not a;
    outputs(8390) <= not b;
    outputs(8391) <= a xor b;
    outputs(8392) <= not b;
    outputs(8393) <= a xor b;
    outputs(8394) <= not b;
    outputs(8395) <= not (a xor b);
    outputs(8396) <= not a;
    outputs(8397) <= not b;
    outputs(8398) <= b;
    outputs(8399) <= not a;
    outputs(8400) <= a xor b;
    outputs(8401) <= b;
    outputs(8402) <= not b;
    outputs(8403) <= not b;
    outputs(8404) <= a xor b;
    outputs(8405) <= not (a xor b);
    outputs(8406) <= not a;
    outputs(8407) <= not b;
    outputs(8408) <= not b;
    outputs(8409) <= not (a or b);
    outputs(8410) <= not a;
    outputs(8411) <= not (a xor b);
    outputs(8412) <= a or b;
    outputs(8413) <= not b;
    outputs(8414) <= a and b;
    outputs(8415) <= a;
    outputs(8416) <= b;
    outputs(8417) <= not b;
    outputs(8418) <= not (a and b);
    outputs(8419) <= not a;
    outputs(8420) <= a;
    outputs(8421) <= a and b;
    outputs(8422) <= not (a xor b);
    outputs(8423) <= not (a and b);
    outputs(8424) <= not a;
    outputs(8425) <= a;
    outputs(8426) <= not (a xor b);
    outputs(8427) <= not b or a;
    outputs(8428) <= b;
    outputs(8429) <= not (a xor b);
    outputs(8430) <= not b or a;
    outputs(8431) <= not (a xor b);
    outputs(8432) <= not (a xor b);
    outputs(8433) <= a;
    outputs(8434) <= a xor b;
    outputs(8435) <= a;
    outputs(8436) <= not a;
    outputs(8437) <= a xor b;
    outputs(8438) <= a xor b;
    outputs(8439) <= a;
    outputs(8440) <= b;
    outputs(8441) <= not a;
    outputs(8442) <= a xor b;
    outputs(8443) <= not a;
    outputs(8444) <= not b;
    outputs(8445) <= not (a xor b);
    outputs(8446) <= not (a and b);
    outputs(8447) <= a xor b;
    outputs(8448) <= a and b;
    outputs(8449) <= not b;
    outputs(8450) <= a xor b;
    outputs(8451) <= a xor b;
    outputs(8452) <= not b or a;
    outputs(8453) <= a;
    outputs(8454) <= b;
    outputs(8455) <= b;
    outputs(8456) <= a;
    outputs(8457) <= b;
    outputs(8458) <= not b;
    outputs(8459) <= a xor b;
    outputs(8460) <= not (a xor b);
    outputs(8461) <= a xor b;
    outputs(8462) <= not a;
    outputs(8463) <= a xor b;
    outputs(8464) <= b;
    outputs(8465) <= not (a xor b);
    outputs(8466) <= a;
    outputs(8467) <= not a;
    outputs(8468) <= not a;
    outputs(8469) <= a xor b;
    outputs(8470) <= a xor b;
    outputs(8471) <= a xor b;
    outputs(8472) <= a and b;
    outputs(8473) <= a;
    outputs(8474) <= a;
    outputs(8475) <= not (a xor b);
    outputs(8476) <= not (a or b);
    outputs(8477) <= a and b;
    outputs(8478) <= not a or b;
    outputs(8479) <= not b or a;
    outputs(8480) <= a xor b;
    outputs(8481) <= a xor b;
    outputs(8482) <= not a;
    outputs(8483) <= a and not b;
    outputs(8484) <= not a;
    outputs(8485) <= a xor b;
    outputs(8486) <= not a;
    outputs(8487) <= not (a and b);
    outputs(8488) <= not a or b;
    outputs(8489) <= b;
    outputs(8490) <= a xor b;
    outputs(8491) <= not b;
    outputs(8492) <= not b;
    outputs(8493) <= a xor b;
    outputs(8494) <= a xor b;
    outputs(8495) <= a;
    outputs(8496) <= a xor b;
    outputs(8497) <= not (a xor b);
    outputs(8498) <= a and b;
    outputs(8499) <= not a;
    outputs(8500) <= not a;
    outputs(8501) <= not a;
    outputs(8502) <= a and not b;
    outputs(8503) <= a xor b;
    outputs(8504) <= a and b;
    outputs(8505) <= a or b;
    outputs(8506) <= a xor b;
    outputs(8507) <= a xor b;
    outputs(8508) <= not b;
    outputs(8509) <= not (a xor b);
    outputs(8510) <= a and b;
    outputs(8511) <= b and not a;
    outputs(8512) <= a and not b;
    outputs(8513) <= a and not b;
    outputs(8514) <= a;
    outputs(8515) <= not a;
    outputs(8516) <= b;
    outputs(8517) <= a and not b;
    outputs(8518) <= a;
    outputs(8519) <= not b or a;
    outputs(8520) <= a and not b;
    outputs(8521) <= a xor b;
    outputs(8522) <= b;
    outputs(8523) <= not b;
    outputs(8524) <= a xor b;
    outputs(8525) <= not a;
    outputs(8526) <= b;
    outputs(8527) <= not a;
    outputs(8528) <= b;
    outputs(8529) <= not b;
    outputs(8530) <= not a;
    outputs(8531) <= not b;
    outputs(8532) <= a xor b;
    outputs(8533) <= not a;
    outputs(8534) <= not b or a;
    outputs(8535) <= b;
    outputs(8536) <= b and not a;
    outputs(8537) <= a or b;
    outputs(8538) <= a;
    outputs(8539) <= not (a xor b);
    outputs(8540) <= a xor b;
    outputs(8541) <= a or b;
    outputs(8542) <= a;
    outputs(8543) <= b and not a;
    outputs(8544) <= not a or b;
    outputs(8545) <= a xor b;
    outputs(8546) <= not (a and b);
    outputs(8547) <= b and not a;
    outputs(8548) <= not b;
    outputs(8549) <= a or b;
    outputs(8550) <= not (a or b);
    outputs(8551) <= not (a xor b);
    outputs(8552) <= a;
    outputs(8553) <= a xor b;
    outputs(8554) <= a xor b;
    outputs(8555) <= a xor b;
    outputs(8556) <= not a;
    outputs(8557) <= a xor b;
    outputs(8558) <= not b or a;
    outputs(8559) <= a xor b;
    outputs(8560) <= a;
    outputs(8561) <= a;
    outputs(8562) <= a or b;
    outputs(8563) <= not (a xor b);
    outputs(8564) <= not (a xor b);
    outputs(8565) <= not b;
    outputs(8566) <= not b or a;
    outputs(8567) <= not b;
    outputs(8568) <= a and not b;
    outputs(8569) <= not b;
    outputs(8570) <= not a;
    outputs(8571) <= a xor b;
    outputs(8572) <= not (a xor b);
    outputs(8573) <= not b;
    outputs(8574) <= a xor b;
    outputs(8575) <= not (a xor b);
    outputs(8576) <= not a;
    outputs(8577) <= not b;
    outputs(8578) <= not a;
    outputs(8579) <= a or b;
    outputs(8580) <= a;
    outputs(8581) <= not b;
    outputs(8582) <= a xor b;
    outputs(8583) <= a;
    outputs(8584) <= a xor b;
    outputs(8585) <= a xor b;
    outputs(8586) <= a;
    outputs(8587) <= not (a and b);
    outputs(8588) <= b;
    outputs(8589) <= a xor b;
    outputs(8590) <= a;
    outputs(8591) <= not (a xor b);
    outputs(8592) <= b;
    outputs(8593) <= a xor b;
    outputs(8594) <= not a or b;
    outputs(8595) <= a xor b;
    outputs(8596) <= not a or b;
    outputs(8597) <= not a;
    outputs(8598) <= b;
    outputs(8599) <= a and not b;
    outputs(8600) <= a;
    outputs(8601) <= not (a xor b);
    outputs(8602) <= a and not b;
    outputs(8603) <= not b;
    outputs(8604) <= not (a xor b);
    outputs(8605) <= a xor b;
    outputs(8606) <= not a;
    outputs(8607) <= a;
    outputs(8608) <= not (a xor b);
    outputs(8609) <= not (a xor b);
    outputs(8610) <= b and not a;
    outputs(8611) <= not b;
    outputs(8612) <= not a;
    outputs(8613) <= not a;
    outputs(8614) <= a;
    outputs(8615) <= not (a xor b);
    outputs(8616) <= not (a xor b);
    outputs(8617) <= b;
    outputs(8618) <= a;
    outputs(8619) <= a;
    outputs(8620) <= b;
    outputs(8621) <= not a;
    outputs(8622) <= a xor b;
    outputs(8623) <= a;
    outputs(8624) <= not (a xor b);
    outputs(8625) <= a xor b;
    outputs(8626) <= a xor b;
    outputs(8627) <= b;
    outputs(8628) <= a xor b;
    outputs(8629) <= b and not a;
    outputs(8630) <= not b;
    outputs(8631) <= a;
    outputs(8632) <= a xor b;
    outputs(8633) <= a;
    outputs(8634) <= b;
    outputs(8635) <= b;
    outputs(8636) <= a;
    outputs(8637) <= not (a xor b);
    outputs(8638) <= a and b;
    outputs(8639) <= not b;
    outputs(8640) <= b;
    outputs(8641) <= a or b;
    outputs(8642) <= not (a xor b);
    outputs(8643) <= not b or a;
    outputs(8644) <= not b or a;
    outputs(8645) <= a;
    outputs(8646) <= not a;
    outputs(8647) <= not b;
    outputs(8648) <= not (a xor b);
    outputs(8649) <= not (a or b);
    outputs(8650) <= not (a and b);
    outputs(8651) <= not (a xor b);
    outputs(8652) <= a;
    outputs(8653) <= not (a xor b);
    outputs(8654) <= b;
    outputs(8655) <= not (a xor b);
    outputs(8656) <= not b;
    outputs(8657) <= b;
    outputs(8658) <= a xor b;
    outputs(8659) <= a;
    outputs(8660) <= a xor b;
    outputs(8661) <= not (a xor b);
    outputs(8662) <= a or b;
    outputs(8663) <= not (a or b);
    outputs(8664) <= b;
    outputs(8665) <= not a or b;
    outputs(8666) <= not b;
    outputs(8667) <= b;
    outputs(8668) <= a;
    outputs(8669) <= not (a xor b);
    outputs(8670) <= b;
    outputs(8671) <= not b or a;
    outputs(8672) <= not (a xor b);
    outputs(8673) <= not (a xor b);
    outputs(8674) <= not a;
    outputs(8675) <= a;
    outputs(8676) <= not a;
    outputs(8677) <= b;
    outputs(8678) <= b;
    outputs(8679) <= a;
    outputs(8680) <= not a;
    outputs(8681) <= a and b;
    outputs(8682) <= not (a xor b);
    outputs(8683) <= not a;
    outputs(8684) <= not a;
    outputs(8685) <= a;
    outputs(8686) <= not a;
    outputs(8687) <= b;
    outputs(8688) <= b;
    outputs(8689) <= a or b;
    outputs(8690) <= b;
    outputs(8691) <= a xor b;
    outputs(8692) <= a and b;
    outputs(8693) <= b;
    outputs(8694) <= not (a and b);
    outputs(8695) <= not b;
    outputs(8696) <= not (a or b);
    outputs(8697) <= not (a xor b);
    outputs(8698) <= not b or a;
    outputs(8699) <= not a;
    outputs(8700) <= not a or b;
    outputs(8701) <= not b;
    outputs(8702) <= a;
    outputs(8703) <= a;
    outputs(8704) <= not (a or b);
    outputs(8705) <= not b;
    outputs(8706) <= a;
    outputs(8707) <= b and not a;
    outputs(8708) <= not (a xor b);
    outputs(8709) <= not (a xor b);
    outputs(8710) <= not a;
    outputs(8711) <= not (a xor b);
    outputs(8712) <= a;
    outputs(8713) <= not a or b;
    outputs(8714) <= a or b;
    outputs(8715) <= not b;
    outputs(8716) <= not (a or b);
    outputs(8717) <= b;
    outputs(8718) <= a;
    outputs(8719) <= a;
    outputs(8720) <= b;
    outputs(8721) <= not (a xor b);
    outputs(8722) <= not b;
    outputs(8723) <= a;
    outputs(8724) <= b;
    outputs(8725) <= not a;
    outputs(8726) <= not a;
    outputs(8727) <= a;
    outputs(8728) <= not (a and b);
    outputs(8729) <= b;
    outputs(8730) <= not b;
    outputs(8731) <= not b;
    outputs(8732) <= a xor b;
    outputs(8733) <= b;
    outputs(8734) <= not (a xor b);
    outputs(8735) <= not (a xor b);
    outputs(8736) <= a or b;
    outputs(8737) <= not b;
    outputs(8738) <= not b;
    outputs(8739) <= a;
    outputs(8740) <= a xor b;
    outputs(8741) <= not b;
    outputs(8742) <= not a or b;
    outputs(8743) <= not (a xor b);
    outputs(8744) <= a;
    outputs(8745) <= not b or a;
    outputs(8746) <= not a;
    outputs(8747) <= not (a xor b);
    outputs(8748) <= not (a xor b);
    outputs(8749) <= b;
    outputs(8750) <= a xor b;
    outputs(8751) <= not (a or b);
    outputs(8752) <= not a;
    outputs(8753) <= not (a and b);
    outputs(8754) <= b;
    outputs(8755) <= not a or b;
    outputs(8756) <= a xor b;
    outputs(8757) <= a;
    outputs(8758) <= a xor b;
    outputs(8759) <= not a;
    outputs(8760) <= a or b;
    outputs(8761) <= a;
    outputs(8762) <= a;
    outputs(8763) <= b;
    outputs(8764) <= not b or a;
    outputs(8765) <= a xor b;
    outputs(8766) <= a xor b;
    outputs(8767) <= a;
    outputs(8768) <= not b or a;
    outputs(8769) <= not (a and b);
    outputs(8770) <= a;
    outputs(8771) <= a;
    outputs(8772) <= not a;
    outputs(8773) <= not (a xor b);
    outputs(8774) <= not a or b;
    outputs(8775) <= a or b;
    outputs(8776) <= a and b;
    outputs(8777) <= a xor b;
    outputs(8778) <= a and b;
    outputs(8779) <= a;
    outputs(8780) <= not (a xor b);
    outputs(8781) <= a and not b;
    outputs(8782) <= a xor b;
    outputs(8783) <= a xor b;
    outputs(8784) <= not b;
    outputs(8785) <= not (a and b);
    outputs(8786) <= b;
    outputs(8787) <= not b or a;
    outputs(8788) <= not b;
    outputs(8789) <= a xor b;
    outputs(8790) <= b;
    outputs(8791) <= not (a xor b);
    outputs(8792) <= b;
    outputs(8793) <= not a;
    outputs(8794) <= not (a xor b);
    outputs(8795) <= a;
    outputs(8796) <= not b;
    outputs(8797) <= b;
    outputs(8798) <= a;
    outputs(8799) <= not (a xor b);
    outputs(8800) <= a xor b;
    outputs(8801) <= not a;
    outputs(8802) <= b;
    outputs(8803) <= not (a xor b);
    outputs(8804) <= not b;
    outputs(8805) <= b and not a;
    outputs(8806) <= a and not b;
    outputs(8807) <= not (a xor b);
    outputs(8808) <= not b;
    outputs(8809) <= a;
    outputs(8810) <= a and b;
    outputs(8811) <= not (a and b);
    outputs(8812) <= a;
    outputs(8813) <= a xor b;
    outputs(8814) <= a;
    outputs(8815) <= not (a xor b);
    outputs(8816) <= a xor b;
    outputs(8817) <= not a;
    outputs(8818) <= a xor b;
    outputs(8819) <= not a;
    outputs(8820) <= a;
    outputs(8821) <= a xor b;
    outputs(8822) <= not (a xor b);
    outputs(8823) <= not (a or b);
    outputs(8824) <= a and b;
    outputs(8825) <= not (a xor b);
    outputs(8826) <= not b;
    outputs(8827) <= a xor b;
    outputs(8828) <= a xor b;
    outputs(8829) <= b;
    outputs(8830) <= a and not b;
    outputs(8831) <= a and b;
    outputs(8832) <= a xor b;
    outputs(8833) <= b;
    outputs(8834) <= not (a xor b);
    outputs(8835) <= not (a or b);
    outputs(8836) <= a xor b;
    outputs(8837) <= not b;
    outputs(8838) <= not (a and b);
    outputs(8839) <= a and b;
    outputs(8840) <= a xor b;
    outputs(8841) <= a xor b;
    outputs(8842) <= not a;
    outputs(8843) <= a and not b;
    outputs(8844) <= b;
    outputs(8845) <= not a;
    outputs(8846) <= not (a xor b);
    outputs(8847) <= a xor b;
    outputs(8848) <= a;
    outputs(8849) <= b;
    outputs(8850) <= not a;
    outputs(8851) <= not a;
    outputs(8852) <= not (a xor b);
    outputs(8853) <= not (a xor b);
    outputs(8854) <= a xor b;
    outputs(8855) <= a xor b;
    outputs(8856) <= not (a or b);
    outputs(8857) <= a;
    outputs(8858) <= not b or a;
    outputs(8859) <= not a or b;
    outputs(8860) <= not b or a;
    outputs(8861) <= a xor b;
    outputs(8862) <= not b;
    outputs(8863) <= a;
    outputs(8864) <= not b;
    outputs(8865) <= a xor b;
    outputs(8866) <= not (a xor b);
    outputs(8867) <= not (a xor b);
    outputs(8868) <= not a;
    outputs(8869) <= not (a xor b);
    outputs(8870) <= not (a xor b);
    outputs(8871) <= a xor b;
    outputs(8872) <= not (a xor b);
    outputs(8873) <= not (a or b);
    outputs(8874) <= not b;
    outputs(8875) <= a;
    outputs(8876) <= not a;
    outputs(8877) <= not a;
    outputs(8878) <= a;
    outputs(8879) <= not (a xor b);
    outputs(8880) <= not b;
    outputs(8881) <= a;
    outputs(8882) <= not b or a;
    outputs(8883) <= not a;
    outputs(8884) <= a xor b;
    outputs(8885) <= not (a xor b);
    outputs(8886) <= not a;
    outputs(8887) <= not (a xor b);
    outputs(8888) <= b;
    outputs(8889) <= not (a xor b);
    outputs(8890) <= b;
    outputs(8891) <= not (a xor b);
    outputs(8892) <= a;
    outputs(8893) <= not b or a;
    outputs(8894) <= a;
    outputs(8895) <= not a;
    outputs(8896) <= a;
    outputs(8897) <= b;
    outputs(8898) <= not (a xor b);
    outputs(8899) <= b;
    outputs(8900) <= b;
    outputs(8901) <= not (a xor b);
    outputs(8902) <= not b or a;
    outputs(8903) <= not (a xor b);
    outputs(8904) <= a xor b;
    outputs(8905) <= not b;
    outputs(8906) <= not a or b;
    outputs(8907) <= a xor b;
    outputs(8908) <= a and b;
    outputs(8909) <= not (a or b);
    outputs(8910) <= a xor b;
    outputs(8911) <= a xor b;
    outputs(8912) <= not (a xor b);
    outputs(8913) <= not (a xor b);
    outputs(8914) <= b;
    outputs(8915) <= a;
    outputs(8916) <= a;
    outputs(8917) <= a xor b;
    outputs(8918) <= not b or a;
    outputs(8919) <= not a;
    outputs(8920) <= a;
    outputs(8921) <= not (a xor b);
    outputs(8922) <= not (a xor b);
    outputs(8923) <= not a;
    outputs(8924) <= a xor b;
    outputs(8925) <= b and not a;
    outputs(8926) <= not b;
    outputs(8927) <= a;
    outputs(8928) <= not a;
    outputs(8929) <= not a;
    outputs(8930) <= not a or b;
    outputs(8931) <= not a;
    outputs(8932) <= a or b;
    outputs(8933) <= a xor b;
    outputs(8934) <= not (a and b);
    outputs(8935) <= b and not a;
    outputs(8936) <= a;
    outputs(8937) <= a xor b;
    outputs(8938) <= a xor b;
    outputs(8939) <= a xor b;
    outputs(8940) <= b;
    outputs(8941) <= not a;
    outputs(8942) <= a xor b;
    outputs(8943) <= not a;
    outputs(8944) <= not a;
    outputs(8945) <= a xor b;
    outputs(8946) <= not (a xor b);
    outputs(8947) <= not a;
    outputs(8948) <= not (a xor b);
    outputs(8949) <= not b;
    outputs(8950) <= not a or b;
    outputs(8951) <= not b or a;
    outputs(8952) <= not b;
    outputs(8953) <= not (a xor b);
    outputs(8954) <= not (a xor b);
    outputs(8955) <= b;
    outputs(8956) <= b;
    outputs(8957) <= a xor b;
    outputs(8958) <= not (a xor b);
    outputs(8959) <= a and not b;
    outputs(8960) <= not a or b;
    outputs(8961) <= a or b;
    outputs(8962) <= not a;
    outputs(8963) <= not (a xor b);
    outputs(8964) <= not a;
    outputs(8965) <= b;
    outputs(8966) <= not (a and b);
    outputs(8967) <= a and b;
    outputs(8968) <= not a;
    outputs(8969) <= a and b;
    outputs(8970) <= b;
    outputs(8971) <= a xor b;
    outputs(8972) <= not a;
    outputs(8973) <= not b;
    outputs(8974) <= not b;
    outputs(8975) <= b and not a;
    outputs(8976) <= a;
    outputs(8977) <= not b;
    outputs(8978) <= not a or b;
    outputs(8979) <= a;
    outputs(8980) <= not b;
    outputs(8981) <= not b;
    outputs(8982) <= not (a xor b);
    outputs(8983) <= a xor b;
    outputs(8984) <= not (a xor b);
    outputs(8985) <= a;
    outputs(8986) <= not b;
    outputs(8987) <= a;
    outputs(8988) <= a xor b;
    outputs(8989) <= a and b;
    outputs(8990) <= a;
    outputs(8991) <= a xor b;
    outputs(8992) <= not (a xor b);
    outputs(8993) <= not a or b;
    outputs(8994) <= a xor b;
    outputs(8995) <= a xor b;
    outputs(8996) <= b;
    outputs(8997) <= not a or b;
    outputs(8998) <= a xor b;
    outputs(8999) <= a xor b;
    outputs(9000) <= not a;
    outputs(9001) <= a xor b;
    outputs(9002) <= not a or b;
    outputs(9003) <= a and b;
    outputs(9004) <= not b;
    outputs(9005) <= b;
    outputs(9006) <= not (a and b);
    outputs(9007) <= not (a xor b);
    outputs(9008) <= not b;
    outputs(9009) <= not (a xor b);
    outputs(9010) <= b;
    outputs(9011) <= not a;
    outputs(9012) <= not (a xor b);
    outputs(9013) <= not b;
    outputs(9014) <= a and not b;
    outputs(9015) <= a;
    outputs(9016) <= not b;
    outputs(9017) <= not (a xor b);
    outputs(9018) <= not b;
    outputs(9019) <= a xor b;
    outputs(9020) <= not b or a;
    outputs(9021) <= b;
    outputs(9022) <= a xor b;
    outputs(9023) <= b;
    outputs(9024) <= not a;
    outputs(9025) <= not a;
    outputs(9026) <= not b;
    outputs(9027) <= not (a or b);
    outputs(9028) <= a and not b;
    outputs(9029) <= a xor b;
    outputs(9030) <= a xor b;
    outputs(9031) <= not (a xor b);
    outputs(9032) <= not a;
    outputs(9033) <= a xor b;
    outputs(9034) <= a or b;
    outputs(9035) <= a or b;
    outputs(9036) <= a and not b;
    outputs(9037) <= b;
    outputs(9038) <= not (a xor b);
    outputs(9039) <= b;
    outputs(9040) <= not b;
    outputs(9041) <= not (a xor b);
    outputs(9042) <= a and not b;
    outputs(9043) <= a xor b;
    outputs(9044) <= a and b;
    outputs(9045) <= not b or a;
    outputs(9046) <= not b or a;
    outputs(9047) <= not (a xor b);
    outputs(9048) <= not (a xor b);
    outputs(9049) <= not (a xor b);
    outputs(9050) <= not b;
    outputs(9051) <= not a;
    outputs(9052) <= a and b;
    outputs(9053) <= not (a xor b);
    outputs(9054) <= not (a xor b);
    outputs(9055) <= not a;
    outputs(9056) <= a xor b;
    outputs(9057) <= a xor b;
    outputs(9058) <= not (a xor b);
    outputs(9059) <= b;
    outputs(9060) <= not b;
    outputs(9061) <= not b;
    outputs(9062) <= a and b;
    outputs(9063) <= not (a xor b);
    outputs(9064) <= a;
    outputs(9065) <= b;
    outputs(9066) <= not b or a;
    outputs(9067) <= a;
    outputs(9068) <= not a;
    outputs(9069) <= b;
    outputs(9070) <= not (a xor b);
    outputs(9071) <= b;
    outputs(9072) <= not b;
    outputs(9073) <= b;
    outputs(9074) <= a and b;
    outputs(9075) <= a;
    outputs(9076) <= not a;
    outputs(9077) <= b;
    outputs(9078) <= a xor b;
    outputs(9079) <= not (a and b);
    outputs(9080) <= a;
    outputs(9081) <= not (a or b);
    outputs(9082) <= not b;
    outputs(9083) <= not a or b;
    outputs(9084) <= b;
    outputs(9085) <= not (a or b);
    outputs(9086) <= not (a and b);
    outputs(9087) <= a xor b;
    outputs(9088) <= not a;
    outputs(9089) <= not (a xor b);
    outputs(9090) <= a;
    outputs(9091) <= not (a xor b);
    outputs(9092) <= not (a and b);
    outputs(9093) <= b and not a;
    outputs(9094) <= a;
    outputs(9095) <= not a;
    outputs(9096) <= not b;
    outputs(9097) <= a xor b;
    outputs(9098) <= not (a xor b);
    outputs(9099) <= not b;
    outputs(9100) <= not (a or b);
    outputs(9101) <= a xor b;
    outputs(9102) <= not (a xor b);
    outputs(9103) <= a;
    outputs(9104) <= not (a xor b);
    outputs(9105) <= not (a and b);
    outputs(9106) <= a and not b;
    outputs(9107) <= b;
    outputs(9108) <= a xor b;
    outputs(9109) <= not b;
    outputs(9110) <= not b or a;
    outputs(9111) <= not b or a;
    outputs(9112) <= b;
    outputs(9113) <= not a or b;
    outputs(9114) <= a and not b;
    outputs(9115) <= not (a xor b);
    outputs(9116) <= a;
    outputs(9117) <= not (a xor b);
    outputs(9118) <= not (a and b);
    outputs(9119) <= a;
    outputs(9120) <= b;
    outputs(9121) <= not (a xor b);
    outputs(9122) <= not (a xor b);
    outputs(9123) <= not b;
    outputs(9124) <= not b;
    outputs(9125) <= not (a xor b);
    outputs(9126) <= b and not a;
    outputs(9127) <= not (a xor b);
    outputs(9128) <= a;
    outputs(9129) <= a xor b;
    outputs(9130) <= a;
    outputs(9131) <= a;
    outputs(9132) <= a xor b;
    outputs(9133) <= a;
    outputs(9134) <= not b;
    outputs(9135) <= not a or b;
    outputs(9136) <= a xor b;
    outputs(9137) <= a;
    outputs(9138) <= a or b;
    outputs(9139) <= not a;
    outputs(9140) <= not a;
    outputs(9141) <= not a;
    outputs(9142) <= not (a xor b);
    outputs(9143) <= a or b;
    outputs(9144) <= not a or b;
    outputs(9145) <= a;
    outputs(9146) <= a or b;
    outputs(9147) <= not a or b;
    outputs(9148) <= b;
    outputs(9149) <= a xor b;
    outputs(9150) <= not a or b;
    outputs(9151) <= a or b;
    outputs(9152) <= b;
    outputs(9153) <= not b;
    outputs(9154) <= a and b;
    outputs(9155) <= not (a xor b);
    outputs(9156) <= not (a or b);
    outputs(9157) <= not a;
    outputs(9158) <= not a;
    outputs(9159) <= a xor b;
    outputs(9160) <= not b;
    outputs(9161) <= not (a xor b);
    outputs(9162) <= not b;
    outputs(9163) <= a xor b;
    outputs(9164) <= a or b;
    outputs(9165) <= a;
    outputs(9166) <= b;
    outputs(9167) <= a xor b;
    outputs(9168) <= not (a xor b);
    outputs(9169) <= not (a xor b);
    outputs(9170) <= a xor b;
    outputs(9171) <= not (a xor b);
    outputs(9172) <= not b;
    outputs(9173) <= not (a xor b);
    outputs(9174) <= not a or b;
    outputs(9175) <= a;
    outputs(9176) <= a;
    outputs(9177) <= not (a xor b);
    outputs(9178) <= not b;
    outputs(9179) <= a;
    outputs(9180) <= a;
    outputs(9181) <= not a or b;
    outputs(9182) <= a;
    outputs(9183) <= b;
    outputs(9184) <= b and not a;
    outputs(9185) <= a xor b;
    outputs(9186) <= a xor b;
    outputs(9187) <= a xor b;
    outputs(9188) <= b;
    outputs(9189) <= b and not a;
    outputs(9190) <= a xor b;
    outputs(9191) <= not (a and b);
    outputs(9192) <= not (a and b);
    outputs(9193) <= a xor b;
    outputs(9194) <= not (a or b);
    outputs(9195) <= not a;
    outputs(9196) <= a and b;
    outputs(9197) <= b;
    outputs(9198) <= not (a and b);
    outputs(9199) <= not a;
    outputs(9200) <= a;
    outputs(9201) <= not a;
    outputs(9202) <= not a or b;
    outputs(9203) <= b;
    outputs(9204) <= a xor b;
    outputs(9205) <= not (a xor b);
    outputs(9206) <= a and b;
    outputs(9207) <= b;
    outputs(9208) <= a xor b;
    outputs(9209) <= not b or a;
    outputs(9210) <= not b;
    outputs(9211) <= not (a xor b);
    outputs(9212) <= not a or b;
    outputs(9213) <= not (a xor b);
    outputs(9214) <= not (a xor b);
    outputs(9215) <= not (a and b);
    outputs(9216) <= not b or a;
    outputs(9217) <= a;
    outputs(9218) <= a;
    outputs(9219) <= not (a and b);
    outputs(9220) <= not b;
    outputs(9221) <= not b;
    outputs(9222) <= b;
    outputs(9223) <= b and not a;
    outputs(9224) <= b;
    outputs(9225) <= b;
    outputs(9226) <= not (a xor b);
    outputs(9227) <= a and b;
    outputs(9228) <= b;
    outputs(9229) <= not (a xor b);
    outputs(9230) <= not a;
    outputs(9231) <= not b;
    outputs(9232) <= not (a xor b);
    outputs(9233) <= not (a xor b);
    outputs(9234) <= not b;
    outputs(9235) <= a xor b;
    outputs(9236) <= not b or a;
    outputs(9237) <= not a;
    outputs(9238) <= not (a xor b);
    outputs(9239) <= not b;
    outputs(9240) <= not (a xor b);
    outputs(9241) <= not b;
    outputs(9242) <= b;
    outputs(9243) <= not a;
    outputs(9244) <= b;
    outputs(9245) <= not (a and b);
    outputs(9246) <= a;
    outputs(9247) <= a xor b;
    outputs(9248) <= not a;
    outputs(9249) <= not (a xor b);
    outputs(9250) <= not (a xor b);
    outputs(9251) <= not (a xor b);
    outputs(9252) <= not b;
    outputs(9253) <= not a;
    outputs(9254) <= not b;
    outputs(9255) <= a xor b;
    outputs(9256) <= not a;
    outputs(9257) <= a;
    outputs(9258) <= not (a xor b);
    outputs(9259) <= a;
    outputs(9260) <= not (a xor b);
    outputs(9261) <= not a;
    outputs(9262) <= a and b;
    outputs(9263) <= not (a xor b);
    outputs(9264) <= not b;
    outputs(9265) <= not (a xor b);
    outputs(9266) <= not b or a;
    outputs(9267) <= not (a xor b);
    outputs(9268) <= a;
    outputs(9269) <= not (a xor b);
    outputs(9270) <= a xor b;
    outputs(9271) <= b;
    outputs(9272) <= a xor b;
    outputs(9273) <= a;
    outputs(9274) <= b;
    outputs(9275) <= a xor b;
    outputs(9276) <= not (a or b);
    outputs(9277) <= a and not b;
    outputs(9278) <= a xor b;
    outputs(9279) <= not b;
    outputs(9280) <= a xor b;
    outputs(9281) <= not (a or b);
    outputs(9282) <= not a;
    outputs(9283) <= a;
    outputs(9284) <= a and b;
    outputs(9285) <= not (a xor b);
    outputs(9286) <= not b;
    outputs(9287) <= not (a xor b);
    outputs(9288) <= a and b;
    outputs(9289) <= not (a xor b);
    outputs(9290) <= not a;
    outputs(9291) <= a xor b;
    outputs(9292) <= not (a xor b);
    outputs(9293) <= not b or a;
    outputs(9294) <= not b;
    outputs(9295) <= b;
    outputs(9296) <= not a or b;
    outputs(9297) <= not a;
    outputs(9298) <= not (a or b);
    outputs(9299) <= a;
    outputs(9300) <= not (a xor b);
    outputs(9301) <= a xor b;
    outputs(9302) <= not b;
    outputs(9303) <= not a or b;
    outputs(9304) <= b and not a;
    outputs(9305) <= a;
    outputs(9306) <= a and b;
    outputs(9307) <= not (a and b);
    outputs(9308) <= a xor b;
    outputs(9309) <= a xor b;
    outputs(9310) <= a and not b;
    outputs(9311) <= a;
    outputs(9312) <= b;
    outputs(9313) <= not b;
    outputs(9314) <= b;
    outputs(9315) <= not (a xor b);
    outputs(9316) <= a and b;
    outputs(9317) <= not a;
    outputs(9318) <= a xor b;
    outputs(9319) <= a xor b;
    outputs(9320) <= not b;
    outputs(9321) <= b and not a;
    outputs(9322) <= a xor b;
    outputs(9323) <= not a;
    outputs(9324) <= not (a xor b);
    outputs(9325) <= not (a and b);
    outputs(9326) <= a;
    outputs(9327) <= not (a xor b);
    outputs(9328) <= not b;
    outputs(9329) <= not b;
    outputs(9330) <= b and not a;
    outputs(9331) <= not a;
    outputs(9332) <= a or b;
    outputs(9333) <= b;
    outputs(9334) <= a xor b;
    outputs(9335) <= b;
    outputs(9336) <= b;
    outputs(9337) <= not a or b;
    outputs(9338) <= not b;
    outputs(9339) <= a and not b;
    outputs(9340) <= a and b;
    outputs(9341) <= b;
    outputs(9342) <= not b or a;
    outputs(9343) <= b;
    outputs(9344) <= not b;
    outputs(9345) <= b;
    outputs(9346) <= a and b;
    outputs(9347) <= not b;
    outputs(9348) <= a and b;
    outputs(9349) <= a and not b;
    outputs(9350) <= a;
    outputs(9351) <= not b;
    outputs(9352) <= a and not b;
    outputs(9353) <= a and not b;
    outputs(9354) <= a xor b;
    outputs(9355) <= a;
    outputs(9356) <= not b;
    outputs(9357) <= not (a xor b);
    outputs(9358) <= a;
    outputs(9359) <= not a;
    outputs(9360) <= a xor b;
    outputs(9361) <= a xor b;
    outputs(9362) <= a and b;
    outputs(9363) <= b and not a;
    outputs(9364) <= not (a or b);
    outputs(9365) <= not (a xor b);
    outputs(9366) <= a and not b;
    outputs(9367) <= a xor b;
    outputs(9368) <= a xor b;
    outputs(9369) <= not b;
    outputs(9370) <= a xor b;
    outputs(9371) <= not (a or b);
    outputs(9372) <= not (a xor b);
    outputs(9373) <= a and not b;
    outputs(9374) <= not (a and b);
    outputs(9375) <= not b;
    outputs(9376) <= b;
    outputs(9377) <= not (a xor b);
    outputs(9378) <= not a;
    outputs(9379) <= not b;
    outputs(9380) <= not (a xor b);
    outputs(9381) <= not b;
    outputs(9382) <= a and b;
    outputs(9383) <= not b or a;
    outputs(9384) <= not a;
    outputs(9385) <= not (a xor b);
    outputs(9386) <= not (a xor b);
    outputs(9387) <= a xor b;
    outputs(9388) <= not (a and b);
    outputs(9389) <= not a;
    outputs(9390) <= b;
    outputs(9391) <= not b or a;
    outputs(9392) <= not (a xor b);
    outputs(9393) <= a xor b;
    outputs(9394) <= a;
    outputs(9395) <= not b;
    outputs(9396) <= b;
    outputs(9397) <= a;
    outputs(9398) <= a and b;
    outputs(9399) <= not a;
    outputs(9400) <= b;
    outputs(9401) <= a xor b;
    outputs(9402) <= not a;
    outputs(9403) <= a and not b;
    outputs(9404) <= b;
    outputs(9405) <= b and not a;
    outputs(9406) <= b;
    outputs(9407) <= a xor b;
    outputs(9408) <= b;
    outputs(9409) <= not (a or b);
    outputs(9410) <= not a;
    outputs(9411) <= not (a xor b);
    outputs(9412) <= a;
    outputs(9413) <= a and not b;
    outputs(9414) <= not a;
    outputs(9415) <= b;
    outputs(9416) <= not (a xor b);
    outputs(9417) <= not (a xor b);
    outputs(9418) <= not (a xor b);
    outputs(9419) <= not a;
    outputs(9420) <= b;
    outputs(9421) <= not a;
    outputs(9422) <= a xor b;
    outputs(9423) <= b and not a;
    outputs(9424) <= not (a xor b);
    outputs(9425) <= not (a xor b);
    outputs(9426) <= a;
    outputs(9427) <= not (a xor b);
    outputs(9428) <= not (a or b);
    outputs(9429) <= b;
    outputs(9430) <= not (a and b);
    outputs(9431) <= not a or b;
    outputs(9432) <= not a;
    outputs(9433) <= a and b;
    outputs(9434) <= a xor b;
    outputs(9435) <= a;
    outputs(9436) <= not b;
    outputs(9437) <= a;
    outputs(9438) <= a and not b;
    outputs(9439) <= a;
    outputs(9440) <= b;
    outputs(9441) <= not b or a;
    outputs(9442) <= a xor b;
    outputs(9443) <= a xor b;
    outputs(9444) <= not (a xor b);
    outputs(9445) <= a;
    outputs(9446) <= not (a xor b);
    outputs(9447) <= not (a xor b);
    outputs(9448) <= not b;
    outputs(9449) <= not b or a;
    outputs(9450) <= a;
    outputs(9451) <= a;
    outputs(9452) <= not b;
    outputs(9453) <= a xor b;
    outputs(9454) <= a xor b;
    outputs(9455) <= not a or b;
    outputs(9456) <= a xor b;
    outputs(9457) <= a;
    outputs(9458) <= a;
    outputs(9459) <= b;
    outputs(9460) <= not (a and b);
    outputs(9461) <= not b;
    outputs(9462) <= not (a and b);
    outputs(9463) <= b and not a;
    outputs(9464) <= a xor b;
    outputs(9465) <= not a;
    outputs(9466) <= a;
    outputs(9467) <= b;
    outputs(9468) <= not b;
    outputs(9469) <= a xor b;
    outputs(9470) <= not b;
    outputs(9471) <= not b;
    outputs(9472) <= a xor b;
    outputs(9473) <= a or b;
    outputs(9474) <= not b;
    outputs(9475) <= b;
    outputs(9476) <= not (a xor b);
    outputs(9477) <= a;
    outputs(9478) <= not (a and b);
    outputs(9479) <= a;
    outputs(9480) <= not b;
    outputs(9481) <= b;
    outputs(9482) <= b;
    outputs(9483) <= b and not a;
    outputs(9484) <= a and not b;
    outputs(9485) <= not a;
    outputs(9486) <= not a;
    outputs(9487) <= not b;
    outputs(9488) <= not b;
    outputs(9489) <= b;
    outputs(9490) <= a and not b;
    outputs(9491) <= not (a or b);
    outputs(9492) <= not (a xor b);
    outputs(9493) <= b and not a;
    outputs(9494) <= not b;
    outputs(9495) <= not (a xor b);
    outputs(9496) <= not a;
    outputs(9497) <= a xor b;
    outputs(9498) <= not b;
    outputs(9499) <= a and not b;
    outputs(9500) <= not (a xor b);
    outputs(9501) <= a;
    outputs(9502) <= not (a xor b);
    outputs(9503) <= not a;
    outputs(9504) <= a;
    outputs(9505) <= b and not a;
    outputs(9506) <= not (a xor b);
    outputs(9507) <= a and not b;
    outputs(9508) <= not (a xor b);
    outputs(9509) <= a;
    outputs(9510) <= not (a or b);
    outputs(9511) <= b;
    outputs(9512) <= a and b;
    outputs(9513) <= not a;
    outputs(9514) <= not a or b;
    outputs(9515) <= not b;
    outputs(9516) <= not (a xor b);
    outputs(9517) <= a and not b;
    outputs(9518) <= not a;
    outputs(9519) <= not (a and b);
    outputs(9520) <= b;
    outputs(9521) <= not (a or b);
    outputs(9522) <= b;
    outputs(9523) <= a xor b;
    outputs(9524) <= b and not a;
    outputs(9525) <= a;
    outputs(9526) <= b;
    outputs(9527) <= not a;
    outputs(9528) <= not b;
    outputs(9529) <= a xor b;
    outputs(9530) <= a xor b;
    outputs(9531) <= b and not a;
    outputs(9532) <= a xor b;
    outputs(9533) <= a xor b;
    outputs(9534) <= b and not a;
    outputs(9535) <= a and b;
    outputs(9536) <= not (a or b);
    outputs(9537) <= a and not b;
    outputs(9538) <= not b;
    outputs(9539) <= not b;
    outputs(9540) <= a xor b;
    outputs(9541) <= a;
    outputs(9542) <= a and b;
    outputs(9543) <= not (a xor b);
    outputs(9544) <= a;
    outputs(9545) <= not (a xor b);
    outputs(9546) <= a xor b;
    outputs(9547) <= not (a xor b);
    outputs(9548) <= not (a or b);
    outputs(9549) <= a and not b;
    outputs(9550) <= a or b;
    outputs(9551) <= b and not a;
    outputs(9552) <= a or b;
    outputs(9553) <= not a or b;
    outputs(9554) <= a or b;
    outputs(9555) <= not b;
    outputs(9556) <= not (a xor b);
    outputs(9557) <= a;
    outputs(9558) <= a;
    outputs(9559) <= not a;
    outputs(9560) <= b;
    outputs(9561) <= b and not a;
    outputs(9562) <= not a;
    outputs(9563) <= a xor b;
    outputs(9564) <= not a;
    outputs(9565) <= not b;
    outputs(9566) <= b;
    outputs(9567) <= b and not a;
    outputs(9568) <= a and b;
    outputs(9569) <= not (a xor b);
    outputs(9570) <= not (a or b);
    outputs(9571) <= not b;
    outputs(9572) <= not b;
    outputs(9573) <= b and not a;
    outputs(9574) <= not a;
    outputs(9575) <= not a;
    outputs(9576) <= not (a or b);
    outputs(9577) <= not a;
    outputs(9578) <= not (a or b);
    outputs(9579) <= not (a or b);
    outputs(9580) <= not b;
    outputs(9581) <= not a or b;
    outputs(9582) <= a xor b;
    outputs(9583) <= not a;
    outputs(9584) <= a xor b;
    outputs(9585) <= a and not b;
    outputs(9586) <= not (a xor b);
    outputs(9587) <= not (a xor b);
    outputs(9588) <= not (a xor b);
    outputs(9589) <= not (a and b);
    outputs(9590) <= a and b;
    outputs(9591) <= b and not a;
    outputs(9592) <= b;
    outputs(9593) <= b and not a;
    outputs(9594) <= a and not b;
    outputs(9595) <= not (a xor b);
    outputs(9596) <= not (a or b);
    outputs(9597) <= a xor b;
    outputs(9598) <= not (a xor b);
    outputs(9599) <= not (a or b);
    outputs(9600) <= a and not b;
    outputs(9601) <= not (a xor b);
    outputs(9602) <= a;
    outputs(9603) <= b;
    outputs(9604) <= not b;
    outputs(9605) <= a;
    outputs(9606) <= not (a xor b);
    outputs(9607) <= not b;
    outputs(9608) <= a or b;
    outputs(9609) <= a xor b;
    outputs(9610) <= not b;
    outputs(9611) <= b;
    outputs(9612) <= not a;
    outputs(9613) <= not (a xor b);
    outputs(9614) <= not (a xor b);
    outputs(9615) <= a and b;
    outputs(9616) <= not b;
    outputs(9617) <= b;
    outputs(9618) <= not (a and b);
    outputs(9619) <= not a;
    outputs(9620) <= a or b;
    outputs(9621) <= not (a and b);
    outputs(9622) <= not a or b;
    outputs(9623) <= a xor b;
    outputs(9624) <= a and b;
    outputs(9625) <= not (a xor b);
    outputs(9626) <= b and not a;
    outputs(9627) <= b;
    outputs(9628) <= not b;
    outputs(9629) <= b and not a;
    outputs(9630) <= a and b;
    outputs(9631) <= a;
    outputs(9632) <= not (a xor b);
    outputs(9633) <= not (a xor b);
    outputs(9634) <= not (a or b);
    outputs(9635) <= a;
    outputs(9636) <= not (a xor b);
    outputs(9637) <= not a;
    outputs(9638) <= not b;
    outputs(9639) <= a or b;
    outputs(9640) <= a;
    outputs(9641) <= b;
    outputs(9642) <= not b;
    outputs(9643) <= a xor b;
    outputs(9644) <= not (a xor b);
    outputs(9645) <= a and b;
    outputs(9646) <= not a;
    outputs(9647) <= not b;
    outputs(9648) <= not (a xor b);
    outputs(9649) <= not b;
    outputs(9650) <= a;
    outputs(9651) <= not a;
    outputs(9652) <= not (a xor b);
    outputs(9653) <= b;
    outputs(9654) <= a and not b;
    outputs(9655) <= b;
    outputs(9656) <= a or b;
    outputs(9657) <= b and not a;
    outputs(9658) <= not a or b;
    outputs(9659) <= not a;
    outputs(9660) <= not (a and b);
    outputs(9661) <= a xor b;
    outputs(9662) <= a xor b;
    outputs(9663) <= not (a xor b);
    outputs(9664) <= b and not a;
    outputs(9665) <= not a;
    outputs(9666) <= not (a or b);
    outputs(9667) <= not a;
    outputs(9668) <= not b;
    outputs(9669) <= b;
    outputs(9670) <= not b or a;
    outputs(9671) <= a;
    outputs(9672) <= a xor b;
    outputs(9673) <= a or b;
    outputs(9674) <= not b;
    outputs(9675) <= not b;
    outputs(9676) <= a xor b;
    outputs(9677) <= a and b;
    outputs(9678) <= not a;
    outputs(9679) <= b and not a;
    outputs(9680) <= not a;
    outputs(9681) <= a xor b;
    outputs(9682) <= a;
    outputs(9683) <= not b or a;
    outputs(9684) <= b and not a;
    outputs(9685) <= b;
    outputs(9686) <= b;
    outputs(9687) <= not (a xor b);
    outputs(9688) <= not (a xor b);
    outputs(9689) <= not (a xor b);
    outputs(9690) <= not (a and b);
    outputs(9691) <= b and not a;
    outputs(9692) <= not (a or b);
    outputs(9693) <= a;
    outputs(9694) <= b and not a;
    outputs(9695) <= not (a xor b);
    outputs(9696) <= not a or b;
    outputs(9697) <= b;
    outputs(9698) <= not a;
    outputs(9699) <= a and not b;
    outputs(9700) <= not a;
    outputs(9701) <= a and not b;
    outputs(9702) <= a;
    outputs(9703) <= a and b;
    outputs(9704) <= b;
    outputs(9705) <= not (a or b);
    outputs(9706) <= a or b;
    outputs(9707) <= not (a or b);
    outputs(9708) <= a xor b;
    outputs(9709) <= not b or a;
    outputs(9710) <= not (a xor b);
    outputs(9711) <= a;
    outputs(9712) <= b;
    outputs(9713) <= b;
    outputs(9714) <= b and not a;
    outputs(9715) <= not (a xor b);
    outputs(9716) <= not (a or b);
    outputs(9717) <= a xor b;
    outputs(9718) <= a or b;
    outputs(9719) <= not (a xor b);
    outputs(9720) <= not a;
    outputs(9721) <= b;
    outputs(9722) <= not b;
    outputs(9723) <= b;
    outputs(9724) <= a and not b;
    outputs(9725) <= not (a xor b);
    outputs(9726) <= not a;
    outputs(9727) <= a;
    outputs(9728) <= b;
    outputs(9729) <= not b;
    outputs(9730) <= a xor b;
    outputs(9731) <= not a;
    outputs(9732) <= not b;
    outputs(9733) <= b;
    outputs(9734) <= a;
    outputs(9735) <= not (a xor b);
    outputs(9736) <= not b or a;
    outputs(9737) <= a;
    outputs(9738) <= a xor b;
    outputs(9739) <= not b or a;
    outputs(9740) <= b and not a;
    outputs(9741) <= a xor b;
    outputs(9742) <= not b;
    outputs(9743) <= a;
    outputs(9744) <= not (a xor b);
    outputs(9745) <= a;
    outputs(9746) <= a;
    outputs(9747) <= b;
    outputs(9748) <= not (a or b);
    outputs(9749) <= not b;
    outputs(9750) <= not (a xor b);
    outputs(9751) <= a or b;
    outputs(9752) <= not a;
    outputs(9753) <= a xor b;
    outputs(9754) <= a;
    outputs(9755) <= not (a xor b);
    outputs(9756) <= a xor b;
    outputs(9757) <= a or b;
    outputs(9758) <= not a;
    outputs(9759) <= not a;
    outputs(9760) <= a xor b;
    outputs(9761) <= b;
    outputs(9762) <= not (a xor b);
    outputs(9763) <= not b or a;
    outputs(9764) <= a and b;
    outputs(9765) <= b;
    outputs(9766) <= a;
    outputs(9767) <= b;
    outputs(9768) <= a xor b;
    outputs(9769) <= a or b;
    outputs(9770) <= b and not a;
    outputs(9771) <= not (a or b);
    outputs(9772) <= not b;
    outputs(9773) <= a xor b;
    outputs(9774) <= not a;
    outputs(9775) <= not a;
    outputs(9776) <= not a;
    outputs(9777) <= a or b;
    outputs(9778) <= not (a and b);
    outputs(9779) <= a;
    outputs(9780) <= b;
    outputs(9781) <= a and b;
    outputs(9782) <= not a;
    outputs(9783) <= a xor b;
    outputs(9784) <= not b;
    outputs(9785) <= not b;
    outputs(9786) <= a xor b;
    outputs(9787) <= not (a or b);
    outputs(9788) <= not b or a;
    outputs(9789) <= not (a or b);
    outputs(9790) <= a xor b;
    outputs(9791) <= a xor b;
    outputs(9792) <= not b;
    outputs(9793) <= not (a xor b);
    outputs(9794) <= b;
    outputs(9795) <= a;
    outputs(9796) <= a;
    outputs(9797) <= not a;
    outputs(9798) <= a xor b;
    outputs(9799) <= not a;
    outputs(9800) <= not b;
    outputs(9801) <= not a;
    outputs(9802) <= not b;
    outputs(9803) <= a xor b;
    outputs(9804) <= a;
    outputs(9805) <= b and not a;
    outputs(9806) <= a xor b;
    outputs(9807) <= b and not a;
    outputs(9808) <= a;
    outputs(9809) <= not b;
    outputs(9810) <= not b;
    outputs(9811) <= not a;
    outputs(9812) <= b;
    outputs(9813) <= a;
    outputs(9814) <= not a;
    outputs(9815) <= b;
    outputs(9816) <= a xor b;
    outputs(9817) <= b;
    outputs(9818) <= a;
    outputs(9819) <= not a;
    outputs(9820) <= b;
    outputs(9821) <= a;
    outputs(9822) <= b;
    outputs(9823) <= a xor b;
    outputs(9824) <= not (a and b);
    outputs(9825) <= b;
    outputs(9826) <= not a;
    outputs(9827) <= not b;
    outputs(9828) <= a and not b;
    outputs(9829) <= a xor b;
    outputs(9830) <= a xor b;
    outputs(9831) <= b;
    outputs(9832) <= a xor b;
    outputs(9833) <= not b or a;
    outputs(9834) <= b;
    outputs(9835) <= not (a xor b);
    outputs(9836) <= not a;
    outputs(9837) <= not (a xor b);
    outputs(9838) <= a xor b;
    outputs(9839) <= b and not a;
    outputs(9840) <= a xor b;
    outputs(9841) <= not a or b;
    outputs(9842) <= not a;
    outputs(9843) <= a;
    outputs(9844) <= not a;
    outputs(9845) <= not b;
    outputs(9846) <= not b;
    outputs(9847) <= not b;
    outputs(9848) <= not a;
    outputs(9849) <= not a;
    outputs(9850) <= a and b;
    outputs(9851) <= a xor b;
    outputs(9852) <= a xor b;
    outputs(9853) <= a and b;
    outputs(9854) <= b and not a;
    outputs(9855) <= a;
    outputs(9856) <= a xor b;
    outputs(9857) <= not (a xor b);
    outputs(9858) <= b and not a;
    outputs(9859) <= a;
    outputs(9860) <= not a;
    outputs(9861) <= not a;
    outputs(9862) <= a and b;
    outputs(9863) <= not (a xor b);
    outputs(9864) <= a xor b;
    outputs(9865) <= a and b;
    outputs(9866) <= a and not b;
    outputs(9867) <= b;
    outputs(9868) <= a and b;
    outputs(9869) <= a;
    outputs(9870) <= b and not a;
    outputs(9871) <= not b;
    outputs(9872) <= a;
    outputs(9873) <= a and not b;
    outputs(9874) <= a xor b;
    outputs(9875) <= b;
    outputs(9876) <= not (a xor b);
    outputs(9877) <= not b;
    outputs(9878) <= a;
    outputs(9879) <= a and not b;
    outputs(9880) <= a or b;
    outputs(9881) <= a;
    outputs(9882) <= a;
    outputs(9883) <= not (a and b);
    outputs(9884) <= a xor b;
    outputs(9885) <= not b;
    outputs(9886) <= a and not b;
    outputs(9887) <= not b;
    outputs(9888) <= a xor b;
    outputs(9889) <= a xor b;
    outputs(9890) <= b;
    outputs(9891) <= not a;
    outputs(9892) <= not b or a;
    outputs(9893) <= not (a xor b);
    outputs(9894) <= a;
    outputs(9895) <= not a;
    outputs(9896) <= a and not b;
    outputs(9897) <= not (a or b);
    outputs(9898) <= a;
    outputs(9899) <= not a;
    outputs(9900) <= not a;
    outputs(9901) <= a and b;
    outputs(9902) <= not (a xor b);
    outputs(9903) <= not (a xor b);
    outputs(9904) <= a;
    outputs(9905) <= not b;
    outputs(9906) <= b;
    outputs(9907) <= a;
    outputs(9908) <= b;
    outputs(9909) <= a and b;
    outputs(9910) <= a and not b;
    outputs(9911) <= not b;
    outputs(9912) <= not (a or b);
    outputs(9913) <= a;
    outputs(9914) <= a;
    outputs(9915) <= a and b;
    outputs(9916) <= a xor b;
    outputs(9917) <= not (a and b);
    outputs(9918) <= not b;
    outputs(9919) <= b;
    outputs(9920) <= b;
    outputs(9921) <= b and not a;
    outputs(9922) <= a and b;
    outputs(9923) <= not a;
    outputs(9924) <= not (a xor b);
    outputs(9925) <= a xor b;
    outputs(9926) <= not b;
    outputs(9927) <= a;
    outputs(9928) <= a xor b;
    outputs(9929) <= b;
    outputs(9930) <= not (a or b);
    outputs(9931) <= b;
    outputs(9932) <= a and not b;
    outputs(9933) <= a xor b;
    outputs(9934) <= a xor b;
    outputs(9935) <= not a;
    outputs(9936) <= not a;
    outputs(9937) <= not a;
    outputs(9938) <= not (a xor b);
    outputs(9939) <= b and not a;
    outputs(9940) <= not b;
    outputs(9941) <= b;
    outputs(9942) <= a xor b;
    outputs(9943) <= not (a or b);
    outputs(9944) <= a xor b;
    outputs(9945) <= not b;
    outputs(9946) <= a;
    outputs(9947) <= not b;
    outputs(9948) <= a xor b;
    outputs(9949) <= b;
    outputs(9950) <= a;
    outputs(9951) <= not b;
    outputs(9952) <= a;
    outputs(9953) <= not (a and b);
    outputs(9954) <= b;
    outputs(9955) <= a or b;
    outputs(9956) <= not (a xor b);
    outputs(9957) <= not b;
    outputs(9958) <= a xor b;
    outputs(9959) <= a and not b;
    outputs(9960) <= a;
    outputs(9961) <= b and not a;
    outputs(9962) <= not (a or b);
    outputs(9963) <= a xor b;
    outputs(9964) <= a and not b;
    outputs(9965) <= a;
    outputs(9966) <= a xor b;
    outputs(9967) <= a or b;
    outputs(9968) <= a;
    outputs(9969) <= not b;
    outputs(9970) <= b;
    outputs(9971) <= b and not a;
    outputs(9972) <= not b;
    outputs(9973) <= not (a xor b);
    outputs(9974) <= not (a xor b);
    outputs(9975) <= a xor b;
    outputs(9976) <= a or b;
    outputs(9977) <= b;
    outputs(9978) <= b;
    outputs(9979) <= not b;
    outputs(9980) <= a and b;
    outputs(9981) <= a and b;
    outputs(9982) <= b;
    outputs(9983) <= not (a xor b);
    outputs(9984) <= b;
    outputs(9985) <= a and b;
    outputs(9986) <= not (a or b);
    outputs(9987) <= a xor b;
    outputs(9988) <= a and b;
    outputs(9989) <= b;
    outputs(9990) <= a;
    outputs(9991) <= a;
    outputs(9992) <= not a;
    outputs(9993) <= not (a xor b);
    outputs(9994) <= not a;
    outputs(9995) <= not a;
    outputs(9996) <= a and not b;
    outputs(9997) <= not b;
    outputs(9998) <= a xor b;
    outputs(9999) <= a xor b;
    outputs(10000) <= a and b;
    outputs(10001) <= b and not a;
    outputs(10002) <= a xor b;
    outputs(10003) <= not a;
    outputs(10004) <= a and b;
    outputs(10005) <= not b;
    outputs(10006) <= not b;
    outputs(10007) <= not a;
    outputs(10008) <= a and not b;
    outputs(10009) <= a xor b;
    outputs(10010) <= b;
    outputs(10011) <= not b;
    outputs(10012) <= not (a xor b);
    outputs(10013) <= b;
    outputs(10014) <= a;
    outputs(10015) <= a xor b;
    outputs(10016) <= not a;
    outputs(10017) <= b;
    outputs(10018) <= not (a xor b);
    outputs(10019) <= b;
    outputs(10020) <= not b;
    outputs(10021) <= a xor b;
    outputs(10022) <= not (a xor b);
    outputs(10023) <= a;
    outputs(10024) <= a;
    outputs(10025) <= not (a xor b);
    outputs(10026) <= not b;
    outputs(10027) <= a xor b;
    outputs(10028) <= a xor b;
    outputs(10029) <= a xor b;
    outputs(10030) <= a xor b;
    outputs(10031) <= not (a xor b);
    outputs(10032) <= not b;
    outputs(10033) <= a xor b;
    outputs(10034) <= not (a and b);
    outputs(10035) <= b;
    outputs(10036) <= not a;
    outputs(10037) <= b and not a;
    outputs(10038) <= not (a and b);
    outputs(10039) <= a and not b;
    outputs(10040) <= not a;
    outputs(10041) <= a and b;
    outputs(10042) <= a and b;
    outputs(10043) <= a;
    outputs(10044) <= a;
    outputs(10045) <= b;
    outputs(10046) <= a xor b;
    outputs(10047) <= a xor b;
    outputs(10048) <= a or b;
    outputs(10049) <= not a;
    outputs(10050) <= not a or b;
    outputs(10051) <= a or b;
    outputs(10052) <= not (a xor b);
    outputs(10053) <= not (a xor b);
    outputs(10054) <= a xor b;
    outputs(10055) <= b;
    outputs(10056) <= b;
    outputs(10057) <= not (a or b);
    outputs(10058) <= not a;
    outputs(10059) <= not a;
    outputs(10060) <= not (a or b);
    outputs(10061) <= not (a xor b);
    outputs(10062) <= a and not b;
    outputs(10063) <= b;
    outputs(10064) <= not a;
    outputs(10065) <= a or b;
    outputs(10066) <= not (a and b);
    outputs(10067) <= a xor b;
    outputs(10068) <= b;
    outputs(10069) <= a;
    outputs(10070) <= a xor b;
    outputs(10071) <= a;
    outputs(10072) <= not (a xor b);
    outputs(10073) <= not (a xor b);
    outputs(10074) <= not (a xor b);
    outputs(10075) <= b;
    outputs(10076) <= not b;
    outputs(10077) <= not (a or b);
    outputs(10078) <= a;
    outputs(10079) <= a and b;
    outputs(10080) <= not (a or b);
    outputs(10081) <= a;
    outputs(10082) <= not b;
    outputs(10083) <= not (a or b);
    outputs(10084) <= a and b;
    outputs(10085) <= not a;
    outputs(10086) <= a and b;
    outputs(10087) <= a xor b;
    outputs(10088) <= not (a xor b);
    outputs(10089) <= not (a xor b);
    outputs(10090) <= a;
    outputs(10091) <= b and not a;
    outputs(10092) <= a xor b;
    outputs(10093) <= b;
    outputs(10094) <= not (a xor b);
    outputs(10095) <= a;
    outputs(10096) <= not (a or b);
    outputs(10097) <= a xor b;
    outputs(10098) <= not (a xor b);
    outputs(10099) <= not b;
    outputs(10100) <= a and not b;
    outputs(10101) <= not b;
    outputs(10102) <= not (a xor b);
    outputs(10103) <= a xor b;
    outputs(10104) <= not (a or b);
    outputs(10105) <= a;
    outputs(10106) <= b;
    outputs(10107) <= not b;
    outputs(10108) <= not a;
    outputs(10109) <= not b;
    outputs(10110) <= not a;
    outputs(10111) <= a or b;
    outputs(10112) <= a and b;
    outputs(10113) <= not (a xor b);
    outputs(10114) <= not b;
    outputs(10115) <= b;
    outputs(10116) <= not a;
    outputs(10117) <= a xor b;
    outputs(10118) <= b;
    outputs(10119) <= a or b;
    outputs(10120) <= not b;
    outputs(10121) <= b;
    outputs(10122) <= b;
    outputs(10123) <= a and b;
    outputs(10124) <= a;
    outputs(10125) <= a xor b;
    outputs(10126) <= a and b;
    outputs(10127) <= not a or b;
    outputs(10128) <= b;
    outputs(10129) <= b;
    outputs(10130) <= b;
    outputs(10131) <= b and not a;
    outputs(10132) <= not (a or b);
    outputs(10133) <= not b;
    outputs(10134) <= b and not a;
    outputs(10135) <= a xor b;
    outputs(10136) <= not (a xor b);
    outputs(10137) <= b;
    outputs(10138) <= a and b;
    outputs(10139) <= not b or a;
    outputs(10140) <= a xor b;
    outputs(10141) <= a or b;
    outputs(10142) <= not (a xor b);
    outputs(10143) <= not a;
    outputs(10144) <= not a;
    outputs(10145) <= not b;
    outputs(10146) <= not b or a;
    outputs(10147) <= a;
    outputs(10148) <= a xor b;
    outputs(10149) <= b;
    outputs(10150) <= b;
    outputs(10151) <= a and b;
    outputs(10152) <= not b or a;
    outputs(10153) <= not a;
    outputs(10154) <= not (a xor b);
    outputs(10155) <= a xor b;
    outputs(10156) <= a xor b;
    outputs(10157) <= not a;
    outputs(10158) <= a xor b;
    outputs(10159) <= not b;
    outputs(10160) <= a xor b;
    outputs(10161) <= a xor b;
    outputs(10162) <= not (a xor b);
    outputs(10163) <= a xor b;
    outputs(10164) <= a;
    outputs(10165) <= a xor b;
    outputs(10166) <= a and not b;
    outputs(10167) <= not (a xor b);
    outputs(10168) <= b;
    outputs(10169) <= a;
    outputs(10170) <= not b;
    outputs(10171) <= not a;
    outputs(10172) <= a xor b;
    outputs(10173) <= a xor b;
    outputs(10174) <= not b;
    outputs(10175) <= not (a xor b);
    outputs(10176) <= a xor b;
    outputs(10177) <= not (a xor b);
    outputs(10178) <= not b;
    outputs(10179) <= not (a xor b);
    outputs(10180) <= a xor b;
    outputs(10181) <= a xor b;
    outputs(10182) <= b;
    outputs(10183) <= not a;
    outputs(10184) <= not (a xor b);
    outputs(10185) <= not (a xor b);
    outputs(10186) <= a or b;
    outputs(10187) <= b;
    outputs(10188) <= a;
    outputs(10189) <= a and b;
    outputs(10190) <= a xor b;
    outputs(10191) <= not (a or b);
    outputs(10192) <= not (a or b);
    outputs(10193) <= not (a xor b);
    outputs(10194) <= b;
    outputs(10195) <= not a;
    outputs(10196) <= b;
    outputs(10197) <= not b;
    outputs(10198) <= not (a xor b);
    outputs(10199) <= not b;
    outputs(10200) <= not b;
    outputs(10201) <= not (a xor b);
    outputs(10202) <= a and not b;
    outputs(10203) <= a xor b;
    outputs(10204) <= a and b;
    outputs(10205) <= a xor b;
    outputs(10206) <= b;
    outputs(10207) <= not (a or b);
    outputs(10208) <= b and not a;
    outputs(10209) <= not a;
    outputs(10210) <= not (a or b);
    outputs(10211) <= a;
    outputs(10212) <= not (a xor b);
    outputs(10213) <= a xor b;
    outputs(10214) <= a;
    outputs(10215) <= not b or a;
    outputs(10216) <= a xor b;
    outputs(10217) <= not b;
    outputs(10218) <= b;
    outputs(10219) <= not b;
    outputs(10220) <= a;
    outputs(10221) <= a xor b;
    outputs(10222) <= a and b;
    outputs(10223) <= not (a xor b);
    outputs(10224) <= not a or b;
    outputs(10225) <= not a;
    outputs(10226) <= not (a and b);
    outputs(10227) <= not b or a;
    outputs(10228) <= a;
    outputs(10229) <= b;
    outputs(10230) <= a or b;
    outputs(10231) <= b;
    outputs(10232) <= not a;
    outputs(10233) <= not (a or b);
    outputs(10234) <= b;
    outputs(10235) <= a xor b;
    outputs(10236) <= a and not b;
    outputs(10237) <= not (a xor b);
    outputs(10238) <= a or b;
    outputs(10239) <= not b;
end Behavioral;
