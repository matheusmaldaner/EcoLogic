module logic_network(
    input wire [1023:0] inputs,
    output wire [9:0] outputs
);

    wire [10239:0] layer0_outputs;

    assign layer0_outputs[0] = ~((inputs[307]) & (inputs[967]));
    assign layer0_outputs[1] = ~((inputs[310]) ^ (inputs[718]));
    assign layer0_outputs[2] = (inputs[217]) & ~(inputs[830]);
    assign layer0_outputs[3] = (inputs[354]) & ~(inputs[904]);
    assign layer0_outputs[4] = ~((inputs[812]) ^ (inputs[875]));
    assign layer0_outputs[5] = ~((inputs[735]) ^ (inputs[126]));
    assign layer0_outputs[6] = inputs[274];
    assign layer0_outputs[7] = ~((inputs[310]) ^ (inputs[544]));
    assign layer0_outputs[8] = (inputs[163]) & ~(inputs[999]);
    assign layer0_outputs[9] = (inputs[487]) & ~(inputs[898]);
    assign layer0_outputs[10] = inputs[500];
    assign layer0_outputs[11] = ~(inputs[851]) | (inputs[62]);
    assign layer0_outputs[12] = (inputs[479]) & ~(inputs[757]);
    assign layer0_outputs[13] = ~(inputs[501]) | (inputs[89]);
    assign layer0_outputs[14] = ~((inputs[826]) & (inputs[1006]));
    assign layer0_outputs[15] = (inputs[590]) | (inputs[916]);
    assign layer0_outputs[16] = ~(inputs[611]);
    assign layer0_outputs[17] = (inputs[674]) ^ (inputs[998]);
    assign layer0_outputs[18] = inputs[265];
    assign layer0_outputs[19] = inputs[558];
    assign layer0_outputs[20] = ~((inputs[337]) ^ (inputs[859]));
    assign layer0_outputs[21] = ~((inputs[222]) | (inputs[362]));
    assign layer0_outputs[22] = (inputs[919]) | (inputs[584]);
    assign layer0_outputs[23] = ~(inputs[814]);
    assign layer0_outputs[24] = ~(inputs[726]) | (inputs[71]);
    assign layer0_outputs[25] = (inputs[858]) & ~(inputs[34]);
    assign layer0_outputs[26] = (inputs[778]) & ~(inputs[162]);
    assign layer0_outputs[27] = ~(inputs[147]) | (inputs[17]);
    assign layer0_outputs[28] = (inputs[968]) | (inputs[567]);
    assign layer0_outputs[29] = (inputs[48]) | (inputs[712]);
    assign layer0_outputs[30] = ~((inputs[265]) | (inputs[31]));
    assign layer0_outputs[31] = ~((inputs[265]) ^ (inputs[158]));
    assign layer0_outputs[32] = (inputs[287]) ^ (inputs[653]);
    assign layer0_outputs[33] = ~(inputs[145]) | (inputs[798]);
    assign layer0_outputs[34] = (inputs[878]) & ~(inputs[491]);
    assign layer0_outputs[35] = ~(inputs[62]);
    assign layer0_outputs[36] = ~((inputs[522]) | (inputs[948]));
    assign layer0_outputs[37] = inputs[1012];
    assign layer0_outputs[38] = (inputs[558]) & (inputs[190]);
    assign layer0_outputs[39] = inputs[306];
    assign layer0_outputs[40] = ~((inputs[180]) | (inputs[1013]));
    assign layer0_outputs[41] = (inputs[197]) & (inputs[968]);
    assign layer0_outputs[42] = ~((inputs[286]) | (inputs[623]));
    assign layer0_outputs[43] = inputs[471];
    assign layer0_outputs[44] = inputs[900];
    assign layer0_outputs[45] = ~(inputs[491]);
    assign layer0_outputs[46] = ~((inputs[300]) ^ (inputs[629]));
    assign layer0_outputs[47] = ~(inputs[903]);
    assign layer0_outputs[48] = ~(inputs[186]);
    assign layer0_outputs[49] = ~((inputs[797]) ^ (inputs[773]));
    assign layer0_outputs[50] = inputs[108];
    assign layer0_outputs[51] = (inputs[615]) | (inputs[342]);
    assign layer0_outputs[52] = inputs[264];
    assign layer0_outputs[53] = (inputs[78]) & ~(inputs[181]);
    assign layer0_outputs[54] = ~((inputs[343]) ^ (inputs[631]));
    assign layer0_outputs[55] = ~((inputs[611]) | (inputs[752]));
    assign layer0_outputs[56] = inputs[190];
    assign layer0_outputs[57] = (inputs[320]) ^ (inputs[91]);
    assign layer0_outputs[58] = (inputs[835]) | (inputs[435]);
    assign layer0_outputs[59] = (inputs[1011]) ^ (inputs[20]);
    assign layer0_outputs[60] = ~(inputs[975]);
    assign layer0_outputs[61] = ~((inputs[248]) | (inputs[425]));
    assign layer0_outputs[62] = (inputs[1017]) & ~(inputs[961]);
    assign layer0_outputs[63] = ~((inputs[364]) ^ (inputs[755]));
    assign layer0_outputs[64] = ~(inputs[895]);
    assign layer0_outputs[65] = (inputs[38]) ^ (inputs[93]);
    assign layer0_outputs[66] = (inputs[306]) & ~(inputs[940]);
    assign layer0_outputs[67] = ~(inputs[346]);
    assign layer0_outputs[68] = (inputs[471]) & ~(inputs[898]);
    assign layer0_outputs[69] = ~((inputs[685]) | (inputs[261]));
    assign layer0_outputs[70] = (inputs[914]) ^ (inputs[818]);
    assign layer0_outputs[71] = ~(inputs[598]);
    assign layer0_outputs[72] = (inputs[343]) & ~(inputs[578]);
    assign layer0_outputs[73] = ~(inputs[672]);
    assign layer0_outputs[74] = ~((inputs[248]) | (inputs[208]));
    assign layer0_outputs[75] = inputs[601];
    assign layer0_outputs[76] = (inputs[377]) & ~(inputs[194]);
    assign layer0_outputs[77] = inputs[578];
    assign layer0_outputs[78] = inputs[525];
    assign layer0_outputs[79] = ~(inputs[750]) | (inputs[614]);
    assign layer0_outputs[80] = inputs[910];
    assign layer0_outputs[81] = ~(inputs[34]) | (inputs[131]);
    assign layer0_outputs[82] = ~((inputs[230]) & (inputs[225]));
    assign layer0_outputs[83] = inputs[581];
    assign layer0_outputs[84] = ~((inputs[664]) ^ (inputs[790]));
    assign layer0_outputs[85] = ~(inputs[344]);
    assign layer0_outputs[86] = ~(inputs[498]) | (inputs[75]);
    assign layer0_outputs[87] = ~((inputs[465]) | (inputs[875]));
    assign layer0_outputs[88] = ~(inputs[406]) | (inputs[901]);
    assign layer0_outputs[89] = ~((inputs[361]) | (inputs[331]));
    assign layer0_outputs[90] = ~((inputs[351]) | (inputs[574]));
    assign layer0_outputs[91] = ~((inputs[992]) ^ (inputs[785]));
    assign layer0_outputs[92] = ~((inputs[722]) | (inputs[84]));
    assign layer0_outputs[93] = ~((inputs[1013]) | (inputs[185]));
    assign layer0_outputs[94] = (inputs[293]) | (inputs[154]);
    assign layer0_outputs[95] = inputs[618];
    assign layer0_outputs[96] = ~((inputs[260]) | (inputs[248]));
    assign layer0_outputs[97] = ~(inputs[462]);
    assign layer0_outputs[98] = (inputs[491]) ^ (inputs[266]);
    assign layer0_outputs[99] = (inputs[398]) | (inputs[879]);
    assign layer0_outputs[100] = ~(inputs[935]) | (inputs[131]);
    assign layer0_outputs[101] = ~((inputs[212]) & (inputs[310]));
    assign layer0_outputs[102] = (inputs[725]) & ~(inputs[387]);
    assign layer0_outputs[103] = ~(inputs[562]);
    assign layer0_outputs[104] = ~((inputs[165]) | (inputs[497]));
    assign layer0_outputs[105] = ~((inputs[865]) | (inputs[344]));
    assign layer0_outputs[106] = ~((inputs[834]) | (inputs[703]));
    assign layer0_outputs[107] = ~((inputs[961]) | (inputs[31]));
    assign layer0_outputs[108] = (inputs[102]) | (inputs[211]);
    assign layer0_outputs[109] = (inputs[291]) | (inputs[884]);
    assign layer0_outputs[110] = inputs[659];
    assign layer0_outputs[111] = ~((inputs[285]) ^ (inputs[455]));
    assign layer0_outputs[112] = (inputs[610]) | (inputs[672]);
    assign layer0_outputs[113] = inputs[270];
    assign layer0_outputs[114] = ~((inputs[935]) | (inputs[331]));
    assign layer0_outputs[115] = (inputs[413]) ^ (inputs[843]);
    assign layer0_outputs[116] = (inputs[798]) & ~(inputs[9]);
    assign layer0_outputs[117] = (inputs[725]) ^ (inputs[291]);
    assign layer0_outputs[118] = ~((inputs[374]) | (inputs[107]));
    assign layer0_outputs[119] = inputs[43];
    assign layer0_outputs[120] = ~((inputs[689]) | (inputs[538]));
    assign layer0_outputs[121] = (inputs[548]) | (inputs[363]);
    assign layer0_outputs[122] = ~((inputs[143]) ^ (inputs[154]));
    assign layer0_outputs[123] = (inputs[316]) | (inputs[986]);
    assign layer0_outputs[124] = ~((inputs[836]) ^ (inputs[810]));
    assign layer0_outputs[125] = inputs[160];
    assign layer0_outputs[126] = (inputs[768]) & ~(inputs[827]);
    assign layer0_outputs[127] = ~((inputs[427]) ^ (inputs[606]));
    assign layer0_outputs[128] = ~((inputs[898]) | (inputs[1001]));
    assign layer0_outputs[129] = inputs[391];
    assign layer0_outputs[130] = ~(inputs[492]);
    assign layer0_outputs[131] = (inputs[391]) & ~(inputs[572]);
    assign layer0_outputs[132] = inputs[871];
    assign layer0_outputs[133] = inputs[423];
    assign layer0_outputs[134] = ~(inputs[537]);
    assign layer0_outputs[135] = ~(inputs[653]);
    assign layer0_outputs[136] = ~(inputs[65]) | (inputs[69]);
    assign layer0_outputs[137] = ~(inputs[115]) | (inputs[898]);
    assign layer0_outputs[138] = ~((inputs[8]) & (inputs[893]));
    assign layer0_outputs[139] = inputs[493];
    assign layer0_outputs[140] = (inputs[684]) | (inputs[986]);
    assign layer0_outputs[141] = ~((inputs[888]) ^ (inputs[788]));
    assign layer0_outputs[142] = ~((inputs[520]) ^ (inputs[2]));
    assign layer0_outputs[143] = ~((inputs[823]) | (inputs[1018]));
    assign layer0_outputs[144] = (inputs[253]) ^ (inputs[1021]);
    assign layer0_outputs[145] = (inputs[841]) & ~(inputs[997]);
    assign layer0_outputs[146] = inputs[624];
    assign layer0_outputs[147] = ~(inputs[727]) | (inputs[422]);
    assign layer0_outputs[148] = (inputs[807]) & ~(inputs[141]);
    assign layer0_outputs[149] = ~(inputs[173]) | (inputs[411]);
    assign layer0_outputs[150] = (inputs[508]) ^ (inputs[115]);
    assign layer0_outputs[151] = (inputs[928]) | (inputs[132]);
    assign layer0_outputs[152] = ~((inputs[175]) ^ (inputs[91]));
    assign layer0_outputs[153] = inputs[372];
    assign layer0_outputs[154] = inputs[912];
    assign layer0_outputs[155] = inputs[1017];
    assign layer0_outputs[156] = ~(inputs[803]);
    assign layer0_outputs[157] = ~((inputs[376]) | (inputs[590]));
    assign layer0_outputs[158] = ~(inputs[612]);
    assign layer0_outputs[159] = (inputs[718]) | (inputs[96]);
    assign layer0_outputs[160] = (inputs[0]) & ~(inputs[1021]);
    assign layer0_outputs[161] = ~(inputs[184]);
    assign layer0_outputs[162] = (inputs[959]) & ~(inputs[886]);
    assign layer0_outputs[163] = inputs[228];
    assign layer0_outputs[164] = (inputs[587]) | (inputs[43]);
    assign layer0_outputs[165] = inputs[222];
    assign layer0_outputs[166] = ~(inputs[341]);
    assign layer0_outputs[167] = (inputs[224]) & (inputs[909]);
    assign layer0_outputs[168] = ~(inputs[471]);
    assign layer0_outputs[169] = (inputs[395]) | (inputs[203]);
    assign layer0_outputs[170] = (inputs[727]) | (inputs[572]);
    assign layer0_outputs[171] = (inputs[890]) | (inputs[284]);
    assign layer0_outputs[172] = (inputs[116]) | (inputs[436]);
    assign layer0_outputs[173] = ~((inputs[778]) | (inputs[259]));
    assign layer0_outputs[174] = ~((inputs[757]) ^ (inputs[329]));
    assign layer0_outputs[175] = inputs[209];
    assign layer0_outputs[176] = inputs[298];
    assign layer0_outputs[177] = ~((inputs[374]) | (inputs[130]));
    assign layer0_outputs[178] = ~((inputs[747]) ^ (inputs[224]));
    assign layer0_outputs[179] = ~((inputs[883]) ^ (inputs[967]));
    assign layer0_outputs[180] = ~(inputs[715]);
    assign layer0_outputs[181] = (inputs[546]) | (inputs[706]);
    assign layer0_outputs[182] = ~(inputs[313]) | (inputs[958]);
    assign layer0_outputs[183] = ~(inputs[722]);
    assign layer0_outputs[184] = (inputs[688]) | (inputs[989]);
    assign layer0_outputs[185] = ~(inputs[782]);
    assign layer0_outputs[186] = inputs[760];
    assign layer0_outputs[187] = ~(inputs[934]);
    assign layer0_outputs[188] = ~((inputs[579]) | (inputs[0]));
    assign layer0_outputs[189] = ~((inputs[1019]) | (inputs[795]));
    assign layer0_outputs[190] = (inputs[743]) & ~(inputs[985]);
    assign layer0_outputs[191] = (inputs[311]) & ~(inputs[554]);
    assign layer0_outputs[192] = (inputs[115]) ^ (inputs[267]);
    assign layer0_outputs[193] = ~(inputs[368]) | (inputs[802]);
    assign layer0_outputs[194] = (inputs[877]) ^ (inputs[1020]);
    assign layer0_outputs[195] = (inputs[595]) | (inputs[332]);
    assign layer0_outputs[196] = ~((inputs[706]) & (inputs[674]));
    assign layer0_outputs[197] = ~(inputs[47]) | (inputs[641]);
    assign layer0_outputs[198] = (inputs[1023]) & (inputs[96]);
    assign layer0_outputs[199] = ~((inputs[215]) | (inputs[806]));
    assign layer0_outputs[200] = ~(inputs[18]) | (inputs[155]);
    assign layer0_outputs[201] = (inputs[877]) & ~(inputs[891]);
    assign layer0_outputs[202] = (inputs[394]) | (inputs[392]);
    assign layer0_outputs[203] = ~(inputs[234]);
    assign layer0_outputs[204] = (inputs[250]) | (inputs[119]);
    assign layer0_outputs[205] = ~(inputs[768]);
    assign layer0_outputs[206] = (inputs[36]) & (inputs[486]);
    assign layer0_outputs[207] = (inputs[238]) | (inputs[258]);
    assign layer0_outputs[208] = ~(inputs[112]);
    assign layer0_outputs[209] = ~(inputs[853]) | (inputs[671]);
    assign layer0_outputs[210] = ~(inputs[843]);
    assign layer0_outputs[211] = (inputs[466]) & ~(inputs[442]);
    assign layer0_outputs[212] = (inputs[367]) ^ (inputs[835]);
    assign layer0_outputs[213] = (inputs[677]) ^ (inputs[296]);
    assign layer0_outputs[214] = (inputs[252]) ^ (inputs[889]);
    assign layer0_outputs[215] = ~((inputs[586]) | (inputs[425]));
    assign layer0_outputs[216] = ~((inputs[793]) & (inputs[123]));
    assign layer0_outputs[217] = (inputs[592]) ^ (inputs[957]);
    assign layer0_outputs[218] = (inputs[919]) ^ (inputs[136]);
    assign layer0_outputs[219] = inputs[852];
    assign layer0_outputs[220] = (inputs[560]) ^ (inputs[291]);
    assign layer0_outputs[221] = inputs[506];
    assign layer0_outputs[222] = (inputs[527]) | (inputs[23]);
    assign layer0_outputs[223] = (inputs[343]) & ~(inputs[97]);
    assign layer0_outputs[224] = ~((inputs[657]) | (inputs[363]));
    assign layer0_outputs[225] = (inputs[404]) & ~(inputs[283]);
    assign layer0_outputs[226] = ~(inputs[839]);
    assign layer0_outputs[227] = ~(inputs[807]);
    assign layer0_outputs[228] = inputs[408];
    assign layer0_outputs[229] = ~(inputs[140]);
    assign layer0_outputs[230] = (inputs[254]) & (inputs[414]);
    assign layer0_outputs[231] = inputs[795];
    assign layer0_outputs[232] = ~(inputs[885]);
    assign layer0_outputs[233] = inputs[558];
    assign layer0_outputs[234] = ~((inputs[283]) & (inputs[376]));
    assign layer0_outputs[235] = inputs[594];
    assign layer0_outputs[236] = (inputs[921]) & ~(inputs[153]);
    assign layer0_outputs[237] = (inputs[995]) & (inputs[670]);
    assign layer0_outputs[238] = (inputs[183]) | (inputs[486]);
    assign layer0_outputs[239] = inputs[243];
    assign layer0_outputs[240] = ~((inputs[804]) | (inputs[851]));
    assign layer0_outputs[241] = (inputs[949]) & ~(inputs[869]);
    assign layer0_outputs[242] = ~(inputs[423]);
    assign layer0_outputs[243] = (inputs[666]) | (inputs[235]);
    assign layer0_outputs[244] = ~((inputs[464]) ^ (inputs[997]));
    assign layer0_outputs[245] = inputs[565];
    assign layer0_outputs[246] = inputs[720];
    assign layer0_outputs[247] = ~((inputs[142]) | (inputs[730]));
    assign layer0_outputs[248] = ~((inputs[510]) | (inputs[219]));
    assign layer0_outputs[249] = ~(inputs[464]) | (inputs[508]);
    assign layer0_outputs[250] = (inputs[904]) & ~(inputs[987]);
    assign layer0_outputs[251] = (inputs[500]) | (inputs[30]);
    assign layer0_outputs[252] = ~((inputs[77]) & (inputs[322]));
    assign layer0_outputs[253] = inputs[430];
    assign layer0_outputs[254] = (inputs[165]) | (inputs[537]);
    assign layer0_outputs[255] = inputs[300];
    assign layer0_outputs[256] = inputs[216];
    assign layer0_outputs[257] = ~(inputs[426]) | (inputs[667]);
    assign layer0_outputs[258] = inputs[252];
    assign layer0_outputs[259] = ~((inputs[584]) | (inputs[793]));
    assign layer0_outputs[260] = ~((inputs[852]) | (inputs[836]));
    assign layer0_outputs[261] = ~(inputs[65]) | (inputs[542]);
    assign layer0_outputs[262] = ~(inputs[749]);
    assign layer0_outputs[263] = ~(inputs[304]);
    assign layer0_outputs[264] = ~(inputs[128]) | (inputs[454]);
    assign layer0_outputs[265] = ~((inputs[960]) | (inputs[8]));
    assign layer0_outputs[266] = (inputs[386]) & (inputs[833]);
    assign layer0_outputs[267] = inputs[569];
    assign layer0_outputs[268] = (inputs[8]) | (inputs[530]);
    assign layer0_outputs[269] = 1'b1;
    assign layer0_outputs[270] = ~(inputs[140]);
    assign layer0_outputs[271] = ~((inputs[138]) | (inputs[509]));
    assign layer0_outputs[272] = ~(inputs[549]) | (inputs[966]);
    assign layer0_outputs[273] = ~((inputs[157]) ^ (inputs[173]));
    assign layer0_outputs[274] = ~((inputs[313]) ^ (inputs[75]));
    assign layer0_outputs[275] = (inputs[774]) | (inputs[462]);
    assign layer0_outputs[276] = ~(inputs[969]) | (inputs[314]);
    assign layer0_outputs[277] = (inputs[902]) | (inputs[278]);
    assign layer0_outputs[278] = (inputs[660]) & ~(inputs[741]);
    assign layer0_outputs[279] = (inputs[842]) & ~(inputs[24]);
    assign layer0_outputs[280] = (inputs[666]) | (inputs[364]);
    assign layer0_outputs[281] = ~(inputs[12]);
    assign layer0_outputs[282] = (inputs[114]) ^ (inputs[790]);
    assign layer0_outputs[283] = ~((inputs[833]) ^ (inputs[1]));
    assign layer0_outputs[284] = ~((inputs[571]) & (inputs[782]));
    assign layer0_outputs[285] = ~((inputs[318]) ^ (inputs[908]));
    assign layer0_outputs[286] = ~(inputs[558]);
    assign layer0_outputs[287] = ~((inputs[765]) ^ (inputs[260]));
    assign layer0_outputs[288] = (inputs[795]) | (inputs[512]);
    assign layer0_outputs[289] = (inputs[709]) | (inputs[733]);
    assign layer0_outputs[290] = (inputs[324]) ^ (inputs[531]);
    assign layer0_outputs[291] = inputs[82];
    assign layer0_outputs[292] = ~((inputs[887]) | (inputs[275]));
    assign layer0_outputs[293] = (inputs[101]) ^ (inputs[934]);
    assign layer0_outputs[294] = ~(inputs[596]);
    assign layer0_outputs[295] = (inputs[377]) | (inputs[65]);
    assign layer0_outputs[296] = (inputs[619]) | (inputs[139]);
    assign layer0_outputs[297] = ~(inputs[529]);
    assign layer0_outputs[298] = ~(inputs[534]) | (inputs[954]);
    assign layer0_outputs[299] = ~(inputs[139]);
    assign layer0_outputs[300] = 1'b1;
    assign layer0_outputs[301] = ~((inputs[874]) ^ (inputs[780]));
    assign layer0_outputs[302] = ~(inputs[501]);
    assign layer0_outputs[303] = (inputs[445]) | (inputs[788]);
    assign layer0_outputs[304] = (inputs[755]) | (inputs[545]);
    assign layer0_outputs[305] = ~(inputs[951]);
    assign layer0_outputs[306] = (inputs[446]) | (inputs[845]);
    assign layer0_outputs[307] = ~(inputs[221]) | (inputs[983]);
    assign layer0_outputs[308] = inputs[26];
    assign layer0_outputs[309] = ~((inputs[957]) ^ (inputs[409]));
    assign layer0_outputs[310] = (inputs[61]) | (inputs[175]);
    assign layer0_outputs[311] = ~(inputs[453]) | (inputs[568]);
    assign layer0_outputs[312] = ~(inputs[931]) | (inputs[45]);
    assign layer0_outputs[313] = 1'b0;
    assign layer0_outputs[314] = (inputs[176]) | (inputs[786]);
    assign layer0_outputs[315] = inputs[883];
    assign layer0_outputs[316] = ~(inputs[137]) | (inputs[226]);
    assign layer0_outputs[317] = ~(inputs[854]);
    assign layer0_outputs[318] = inputs[101];
    assign layer0_outputs[319] = ~((inputs[29]) | (inputs[512]));
    assign layer0_outputs[320] = (inputs[527]) & ~(inputs[70]);
    assign layer0_outputs[321] = ~((inputs[479]) | (inputs[401]));
    assign layer0_outputs[322] = (inputs[575]) ^ (inputs[731]);
    assign layer0_outputs[323] = ~(inputs[353]);
    assign layer0_outputs[324] = (inputs[863]) & (inputs[148]);
    assign layer0_outputs[325] = ~((inputs[674]) | (inputs[632]));
    assign layer0_outputs[326] = inputs[559];
    assign layer0_outputs[327] = ~(inputs[540]) | (inputs[46]);
    assign layer0_outputs[328] = ~(inputs[644]);
    assign layer0_outputs[329] = (inputs[54]) | (inputs[113]);
    assign layer0_outputs[330] = inputs[706];
    assign layer0_outputs[331] = ~((inputs[243]) | (inputs[526]));
    assign layer0_outputs[332] = ~((inputs[140]) | (inputs[651]));
    assign layer0_outputs[333] = ~((inputs[540]) ^ (inputs[2]));
    assign layer0_outputs[334] = (inputs[468]) ^ (inputs[663]);
    assign layer0_outputs[335] = 1'b0;
    assign layer0_outputs[336] = (inputs[363]) | (inputs[671]);
    assign layer0_outputs[337] = ~((inputs[410]) | (inputs[553]));
    assign layer0_outputs[338] = ~(inputs[232]) | (inputs[516]);
    assign layer0_outputs[339] = ~(inputs[567]);
    assign layer0_outputs[340] = ~(inputs[715]);
    assign layer0_outputs[341] = inputs[94];
    assign layer0_outputs[342] = ~(inputs[398]) | (inputs[831]);
    assign layer0_outputs[343] = (inputs[242]) & ~(inputs[508]);
    assign layer0_outputs[344] = inputs[493];
    assign layer0_outputs[345] = (inputs[811]) | (inputs[702]);
    assign layer0_outputs[346] = ~(inputs[595]) | (inputs[693]);
    assign layer0_outputs[347] = (inputs[788]) | (inputs[105]);
    assign layer0_outputs[348] = inputs[725];
    assign layer0_outputs[349] = (inputs[480]) | (inputs[915]);
    assign layer0_outputs[350] = ~(inputs[189]);
    assign layer0_outputs[351] = ~((inputs[938]) ^ (inputs[380]));
    assign layer0_outputs[352] = inputs[396];
    assign layer0_outputs[353] = (inputs[585]) & ~(inputs[858]);
    assign layer0_outputs[354] = (inputs[343]) | (inputs[478]);
    assign layer0_outputs[355] = (inputs[824]) | (inputs[643]);
    assign layer0_outputs[356] = (inputs[779]) ^ (inputs[903]);
    assign layer0_outputs[357] = 1'b0;
    assign layer0_outputs[358] = (inputs[744]) & ~(inputs[958]);
    assign layer0_outputs[359] = ~((inputs[445]) | (inputs[601]));
    assign layer0_outputs[360] = ~(inputs[389]);
    assign layer0_outputs[361] = ~((inputs[824]) | (inputs[251]));
    assign layer0_outputs[362] = ~((inputs[146]) | (inputs[729]));
    assign layer0_outputs[363] = (inputs[914]) & ~(inputs[808]);
    assign layer0_outputs[364] = ~(inputs[603]) | (inputs[741]);
    assign layer0_outputs[365] = ~(inputs[759]);
    assign layer0_outputs[366] = ~(inputs[395]) | (inputs[739]);
    assign layer0_outputs[367] = ~(inputs[758]) | (inputs[439]);
    assign layer0_outputs[368] = ~((inputs[315]) | (inputs[334]));
    assign layer0_outputs[369] = (inputs[505]) & ~(inputs[993]);
    assign layer0_outputs[370] = 1'b0;
    assign layer0_outputs[371] = ~((inputs[1019]) | (inputs[923]));
    assign layer0_outputs[372] = ~((inputs[976]) ^ (inputs[838]));
    assign layer0_outputs[373] = ~(inputs[160]) | (inputs[481]);
    assign layer0_outputs[374] = (inputs[882]) ^ (inputs[971]);
    assign layer0_outputs[375] = (inputs[151]) & ~(inputs[989]);
    assign layer0_outputs[376] = ~((inputs[28]) | (inputs[100]));
    assign layer0_outputs[377] = ~(inputs[364]) | (inputs[142]);
    assign layer0_outputs[378] = ~((inputs[148]) | (inputs[146]));
    assign layer0_outputs[379] = ~(inputs[958]);
    assign layer0_outputs[380] = (inputs[90]) ^ (inputs[648]);
    assign layer0_outputs[381] = ~(inputs[676]) | (inputs[67]);
    assign layer0_outputs[382] = ~(inputs[972]) | (inputs[271]);
    assign layer0_outputs[383] = ~(inputs[50]) | (inputs[769]);
    assign layer0_outputs[384] = ~(inputs[233]);
    assign layer0_outputs[385] = inputs[590];
    assign layer0_outputs[386] = (inputs[219]) & ~(inputs[92]);
    assign layer0_outputs[387] = ~(inputs[460]) | (inputs[102]);
    assign layer0_outputs[388] = ~((inputs[276]) | (inputs[374]));
    assign layer0_outputs[389] = ~(inputs[710]) | (inputs[946]);
    assign layer0_outputs[390] = ~(inputs[896]) | (inputs[501]);
    assign layer0_outputs[391] = ~((inputs[122]) ^ (inputs[440]));
    assign layer0_outputs[392] = (inputs[219]) & ~(inputs[606]);
    assign layer0_outputs[393] = (inputs[472]) & ~(inputs[35]);
    assign layer0_outputs[394] = (inputs[133]) ^ (inputs[264]);
    assign layer0_outputs[395] = ~(inputs[653]);
    assign layer0_outputs[396] = inputs[465];
    assign layer0_outputs[397] = (inputs[555]) ^ (inputs[992]);
    assign layer0_outputs[398] = inputs[661];
    assign layer0_outputs[399] = ~((inputs[247]) | (inputs[985]));
    assign layer0_outputs[400] = 1'b0;
    assign layer0_outputs[401] = (inputs[437]) & (inputs[557]);
    assign layer0_outputs[402] = inputs[793];
    assign layer0_outputs[403] = ~(inputs[694]) | (inputs[224]);
    assign layer0_outputs[404] = ~(inputs[211]);
    assign layer0_outputs[405] = ~((inputs[677]) ^ (inputs[96]));
    assign layer0_outputs[406] = (inputs[172]) & ~(inputs[547]);
    assign layer0_outputs[407] = (inputs[342]) & ~(inputs[82]);
    assign layer0_outputs[408] = (inputs[100]) ^ (inputs[951]);
    assign layer0_outputs[409] = (inputs[174]) | (inputs[452]);
    assign layer0_outputs[410] = inputs[717];
    assign layer0_outputs[411] = ~((inputs[901]) & (inputs[285]));
    assign layer0_outputs[412] = ~(inputs[63]) | (inputs[802]);
    assign layer0_outputs[413] = ~((inputs[619]) | (inputs[245]));
    assign layer0_outputs[414] = (inputs[428]) & ~(inputs[944]);
    assign layer0_outputs[415] = ~(inputs[435]) | (inputs[925]);
    assign layer0_outputs[416] = ~((inputs[711]) | (inputs[205]));
    assign layer0_outputs[417] = ~(inputs[802]) | (inputs[972]);
    assign layer0_outputs[418] = ~(inputs[953]) | (inputs[900]);
    assign layer0_outputs[419] = ~(inputs[74]) | (inputs[611]);
    assign layer0_outputs[420] = ~((inputs[767]) ^ (inputs[221]));
    assign layer0_outputs[421] = (inputs[73]) | (inputs[726]);
    assign layer0_outputs[422] = inputs[867];
    assign layer0_outputs[423] = ~(inputs[91]) | (inputs[204]);
    assign layer0_outputs[424] = (inputs[11]) | (inputs[751]);
    assign layer0_outputs[425] = inputs[53];
    assign layer0_outputs[426] = ~(inputs[504]);
    assign layer0_outputs[427] = inputs[57];
    assign layer0_outputs[428] = 1'b0;
    assign layer0_outputs[429] = ~(inputs[995]);
    assign layer0_outputs[430] = ~((inputs[593]) ^ (inputs[229]));
    assign layer0_outputs[431] = ~(inputs[916]) | (inputs[645]);
    assign layer0_outputs[432] = (inputs[896]) & (inputs[1004]);
    assign layer0_outputs[433] = ~(inputs[443]) | (inputs[954]);
    assign layer0_outputs[434] = ~(inputs[920]);
    assign layer0_outputs[435] = (inputs[596]) & ~(inputs[117]);
    assign layer0_outputs[436] = ~(inputs[275]) | (inputs[466]);
    assign layer0_outputs[437] = (inputs[937]) | (inputs[624]);
    assign layer0_outputs[438] = (inputs[341]) & ~(inputs[76]);
    assign layer0_outputs[439] = (inputs[818]) | (inputs[677]);
    assign layer0_outputs[440] = inputs[170];
    assign layer0_outputs[441] = ~(inputs[81]) | (inputs[392]);
    assign layer0_outputs[442] = ~((inputs[109]) ^ (inputs[17]));
    assign layer0_outputs[443] = ~((inputs[937]) | (inputs[119]));
    assign layer0_outputs[444] = ~((inputs[842]) | (inputs[940]));
    assign layer0_outputs[445] = ~((inputs[729]) ^ (inputs[861]));
    assign layer0_outputs[446] = 1'b0;
    assign layer0_outputs[447] = (inputs[146]) ^ (inputs[955]);
    assign layer0_outputs[448] = ~(inputs[446]) | (inputs[577]);
    assign layer0_outputs[449] = (inputs[663]) & ~(inputs[518]);
    assign layer0_outputs[450] = ~((inputs[971]) ^ (inputs[92]));
    assign layer0_outputs[451] = ~(inputs[487]);
    assign layer0_outputs[452] = inputs[565];
    assign layer0_outputs[453] = (inputs[802]) | (inputs[585]);
    assign layer0_outputs[454] = ~(inputs[463]);
    assign layer0_outputs[455] = inputs[338];
    assign layer0_outputs[456] = (inputs[125]) ^ (inputs[914]);
    assign layer0_outputs[457] = ~((inputs[176]) | (inputs[647]));
    assign layer0_outputs[458] = ~(inputs[428]) | (inputs[912]);
    assign layer0_outputs[459] = ~((inputs[934]) | (inputs[724]));
    assign layer0_outputs[460] = inputs[940];
    assign layer0_outputs[461] = (inputs[783]) & ~(inputs[515]);
    assign layer0_outputs[462] = ~(inputs[450]);
    assign layer0_outputs[463] = inputs[393];
    assign layer0_outputs[464] = ~((inputs[772]) ^ (inputs[730]));
    assign layer0_outputs[465] = 1'b1;
    assign layer0_outputs[466] = ~(inputs[334]) | (inputs[643]);
    assign layer0_outputs[467] = 1'b0;
    assign layer0_outputs[468] = ~(inputs[386]) | (inputs[445]);
    assign layer0_outputs[469] = ~(inputs[517]);
    assign layer0_outputs[470] = (inputs[211]) ^ (inputs[713]);
    assign layer0_outputs[471] = ~(inputs[915]);
    assign layer0_outputs[472] = (inputs[110]) | (inputs[956]);
    assign layer0_outputs[473] = (inputs[1010]) ^ (inputs[800]);
    assign layer0_outputs[474] = (inputs[469]) & ~(inputs[170]);
    assign layer0_outputs[475] = (inputs[347]) ^ (inputs[833]);
    assign layer0_outputs[476] = ~((inputs[680]) | (inputs[743]));
    assign layer0_outputs[477] = ~((inputs[988]) & (inputs[979]));
    assign layer0_outputs[478] = (inputs[370]) | (inputs[765]);
    assign layer0_outputs[479] = (inputs[118]) & (inputs[256]);
    assign layer0_outputs[480] = inputs[715];
    assign layer0_outputs[481] = ~((inputs[264]) | (inputs[880]));
    assign layer0_outputs[482] = inputs[533];
    assign layer0_outputs[483] = ~((inputs[600]) ^ (inputs[648]));
    assign layer0_outputs[484] = ~(inputs[691]);
    assign layer0_outputs[485] = ~(inputs[701]);
    assign layer0_outputs[486] = ~((inputs[791]) | (inputs[718]));
    assign layer0_outputs[487] = (inputs[620]) & ~(inputs[16]);
    assign layer0_outputs[488] = (inputs[197]) ^ (inputs[632]);
    assign layer0_outputs[489] = ~((inputs[987]) ^ (inputs[225]));
    assign layer0_outputs[490] = ~(inputs[373]) | (inputs[194]);
    assign layer0_outputs[491] = ~(inputs[371]);
    assign layer0_outputs[492] = ~((inputs[378]) ^ (inputs[373]));
    assign layer0_outputs[493] = ~((inputs[323]) | (inputs[171]));
    assign layer0_outputs[494] = (inputs[1]) | (inputs[33]);
    assign layer0_outputs[495] = ~((inputs[620]) | (inputs[830]));
    assign layer0_outputs[496] = inputs[538];
    assign layer0_outputs[497] = ~(inputs[468]) | (inputs[663]);
    assign layer0_outputs[498] = ~(inputs[808]) | (inputs[291]);
    assign layer0_outputs[499] = (inputs[878]) & ~(inputs[144]);
    assign layer0_outputs[500] = ~((inputs[801]) ^ (inputs[812]));
    assign layer0_outputs[501] = (inputs[937]) & ~(inputs[199]);
    assign layer0_outputs[502] = (inputs[79]) & ~(inputs[993]);
    assign layer0_outputs[503] = (inputs[249]) & ~(inputs[32]);
    assign layer0_outputs[504] = 1'b0;
    assign layer0_outputs[505] = (inputs[156]) & ~(inputs[583]);
    assign layer0_outputs[506] = ~(inputs[720]);
    assign layer0_outputs[507] = ~((inputs[985]) ^ (inputs[458]));
    assign layer0_outputs[508] = (inputs[580]) ^ (inputs[565]);
    assign layer0_outputs[509] = inputs[942];
    assign layer0_outputs[510] = inputs[877];
    assign layer0_outputs[511] = (inputs[319]) & ~(inputs[0]);
    assign layer0_outputs[512] = ~(inputs[940]) | (inputs[444]);
    assign layer0_outputs[513] = (inputs[499]) & ~(inputs[155]);
    assign layer0_outputs[514] = (inputs[115]) & ~(inputs[701]);
    assign layer0_outputs[515] = (inputs[811]) ^ (inputs[854]);
    assign layer0_outputs[516] = inputs[560];
    assign layer0_outputs[517] = ~(inputs[413]);
    assign layer0_outputs[518] = (inputs[76]) & (inputs[707]);
    assign layer0_outputs[519] = ~((inputs[194]) ^ (inputs[403]));
    assign layer0_outputs[520] = ~(inputs[645]);
    assign layer0_outputs[521] = (inputs[44]) | (inputs[726]);
    assign layer0_outputs[522] = ~((inputs[957]) & (inputs[67]));
    assign layer0_outputs[523] = (inputs[68]) | (inputs[284]);
    assign layer0_outputs[524] = inputs[552];
    assign layer0_outputs[525] = ~(inputs[886]);
    assign layer0_outputs[526] = (inputs[846]) & ~(inputs[36]);
    assign layer0_outputs[527] = (inputs[500]) | (inputs[387]);
    assign layer0_outputs[528] = (inputs[708]) | (inputs[684]);
    assign layer0_outputs[529] = ~(inputs[626]) | (inputs[894]);
    assign layer0_outputs[530] = ~((inputs[958]) ^ (inputs[537]));
    assign layer0_outputs[531] = (inputs[170]) | (inputs[818]);
    assign layer0_outputs[532] = (inputs[366]) ^ (inputs[666]);
    assign layer0_outputs[533] = ~((inputs[39]) ^ (inputs[165]));
    assign layer0_outputs[534] = (inputs[641]) ^ (inputs[311]);
    assign layer0_outputs[535] = (inputs[924]) ^ (inputs[777]);
    assign layer0_outputs[536] = ~((inputs[918]) ^ (inputs[445]));
    assign layer0_outputs[537] = ~((inputs[353]) ^ (inputs[693]));
    assign layer0_outputs[538] = ~(inputs[424]);
    assign layer0_outputs[539] = 1'b0;
    assign layer0_outputs[540] = ~((inputs[11]) | (inputs[643]));
    assign layer0_outputs[541] = ~(inputs[709]) | (inputs[518]);
    assign layer0_outputs[542] = ~(inputs[589]) | (inputs[770]);
    assign layer0_outputs[543] = ~((inputs[404]) | (inputs[230]));
    assign layer0_outputs[544] = (inputs[631]) & ~(inputs[853]);
    assign layer0_outputs[545] = inputs[653];
    assign layer0_outputs[546] = ~((inputs[1005]) ^ (inputs[959]));
    assign layer0_outputs[547] = ~((inputs[226]) ^ (inputs[109]));
    assign layer0_outputs[548] = ~((inputs[176]) | (inputs[822]));
    assign layer0_outputs[549] = ~((inputs[923]) | (inputs[407]));
    assign layer0_outputs[550] = (inputs[626]) & ~(inputs[204]);
    assign layer0_outputs[551] = ~((inputs[5]) & (inputs[823]));
    assign layer0_outputs[552] = 1'b0;
    assign layer0_outputs[553] = ~(inputs[349]);
    assign layer0_outputs[554] = ~(inputs[489]) | (inputs[327]);
    assign layer0_outputs[555] = ~(inputs[578]) | (inputs[997]);
    assign layer0_outputs[556] = 1'b1;
    assign layer0_outputs[557] = ~((inputs[999]) | (inputs[461]));
    assign layer0_outputs[558] = ~(inputs[302]) | (inputs[458]);
    assign layer0_outputs[559] = ~(inputs[652]) | (inputs[1002]);
    assign layer0_outputs[560] = (inputs[601]) | (inputs[38]);
    assign layer0_outputs[561] = ~(inputs[713]) | (inputs[900]);
    assign layer0_outputs[562] = (inputs[654]) | (inputs[261]);
    assign layer0_outputs[563] = 1'b0;
    assign layer0_outputs[564] = inputs[781];
    assign layer0_outputs[565] = (inputs[425]) | (inputs[376]);
    assign layer0_outputs[566] = inputs[549];
    assign layer0_outputs[567] = (inputs[742]) & ~(inputs[94]);
    assign layer0_outputs[568] = ~(inputs[338]);
    assign layer0_outputs[569] = (inputs[561]) & ~(inputs[486]);
    assign layer0_outputs[570] = (inputs[58]) ^ (inputs[494]);
    assign layer0_outputs[571] = ~(inputs[733]);
    assign layer0_outputs[572] = (inputs[388]) & ~(inputs[800]);
    assign layer0_outputs[573] = (inputs[754]) & ~(inputs[358]);
    assign layer0_outputs[574] = inputs[772];
    assign layer0_outputs[575] = (inputs[1008]) & ~(inputs[1017]);
    assign layer0_outputs[576] = (inputs[963]) & (inputs[68]);
    assign layer0_outputs[577] = ~(inputs[278]);
    assign layer0_outputs[578] = ~((inputs[711]) ^ (inputs[228]));
    assign layer0_outputs[579] = ~(inputs[538]) | (inputs[201]);
    assign layer0_outputs[580] = ~((inputs[85]) | (inputs[1002]));
    assign layer0_outputs[581] = ~(inputs[115]);
    assign layer0_outputs[582] = ~(inputs[653]) | (inputs[357]);
    assign layer0_outputs[583] = ~((inputs[374]) | (inputs[356]));
    assign layer0_outputs[584] = (inputs[992]) | (inputs[697]);
    assign layer0_outputs[585] = (inputs[886]) & (inputs[768]);
    assign layer0_outputs[586] = (inputs[361]) ^ (inputs[430]);
    assign layer0_outputs[587] = ~(inputs[715]);
    assign layer0_outputs[588] = inputs[692];
    assign layer0_outputs[589] = inputs[920];
    assign layer0_outputs[590] = inputs[24];
    assign layer0_outputs[591] = inputs[408];
    assign layer0_outputs[592] = ~(inputs[996]) | (inputs[82]);
    assign layer0_outputs[593] = ~((inputs[908]) ^ (inputs[910]));
    assign layer0_outputs[594] = inputs[304];
    assign layer0_outputs[595] = ~(inputs[808]) | (inputs[155]);
    assign layer0_outputs[596] = ~((inputs[589]) | (inputs[446]));
    assign layer0_outputs[597] = (inputs[269]) | (inputs[589]);
    assign layer0_outputs[598] = (inputs[80]) & (inputs[280]);
    assign layer0_outputs[599] = (inputs[289]) & (inputs[320]);
    assign layer0_outputs[600] = inputs[901];
    assign layer0_outputs[601] = ~(inputs[606]) | (inputs[10]);
    assign layer0_outputs[602] = inputs[129];
    assign layer0_outputs[603] = ~((inputs[30]) | (inputs[655]));
    assign layer0_outputs[604] = (inputs[897]) & ~(inputs[24]);
    assign layer0_outputs[605] = ~(inputs[54]);
    assign layer0_outputs[606] = inputs[619];
    assign layer0_outputs[607] = (inputs[640]) | (inputs[518]);
    assign layer0_outputs[608] = (inputs[406]) ^ (inputs[961]);
    assign layer0_outputs[609] = ~((inputs[827]) ^ (inputs[73]));
    assign layer0_outputs[610] = ~(inputs[601]);
    assign layer0_outputs[611] = ~((inputs[649]) ^ (inputs[780]));
    assign layer0_outputs[612] = (inputs[944]) | (inputs[983]);
    assign layer0_outputs[613] = ~((inputs[262]) ^ (inputs[707]));
    assign layer0_outputs[614] = ~((inputs[995]) | (inputs[469]));
    assign layer0_outputs[615] = (inputs[362]) & ~(inputs[117]);
    assign layer0_outputs[616] = (inputs[246]) & (inputs[1002]);
    assign layer0_outputs[617] = (inputs[424]) & ~(inputs[383]);
    assign layer0_outputs[618] = ~((inputs[847]) ^ (inputs[968]));
    assign layer0_outputs[619] = (inputs[432]) & ~(inputs[389]);
    assign layer0_outputs[620] = (inputs[592]) | (inputs[540]);
    assign layer0_outputs[621] = 1'b1;
    assign layer0_outputs[622] = inputs[471];
    assign layer0_outputs[623] = ~((inputs[728]) & (inputs[634]));
    assign layer0_outputs[624] = (inputs[998]) ^ (inputs[457]);
    assign layer0_outputs[625] = ~((inputs[795]) | (inputs[16]));
    assign layer0_outputs[626] = ~(inputs[956]) | (inputs[419]);
    assign layer0_outputs[627] = (inputs[208]) ^ (inputs[135]);
    assign layer0_outputs[628] = ~(inputs[736]);
    assign layer0_outputs[629] = (inputs[621]) | (inputs[145]);
    assign layer0_outputs[630] = ~((inputs[337]) | (inputs[739]));
    assign layer0_outputs[631] = (inputs[577]) & (inputs[858]);
    assign layer0_outputs[632] = (inputs[175]) & ~(inputs[356]);
    assign layer0_outputs[633] = ~(inputs[947]);
    assign layer0_outputs[634] = inputs[883];
    assign layer0_outputs[635] = ~(inputs[1023]) | (inputs[186]);
    assign layer0_outputs[636] = inputs[321];
    assign layer0_outputs[637] = inputs[850];
    assign layer0_outputs[638] = (inputs[389]) ^ (inputs[137]);
    assign layer0_outputs[639] = inputs[592];
    assign layer0_outputs[640] = ~((inputs[379]) ^ (inputs[151]));
    assign layer0_outputs[641] = ~((inputs[663]) ^ (inputs[201]));
    assign layer0_outputs[642] = (inputs[801]) ^ (inputs[743]);
    assign layer0_outputs[643] = (inputs[632]) | (inputs[210]);
    assign layer0_outputs[644] = inputs[659];
    assign layer0_outputs[645] = (inputs[686]) ^ (inputs[830]);
    assign layer0_outputs[646] = (inputs[764]) | (inputs[175]);
    assign layer0_outputs[647] = inputs[429];
    assign layer0_outputs[648] = ~((inputs[285]) | (inputs[430]));
    assign layer0_outputs[649] = ~(inputs[849]) | (inputs[201]);
    assign layer0_outputs[650] = ~(inputs[224]) | (inputs[483]);
    assign layer0_outputs[651] = (inputs[809]) & ~(inputs[865]);
    assign layer0_outputs[652] = (inputs[221]) ^ (inputs[496]);
    assign layer0_outputs[653] = (inputs[292]) | (inputs[989]);
    assign layer0_outputs[654] = (inputs[644]) & (inputs[610]);
    assign layer0_outputs[655] = (inputs[342]) & (inputs[297]);
    assign layer0_outputs[656] = ~((inputs[290]) & (inputs[13]));
    assign layer0_outputs[657] = 1'b1;
    assign layer0_outputs[658] = ~(inputs[593]) | (inputs[364]);
    assign layer0_outputs[659] = ~((inputs[694]) | (inputs[116]));
    assign layer0_outputs[660] = 1'b0;
    assign layer0_outputs[661] = (inputs[688]) & ~(inputs[677]);
    assign layer0_outputs[662] = ~(inputs[820]) | (inputs[30]);
    assign layer0_outputs[663] = ~((inputs[577]) | (inputs[272]));
    assign layer0_outputs[664] = (inputs[676]) ^ (inputs[809]);
    assign layer0_outputs[665] = (inputs[134]) | (inputs[211]);
    assign layer0_outputs[666] = (inputs[759]) ^ (inputs[522]);
    assign layer0_outputs[667] = inputs[617];
    assign layer0_outputs[668] = (inputs[502]) & ~(inputs[770]);
    assign layer0_outputs[669] = ~(inputs[406]);
    assign layer0_outputs[670] = inputs[460];
    assign layer0_outputs[671] = ~(inputs[691]);
    assign layer0_outputs[672] = 1'b0;
    assign layer0_outputs[673] = (inputs[517]) | (inputs[656]);
    assign layer0_outputs[674] = inputs[459];
    assign layer0_outputs[675] = ~(inputs[35]);
    assign layer0_outputs[676] = (inputs[536]) & ~(inputs[997]);
    assign layer0_outputs[677] = inputs[267];
    assign layer0_outputs[678] = (inputs[580]) ^ (inputs[351]);
    assign layer0_outputs[679] = ~((inputs[672]) ^ (inputs[573]));
    assign layer0_outputs[680] = ~((inputs[682]) | (inputs[636]));
    assign layer0_outputs[681] = ~(inputs[981]) | (inputs[255]);
    assign layer0_outputs[682] = (inputs[820]) & ~(inputs[144]);
    assign layer0_outputs[683] = (inputs[517]) ^ (inputs[756]);
    assign layer0_outputs[684] = ~(inputs[39]);
    assign layer0_outputs[685] = inputs[915];
    assign layer0_outputs[686] = ~((inputs[115]) & (inputs[939]));
    assign layer0_outputs[687] = (inputs[679]) & ~(inputs[61]);
    assign layer0_outputs[688] = ~(inputs[272]) | (inputs[615]);
    assign layer0_outputs[689] = ~((inputs[429]) | (inputs[555]));
    assign layer0_outputs[690] = ~(inputs[519]);
    assign layer0_outputs[691] = (inputs[219]) & ~(inputs[930]);
    assign layer0_outputs[692] = (inputs[428]) & ~(inputs[677]);
    assign layer0_outputs[693] = inputs[390];
    assign layer0_outputs[694] = (inputs[878]) | (inputs[942]);
    assign layer0_outputs[695] = ~((inputs[201]) & (inputs[356]));
    assign layer0_outputs[696] = ~((inputs[686]) | (inputs[710]));
    assign layer0_outputs[697] = inputs[498];
    assign layer0_outputs[698] = (inputs[206]) & ~(inputs[566]);
    assign layer0_outputs[699] = ~(inputs[141]) | (inputs[19]);
    assign layer0_outputs[700] = ~((inputs[413]) ^ (inputs[833]));
    assign layer0_outputs[701] = ~(inputs[749]);
    assign layer0_outputs[702] = (inputs[488]) | (inputs[47]);
    assign layer0_outputs[703] = ~(inputs[649]) | (inputs[671]);
    assign layer0_outputs[704] = ~(inputs[942]) | (inputs[148]);
    assign layer0_outputs[705] = 1'b0;
    assign layer0_outputs[706] = ~(inputs[3]) | (inputs[698]);
    assign layer0_outputs[707] = (inputs[9]) & ~(inputs[703]);
    assign layer0_outputs[708] = ~((inputs[966]) & (inputs[887]));
    assign layer0_outputs[709] = (inputs[662]) | (inputs[632]);
    assign layer0_outputs[710] = (inputs[979]) | (inputs[909]);
    assign layer0_outputs[711] = ~(inputs[604]);
    assign layer0_outputs[712] = (inputs[276]) & ~(inputs[770]);
    assign layer0_outputs[713] = inputs[495];
    assign layer0_outputs[714] = ~(inputs[821]) | (inputs[385]);
    assign layer0_outputs[715] = ~(inputs[749]);
    assign layer0_outputs[716] = ~((inputs[607]) ^ (inputs[205]));
    assign layer0_outputs[717] = (inputs[315]) ^ (inputs[64]);
    assign layer0_outputs[718] = ~(inputs[459]);
    assign layer0_outputs[719] = ~(inputs[436]);
    assign layer0_outputs[720] = ~(inputs[585]);
    assign layer0_outputs[721] = inputs[309];
    assign layer0_outputs[722] = ~(inputs[599]) | (inputs[281]);
    assign layer0_outputs[723] = (inputs[686]) & ~(inputs[381]);
    assign layer0_outputs[724] = inputs[347];
    assign layer0_outputs[725] = inputs[740];
    assign layer0_outputs[726] = 1'b1;
    assign layer0_outputs[727] = ~((inputs[324]) ^ (inputs[540]));
    assign layer0_outputs[728] = ~((inputs[484]) & (inputs[355]));
    assign layer0_outputs[729] = (inputs[962]) | (inputs[354]);
    assign layer0_outputs[730] = (inputs[40]) ^ (inputs[443]);
    assign layer0_outputs[731] = ~((inputs[807]) ^ (inputs[529]));
    assign layer0_outputs[732] = (inputs[499]) & ~(inputs[888]);
    assign layer0_outputs[733] = inputs[531];
    assign layer0_outputs[734] = ~(inputs[861]) | (inputs[50]);
    assign layer0_outputs[735] = ~((inputs[924]) & (inputs[162]));
    assign layer0_outputs[736] = ~(inputs[824]);
    assign layer0_outputs[737] = (inputs[504]) | (inputs[344]);
    assign layer0_outputs[738] = ~((inputs[686]) | (inputs[444]));
    assign layer0_outputs[739] = (inputs[382]) & ~(inputs[820]);
    assign layer0_outputs[740] = ~((inputs[871]) & (inputs[79]));
    assign layer0_outputs[741] = 1'b1;
    assign layer0_outputs[742] = ~((inputs[603]) ^ (inputs[980]));
    assign layer0_outputs[743] = (inputs[984]) | (inputs[745]);
    assign layer0_outputs[744] = (inputs[978]) ^ (inputs[319]);
    assign layer0_outputs[745] = (inputs[358]) & (inputs[367]);
    assign layer0_outputs[746] = (inputs[43]) | (inputs[1010]);
    assign layer0_outputs[747] = inputs[787];
    assign layer0_outputs[748] = (inputs[943]) | (inputs[630]);
    assign layer0_outputs[749] = (inputs[257]) ^ (inputs[775]);
    assign layer0_outputs[750] = (inputs[257]) ^ (inputs[21]);
    assign layer0_outputs[751] = (inputs[386]) ^ (inputs[813]);
    assign layer0_outputs[752] = ~((inputs[185]) | (inputs[725]));
    assign layer0_outputs[753] = (inputs[171]) & ~(inputs[968]);
    assign layer0_outputs[754] = ~((inputs[524]) ^ (inputs[817]));
    assign layer0_outputs[755] = (inputs[66]) & (inputs[23]);
    assign layer0_outputs[756] = ~((inputs[2]) | (inputs[338]));
    assign layer0_outputs[757] = ~((inputs[843]) & (inputs[424]));
    assign layer0_outputs[758] = ~((inputs[529]) | (inputs[982]));
    assign layer0_outputs[759] = ~((inputs[803]) ^ (inputs[849]));
    assign layer0_outputs[760] = (inputs[193]) & (inputs[387]);
    assign layer0_outputs[761] = ~(inputs[478]);
    assign layer0_outputs[762] = ~((inputs[560]) | (inputs[225]));
    assign layer0_outputs[763] = inputs[270];
    assign layer0_outputs[764] = 1'b1;
    assign layer0_outputs[765] = (inputs[536]) & ~(inputs[718]);
    assign layer0_outputs[766] = ~(inputs[936]);
    assign layer0_outputs[767] = ~((inputs[662]) | (inputs[58]));
    assign layer0_outputs[768] = 1'b1;
    assign layer0_outputs[769] = ~((inputs[973]) ^ (inputs[522]));
    assign layer0_outputs[770] = inputs[498];
    assign layer0_outputs[771] = (inputs[571]) | (inputs[574]);
    assign layer0_outputs[772] = ~(inputs[981]) | (inputs[95]);
    assign layer0_outputs[773] = inputs[59];
    assign layer0_outputs[774] = (inputs[1020]) & ~(inputs[766]);
    assign layer0_outputs[775] = inputs[571];
    assign layer0_outputs[776] = (inputs[53]) ^ (inputs[628]);
    assign layer0_outputs[777] = (inputs[42]) | (inputs[401]);
    assign layer0_outputs[778] = ~((inputs[972]) ^ (inputs[770]));
    assign layer0_outputs[779] = (inputs[357]) | (inputs[729]);
    assign layer0_outputs[780] = inputs[225];
    assign layer0_outputs[781] = inputs[297];
    assign layer0_outputs[782] = inputs[176];
    assign layer0_outputs[783] = (inputs[927]) & (inputs[22]);
    assign layer0_outputs[784] = (inputs[334]) & ~(inputs[161]);
    assign layer0_outputs[785] = (inputs[498]) & (inputs[661]);
    assign layer0_outputs[786] = ~((inputs[666]) | (inputs[50]));
    assign layer0_outputs[787] = ~((inputs[333]) ^ (inputs[576]));
    assign layer0_outputs[788] = ~(inputs[333]);
    assign layer0_outputs[789] = ~((inputs[800]) | (inputs[659]));
    assign layer0_outputs[790] = (inputs[127]) ^ (inputs[763]);
    assign layer0_outputs[791] = ~((inputs[633]) | (inputs[134]));
    assign layer0_outputs[792] = (inputs[650]) | (inputs[322]);
    assign layer0_outputs[793] = ~((inputs[16]) ^ (inputs[588]));
    assign layer0_outputs[794] = ~((inputs[476]) | (inputs[722]));
    assign layer0_outputs[795] = (inputs[103]) & (inputs[188]);
    assign layer0_outputs[796] = (inputs[943]) & ~(inputs[260]);
    assign layer0_outputs[797] = ~((inputs[552]) ^ (inputs[490]));
    assign layer0_outputs[798] = ~(inputs[370]) | (inputs[299]);
    assign layer0_outputs[799] = ~(inputs[490]) | (inputs[250]);
    assign layer0_outputs[800] = (inputs[787]) ^ (inputs[191]);
    assign layer0_outputs[801] = (inputs[219]) & (inputs[8]);
    assign layer0_outputs[802] = (inputs[595]) & ~(inputs[780]);
    assign layer0_outputs[803] = ~((inputs[121]) | (inputs[437]));
    assign layer0_outputs[804] = inputs[627];
    assign layer0_outputs[805] = inputs[322];
    assign layer0_outputs[806] = ~(inputs[555]);
    assign layer0_outputs[807] = ~((inputs[982]) & (inputs[450]));
    assign layer0_outputs[808] = ~(inputs[533]);
    assign layer0_outputs[809] = 1'b0;
    assign layer0_outputs[810] = (inputs[116]) & (inputs[119]);
    assign layer0_outputs[811] = ~(inputs[308]);
    assign layer0_outputs[812] = (inputs[342]) | (inputs[79]);
    assign layer0_outputs[813] = ~((inputs[93]) ^ (inputs[350]));
    assign layer0_outputs[814] = ~(inputs[264]);
    assign layer0_outputs[815] = inputs[740];
    assign layer0_outputs[816] = ~(inputs[1009]);
    assign layer0_outputs[817] = inputs[879];
    assign layer0_outputs[818] = (inputs[312]) & (inputs[40]);
    assign layer0_outputs[819] = ~(inputs[635]) | (inputs[435]);
    assign layer0_outputs[820] = (inputs[840]) ^ (inputs[990]);
    assign layer0_outputs[821] = ~(inputs[790]);
    assign layer0_outputs[822] = ~((inputs[491]) & (inputs[429]));
    assign layer0_outputs[823] = ~((inputs[162]) & (inputs[102]));
    assign layer0_outputs[824] = inputs[720];
    assign layer0_outputs[825] = (inputs[411]) ^ (inputs[517]);
    assign layer0_outputs[826] = ~(inputs[902]) | (inputs[1008]);
    assign layer0_outputs[827] = 1'b1;
    assign layer0_outputs[828] = (inputs[348]) & ~(inputs[633]);
    assign layer0_outputs[829] = ~(inputs[569]);
    assign layer0_outputs[830] = (inputs[920]) & ~(inputs[325]);
    assign layer0_outputs[831] = ~(inputs[196]);
    assign layer0_outputs[832] = ~((inputs[966]) ^ (inputs[825]));
    assign layer0_outputs[833] = ~(inputs[497]);
    assign layer0_outputs[834] = ~((inputs[398]) ^ (inputs[976]));
    assign layer0_outputs[835] = ~(inputs[1022]) | (inputs[796]);
    assign layer0_outputs[836] = ~(inputs[594]);
    assign layer0_outputs[837] = (inputs[336]) & ~(inputs[867]);
    assign layer0_outputs[838] = (inputs[397]) ^ (inputs[164]);
    assign layer0_outputs[839] = ~(inputs[327]);
    assign layer0_outputs[840] = (inputs[215]) ^ (inputs[747]);
    assign layer0_outputs[841] = ~((inputs[846]) | (inputs[251]));
    assign layer0_outputs[842] = (inputs[690]) & ~(inputs[840]);
    assign layer0_outputs[843] = (inputs[236]) | (inputs[172]);
    assign layer0_outputs[844] = (inputs[335]) ^ (inputs[2]);
    assign layer0_outputs[845] = ~(inputs[584]);
    assign layer0_outputs[846] = 1'b0;
    assign layer0_outputs[847] = (inputs[855]) ^ (inputs[819]);
    assign layer0_outputs[848] = (inputs[775]) | (inputs[692]);
    assign layer0_outputs[849] = ~(inputs[362]);
    assign layer0_outputs[850] = ~((inputs[576]) | (inputs[318]));
    assign layer0_outputs[851] = ~(inputs[555]) | (inputs[254]);
    assign layer0_outputs[852] = ~(inputs[148]) | (inputs[962]);
    assign layer0_outputs[853] = (inputs[348]) & (inputs[742]);
    assign layer0_outputs[854] = ~((inputs[729]) ^ (inputs[334]));
    assign layer0_outputs[855] = ~((inputs[59]) | (inputs[432]));
    assign layer0_outputs[856] = ~(inputs[786]) | (inputs[576]);
    assign layer0_outputs[857] = (inputs[180]) & ~(inputs[2]);
    assign layer0_outputs[858] = (inputs[322]) & ~(inputs[520]);
    assign layer0_outputs[859] = (inputs[10]) & ~(inputs[163]);
    assign layer0_outputs[860] = inputs[613];
    assign layer0_outputs[861] = ~(inputs[307]) | (inputs[384]);
    assign layer0_outputs[862] = ~((inputs[51]) ^ (inputs[57]));
    assign layer0_outputs[863] = ~(inputs[715]) | (inputs[184]);
    assign layer0_outputs[864] = ~(inputs[637]) | (inputs[638]);
    assign layer0_outputs[865] = ~(inputs[436]);
    assign layer0_outputs[866] = ~(inputs[669]) | (inputs[628]);
    assign layer0_outputs[867] = ~((inputs[977]) ^ (inputs[234]));
    assign layer0_outputs[868] = inputs[949];
    assign layer0_outputs[869] = ~((inputs[790]) | (inputs[683]));
    assign layer0_outputs[870] = ~(inputs[420]) | (inputs[420]);
    assign layer0_outputs[871] = ~((inputs[424]) ^ (inputs[381]));
    assign layer0_outputs[872] = (inputs[870]) & ~(inputs[801]);
    assign layer0_outputs[873] = ~(inputs[577]) | (inputs[827]);
    assign layer0_outputs[874] = ~(inputs[322]);
    assign layer0_outputs[875] = (inputs[622]) | (inputs[617]);
    assign layer0_outputs[876] = inputs[62];
    assign layer0_outputs[877] = ~((inputs[941]) ^ (inputs[257]));
    assign layer0_outputs[878] = ~(inputs[211]);
    assign layer0_outputs[879] = (inputs[602]) ^ (inputs[100]);
    assign layer0_outputs[880] = inputs[134];
    assign layer0_outputs[881] = (inputs[473]) | (inputs[944]);
    assign layer0_outputs[882] = inputs[1004];
    assign layer0_outputs[883] = (inputs[907]) | (inputs[526]);
    assign layer0_outputs[884] = (inputs[475]) & ~(inputs[828]);
    assign layer0_outputs[885] = (inputs[654]) & ~(inputs[288]);
    assign layer0_outputs[886] = (inputs[304]) ^ (inputs[815]);
    assign layer0_outputs[887] = (inputs[875]) & ~(inputs[257]);
    assign layer0_outputs[888] = ~((inputs[69]) ^ (inputs[358]));
    assign layer0_outputs[889] = ~((inputs[969]) ^ (inputs[206]));
    assign layer0_outputs[890] = ~(inputs[431]) | (inputs[888]);
    assign layer0_outputs[891] = ~((inputs[525]) | (inputs[927]));
    assign layer0_outputs[892] = (inputs[296]) | (inputs[94]);
    assign layer0_outputs[893] = ~((inputs[878]) ^ (inputs[895]));
    assign layer0_outputs[894] = ~((inputs[965]) ^ (inputs[708]));
    assign layer0_outputs[895] = ~(inputs[52]);
    assign layer0_outputs[896] = ~(inputs[435]) | (inputs[47]);
    assign layer0_outputs[897] = (inputs[251]) ^ (inputs[774]);
    assign layer0_outputs[898] = ~((inputs[917]) ^ (inputs[315]));
    assign layer0_outputs[899] = ~((inputs[559]) ^ (inputs[998]));
    assign layer0_outputs[900] = (inputs[702]) ^ (inputs[744]);
    assign layer0_outputs[901] = (inputs[587]) ^ (inputs[735]);
    assign layer0_outputs[902] = ~((inputs[138]) | (inputs[697]));
    assign layer0_outputs[903] = (inputs[1]) & (inputs[532]);
    assign layer0_outputs[904] = (inputs[8]) & ~(inputs[476]);
    assign layer0_outputs[905] = ~((inputs[561]) | (inputs[413]));
    assign layer0_outputs[906] = (inputs[769]) | (inputs[582]);
    assign layer0_outputs[907] = (inputs[635]) & ~(inputs[829]);
    assign layer0_outputs[908] = ~(inputs[96]) | (inputs[222]);
    assign layer0_outputs[909] = inputs[563];
    assign layer0_outputs[910] = ~((inputs[56]) | (inputs[623]));
    assign layer0_outputs[911] = ~((inputs[995]) & (inputs[744]));
    assign layer0_outputs[912] = ~(inputs[758]) | (inputs[454]);
    assign layer0_outputs[913] = ~(inputs[638]) | (inputs[875]);
    assign layer0_outputs[914] = (inputs[902]) | (inputs[8]);
    assign layer0_outputs[915] = 1'b1;
    assign layer0_outputs[916] = ~(inputs[377]);
    assign layer0_outputs[917] = inputs[679];
    assign layer0_outputs[918] = ~((inputs[870]) | (inputs[268]));
    assign layer0_outputs[919] = 1'b1;
    assign layer0_outputs[920] = inputs[683];
    assign layer0_outputs[921] = ~(inputs[332]) | (inputs[743]);
    assign layer0_outputs[922] = inputs[847];
    assign layer0_outputs[923] = (inputs[935]) & ~(inputs[888]);
    assign layer0_outputs[924] = ~(inputs[893]) | (inputs[965]);
    assign layer0_outputs[925] = ~(inputs[702]) | (inputs[919]);
    assign layer0_outputs[926] = inputs[478];
    assign layer0_outputs[927] = (inputs[624]) ^ (inputs[63]);
    assign layer0_outputs[928] = ~(inputs[313]) | (inputs[997]);
    assign layer0_outputs[929] = (inputs[190]) & ~(inputs[231]);
    assign layer0_outputs[930] = (inputs[809]) & ~(inputs[419]);
    assign layer0_outputs[931] = inputs[320];
    assign layer0_outputs[932] = 1'b0;
    assign layer0_outputs[933] = inputs[264];
    assign layer0_outputs[934] = ~(inputs[877]);
    assign layer0_outputs[935] = ~(inputs[498]) | (inputs[696]);
    assign layer0_outputs[936] = ~((inputs[682]) ^ (inputs[399]));
    assign layer0_outputs[937] = (inputs[941]) | (inputs[324]);
    assign layer0_outputs[938] = ~((inputs[502]) ^ (inputs[399]));
    assign layer0_outputs[939] = (inputs[549]) & ~(inputs[1015]);
    assign layer0_outputs[940] = ~(inputs[712]) | (inputs[917]);
    assign layer0_outputs[941] = ~(inputs[453]) | (inputs[384]);
    assign layer0_outputs[942] = ~((inputs[669]) | (inputs[855]));
    assign layer0_outputs[943] = inputs[395];
    assign layer0_outputs[944] = (inputs[659]) & (inputs[82]);
    assign layer0_outputs[945] = ~(inputs[711]);
    assign layer0_outputs[946] = (inputs[49]) | (inputs[531]);
    assign layer0_outputs[947] = ~(inputs[266]) | (inputs[536]);
    assign layer0_outputs[948] = (inputs[524]) | (inputs[458]);
    assign layer0_outputs[949] = ~(inputs[722]) | (inputs[34]);
    assign layer0_outputs[950] = ~(inputs[890]);
    assign layer0_outputs[951] = (inputs[533]) | (inputs[506]);
    assign layer0_outputs[952] = (inputs[114]) | (inputs[402]);
    assign layer0_outputs[953] = inputs[233];
    assign layer0_outputs[954] = ~((inputs[115]) ^ (inputs[868]));
    assign layer0_outputs[955] = (inputs[225]) | (inputs[630]);
    assign layer0_outputs[956] = (inputs[490]) & ~(inputs[609]);
    assign layer0_outputs[957] = (inputs[145]) ^ (inputs[291]);
    assign layer0_outputs[958] = (inputs[866]) | (inputs[292]);
    assign layer0_outputs[959] = (inputs[857]) & ~(inputs[104]);
    assign layer0_outputs[960] = ~((inputs[821]) ^ (inputs[44]));
    assign layer0_outputs[961] = inputs[612];
    assign layer0_outputs[962] = inputs[89];
    assign layer0_outputs[963] = ~((inputs[627]) ^ (inputs[932]));
    assign layer0_outputs[964] = (inputs[284]) | (inputs[240]);
    assign layer0_outputs[965] = ~(inputs[601]);
    assign layer0_outputs[966] = (inputs[334]) | (inputs[941]);
    assign layer0_outputs[967] = inputs[523];
    assign layer0_outputs[968] = ~(inputs[341]);
    assign layer0_outputs[969] = ~(inputs[628]);
    assign layer0_outputs[970] = ~((inputs[579]) | (inputs[344]));
    assign layer0_outputs[971] = ~((inputs[184]) | (inputs[952]));
    assign layer0_outputs[972] = ~(inputs[706]) | (inputs[959]);
    assign layer0_outputs[973] = inputs[754];
    assign layer0_outputs[974] = (inputs[247]) | (inputs[904]);
    assign layer0_outputs[975] = ~(inputs[783]);
    assign layer0_outputs[976] = ~(inputs[505]);
    assign layer0_outputs[977] = ~((inputs[184]) | (inputs[362]));
    assign layer0_outputs[978] = (inputs[519]) & ~(inputs[982]);
    assign layer0_outputs[979] = ~(inputs[150]) | (inputs[47]);
    assign layer0_outputs[980] = (inputs[48]) & ~(inputs[796]);
    assign layer0_outputs[981] = ~(inputs[682]);
    assign layer0_outputs[982] = inputs[398];
    assign layer0_outputs[983] = (inputs[380]) ^ (inputs[183]);
    assign layer0_outputs[984] = ~((inputs[288]) & (inputs[1009]));
    assign layer0_outputs[985] = ~((inputs[191]) & (inputs[988]));
    assign layer0_outputs[986] = inputs[459];
    assign layer0_outputs[987] = ~((inputs[462]) ^ (inputs[557]));
    assign layer0_outputs[988] = inputs[825];
    assign layer0_outputs[989] = (inputs[574]) ^ (inputs[1000]);
    assign layer0_outputs[990] = (inputs[743]) | (inputs[711]);
    assign layer0_outputs[991] = (inputs[920]) & (inputs[640]);
    assign layer0_outputs[992] = inputs[218];
    assign layer0_outputs[993] = (inputs[18]) | (inputs[128]);
    assign layer0_outputs[994] = ~((inputs[538]) | (inputs[844]));
    assign layer0_outputs[995] = ~((inputs[474]) ^ (inputs[775]));
    assign layer0_outputs[996] = ~(inputs[329]);
    assign layer0_outputs[997] = ~((inputs[714]) | (inputs[486]));
    assign layer0_outputs[998] = ~(inputs[254]);
    assign layer0_outputs[999] = ~(inputs[500]);
    assign layer0_outputs[1000] = ~((inputs[878]) | (inputs[139]));
    assign layer0_outputs[1001] = ~(inputs[744]);
    assign layer0_outputs[1002] = (inputs[80]) & ~(inputs[642]);
    assign layer0_outputs[1003] = ~(inputs[815]) | (inputs[195]);
    assign layer0_outputs[1004] = (inputs[217]) & ~(inputs[507]);
    assign layer0_outputs[1005] = (inputs[51]) | (inputs[318]);
    assign layer0_outputs[1006] = ~(inputs[442]) | (inputs[797]);
    assign layer0_outputs[1007] = inputs[382];
    assign layer0_outputs[1008] = (inputs[85]) & ~(inputs[53]);
    assign layer0_outputs[1009] = inputs[680];
    assign layer0_outputs[1010] = ~((inputs[173]) ^ (inputs[480]));
    assign layer0_outputs[1011] = (inputs[72]) ^ (inputs[408]);
    assign layer0_outputs[1012] = (inputs[870]) | (inputs[404]);
    assign layer0_outputs[1013] = ~((inputs[647]) ^ (inputs[205]));
    assign layer0_outputs[1014] = ~((inputs[237]) | (inputs[680]));
    assign layer0_outputs[1015] = (inputs[835]) | (inputs[34]);
    assign layer0_outputs[1016] = ~(inputs[777]);
    assign layer0_outputs[1017] = ~(inputs[296]) | (inputs[930]);
    assign layer0_outputs[1018] = ~(inputs[719]);
    assign layer0_outputs[1019] = 1'b0;
    assign layer0_outputs[1020] = (inputs[0]) & ~(inputs[831]);
    assign layer0_outputs[1021] = ~(inputs[884]);
    assign layer0_outputs[1022] = (inputs[774]) & ~(inputs[192]);
    assign layer0_outputs[1023] = inputs[554];
    assign layer0_outputs[1024] = inputs[325];
    assign layer0_outputs[1025] = (inputs[236]) & ~(inputs[163]);
    assign layer0_outputs[1026] = 1'b0;
    assign layer0_outputs[1027] = (inputs[827]) ^ (inputs[716]);
    assign layer0_outputs[1028] = ~(inputs[850]) | (inputs[638]);
    assign layer0_outputs[1029] = ~(inputs[730]);
    assign layer0_outputs[1030] = ~((inputs[60]) ^ (inputs[464]));
    assign layer0_outputs[1031] = ~((inputs[875]) ^ (inputs[259]));
    assign layer0_outputs[1032] = ~((inputs[602]) | (inputs[586]));
    assign layer0_outputs[1033] = ~(inputs[822]) | (inputs[921]);
    assign layer0_outputs[1034] = inputs[92];
    assign layer0_outputs[1035] = (inputs[1]) ^ (inputs[379]);
    assign layer0_outputs[1036] = ~((inputs[550]) | (inputs[155]));
    assign layer0_outputs[1037] = (inputs[274]) & ~(inputs[153]);
    assign layer0_outputs[1038] = ~(inputs[834]);
    assign layer0_outputs[1039] = (inputs[682]) & ~(inputs[675]);
    assign layer0_outputs[1040] = inputs[546];
    assign layer0_outputs[1041] = inputs[303];
    assign layer0_outputs[1042] = ~(inputs[906]);
    assign layer0_outputs[1043] = ~(inputs[338]) | (inputs[866]);
    assign layer0_outputs[1044] = ~(inputs[587]);
    assign layer0_outputs[1045] = 1'b0;
    assign layer0_outputs[1046] = ~((inputs[574]) & (inputs[229]));
    assign layer0_outputs[1047] = (inputs[1023]) & ~(inputs[1009]);
    assign layer0_outputs[1048] = ~(inputs[942]) | (inputs[646]);
    assign layer0_outputs[1049] = 1'b1;
    assign layer0_outputs[1050] = ~(inputs[266]);
    assign layer0_outputs[1051] = ~(inputs[567]) | (inputs[309]);
    assign layer0_outputs[1052] = (inputs[273]) ^ (inputs[126]);
    assign layer0_outputs[1053] = 1'b0;
    assign layer0_outputs[1054] = (inputs[971]) | (inputs[141]);
    assign layer0_outputs[1055] = ~(inputs[32]) | (inputs[834]);
    assign layer0_outputs[1056] = ~(inputs[317]);
    assign layer0_outputs[1057] = ~(inputs[193]);
    assign layer0_outputs[1058] = ~((inputs[576]) & (inputs[145]));
    assign layer0_outputs[1059] = ~((inputs[66]) ^ (inputs[438]));
    assign layer0_outputs[1060] = ~(inputs[639]);
    assign layer0_outputs[1061] = ~(inputs[824]);
    assign layer0_outputs[1062] = (inputs[653]) & ~(inputs[263]);
    assign layer0_outputs[1063] = (inputs[905]) & ~(inputs[140]);
    assign layer0_outputs[1064] = ~(inputs[613]);
    assign layer0_outputs[1065] = 1'b1;
    assign layer0_outputs[1066] = ~(inputs[633]);
    assign layer0_outputs[1067] = 1'b0;
    assign layer0_outputs[1068] = (inputs[169]) & ~(inputs[771]);
    assign layer0_outputs[1069] = (inputs[587]) & ~(inputs[899]);
    assign layer0_outputs[1070] = ~((inputs[521]) | (inputs[903]));
    assign layer0_outputs[1071] = (inputs[652]) | (inputs[5]);
    assign layer0_outputs[1072] = 1'b1;
    assign layer0_outputs[1073] = (inputs[958]) | (inputs[43]);
    assign layer0_outputs[1074] = ~((inputs[603]) | (inputs[160]));
    assign layer0_outputs[1075] = ~(inputs[32]);
    assign layer0_outputs[1076] = ~(inputs[136]);
    assign layer0_outputs[1077] = (inputs[701]) ^ (inputs[284]);
    assign layer0_outputs[1078] = inputs[867];
    assign layer0_outputs[1079] = ~((inputs[644]) | (inputs[410]));
    assign layer0_outputs[1080] = (inputs[800]) ^ (inputs[740]);
    assign layer0_outputs[1081] = ~((inputs[183]) ^ (inputs[310]));
    assign layer0_outputs[1082] = ~(inputs[175]) | (inputs[313]);
    assign layer0_outputs[1083] = ~(inputs[289]);
    assign layer0_outputs[1084] = (inputs[525]) & ~(inputs[957]);
    assign layer0_outputs[1085] = inputs[812];
    assign layer0_outputs[1086] = inputs[925];
    assign layer0_outputs[1087] = ~((inputs[879]) | (inputs[398]));
    assign layer0_outputs[1088] = ~(inputs[620]);
    assign layer0_outputs[1089] = inputs[397];
    assign layer0_outputs[1090] = ~((inputs[11]) | (inputs[54]));
    assign layer0_outputs[1091] = ~((inputs[609]) ^ (inputs[12]));
    assign layer0_outputs[1092] = (inputs[551]) ^ (inputs[495]);
    assign layer0_outputs[1093] = ~(inputs[668]) | (inputs[449]);
    assign layer0_outputs[1094] = inputs[626];
    assign layer0_outputs[1095] = (inputs[379]) & ~(inputs[273]);
    assign layer0_outputs[1096] = ~((inputs[699]) | (inputs[165]));
    assign layer0_outputs[1097] = inputs[798];
    assign layer0_outputs[1098] = ~(inputs[349]);
    assign layer0_outputs[1099] = (inputs[526]) | (inputs[352]);
    assign layer0_outputs[1100] = ~((inputs[46]) ^ (inputs[636]));
    assign layer0_outputs[1101] = (inputs[751]) ^ (inputs[191]);
    assign layer0_outputs[1102] = (inputs[425]) & ~(inputs[832]);
    assign layer0_outputs[1103] = ~(inputs[387]) | (inputs[99]);
    assign layer0_outputs[1104] = (inputs[88]) | (inputs[461]);
    assign layer0_outputs[1105] = ~(inputs[141]);
    assign layer0_outputs[1106] = (inputs[564]) ^ (inputs[550]);
    assign layer0_outputs[1107] = (inputs[346]) | (inputs[852]);
    assign layer0_outputs[1108] = (inputs[304]) & ~(inputs[351]);
    assign layer0_outputs[1109] = ~((inputs[831]) & (inputs[868]));
    assign layer0_outputs[1110] = inputs[491];
    assign layer0_outputs[1111] = ~((inputs[143]) ^ (inputs[249]));
    assign layer0_outputs[1112] = inputs[1003];
    assign layer0_outputs[1113] = ~(inputs[653]);
    assign layer0_outputs[1114] = ~((inputs[466]) & (inputs[809]));
    assign layer0_outputs[1115] = (inputs[71]) ^ (inputs[108]);
    assign layer0_outputs[1116] = (inputs[178]) & ~(inputs[487]);
    assign layer0_outputs[1117] = (inputs[230]) | (inputs[617]);
    assign layer0_outputs[1118] = ~(inputs[51]);
    assign layer0_outputs[1119] = ~((inputs[627]) ^ (inputs[807]));
    assign layer0_outputs[1120] = ~((inputs[608]) ^ (inputs[963]));
    assign layer0_outputs[1121] = ~((inputs[578]) & (inputs[354]));
    assign layer0_outputs[1122] = (inputs[170]) ^ (inputs[54]);
    assign layer0_outputs[1123] = (inputs[391]) | (inputs[831]);
    assign layer0_outputs[1124] = ~((inputs[936]) | (inputs[770]));
    assign layer0_outputs[1125] = inputs[867];
    assign layer0_outputs[1126] = (inputs[30]) & ~(inputs[33]);
    assign layer0_outputs[1127] = (inputs[847]) | (inputs[425]);
    assign layer0_outputs[1128] = (inputs[252]) | (inputs[455]);
    assign layer0_outputs[1129] = inputs[603];
    assign layer0_outputs[1130] = inputs[358];
    assign layer0_outputs[1131] = inputs[183];
    assign layer0_outputs[1132] = ~((inputs[982]) | (inputs[802]));
    assign layer0_outputs[1133] = ~(inputs[549]);
    assign layer0_outputs[1134] = ~(inputs[625]);
    assign layer0_outputs[1135] = (inputs[368]) ^ (inputs[119]);
    assign layer0_outputs[1136] = ~(inputs[648]);
    assign layer0_outputs[1137] = inputs[177];
    assign layer0_outputs[1138] = (inputs[17]) ^ (inputs[333]);
    assign layer0_outputs[1139] = 1'b1;
    assign layer0_outputs[1140] = ~((inputs[810]) & (inputs[815]));
    assign layer0_outputs[1141] = ~((inputs[937]) ^ (inputs[598]));
    assign layer0_outputs[1142] = ~(inputs[568]) | (inputs[550]);
    assign layer0_outputs[1143] = ~(inputs[342]) | (inputs[170]);
    assign layer0_outputs[1144] = (inputs[414]) & (inputs[963]);
    assign layer0_outputs[1145] = inputs[803];
    assign layer0_outputs[1146] = 1'b0;
    assign layer0_outputs[1147] = (inputs[629]) ^ (inputs[431]);
    assign layer0_outputs[1148] = ~((inputs[369]) | (inputs[326]));
    assign layer0_outputs[1149] = ~((inputs[304]) | (inputs[18]));
    assign layer0_outputs[1150] = (inputs[276]) & ~(inputs[779]);
    assign layer0_outputs[1151] = ~(inputs[750]);
    assign layer0_outputs[1152] = ~(inputs[586]);
    assign layer0_outputs[1153] = (inputs[622]) ^ (inputs[51]);
    assign layer0_outputs[1154] = (inputs[544]) & ~(inputs[928]);
    assign layer0_outputs[1155] = inputs[659];
    assign layer0_outputs[1156] = 1'b1;
    assign layer0_outputs[1157] = ~((inputs[794]) | (inputs[774]));
    assign layer0_outputs[1158] = ~(inputs[95]);
    assign layer0_outputs[1159] = ~(inputs[500]);
    assign layer0_outputs[1160] = (inputs[185]) & ~(inputs[950]);
    assign layer0_outputs[1161] = ~((inputs[648]) | (inputs[885]));
    assign layer0_outputs[1162] = (inputs[717]) ^ (inputs[436]);
    assign layer0_outputs[1163] = ~((inputs[326]) | (inputs[805]));
    assign layer0_outputs[1164] = (inputs[717]) & ~(inputs[259]);
    assign layer0_outputs[1165] = ~((inputs[220]) ^ (inputs[636]));
    assign layer0_outputs[1166] = (inputs[739]) & ~(inputs[647]);
    assign layer0_outputs[1167] = ~(inputs[778]) | (inputs[162]);
    assign layer0_outputs[1168] = (inputs[956]) ^ (inputs[497]);
    assign layer0_outputs[1169] = inputs[217];
    assign layer0_outputs[1170] = ~((inputs[853]) ^ (inputs[739]));
    assign layer0_outputs[1171] = ~(inputs[312]) | (inputs[172]);
    assign layer0_outputs[1172] = ~(inputs[551]) | (inputs[230]);
    assign layer0_outputs[1173] = (inputs[854]) | (inputs[392]);
    assign layer0_outputs[1174] = ~((inputs[700]) | (inputs[736]));
    assign layer0_outputs[1175] = ~((inputs[539]) ^ (inputs[655]));
    assign layer0_outputs[1176] = inputs[347];
    assign layer0_outputs[1177] = ~((inputs[767]) | (inputs[951]));
    assign layer0_outputs[1178] = (inputs[300]) & ~(inputs[599]);
    assign layer0_outputs[1179] = inputs[694];
    assign layer0_outputs[1180] = (inputs[452]) | (inputs[128]);
    assign layer0_outputs[1181] = (inputs[349]) | (inputs[603]);
    assign layer0_outputs[1182] = ~(inputs[781]) | (inputs[803]);
    assign layer0_outputs[1183] = (inputs[452]) ^ (inputs[264]);
    assign layer0_outputs[1184] = (inputs[406]) | (inputs[912]);
    assign layer0_outputs[1185] = ~(inputs[563]) | (inputs[781]);
    assign layer0_outputs[1186] = (inputs[444]) & ~(inputs[287]);
    assign layer0_outputs[1187] = ~((inputs[8]) ^ (inputs[60]));
    assign layer0_outputs[1188] = ~((inputs[271]) ^ (inputs[144]));
    assign layer0_outputs[1189] = 1'b0;
    assign layer0_outputs[1190] = ~(inputs[541]) | (inputs[956]);
    assign layer0_outputs[1191] = ~((inputs[640]) | (inputs[439]));
    assign layer0_outputs[1192] = ~(inputs[429]);
    assign layer0_outputs[1193] = ~(inputs[763]);
    assign layer0_outputs[1194] = (inputs[124]) & ~(inputs[566]);
    assign layer0_outputs[1195] = (inputs[769]) ^ (inputs[844]);
    assign layer0_outputs[1196] = ~(inputs[535]) | (inputs[729]);
    assign layer0_outputs[1197] = (inputs[117]) & ~(inputs[714]);
    assign layer0_outputs[1198] = ~(inputs[556]) | (inputs[266]);
    assign layer0_outputs[1199] = ~(inputs[660]) | (inputs[871]);
    assign layer0_outputs[1200] = (inputs[927]) & (inputs[66]);
    assign layer0_outputs[1201] = (inputs[680]) & ~(inputs[285]);
    assign layer0_outputs[1202] = ~((inputs[810]) | (inputs[779]));
    assign layer0_outputs[1203] = (inputs[792]) & ~(inputs[224]);
    assign layer0_outputs[1204] = (inputs[619]) ^ (inputs[650]);
    assign layer0_outputs[1205] = ~(inputs[881]) | (inputs[200]);
    assign layer0_outputs[1206] = (inputs[238]) | (inputs[142]);
    assign layer0_outputs[1207] = (inputs[828]) & ~(inputs[789]);
    assign layer0_outputs[1208] = ~(inputs[58]) | (inputs[154]);
    assign layer0_outputs[1209] = ~(inputs[307]) | (inputs[324]);
    assign layer0_outputs[1210] = (inputs[748]) | (inputs[369]);
    assign layer0_outputs[1211] = ~(inputs[307]) | (inputs[9]);
    assign layer0_outputs[1212] = inputs[628];
    assign layer0_outputs[1213] = (inputs[894]) ^ (inputs[35]);
    assign layer0_outputs[1214] = ~(inputs[396]);
    assign layer0_outputs[1215] = ~((inputs[614]) | (inputs[382]));
    assign layer0_outputs[1216] = inputs[555];
    assign layer0_outputs[1217] = ~(inputs[525]) | (inputs[859]);
    assign layer0_outputs[1218] = ~(inputs[55]) | (inputs[1023]);
    assign layer0_outputs[1219] = ~(inputs[745]);
    assign layer0_outputs[1220] = ~((inputs[616]) ^ (inputs[140]));
    assign layer0_outputs[1221] = ~(inputs[431]);
    assign layer0_outputs[1222] = (inputs[478]) & (inputs[480]);
    assign layer0_outputs[1223] = ~(inputs[428]);
    assign layer0_outputs[1224] = ~(inputs[248]) | (inputs[958]);
    assign layer0_outputs[1225] = ~(inputs[620]);
    assign layer0_outputs[1226] = (inputs[776]) & ~(inputs[732]);
    assign layer0_outputs[1227] = ~(inputs[822]) | (inputs[1014]);
    assign layer0_outputs[1228] = 1'b0;
    assign layer0_outputs[1229] = (inputs[899]) ^ (inputs[538]);
    assign layer0_outputs[1230] = ~((inputs[453]) & (inputs[296]));
    assign layer0_outputs[1231] = inputs[782];
    assign layer0_outputs[1232] = (inputs[953]) | (inputs[267]);
    assign layer0_outputs[1233] = (inputs[440]) | (inputs[972]);
    assign layer0_outputs[1234] = ~((inputs[307]) | (inputs[90]));
    assign layer0_outputs[1235] = ~((inputs[110]) ^ (inputs[706]));
    assign layer0_outputs[1236] = (inputs[519]) | (inputs[845]);
    assign layer0_outputs[1237] = ~((inputs[534]) | (inputs[892]));
    assign layer0_outputs[1238] = (inputs[872]) ^ (inputs[325]);
    assign layer0_outputs[1239] = (inputs[1001]) ^ (inputs[77]);
    assign layer0_outputs[1240] = (inputs[498]) & ~(inputs[101]);
    assign layer0_outputs[1241] = (inputs[363]) & ~(inputs[133]);
    assign layer0_outputs[1242] = (inputs[657]) | (inputs[979]);
    assign layer0_outputs[1243] = ~(inputs[94]);
    assign layer0_outputs[1244] = ~(inputs[16]);
    assign layer0_outputs[1245] = inputs[252];
    assign layer0_outputs[1246] = (inputs[622]) & ~(inputs[93]);
    assign layer0_outputs[1247] = (inputs[701]) | (inputs[177]);
    assign layer0_outputs[1248] = inputs[399];
    assign layer0_outputs[1249] = ~((inputs[951]) | (inputs[949]));
    assign layer0_outputs[1250] = inputs[810];
    assign layer0_outputs[1251] = ~(inputs[422]);
    assign layer0_outputs[1252] = inputs[691];
    assign layer0_outputs[1253] = (inputs[1015]) & (inputs[166]);
    assign layer0_outputs[1254] = (inputs[630]) | (inputs[745]);
    assign layer0_outputs[1255] = ~(inputs[314]);
    assign layer0_outputs[1256] = inputs[712];
    assign layer0_outputs[1257] = ~(inputs[209]);
    assign layer0_outputs[1258] = ~((inputs[827]) & (inputs[638]));
    assign layer0_outputs[1259] = (inputs[148]) ^ (inputs[357]);
    assign layer0_outputs[1260] = inputs[577];
    assign layer0_outputs[1261] = ~(inputs[402]) | (inputs[544]);
    assign layer0_outputs[1262] = (inputs[32]) | (inputs[821]);
    assign layer0_outputs[1263] = (inputs[665]) | (inputs[236]);
    assign layer0_outputs[1264] = ~(inputs[886]) | (inputs[738]);
    assign layer0_outputs[1265] = ~((inputs[97]) | (inputs[909]));
    assign layer0_outputs[1266] = (inputs[762]) & ~(inputs[75]);
    assign layer0_outputs[1267] = ~(inputs[894]);
    assign layer0_outputs[1268] = (inputs[147]) ^ (inputs[82]);
    assign layer0_outputs[1269] = (inputs[841]) ^ (inputs[324]);
    assign layer0_outputs[1270] = ~((inputs[255]) & (inputs[1016]));
    assign layer0_outputs[1271] = (inputs[855]) & ~(inputs[352]);
    assign layer0_outputs[1272] = (inputs[393]) & ~(inputs[14]);
    assign layer0_outputs[1273] = (inputs[527]) & ~(inputs[354]);
    assign layer0_outputs[1274] = ~(inputs[842]) | (inputs[931]);
    assign layer0_outputs[1275] = ~(inputs[914]);
    assign layer0_outputs[1276] = (inputs[998]) | (inputs[466]);
    assign layer0_outputs[1277] = ~((inputs[643]) & (inputs[484]));
    assign layer0_outputs[1278] = ~((inputs[618]) | (inputs[579]));
    assign layer0_outputs[1279] = ~(inputs[522]) | (inputs[663]);
    assign layer0_outputs[1280] = ~(inputs[817]);
    assign layer0_outputs[1281] = (inputs[519]) ^ (inputs[167]);
    assign layer0_outputs[1282] = ~((inputs[86]) ^ (inputs[977]));
    assign layer0_outputs[1283] = ~(inputs[463]) | (inputs[479]);
    assign layer0_outputs[1284] = ~(inputs[428]);
    assign layer0_outputs[1285] = ~((inputs[46]) ^ (inputs[387]));
    assign layer0_outputs[1286] = ~(inputs[336]);
    assign layer0_outputs[1287] = ~(inputs[595]) | (inputs[641]);
    assign layer0_outputs[1288] = ~(inputs[758]);
    assign layer0_outputs[1289] = ~(inputs[393]);
    assign layer0_outputs[1290] = ~(inputs[585]) | (inputs[1000]);
    assign layer0_outputs[1291] = ~((inputs[901]) & (inputs[39]));
    assign layer0_outputs[1292] = 1'b0;
    assign layer0_outputs[1293] = ~(inputs[845]);
    assign layer0_outputs[1294] = (inputs[206]) ^ (inputs[269]);
    assign layer0_outputs[1295] = (inputs[501]) & ~(inputs[137]);
    assign layer0_outputs[1296] = ~(inputs[494]) | (inputs[10]);
    assign layer0_outputs[1297] = ~((inputs[504]) | (inputs[847]));
    assign layer0_outputs[1298] = inputs[507];
    assign layer0_outputs[1299] = ~(inputs[941]);
    assign layer0_outputs[1300] = inputs[330];
    assign layer0_outputs[1301] = ~((inputs[378]) | (inputs[642]));
    assign layer0_outputs[1302] = ~(inputs[205]) | (inputs[222]);
    assign layer0_outputs[1303] = ~((inputs[77]) | (inputs[295]));
    assign layer0_outputs[1304] = (inputs[955]) | (inputs[998]);
    assign layer0_outputs[1305] = ~(inputs[688]);
    assign layer0_outputs[1306] = (inputs[148]) & ~(inputs[607]);
    assign layer0_outputs[1307] = ~((inputs[701]) ^ (inputs[317]));
    assign layer0_outputs[1308] = ~((inputs[162]) | (inputs[272]));
    assign layer0_outputs[1309] = (inputs[841]) & ~(inputs[572]);
    assign layer0_outputs[1310] = ~((inputs[586]) ^ (inputs[652]));
    assign layer0_outputs[1311] = (inputs[779]) & ~(inputs[923]);
    assign layer0_outputs[1312] = (inputs[194]) ^ (inputs[39]);
    assign layer0_outputs[1313] = ~(inputs[500]) | (inputs[987]);
    assign layer0_outputs[1314] = inputs[984];
    assign layer0_outputs[1315] = ~((inputs[524]) ^ (inputs[484]));
    assign layer0_outputs[1316] = inputs[187];
    assign layer0_outputs[1317] = ~((inputs[999]) ^ (inputs[219]));
    assign layer0_outputs[1318] = ~(inputs[401]);
    assign layer0_outputs[1319] = (inputs[302]) | (inputs[15]);
    assign layer0_outputs[1320] = (inputs[656]) ^ (inputs[738]);
    assign layer0_outputs[1321] = ~(inputs[361]);
    assign layer0_outputs[1322] = (inputs[791]) ^ (inputs[137]);
    assign layer0_outputs[1323] = ~(inputs[224]) | (inputs[75]);
    assign layer0_outputs[1324] = (inputs[533]) & ~(inputs[81]);
    assign layer0_outputs[1325] = ~(inputs[225]) | (inputs[546]);
    assign layer0_outputs[1326] = ~((inputs[170]) | (inputs[448]));
    assign layer0_outputs[1327] = 1'b0;
    assign layer0_outputs[1328] = (inputs[975]) | (inputs[807]);
    assign layer0_outputs[1329] = (inputs[973]) | (inputs[518]);
    assign layer0_outputs[1330] = ~(inputs[370]);
    assign layer0_outputs[1331] = (inputs[621]) & ~(inputs[937]);
    assign layer0_outputs[1332] = (inputs[10]) | (inputs[98]);
    assign layer0_outputs[1333] = (inputs[517]) | (inputs[392]);
    assign layer0_outputs[1334] = inputs[598];
    assign layer0_outputs[1335] = (inputs[237]) ^ (inputs[458]);
    assign layer0_outputs[1336] = (inputs[541]) | (inputs[374]);
    assign layer0_outputs[1337] = ~(inputs[316]);
    assign layer0_outputs[1338] = (inputs[532]) ^ (inputs[708]);
    assign layer0_outputs[1339] = ~((inputs[936]) & (inputs[1016]));
    assign layer0_outputs[1340] = ~((inputs[689]) & (inputs[1012]));
    assign layer0_outputs[1341] = ~(inputs[552]) | (inputs[796]);
    assign layer0_outputs[1342] = ~((inputs[218]) | (inputs[215]));
    assign layer0_outputs[1343] = ~((inputs[436]) | (inputs[1022]));
    assign layer0_outputs[1344] = inputs[301];
    assign layer0_outputs[1345] = (inputs[665]) | (inputs[191]);
    assign layer0_outputs[1346] = ~(inputs[161]);
    assign layer0_outputs[1347] = (inputs[394]) & ~(inputs[833]);
    assign layer0_outputs[1348] = (inputs[558]) & ~(inputs[857]);
    assign layer0_outputs[1349] = (inputs[382]) | (inputs[818]);
    assign layer0_outputs[1350] = (inputs[569]) & ~(inputs[952]);
    assign layer0_outputs[1351] = (inputs[805]) & ~(inputs[709]);
    assign layer0_outputs[1352] = (inputs[617]) ^ (inputs[257]);
    assign layer0_outputs[1353] = (inputs[599]) & ~(inputs[855]);
    assign layer0_outputs[1354] = ~(inputs[622]) | (inputs[136]);
    assign layer0_outputs[1355] = (inputs[312]) & ~(inputs[97]);
    assign layer0_outputs[1356] = (inputs[35]) & ~(inputs[642]);
    assign layer0_outputs[1357] = ~(inputs[713]) | (inputs[978]);
    assign layer0_outputs[1358] = (inputs[877]) & ~(inputs[858]);
    assign layer0_outputs[1359] = (inputs[624]) & ~(inputs[347]);
    assign layer0_outputs[1360] = ~((inputs[169]) | (inputs[372]));
    assign layer0_outputs[1361] = (inputs[91]) ^ (inputs[488]);
    assign layer0_outputs[1362] = (inputs[180]) ^ (inputs[904]);
    assign layer0_outputs[1363] = ~(inputs[550]) | (inputs[31]);
    assign layer0_outputs[1364] = (inputs[693]) & ~(inputs[221]);
    assign layer0_outputs[1365] = ~(inputs[493]) | (inputs[844]);
    assign layer0_outputs[1366] = inputs[1004];
    assign layer0_outputs[1367] = (inputs[327]) | (inputs[1012]);
    assign layer0_outputs[1368] = ~((inputs[748]) | (inputs[552]));
    assign layer0_outputs[1369] = inputs[905];
    assign layer0_outputs[1370] = (inputs[520]) & (inputs[783]);
    assign layer0_outputs[1371] = inputs[757];
    assign layer0_outputs[1372] = (inputs[300]) ^ (inputs[754]);
    assign layer0_outputs[1373] = (inputs[867]) | (inputs[321]);
    assign layer0_outputs[1374] = ~(inputs[559]) | (inputs[27]);
    assign layer0_outputs[1375] = (inputs[275]) & ~(inputs[1005]);
    assign layer0_outputs[1376] = inputs[707];
    assign layer0_outputs[1377] = ~((inputs[280]) ^ (inputs[770]));
    assign layer0_outputs[1378] = (inputs[279]) ^ (inputs[949]);
    assign layer0_outputs[1379] = ~(inputs[66]) | (inputs[921]);
    assign layer0_outputs[1380] = ~((inputs[311]) | (inputs[813]));
    assign layer0_outputs[1381] = ~((inputs[18]) | (inputs[656]));
    assign layer0_outputs[1382] = ~((inputs[434]) ^ (inputs[890]));
    assign layer0_outputs[1383] = (inputs[798]) ^ (inputs[40]);
    assign layer0_outputs[1384] = ~(inputs[935]) | (inputs[160]);
    assign layer0_outputs[1385] = ~((inputs[703]) | (inputs[1014]));
    assign layer0_outputs[1386] = ~((inputs[872]) | (inputs[716]));
    assign layer0_outputs[1387] = ~(inputs[969]) | (inputs[851]);
    assign layer0_outputs[1388] = ~(inputs[284]) | (inputs[4]);
    assign layer0_outputs[1389] = ~((inputs[69]) | (inputs[878]));
    assign layer0_outputs[1390] = (inputs[638]) & (inputs[511]);
    assign layer0_outputs[1391] = ~(inputs[722]) | (inputs[347]);
    assign layer0_outputs[1392] = (inputs[660]) & ~(inputs[733]);
    assign layer0_outputs[1393] = ~((inputs[158]) | (inputs[1016]));
    assign layer0_outputs[1394] = ~((inputs[759]) ^ (inputs[523]));
    assign layer0_outputs[1395] = (inputs[813]) ^ (inputs[928]);
    assign layer0_outputs[1396] = inputs[280];
    assign layer0_outputs[1397] = ~(inputs[570]);
    assign layer0_outputs[1398] = (inputs[116]) & ~(inputs[261]);
    assign layer0_outputs[1399] = ~(inputs[402]) | (inputs[156]);
    assign layer0_outputs[1400] = (inputs[639]) | (inputs[519]);
    assign layer0_outputs[1401] = inputs[212];
    assign layer0_outputs[1402] = ~(inputs[463]);
    assign layer0_outputs[1403] = ~((inputs[346]) | (inputs[494]));
    assign layer0_outputs[1404] = ~(inputs[432]) | (inputs[566]);
    assign layer0_outputs[1405] = ~(inputs[465]) | (inputs[107]);
    assign layer0_outputs[1406] = (inputs[72]) ^ (inputs[639]);
    assign layer0_outputs[1407] = (inputs[40]) & ~(inputs[81]);
    assign layer0_outputs[1408] = inputs[905];
    assign layer0_outputs[1409] = (inputs[247]) | (inputs[513]);
    assign layer0_outputs[1410] = (inputs[222]) & ~(inputs[1011]);
    assign layer0_outputs[1411] = ~((inputs[449]) & (inputs[58]));
    assign layer0_outputs[1412] = (inputs[683]) | (inputs[961]);
    assign layer0_outputs[1413] = ~(inputs[29]);
    assign layer0_outputs[1414] = (inputs[780]) & ~(inputs[409]);
    assign layer0_outputs[1415] = ~((inputs[323]) ^ (inputs[444]));
    assign layer0_outputs[1416] = ~((inputs[414]) | (inputs[664]));
    assign layer0_outputs[1417] = (inputs[280]) | (inputs[996]);
    assign layer0_outputs[1418] = (inputs[543]) & ~(inputs[392]);
    assign layer0_outputs[1419] = (inputs[549]) ^ (inputs[204]);
    assign layer0_outputs[1420] = (inputs[968]) | (inputs[537]);
    assign layer0_outputs[1421] = ~((inputs[279]) | (inputs[36]));
    assign layer0_outputs[1422] = (inputs[217]) ^ (inputs[704]);
    assign layer0_outputs[1423] = (inputs[671]) ^ (inputs[700]);
    assign layer0_outputs[1424] = (inputs[227]) ^ (inputs[829]);
    assign layer0_outputs[1425] = ~((inputs[706]) ^ (inputs[538]));
    assign layer0_outputs[1426] = (inputs[732]) ^ (inputs[506]);
    assign layer0_outputs[1427] = inputs[838];
    assign layer0_outputs[1428] = ~(inputs[258]);
    assign layer0_outputs[1429] = ~(inputs[653]);
    assign layer0_outputs[1430] = ~(inputs[828]);
    assign layer0_outputs[1431] = ~(inputs[631]);
    assign layer0_outputs[1432] = (inputs[752]) & ~(inputs[252]);
    assign layer0_outputs[1433] = 1'b1;
    assign layer0_outputs[1434] = ~(inputs[187]) | (inputs[299]);
    assign layer0_outputs[1435] = ~(inputs[439]);
    assign layer0_outputs[1436] = ~((inputs[779]) ^ (inputs[537]));
    assign layer0_outputs[1437] = ~((inputs[945]) ^ (inputs[560]));
    assign layer0_outputs[1438] = (inputs[164]) & ~(inputs[194]);
    assign layer0_outputs[1439] = ~(inputs[202]);
    assign layer0_outputs[1440] = (inputs[257]) ^ (inputs[332]);
    assign layer0_outputs[1441] = inputs[643];
    assign layer0_outputs[1442] = 1'b0;
    assign layer0_outputs[1443] = (inputs[750]) & ~(inputs[982]);
    assign layer0_outputs[1444] = ~((inputs[793]) | (inputs[906]));
    assign layer0_outputs[1445] = (inputs[635]) & ~(inputs[35]);
    assign layer0_outputs[1446] = (inputs[840]) & (inputs[385]);
    assign layer0_outputs[1447] = inputs[654];
    assign layer0_outputs[1448] = ~((inputs[700]) | (inputs[566]));
    assign layer0_outputs[1449] = ~((inputs[111]) ^ (inputs[233]));
    assign layer0_outputs[1450] = inputs[473];
    assign layer0_outputs[1451] = ~((inputs[203]) | (inputs[621]));
    assign layer0_outputs[1452] = ~(inputs[192]);
    assign layer0_outputs[1453] = (inputs[485]) & ~(inputs[350]);
    assign layer0_outputs[1454] = ~(inputs[711]);
    assign layer0_outputs[1455] = inputs[9];
    assign layer0_outputs[1456] = (inputs[478]) | (inputs[681]);
    assign layer0_outputs[1457] = inputs[717];
    assign layer0_outputs[1458] = ~((inputs[836]) & (inputs[969]));
    assign layer0_outputs[1459] = ~(inputs[298]) | (inputs[475]);
    assign layer0_outputs[1460] = inputs[446];
    assign layer0_outputs[1461] = (inputs[469]) & ~(inputs[691]);
    assign layer0_outputs[1462] = ~(inputs[367]) | (inputs[996]);
    assign layer0_outputs[1463] = ~((inputs[267]) | (inputs[785]));
    assign layer0_outputs[1464] = ~(inputs[487]) | (inputs[255]);
    assign layer0_outputs[1465] = (inputs[77]) ^ (inputs[779]);
    assign layer0_outputs[1466] = ~(inputs[279]);
    assign layer0_outputs[1467] = (inputs[412]) & (inputs[927]);
    assign layer0_outputs[1468] = (inputs[547]) | (inputs[329]);
    assign layer0_outputs[1469] = ~(inputs[91]) | (inputs[1010]);
    assign layer0_outputs[1470] = ~(inputs[1023]);
    assign layer0_outputs[1471] = ~((inputs[669]) | (inputs[152]));
    assign layer0_outputs[1472] = (inputs[946]) | (inputs[104]);
    assign layer0_outputs[1473] = (inputs[296]) & ~(inputs[988]);
    assign layer0_outputs[1474] = ~((inputs[670]) | (inputs[696]));
    assign layer0_outputs[1475] = ~(inputs[559]) | (inputs[78]);
    assign layer0_outputs[1476] = inputs[203];
    assign layer0_outputs[1477] = (inputs[476]) | (inputs[307]);
    assign layer0_outputs[1478] = (inputs[408]) | (inputs[116]);
    assign layer0_outputs[1479] = ~((inputs[393]) | (inputs[564]));
    assign layer0_outputs[1480] = inputs[330];
    assign layer0_outputs[1481] = ~((inputs[373]) ^ (inputs[816]));
    assign layer0_outputs[1482] = inputs[693];
    assign layer0_outputs[1483] = inputs[534];
    assign layer0_outputs[1484] = (inputs[111]) ^ (inputs[559]);
    assign layer0_outputs[1485] = (inputs[476]) & ~(inputs[192]);
    assign layer0_outputs[1486] = ~(inputs[726]);
    assign layer0_outputs[1487] = (inputs[587]) & ~(inputs[814]);
    assign layer0_outputs[1488] = ~((inputs[221]) ^ (inputs[198]));
    assign layer0_outputs[1489] = (inputs[175]) & ~(inputs[283]);
    assign layer0_outputs[1490] = ~((inputs[246]) ^ (inputs[343]));
    assign layer0_outputs[1491] = ~(inputs[488]) | (inputs[699]);
    assign layer0_outputs[1492] = ~((inputs[33]) | (inputs[621]));
    assign layer0_outputs[1493] = inputs[626];
    assign layer0_outputs[1494] = (inputs[420]) ^ (inputs[318]);
    assign layer0_outputs[1495] = ~(inputs[23]);
    assign layer0_outputs[1496] = (inputs[367]) | (inputs[603]);
    assign layer0_outputs[1497] = ~(inputs[874]) | (inputs[139]);
    assign layer0_outputs[1498] = inputs[724];
    assign layer0_outputs[1499] = (inputs[374]) & ~(inputs[667]);
    assign layer0_outputs[1500] = 1'b0;
    assign layer0_outputs[1501] = (inputs[50]) ^ (inputs[798]);
    assign layer0_outputs[1502] = ~(inputs[621]) | (inputs[115]);
    assign layer0_outputs[1503] = ~(inputs[870]) | (inputs[27]);
    assign layer0_outputs[1504] = (inputs[715]) & ~(inputs[133]);
    assign layer0_outputs[1505] = ~((inputs[413]) | (inputs[510]));
    assign layer0_outputs[1506] = ~((inputs[448]) | (inputs[210]));
    assign layer0_outputs[1507] = ~(inputs[493]) | (inputs[1022]);
    assign layer0_outputs[1508] = (inputs[955]) & ~(inputs[945]);
    assign layer0_outputs[1509] = ~((inputs[341]) ^ (inputs[716]));
    assign layer0_outputs[1510] = ~(inputs[794]) | (inputs[31]);
    assign layer0_outputs[1511] = (inputs[687]) | (inputs[311]);
    assign layer0_outputs[1512] = ~(inputs[965]) | (inputs[51]);
    assign layer0_outputs[1513] = ~((inputs[765]) & (inputs[630]));
    assign layer0_outputs[1514] = (inputs[180]) ^ (inputs[695]);
    assign layer0_outputs[1515] = ~(inputs[125]) | (inputs[837]);
    assign layer0_outputs[1516] = ~(inputs[435]);
    assign layer0_outputs[1517] = (inputs[181]) ^ (inputs[516]);
    assign layer0_outputs[1518] = (inputs[471]) ^ (inputs[597]);
    assign layer0_outputs[1519] = (inputs[443]) | (inputs[401]);
    assign layer0_outputs[1520] = inputs[464];
    assign layer0_outputs[1521] = (inputs[713]) & ~(inputs[517]);
    assign layer0_outputs[1522] = (inputs[713]) ^ (inputs[146]);
    assign layer0_outputs[1523] = ~((inputs[396]) & (inputs[521]));
    assign layer0_outputs[1524] = ~(inputs[468]) | (inputs[255]);
    assign layer0_outputs[1525] = ~(inputs[999]);
    assign layer0_outputs[1526] = (inputs[17]) & (inputs[926]);
    assign layer0_outputs[1527] = ~((inputs[106]) | (inputs[635]));
    assign layer0_outputs[1528] = ~(inputs[271]);
    assign layer0_outputs[1529] = ~(inputs[626]);
    assign layer0_outputs[1530] = (inputs[984]) & ~(inputs[609]);
    assign layer0_outputs[1531] = ~(inputs[764]) | (inputs[821]);
    assign layer0_outputs[1532] = ~(inputs[936]);
    assign layer0_outputs[1533] = inputs[488];
    assign layer0_outputs[1534] = 1'b1;
    assign layer0_outputs[1535] = ~(inputs[242]);
    assign layer0_outputs[1536] = (inputs[415]) ^ (inputs[916]);
    assign layer0_outputs[1537] = (inputs[851]) ^ (inputs[1007]);
    assign layer0_outputs[1538] = ~(inputs[298]);
    assign layer0_outputs[1539] = 1'b1;
    assign layer0_outputs[1540] = (inputs[622]) & ~(inputs[668]);
    assign layer0_outputs[1541] = inputs[613];
    assign layer0_outputs[1542] = 1'b1;
    assign layer0_outputs[1543] = ~((inputs[927]) & (inputs[833]));
    assign layer0_outputs[1544] = ~((inputs[520]) ^ (inputs[521]));
    assign layer0_outputs[1545] = ~(inputs[247]);
    assign layer0_outputs[1546] = ~(inputs[711]) | (inputs[926]);
    assign layer0_outputs[1547] = (inputs[554]) & ~(inputs[780]);
    assign layer0_outputs[1548] = ~((inputs[899]) | (inputs[643]));
    assign layer0_outputs[1549] = (inputs[842]) & ~(inputs[902]);
    assign layer0_outputs[1550] = ~((inputs[40]) & (inputs[349]));
    assign layer0_outputs[1551] = ~(inputs[193]) | (inputs[122]);
    assign layer0_outputs[1552] = ~((inputs[859]) ^ (inputs[138]));
    assign layer0_outputs[1553] = inputs[272];
    assign layer0_outputs[1554] = (inputs[155]) | (inputs[865]);
    assign layer0_outputs[1555] = ~((inputs[425]) | (inputs[462]));
    assign layer0_outputs[1556] = (inputs[204]) | (inputs[725]);
    assign layer0_outputs[1557] = ~(inputs[36]) | (inputs[959]);
    assign layer0_outputs[1558] = 1'b0;
    assign layer0_outputs[1559] = ~(inputs[292]) | (inputs[722]);
    assign layer0_outputs[1560] = ~(inputs[848]);
    assign layer0_outputs[1561] = inputs[837];
    assign layer0_outputs[1562] = ~(inputs[86]) | (inputs[925]);
    assign layer0_outputs[1563] = (inputs[484]) | (inputs[401]);
    assign layer0_outputs[1564] = inputs[473];
    assign layer0_outputs[1565] = inputs[215];
    assign layer0_outputs[1566] = ~(inputs[570]) | (inputs[135]);
    assign layer0_outputs[1567] = ~(inputs[9]);
    assign layer0_outputs[1568] = inputs[124];
    assign layer0_outputs[1569] = (inputs[529]) & ~(inputs[172]);
    assign layer0_outputs[1570] = ~(inputs[846]) | (inputs[200]);
    assign layer0_outputs[1571] = ~(inputs[664]) | (inputs[739]);
    assign layer0_outputs[1572] = ~(inputs[594]);
    assign layer0_outputs[1573] = ~(inputs[224]) | (inputs[50]);
    assign layer0_outputs[1574] = ~(inputs[680]);
    assign layer0_outputs[1575] = ~((inputs[114]) & (inputs[678]));
    assign layer0_outputs[1576] = ~(inputs[525]);
    assign layer0_outputs[1577] = ~((inputs[963]) | (inputs[549]));
    assign layer0_outputs[1578] = ~(inputs[183]);
    assign layer0_outputs[1579] = (inputs[545]) ^ (inputs[352]);
    assign layer0_outputs[1580] = ~((inputs[954]) ^ (inputs[958]));
    assign layer0_outputs[1581] = ~(inputs[256]);
    assign layer0_outputs[1582] = (inputs[279]) & ~(inputs[476]);
    assign layer0_outputs[1583] = ~(inputs[328]) | (inputs[126]);
    assign layer0_outputs[1584] = ~(inputs[977]);
    assign layer0_outputs[1585] = 1'b0;
    assign layer0_outputs[1586] = ~(inputs[562]);
    assign layer0_outputs[1587] = ~((inputs[252]) ^ (inputs[451]));
    assign layer0_outputs[1588] = (inputs[98]) & ~(inputs[295]);
    assign layer0_outputs[1589] = ~(inputs[630]) | (inputs[446]);
    assign layer0_outputs[1590] = (inputs[819]) | (inputs[762]);
    assign layer0_outputs[1591] = (inputs[509]) & ~(inputs[675]);
    assign layer0_outputs[1592] = ~((inputs[548]) ^ (inputs[491]));
    assign layer0_outputs[1593] = (inputs[93]) | (inputs[369]);
    assign layer0_outputs[1594] = (inputs[281]) | (inputs[197]);
    assign layer0_outputs[1595] = (inputs[460]) & ~(inputs[977]);
    assign layer0_outputs[1596] = ~((inputs[1]) | (inputs[734]));
    assign layer0_outputs[1597] = (inputs[492]) & ~(inputs[897]);
    assign layer0_outputs[1598] = ~((inputs[584]) | (inputs[218]));
    assign layer0_outputs[1599] = ~(inputs[730]) | (inputs[11]);
    assign layer0_outputs[1600] = ~(inputs[103]);
    assign layer0_outputs[1601] = (inputs[1016]) | (inputs[677]);
    assign layer0_outputs[1602] = ~(inputs[281]) | (inputs[173]);
    assign layer0_outputs[1603] = ~((inputs[466]) | (inputs[694]));
    assign layer0_outputs[1604] = ~(inputs[153]);
    assign layer0_outputs[1605] = ~((inputs[843]) ^ (inputs[10]));
    assign layer0_outputs[1606] = ~((inputs[568]) ^ (inputs[208]));
    assign layer0_outputs[1607] = ~(inputs[457]);
    assign layer0_outputs[1608] = (inputs[858]) ^ (inputs[878]);
    assign layer0_outputs[1609] = ~(inputs[634]);
    assign layer0_outputs[1610] = ~((inputs[304]) | (inputs[893]));
    assign layer0_outputs[1611] = (inputs[633]) & ~(inputs[868]);
    assign layer0_outputs[1612] = ~((inputs[962]) | (inputs[993]));
    assign layer0_outputs[1613] = (inputs[71]) & (inputs[252]);
    assign layer0_outputs[1614] = (inputs[867]) & ~(inputs[23]);
    assign layer0_outputs[1615] = inputs[779];
    assign layer0_outputs[1616] = ~(inputs[823]);
    assign layer0_outputs[1617] = ~(inputs[763]);
    assign layer0_outputs[1618] = inputs[890];
    assign layer0_outputs[1619] = (inputs[509]) & (inputs[578]);
    assign layer0_outputs[1620] = (inputs[295]) ^ (inputs[964]);
    assign layer0_outputs[1621] = (inputs[335]) | (inputs[608]);
    assign layer0_outputs[1622] = ~(inputs[300]);
    assign layer0_outputs[1623] = (inputs[519]) & ~(inputs[980]);
    assign layer0_outputs[1624] = (inputs[571]) | (inputs[564]);
    assign layer0_outputs[1625] = (inputs[879]) | (inputs[894]);
    assign layer0_outputs[1626] = (inputs[835]) & ~(inputs[973]);
    assign layer0_outputs[1627] = (inputs[113]) | (inputs[237]);
    assign layer0_outputs[1628] = ~((inputs[314]) ^ (inputs[128]));
    assign layer0_outputs[1629] = (inputs[544]) ^ (inputs[82]);
    assign layer0_outputs[1630] = inputs[411];
    assign layer0_outputs[1631] = inputs[572];
    assign layer0_outputs[1632] = ~((inputs[484]) | (inputs[932]));
    assign layer0_outputs[1633] = ~((inputs[67]) ^ (inputs[972]));
    assign layer0_outputs[1634] = ~(inputs[817]) | (inputs[70]);
    assign layer0_outputs[1635] = ~(inputs[777]);
    assign layer0_outputs[1636] = ~((inputs[379]) | (inputs[580]));
    assign layer0_outputs[1637] = ~(inputs[430]);
    assign layer0_outputs[1638] = ~(inputs[458]);
    assign layer0_outputs[1639] = ~(inputs[303]);
    assign layer0_outputs[1640] = (inputs[378]) ^ (inputs[299]);
    assign layer0_outputs[1641] = inputs[608];
    assign layer0_outputs[1642] = 1'b0;
    assign layer0_outputs[1643] = (inputs[553]) & ~(inputs[945]);
    assign layer0_outputs[1644] = (inputs[831]) ^ (inputs[490]);
    assign layer0_outputs[1645] = inputs[183];
    assign layer0_outputs[1646] = (inputs[663]) | (inputs[66]);
    assign layer0_outputs[1647] = (inputs[525]) ^ (inputs[536]);
    assign layer0_outputs[1648] = (inputs[598]) & ~(inputs[611]);
    assign layer0_outputs[1649] = ~((inputs[332]) | (inputs[916]));
    assign layer0_outputs[1650] = (inputs[716]) | (inputs[605]);
    assign layer0_outputs[1651] = ~((inputs[721]) ^ (inputs[130]));
    assign layer0_outputs[1652] = (inputs[474]) | (inputs[158]);
    assign layer0_outputs[1653] = inputs[650];
    assign layer0_outputs[1654] = (inputs[759]) | (inputs[980]);
    assign layer0_outputs[1655] = (inputs[774]) & ~(inputs[4]);
    assign layer0_outputs[1656] = (inputs[647]) & ~(inputs[154]);
    assign layer0_outputs[1657] = ~(inputs[499]) | (inputs[959]);
    assign layer0_outputs[1658] = ~((inputs[945]) | (inputs[485]));
    assign layer0_outputs[1659] = ~((inputs[796]) ^ (inputs[340]));
    assign layer0_outputs[1660] = (inputs[100]) | (inputs[618]);
    assign layer0_outputs[1661] = ~((inputs[447]) | (inputs[806]));
    assign layer0_outputs[1662] = ~((inputs[917]) ^ (inputs[66]));
    assign layer0_outputs[1663] = ~((inputs[516]) | (inputs[157]));
    assign layer0_outputs[1664] = inputs[16];
    assign layer0_outputs[1665] = ~(inputs[462]) | (inputs[911]);
    assign layer0_outputs[1666] = ~((inputs[872]) & (inputs[186]));
    assign layer0_outputs[1667] = (inputs[794]) ^ (inputs[104]);
    assign layer0_outputs[1668] = inputs[846];
    assign layer0_outputs[1669] = ~(inputs[282]) | (inputs[681]);
    assign layer0_outputs[1670] = 1'b0;
    assign layer0_outputs[1671] = (inputs[383]) & (inputs[189]);
    assign layer0_outputs[1672] = ~(inputs[947]);
    assign layer0_outputs[1673] = (inputs[163]) | (inputs[65]);
    assign layer0_outputs[1674] = 1'b1;
    assign layer0_outputs[1675] = (inputs[194]) & ~(inputs[1001]);
    assign layer0_outputs[1676] = ~((inputs[235]) ^ (inputs[718]));
    assign layer0_outputs[1677] = (inputs[341]) & ~(inputs[49]);
    assign layer0_outputs[1678] = (inputs[729]) ^ (inputs[233]);
    assign layer0_outputs[1679] = (inputs[742]) | (inputs[817]);
    assign layer0_outputs[1680] = ~(inputs[337]) | (inputs[605]);
    assign layer0_outputs[1681] = inputs[750];
    assign layer0_outputs[1682] = 1'b1;
    assign layer0_outputs[1683] = ~(inputs[427]);
    assign layer0_outputs[1684] = (inputs[148]) & ~(inputs[40]);
    assign layer0_outputs[1685] = (inputs[689]) & ~(inputs[765]);
    assign layer0_outputs[1686] = inputs[403];
    assign layer0_outputs[1687] = ~(inputs[625]) | (inputs[394]);
    assign layer0_outputs[1688] = 1'b1;
    assign layer0_outputs[1689] = ~(inputs[408]) | (inputs[928]);
    assign layer0_outputs[1690] = (inputs[113]) & ~(inputs[987]);
    assign layer0_outputs[1691] = ~(inputs[492]);
    assign layer0_outputs[1692] = ~(inputs[621]);
    assign layer0_outputs[1693] = ~((inputs[828]) | (inputs[561]));
    assign layer0_outputs[1694] = ~((inputs[391]) | (inputs[228]));
    assign layer0_outputs[1695] = ~(inputs[757]);
    assign layer0_outputs[1696] = (inputs[177]) ^ (inputs[922]);
    assign layer0_outputs[1697] = (inputs[819]) & ~(inputs[645]);
    assign layer0_outputs[1698] = ~(inputs[494]);
    assign layer0_outputs[1699] = ~((inputs[306]) | (inputs[406]));
    assign layer0_outputs[1700] = inputs[278];
    assign layer0_outputs[1701] = (inputs[49]) | (inputs[86]);
    assign layer0_outputs[1702] = (inputs[209]) | (inputs[54]);
    assign layer0_outputs[1703] = (inputs[731]) & ~(inputs[160]);
    assign layer0_outputs[1704] = (inputs[754]) ^ (inputs[819]);
    assign layer0_outputs[1705] = (inputs[265]) | (inputs[757]);
    assign layer0_outputs[1706] = ~((inputs[910]) ^ (inputs[903]));
    assign layer0_outputs[1707] = (inputs[946]) | (inputs[153]);
    assign layer0_outputs[1708] = 1'b0;
    assign layer0_outputs[1709] = ~((inputs[198]) ^ (inputs[311]));
    assign layer0_outputs[1710] = ~((inputs[507]) ^ (inputs[693]));
    assign layer0_outputs[1711] = (inputs[334]) | (inputs[61]);
    assign layer0_outputs[1712] = inputs[215];
    assign layer0_outputs[1713] = (inputs[298]) ^ (inputs[38]);
    assign layer0_outputs[1714] = ~((inputs[216]) ^ (inputs[719]));
    assign layer0_outputs[1715] = ~((inputs[404]) | (inputs[417]));
    assign layer0_outputs[1716] = (inputs[660]) | (inputs[105]);
    assign layer0_outputs[1717] = (inputs[942]) & ~(inputs[74]);
    assign layer0_outputs[1718] = (inputs[782]) ^ (inputs[201]);
    assign layer0_outputs[1719] = ~(inputs[297]);
    assign layer0_outputs[1720] = ~(inputs[492]);
    assign layer0_outputs[1721] = ~(inputs[700]);
    assign layer0_outputs[1722] = ~(inputs[590]) | (inputs[547]);
    assign layer0_outputs[1723] = inputs[661];
    assign layer0_outputs[1724] = ~(inputs[859]);
    assign layer0_outputs[1725] = inputs[247];
    assign layer0_outputs[1726] = ~(inputs[936]) | (inputs[71]);
    assign layer0_outputs[1727] = (inputs[242]) & ~(inputs[151]);
    assign layer0_outputs[1728] = inputs[428];
    assign layer0_outputs[1729] = ~(inputs[653]) | (inputs[687]);
    assign layer0_outputs[1730] = (inputs[565]) & ~(inputs[212]);
    assign layer0_outputs[1731] = (inputs[770]) & ~(inputs[230]);
    assign layer0_outputs[1732] = inputs[818];
    assign layer0_outputs[1733] = (inputs[806]) & ~(inputs[1007]);
    assign layer0_outputs[1734] = (inputs[628]) ^ (inputs[761]);
    assign layer0_outputs[1735] = (inputs[18]) ^ (inputs[698]);
    assign layer0_outputs[1736] = ~(inputs[847]);
    assign layer0_outputs[1737] = ~((inputs[496]) | (inputs[912]));
    assign layer0_outputs[1738] = (inputs[831]) & ~(inputs[124]);
    assign layer0_outputs[1739] = (inputs[351]) & ~(inputs[160]);
    assign layer0_outputs[1740] = (inputs[667]) ^ (inputs[383]);
    assign layer0_outputs[1741] = (inputs[82]) ^ (inputs[203]);
    assign layer0_outputs[1742] = ~(inputs[910]);
    assign layer0_outputs[1743] = (inputs[531]) | (inputs[19]);
    assign layer0_outputs[1744] = inputs[94];
    assign layer0_outputs[1745] = inputs[538];
    assign layer0_outputs[1746] = inputs[551];
    assign layer0_outputs[1747] = ~(inputs[827]) | (inputs[388]);
    assign layer0_outputs[1748] = inputs[720];
    assign layer0_outputs[1749] = ~((inputs[924]) & (inputs[309]));
    assign layer0_outputs[1750] = inputs[919];
    assign layer0_outputs[1751] = ~(inputs[491]) | (inputs[572]);
    assign layer0_outputs[1752] = ~((inputs[177]) | (inputs[601]));
    assign layer0_outputs[1753] = ~((inputs[604]) | (inputs[303]));
    assign layer0_outputs[1754] = 1'b1;
    assign layer0_outputs[1755] = ~((inputs[770]) & (inputs[372]));
    assign layer0_outputs[1756] = ~((inputs[130]) ^ (inputs[776]));
    assign layer0_outputs[1757] = ~(inputs[601]);
    assign layer0_outputs[1758] = inputs[854];
    assign layer0_outputs[1759] = ~((inputs[897]) | (inputs[433]));
    assign layer0_outputs[1760] = (inputs[289]) ^ (inputs[453]);
    assign layer0_outputs[1761] = inputs[656];
    assign layer0_outputs[1762] = ~(inputs[269]);
    assign layer0_outputs[1763] = (inputs[842]) & ~(inputs[766]);
    assign layer0_outputs[1764] = inputs[776];
    assign layer0_outputs[1765] = (inputs[756]) ^ (inputs[380]);
    assign layer0_outputs[1766] = 1'b0;
    assign layer0_outputs[1767] = ~((inputs[258]) | (inputs[926]));
    assign layer0_outputs[1768] = ~(inputs[908]) | (inputs[414]);
    assign layer0_outputs[1769] = ~((inputs[580]) | (inputs[821]));
    assign layer0_outputs[1770] = (inputs[503]) ^ (inputs[667]);
    assign layer0_outputs[1771] = (inputs[473]) | (inputs[159]);
    assign layer0_outputs[1772] = ~((inputs[138]) | (inputs[647]));
    assign layer0_outputs[1773] = (inputs[824]) & ~(inputs[117]);
    assign layer0_outputs[1774] = ~((inputs[171]) | (inputs[716]));
    assign layer0_outputs[1775] = (inputs[970]) | (inputs[306]);
    assign layer0_outputs[1776] = ~(inputs[469]) | (inputs[87]);
    assign layer0_outputs[1777] = ~(inputs[245]);
    assign layer0_outputs[1778] = (inputs[553]) | (inputs[569]);
    assign layer0_outputs[1779] = ~(inputs[848]) | (inputs[126]);
    assign layer0_outputs[1780] = ~(inputs[239]);
    assign layer0_outputs[1781] = ~(inputs[775]) | (inputs[923]);
    assign layer0_outputs[1782] = ~(inputs[239]) | (inputs[95]);
    assign layer0_outputs[1783] = inputs[178];
    assign layer0_outputs[1784] = ~(inputs[536]) | (inputs[44]);
    assign layer0_outputs[1785] = (inputs[462]) & ~(inputs[566]);
    assign layer0_outputs[1786] = ~((inputs[951]) ^ (inputs[1007]));
    assign layer0_outputs[1787] = (inputs[831]) | (inputs[334]);
    assign layer0_outputs[1788] = inputs[576];
    assign layer0_outputs[1789] = ~(inputs[463]) | (inputs[488]);
    assign layer0_outputs[1790] = (inputs[955]) & (inputs[1017]);
    assign layer0_outputs[1791] = ~(inputs[247]);
    assign layer0_outputs[1792] = ~((inputs[426]) | (inputs[721]));
    assign layer0_outputs[1793] = (inputs[721]) | (inputs[785]);
    assign layer0_outputs[1794] = (inputs[38]) ^ (inputs[477]);
    assign layer0_outputs[1795] = inputs[362];
    assign layer0_outputs[1796] = inputs[188];
    assign layer0_outputs[1797] = ~(inputs[293]);
    assign layer0_outputs[1798] = inputs[811];
    assign layer0_outputs[1799] = ~(inputs[712]);
    assign layer0_outputs[1800] = ~(inputs[212]) | (inputs[539]);
    assign layer0_outputs[1801] = ~(inputs[561]) | (inputs[665]);
    assign layer0_outputs[1802] = ~((inputs[984]) ^ (inputs[165]));
    assign layer0_outputs[1803] = (inputs[581]) | (inputs[104]);
    assign layer0_outputs[1804] = ~((inputs[842]) | (inputs[23]));
    assign layer0_outputs[1805] = (inputs[73]) | (inputs[345]);
    assign layer0_outputs[1806] = (inputs[863]) & ~(inputs[868]);
    assign layer0_outputs[1807] = inputs[386];
    assign layer0_outputs[1808] = (inputs[687]) | (inputs[204]);
    assign layer0_outputs[1809] = inputs[805];
    assign layer0_outputs[1810] = ~(inputs[501]) | (inputs[917]);
    assign layer0_outputs[1811] = 1'b1;
    assign layer0_outputs[1812] = (inputs[395]) & ~(inputs[738]);
    assign layer0_outputs[1813] = ~(inputs[42]);
    assign layer0_outputs[1814] = (inputs[497]) ^ (inputs[321]);
    assign layer0_outputs[1815] = inputs[1000];
    assign layer0_outputs[1816] = (inputs[251]) & ~(inputs[174]);
    assign layer0_outputs[1817] = ~(inputs[651]) | (inputs[69]);
    assign layer0_outputs[1818] = ~(inputs[506]) | (inputs[524]);
    assign layer0_outputs[1819] = ~((inputs[5]) | (inputs[210]));
    assign layer0_outputs[1820] = ~((inputs[766]) ^ (inputs[371]));
    assign layer0_outputs[1821] = ~(inputs[308]);
    assign layer0_outputs[1822] = (inputs[307]) & ~(inputs[130]);
    assign layer0_outputs[1823] = ~(inputs[10]);
    assign layer0_outputs[1824] = 1'b1;
    assign layer0_outputs[1825] = ~(inputs[557]);
    assign layer0_outputs[1826] = ~((inputs[833]) & (inputs[703]));
    assign layer0_outputs[1827] = (inputs[799]) & ~(inputs[571]);
    assign layer0_outputs[1828] = (inputs[541]) & ~(inputs[920]);
    assign layer0_outputs[1829] = 1'b0;
    assign layer0_outputs[1830] = ~(inputs[279]);
    assign layer0_outputs[1831] = ~(inputs[875]) | (inputs[666]);
    assign layer0_outputs[1832] = ~(inputs[250]) | (inputs[702]);
    assign layer0_outputs[1833] = ~(inputs[408]) | (inputs[919]);
    assign layer0_outputs[1834] = ~((inputs[375]) ^ (inputs[596]));
    assign layer0_outputs[1835] = inputs[930];
    assign layer0_outputs[1836] = ~(inputs[563]);
    assign layer0_outputs[1837] = ~((inputs[950]) & (inputs[287]));
    assign layer0_outputs[1838] = inputs[400];
    assign layer0_outputs[1839] = inputs[156];
    assign layer0_outputs[1840] = ~((inputs[263]) | (inputs[683]));
    assign layer0_outputs[1841] = inputs[1];
    assign layer0_outputs[1842] = ~((inputs[668]) | (inputs[652]));
    assign layer0_outputs[1843] = ~(inputs[497]);
    assign layer0_outputs[1844] = inputs[434];
    assign layer0_outputs[1845] = ~(inputs[283]);
    assign layer0_outputs[1846] = ~((inputs[978]) & (inputs[640]));
    assign layer0_outputs[1847] = ~(inputs[136]);
    assign layer0_outputs[1848] = ~((inputs[1004]) ^ (inputs[333]));
    assign layer0_outputs[1849] = (inputs[209]) ^ (inputs[368]);
    assign layer0_outputs[1850] = ~((inputs[239]) & (inputs[199]));
    assign layer0_outputs[1851] = ~(inputs[914]) | (inputs[280]);
    assign layer0_outputs[1852] = (inputs[276]) & ~(inputs[87]);
    assign layer0_outputs[1853] = (inputs[473]) | (inputs[853]);
    assign layer0_outputs[1854] = 1'b0;
    assign layer0_outputs[1855] = (inputs[985]) | (inputs[388]);
    assign layer0_outputs[1856] = ~(inputs[915]);
    assign layer0_outputs[1857] = 1'b0;
    assign layer0_outputs[1858] = (inputs[466]) & ~(inputs[923]);
    assign layer0_outputs[1859] = ~((inputs[839]) | (inputs[63]));
    assign layer0_outputs[1860] = (inputs[48]) & ~(inputs[92]);
    assign layer0_outputs[1861] = ~((inputs[186]) ^ (inputs[487]));
    assign layer0_outputs[1862] = (inputs[849]) & ~(inputs[263]);
    assign layer0_outputs[1863] = ~(inputs[335]) | (inputs[911]);
    assign layer0_outputs[1864] = (inputs[34]) & ~(inputs[936]);
    assign layer0_outputs[1865] = ~(inputs[33]);
    assign layer0_outputs[1866] = (inputs[488]) & ~(inputs[260]);
    assign layer0_outputs[1867] = ~(inputs[619]);
    assign layer0_outputs[1868] = ~((inputs[888]) | (inputs[495]));
    assign layer0_outputs[1869] = (inputs[632]) & ~(inputs[823]);
    assign layer0_outputs[1870] = ~((inputs[435]) | (inputs[967]));
    assign layer0_outputs[1871] = ~(inputs[907]) | (inputs[1012]);
    assign layer0_outputs[1872] = ~(inputs[718]);
    assign layer0_outputs[1873] = inputs[520];
    assign layer0_outputs[1874] = ~(inputs[402]);
    assign layer0_outputs[1875] = inputs[219];
    assign layer0_outputs[1876] = (inputs[377]) & ~(inputs[626]);
    assign layer0_outputs[1877] = 1'b1;
    assign layer0_outputs[1878] = (inputs[936]) | (inputs[337]);
    assign layer0_outputs[1879] = (inputs[179]) ^ (inputs[189]);
    assign layer0_outputs[1880] = (inputs[156]) & (inputs[31]);
    assign layer0_outputs[1881] = ~(inputs[819]) | (inputs[973]);
    assign layer0_outputs[1882] = ~((inputs[459]) ^ (inputs[382]));
    assign layer0_outputs[1883] = inputs[526];
    assign layer0_outputs[1884] = (inputs[672]) | (inputs[632]);
    assign layer0_outputs[1885] = ~((inputs[209]) | (inputs[150]));
    assign layer0_outputs[1886] = ~(inputs[491]);
    assign layer0_outputs[1887] = (inputs[171]) ^ (inputs[951]);
    assign layer0_outputs[1888] = ~((inputs[23]) ^ (inputs[190]));
    assign layer0_outputs[1889] = ~(inputs[116]) | (inputs[110]);
    assign layer0_outputs[1890] = ~((inputs[367]) | (inputs[405]));
    assign layer0_outputs[1891] = ~(inputs[495]);
    assign layer0_outputs[1892] = ~(inputs[294]) | (inputs[512]);
    assign layer0_outputs[1893] = ~((inputs[453]) | (inputs[244]));
    assign layer0_outputs[1894] = (inputs[336]) & ~(inputs[853]);
    assign layer0_outputs[1895] = ~((inputs[125]) & (inputs[293]));
    assign layer0_outputs[1896] = inputs[995];
    assign layer0_outputs[1897] = (inputs[272]) & ~(inputs[865]);
    assign layer0_outputs[1898] = ~(inputs[453]) | (inputs[45]);
    assign layer0_outputs[1899] = ~(inputs[999]) | (inputs[61]);
    assign layer0_outputs[1900] = (inputs[748]) & ~(inputs[901]);
    assign layer0_outputs[1901] = ~(inputs[785]);
    assign layer0_outputs[1902] = (inputs[405]) ^ (inputs[448]);
    assign layer0_outputs[1903] = ~((inputs[401]) ^ (inputs[374]));
    assign layer0_outputs[1904] = ~((inputs[784]) | (inputs[828]));
    assign layer0_outputs[1905] = (inputs[268]) | (inputs[910]);
    assign layer0_outputs[1906] = (inputs[187]) | (inputs[626]);
    assign layer0_outputs[1907] = ~(inputs[562]);
    assign layer0_outputs[1908] = ~(inputs[562]);
    assign layer0_outputs[1909] = 1'b0;
    assign layer0_outputs[1910] = 1'b1;
    assign layer0_outputs[1911] = ~(inputs[896]) | (inputs[697]);
    assign layer0_outputs[1912] = ~((inputs[126]) | (inputs[379]));
    assign layer0_outputs[1913] = ~(inputs[418]) | (inputs[484]);
    assign layer0_outputs[1914] = inputs[253];
    assign layer0_outputs[1915] = ~((inputs[154]) | (inputs[396]));
    assign layer0_outputs[1916] = (inputs[435]) & ~(inputs[110]);
    assign layer0_outputs[1917] = ~((inputs[673]) ^ (inputs[368]));
    assign layer0_outputs[1918] = (inputs[299]) & ~(inputs[19]);
    assign layer0_outputs[1919] = inputs[822];
    assign layer0_outputs[1920] = (inputs[196]) ^ (inputs[724]);
    assign layer0_outputs[1921] = ~(inputs[534]);
    assign layer0_outputs[1922] = (inputs[261]) | (inputs[313]);
    assign layer0_outputs[1923] = inputs[323];
    assign layer0_outputs[1924] = inputs[423];
    assign layer0_outputs[1925] = ~(inputs[253]) | (inputs[41]);
    assign layer0_outputs[1926] = (inputs[942]) & ~(inputs[92]);
    assign layer0_outputs[1927] = (inputs[400]) | (inputs[192]);
    assign layer0_outputs[1928] = ~((inputs[133]) | (inputs[18]));
    assign layer0_outputs[1929] = inputs[837];
    assign layer0_outputs[1930] = (inputs[723]) & ~(inputs[538]);
    assign layer0_outputs[1931] = (inputs[599]) | (inputs[155]);
    assign layer0_outputs[1932] = inputs[593];
    assign layer0_outputs[1933] = ~((inputs[453]) | (inputs[246]));
    assign layer0_outputs[1934] = inputs[726];
    assign layer0_outputs[1935] = ~(inputs[12]) | (inputs[667]);
    assign layer0_outputs[1936] = (inputs[627]) & ~(inputs[380]);
    assign layer0_outputs[1937] = ~(inputs[537]);
    assign layer0_outputs[1938] = (inputs[585]) & ~(inputs[572]);
    assign layer0_outputs[1939] = 1'b0;
    assign layer0_outputs[1940] = ~((inputs[1021]) | (inputs[957]));
    assign layer0_outputs[1941] = ~((inputs[739]) ^ (inputs[354]));
    assign layer0_outputs[1942] = (inputs[625]) & ~(inputs[983]);
    assign layer0_outputs[1943] = inputs[799];
    assign layer0_outputs[1944] = (inputs[491]) | (inputs[22]);
    assign layer0_outputs[1945] = ~(inputs[48]) | (inputs[767]);
    assign layer0_outputs[1946] = (inputs[274]) | (inputs[13]);
    assign layer0_outputs[1947] = (inputs[239]) & ~(inputs[615]);
    assign layer0_outputs[1948] = inputs[666];
    assign layer0_outputs[1949] = ~(inputs[623]);
    assign layer0_outputs[1950] = (inputs[692]) | (inputs[215]);
    assign layer0_outputs[1951] = (inputs[727]) & ~(inputs[928]);
    assign layer0_outputs[1952] = ~((inputs[338]) | (inputs[637]));
    assign layer0_outputs[1953] = (inputs[163]) ^ (inputs[504]);
    assign layer0_outputs[1954] = (inputs[806]) ^ (inputs[726]);
    assign layer0_outputs[1955] = (inputs[453]) & ~(inputs[419]);
    assign layer0_outputs[1956] = ~(inputs[902]) | (inputs[513]);
    assign layer0_outputs[1957] = 1'b0;
    assign layer0_outputs[1958] = (inputs[694]) & ~(inputs[689]);
    assign layer0_outputs[1959] = (inputs[525]) | (inputs[994]);
    assign layer0_outputs[1960] = ~((inputs[583]) | (inputs[604]));
    assign layer0_outputs[1961] = (inputs[627]) & ~(inputs[284]);
    assign layer0_outputs[1962] = inputs[262];
    assign layer0_outputs[1963] = inputs[434];
    assign layer0_outputs[1964] = (inputs[296]) ^ (inputs[83]);
    assign layer0_outputs[1965] = (inputs[498]) & ~(inputs[771]);
    assign layer0_outputs[1966] = 1'b0;
    assign layer0_outputs[1967] = (inputs[213]) & ~(inputs[165]);
    assign layer0_outputs[1968] = ~((inputs[634]) | (inputs[192]));
    assign layer0_outputs[1969] = ~(inputs[1006]);
    assign layer0_outputs[1970] = (inputs[742]) & (inputs[139]);
    assign layer0_outputs[1971] = (inputs[417]) & (inputs[191]);
    assign layer0_outputs[1972] = (inputs[658]) & ~(inputs[9]);
    assign layer0_outputs[1973] = (inputs[206]) & ~(inputs[901]);
    assign layer0_outputs[1974] = ~(inputs[245]);
    assign layer0_outputs[1975] = inputs[539];
    assign layer0_outputs[1976] = ~(inputs[819]) | (inputs[51]);
    assign layer0_outputs[1977] = inputs[530];
    assign layer0_outputs[1978] = ~(inputs[1008]) | (inputs[635]);
    assign layer0_outputs[1979] = ~(inputs[177]) | (inputs[939]);
    assign layer0_outputs[1980] = ~(inputs[716]);
    assign layer0_outputs[1981] = inputs[906];
    assign layer0_outputs[1982] = inputs[901];
    assign layer0_outputs[1983] = ~((inputs[244]) & (inputs[375]));
    assign layer0_outputs[1984] = ~(inputs[364]);
    assign layer0_outputs[1985] = ~(inputs[753]);
    assign layer0_outputs[1986] = (inputs[956]) | (inputs[504]);
    assign layer0_outputs[1987] = (inputs[339]) ^ (inputs[888]);
    assign layer0_outputs[1988] = (inputs[887]) & ~(inputs[905]);
    assign layer0_outputs[1989] = (inputs[729]) | (inputs[723]);
    assign layer0_outputs[1990] = ~((inputs[230]) | (inputs[963]));
    assign layer0_outputs[1991] = ~(inputs[943]);
    assign layer0_outputs[1992] = ~(inputs[422]) | (inputs[546]);
    assign layer0_outputs[1993] = ~(inputs[500]);
    assign layer0_outputs[1994] = ~((inputs[308]) ^ (inputs[51]));
    assign layer0_outputs[1995] = ~(inputs[472]);
    assign layer0_outputs[1996] = (inputs[746]) & ~(inputs[227]);
    assign layer0_outputs[1997] = inputs[809];
    assign layer0_outputs[1998] = (inputs[351]) & ~(inputs[893]);
    assign layer0_outputs[1999] = ~((inputs[946]) | (inputs[833]));
    assign layer0_outputs[2000] = inputs[104];
    assign layer0_outputs[2001] = ~(inputs[555]) | (inputs[545]);
    assign layer0_outputs[2002] = ~((inputs[998]) ^ (inputs[811]));
    assign layer0_outputs[2003] = ~((inputs[576]) | (inputs[820]));
    assign layer0_outputs[2004] = ~((inputs[159]) & (inputs[161]));
    assign layer0_outputs[2005] = ~((inputs[763]) | (inputs[373]));
    assign layer0_outputs[2006] = ~(inputs[526]);
    assign layer0_outputs[2007] = inputs[383];
    assign layer0_outputs[2008] = (inputs[104]) & ~(inputs[34]);
    assign layer0_outputs[2009] = ~((inputs[211]) | (inputs[212]));
    assign layer0_outputs[2010] = ~((inputs[665]) ^ (inputs[318]));
    assign layer0_outputs[2011] = (inputs[841]) & ~(inputs[1001]);
    assign layer0_outputs[2012] = ~((inputs[337]) | (inputs[73]));
    assign layer0_outputs[2013] = (inputs[909]) & ~(inputs[288]);
    assign layer0_outputs[2014] = ~(inputs[653]);
    assign layer0_outputs[2015] = inputs[409];
    assign layer0_outputs[2016] = ~(inputs[944]);
    assign layer0_outputs[2017] = (inputs[367]) | (inputs[411]);
    assign layer0_outputs[2018] = ~(inputs[59]) | (inputs[66]);
    assign layer0_outputs[2019] = (inputs[469]) & ~(inputs[158]);
    assign layer0_outputs[2020] = (inputs[569]) ^ (inputs[219]);
    assign layer0_outputs[2021] = (inputs[137]) ^ (inputs[208]);
    assign layer0_outputs[2022] = ~(inputs[913]);
    assign layer0_outputs[2023] = inputs[708];
    assign layer0_outputs[2024] = ~(inputs[120]) | (inputs[956]);
    assign layer0_outputs[2025] = ~(inputs[744]);
    assign layer0_outputs[2026] = inputs[449];
    assign layer0_outputs[2027] = inputs[305];
    assign layer0_outputs[2028] = ~(inputs[203]) | (inputs[332]);
    assign layer0_outputs[2029] = inputs[1001];
    assign layer0_outputs[2030] = 1'b1;
    assign layer0_outputs[2031] = inputs[649];
    assign layer0_outputs[2032] = (inputs[520]) | (inputs[132]);
    assign layer0_outputs[2033] = ~(inputs[650]);
    assign layer0_outputs[2034] = ~(inputs[1012]);
    assign layer0_outputs[2035] = ~((inputs[588]) ^ (inputs[830]));
    assign layer0_outputs[2036] = 1'b1;
    assign layer0_outputs[2037] = inputs[694];
    assign layer0_outputs[2038] = (inputs[528]) | (inputs[450]);
    assign layer0_outputs[2039] = (inputs[433]) & ~(inputs[28]);
    assign layer0_outputs[2040] = inputs[159];
    assign layer0_outputs[2041] = ~((inputs[86]) | (inputs[98]));
    assign layer0_outputs[2042] = (inputs[460]) & ~(inputs[448]);
    assign layer0_outputs[2043] = ~((inputs[788]) | (inputs[268]));
    assign layer0_outputs[2044] = (inputs[440]) & ~(inputs[795]);
    assign layer0_outputs[2045] = ~((inputs[699]) | (inputs[417]));
    assign layer0_outputs[2046] = ~(inputs[986]) | (inputs[354]);
    assign layer0_outputs[2047] = ~(inputs[249]);
    assign layer0_outputs[2048] = (inputs[485]) & ~(inputs[731]);
    assign layer0_outputs[2049] = ~((inputs[310]) | (inputs[989]));
    assign layer0_outputs[2050] = inputs[461];
    assign layer0_outputs[2051] = ~(inputs[523]) | (inputs[1001]);
    assign layer0_outputs[2052] = ~(inputs[305]);
    assign layer0_outputs[2053] = ~(inputs[274]);
    assign layer0_outputs[2054] = (inputs[470]) | (inputs[143]);
    assign layer0_outputs[2055] = ~((inputs[592]) | (inputs[82]));
    assign layer0_outputs[2056] = ~(inputs[896]) | (inputs[672]);
    assign layer0_outputs[2057] = ~(inputs[289]);
    assign layer0_outputs[2058] = ~(inputs[716]);
    assign layer0_outputs[2059] = ~((inputs[956]) | (inputs[878]));
    assign layer0_outputs[2060] = inputs[932];
    assign layer0_outputs[2061] = (inputs[952]) & ~(inputs[29]);
    assign layer0_outputs[2062] = (inputs[505]) | (inputs[220]);
    assign layer0_outputs[2063] = ~((inputs[573]) ^ (inputs[554]));
    assign layer0_outputs[2064] = inputs[56];
    assign layer0_outputs[2065] = (inputs[375]) | (inputs[930]);
    assign layer0_outputs[2066] = 1'b0;
    assign layer0_outputs[2067] = ~(inputs[320]) | (inputs[851]);
    assign layer0_outputs[2068] = ~((inputs[5]) ^ (inputs[467]));
    assign layer0_outputs[2069] = (inputs[226]) & (inputs[44]);
    assign layer0_outputs[2070] = inputs[1010];
    assign layer0_outputs[2071] = ~(inputs[357]) | (inputs[414]);
    assign layer0_outputs[2072] = (inputs[938]) ^ (inputs[575]);
    assign layer0_outputs[2073] = ~((inputs[981]) | (inputs[921]));
    assign layer0_outputs[2074] = ~((inputs[860]) | (inputs[501]));
    assign layer0_outputs[2075] = ~(inputs[145]);
    assign layer0_outputs[2076] = ~((inputs[429]) | (inputs[512]));
    assign layer0_outputs[2077] = ~(inputs[562]);
    assign layer0_outputs[2078] = ~(inputs[310]);
    assign layer0_outputs[2079] = ~(inputs[499]) | (inputs[432]);
    assign layer0_outputs[2080] = (inputs[285]) & ~(inputs[764]);
    assign layer0_outputs[2081] = inputs[779];
    assign layer0_outputs[2082] = ~(inputs[703]);
    assign layer0_outputs[2083] = inputs[589];
    assign layer0_outputs[2084] = ~((inputs[401]) | (inputs[642]));
    assign layer0_outputs[2085] = inputs[317];
    assign layer0_outputs[2086] = ~(inputs[172]) | (inputs[3]);
    assign layer0_outputs[2087] = 1'b1;
    assign layer0_outputs[2088] = 1'b1;
    assign layer0_outputs[2089] = ~(inputs[498]) | (inputs[985]);
    assign layer0_outputs[2090] = ~((inputs[366]) & (inputs[90]));
    assign layer0_outputs[2091] = (inputs[78]) ^ (inputs[208]);
    assign layer0_outputs[2092] = ~(inputs[16]);
    assign layer0_outputs[2093] = ~(inputs[282]) | (inputs[189]);
    assign layer0_outputs[2094] = inputs[278];
    assign layer0_outputs[2095] = (inputs[279]) ^ (inputs[989]);
    assign layer0_outputs[2096] = ~(inputs[634]) | (inputs[881]);
    assign layer0_outputs[2097] = (inputs[708]) | (inputs[678]);
    assign layer0_outputs[2098] = inputs[507];
    assign layer0_outputs[2099] = ~(inputs[540]) | (inputs[69]);
    assign layer0_outputs[2100] = ~(inputs[614]) | (inputs[514]);
    assign layer0_outputs[2101] = ~((inputs[354]) | (inputs[5]));
    assign layer0_outputs[2102] = (inputs[568]) & ~(inputs[826]);
    assign layer0_outputs[2103] = (inputs[375]) & ~(inputs[355]);
    assign layer0_outputs[2104] = ~(inputs[974]);
    assign layer0_outputs[2105] = ~((inputs[646]) ^ (inputs[251]));
    assign layer0_outputs[2106] = ~((inputs[621]) | (inputs[232]));
    assign layer0_outputs[2107] = (inputs[740]) & (inputs[73]);
    assign layer0_outputs[2108] = (inputs[798]) & (inputs[670]);
    assign layer0_outputs[2109] = ~((inputs[515]) ^ (inputs[159]));
    assign layer0_outputs[2110] = (inputs[373]) & ~(inputs[39]);
    assign layer0_outputs[2111] = (inputs[719]) | (inputs[730]);
    assign layer0_outputs[2112] = (inputs[403]) | (inputs[298]);
    assign layer0_outputs[2113] = inputs[756];
    assign layer0_outputs[2114] = ~((inputs[7]) ^ (inputs[554]));
    assign layer0_outputs[2115] = (inputs[757]) ^ (inputs[1003]);
    assign layer0_outputs[2116] = ~(inputs[1007]) | (inputs[321]);
    assign layer0_outputs[2117] = ~((inputs[664]) ^ (inputs[796]));
    assign layer0_outputs[2118] = ~((inputs[296]) ^ (inputs[805]));
    assign layer0_outputs[2119] = (inputs[978]) & ~(inputs[411]);
    assign layer0_outputs[2120] = ~(inputs[471]) | (inputs[87]);
    assign layer0_outputs[2121] = (inputs[691]) & ~(inputs[837]);
    assign layer0_outputs[2122] = (inputs[458]) ^ (inputs[489]);
    assign layer0_outputs[2123] = (inputs[92]) & ~(inputs[772]);
    assign layer0_outputs[2124] = ~(inputs[776]) | (inputs[900]);
    assign layer0_outputs[2125] = ~(inputs[373]);
    assign layer0_outputs[2126] = inputs[622];
    assign layer0_outputs[2127] = ~((inputs[993]) & (inputs[893]));
    assign layer0_outputs[2128] = inputs[955];
    assign layer0_outputs[2129] = ~(inputs[671]) | (inputs[284]);
    assign layer0_outputs[2130] = ~(inputs[866]);
    assign layer0_outputs[2131] = 1'b1;
    assign layer0_outputs[2132] = (inputs[900]) | (inputs[213]);
    assign layer0_outputs[2133] = (inputs[333]) ^ (inputs[707]);
    assign layer0_outputs[2134] = ~(inputs[721]) | (inputs[871]);
    assign layer0_outputs[2135] = ~((inputs[348]) | (inputs[627]));
    assign layer0_outputs[2136] = (inputs[286]) ^ (inputs[426]);
    assign layer0_outputs[2137] = ~(inputs[491]);
    assign layer0_outputs[2138] = ~(inputs[459]);
    assign layer0_outputs[2139] = (inputs[405]) | (inputs[730]);
    assign layer0_outputs[2140] = ~((inputs[802]) | (inputs[562]));
    assign layer0_outputs[2141] = inputs[459];
    assign layer0_outputs[2142] = ~(inputs[315]);
    assign layer0_outputs[2143] = ~(inputs[251]);
    assign layer0_outputs[2144] = ~((inputs[196]) ^ (inputs[676]));
    assign layer0_outputs[2145] = ~((inputs[896]) ^ (inputs[645]));
    assign layer0_outputs[2146] = (inputs[768]) | (inputs[992]);
    assign layer0_outputs[2147] = (inputs[464]) & ~(inputs[993]);
    assign layer0_outputs[2148] = ~(inputs[184]) | (inputs[358]);
    assign layer0_outputs[2149] = (inputs[60]) | (inputs[648]);
    assign layer0_outputs[2150] = ~(inputs[398]) | (inputs[892]);
    assign layer0_outputs[2151] = ~((inputs[672]) | (inputs[67]));
    assign layer0_outputs[2152] = (inputs[687]) ^ (inputs[194]);
    assign layer0_outputs[2153] = (inputs[870]) & ~(inputs[85]);
    assign layer0_outputs[2154] = (inputs[817]) & ~(inputs[934]);
    assign layer0_outputs[2155] = (inputs[531]) ^ (inputs[759]);
    assign layer0_outputs[2156] = (inputs[666]) ^ (inputs[397]);
    assign layer0_outputs[2157] = (inputs[520]) & ~(inputs[688]);
    assign layer0_outputs[2158] = inputs[406];
    assign layer0_outputs[2159] = 1'b1;
    assign layer0_outputs[2160] = (inputs[663]) ^ (inputs[412]);
    assign layer0_outputs[2161] = (inputs[943]) & (inputs[965]);
    assign layer0_outputs[2162] = (inputs[898]) | (inputs[863]);
    assign layer0_outputs[2163] = 1'b1;
    assign layer0_outputs[2164] = ~((inputs[645]) | (inputs[553]));
    assign layer0_outputs[2165] = ~(inputs[462]);
    assign layer0_outputs[2166] = (inputs[960]) | (inputs[886]);
    assign layer0_outputs[2167] = (inputs[306]) & ~(inputs[263]);
    assign layer0_outputs[2168] = (inputs[372]) ^ (inputs[994]);
    assign layer0_outputs[2169] = inputs[496];
    assign layer0_outputs[2170] = ~(inputs[881]);
    assign layer0_outputs[2171] = (inputs[863]) | (inputs[905]);
    assign layer0_outputs[2172] = inputs[408];
    assign layer0_outputs[2173] = inputs[137];
    assign layer0_outputs[2174] = ~(inputs[127]);
    assign layer0_outputs[2175] = ~(inputs[716]) | (inputs[580]);
    assign layer0_outputs[2176] = ~((inputs[157]) ^ (inputs[852]));
    assign layer0_outputs[2177] = ~(inputs[811]) | (inputs[451]);
    assign layer0_outputs[2178] = ~((inputs[213]) | (inputs[179]));
    assign layer0_outputs[2179] = ~(inputs[400]) | (inputs[832]);
    assign layer0_outputs[2180] = (inputs[430]) & ~(inputs[53]);
    assign layer0_outputs[2181] = ~(inputs[784]);
    assign layer0_outputs[2182] = 1'b1;
    assign layer0_outputs[2183] = ~((inputs[824]) | (inputs[17]));
    assign layer0_outputs[2184] = ~((inputs[375]) | (inputs[186]));
    assign layer0_outputs[2185] = (inputs[624]) ^ (inputs[248]);
    assign layer0_outputs[2186] = (inputs[242]) | (inputs[133]);
    assign layer0_outputs[2187] = ~((inputs[520]) | (inputs[236]));
    assign layer0_outputs[2188] = ~((inputs[900]) & (inputs[1014]));
    assign layer0_outputs[2189] = ~(inputs[619]);
    assign layer0_outputs[2190] = ~((inputs[508]) | (inputs[726]));
    assign layer0_outputs[2191] = ~((inputs[896]) | (inputs[384]));
    assign layer0_outputs[2192] = 1'b1;
    assign layer0_outputs[2193] = ~((inputs[648]) ^ (inputs[616]));
    assign layer0_outputs[2194] = ~(inputs[459]) | (inputs[49]);
    assign layer0_outputs[2195] = (inputs[705]) ^ (inputs[396]);
    assign layer0_outputs[2196] = (inputs[230]) ^ (inputs[692]);
    assign layer0_outputs[2197] = (inputs[144]) ^ (inputs[960]);
    assign layer0_outputs[2198] = ~((inputs[973]) | (inputs[888]));
    assign layer0_outputs[2199] = ~((inputs[983]) & (inputs[184]));
    assign layer0_outputs[2200] = 1'b1;
    assign layer0_outputs[2201] = inputs[808];
    assign layer0_outputs[2202] = ~(inputs[492]);
    assign layer0_outputs[2203] = inputs[306];
    assign layer0_outputs[2204] = (inputs[563]) & ~(inputs[349]);
    assign layer0_outputs[2205] = ~(inputs[54]);
    assign layer0_outputs[2206] = (inputs[140]) & (inputs[296]);
    assign layer0_outputs[2207] = ~(inputs[652]);
    assign layer0_outputs[2208] = ~((inputs[31]) & (inputs[1022]));
    assign layer0_outputs[2209] = ~(inputs[476]);
    assign layer0_outputs[2210] = (inputs[474]) | (inputs[568]);
    assign layer0_outputs[2211] = ~((inputs[934]) | (inputs[77]));
    assign layer0_outputs[2212] = inputs[633];
    assign layer0_outputs[2213] = inputs[814];
    assign layer0_outputs[2214] = inputs[66];
    assign layer0_outputs[2215] = (inputs[810]) & (inputs[813]);
    assign layer0_outputs[2216] = (inputs[752]) & ~(inputs[899]);
    assign layer0_outputs[2217] = inputs[649];
    assign layer0_outputs[2218] = (inputs[675]) & ~(inputs[938]);
    assign layer0_outputs[2219] = ~(inputs[270]);
    assign layer0_outputs[2220] = (inputs[358]) ^ (inputs[801]);
    assign layer0_outputs[2221] = ~(inputs[215]);
    assign layer0_outputs[2222] = (inputs[949]) | (inputs[233]);
    assign layer0_outputs[2223] = ~(inputs[282]);
    assign layer0_outputs[2224] = ~((inputs[254]) | (inputs[546]));
    assign layer0_outputs[2225] = (inputs[107]) ^ (inputs[119]);
    assign layer0_outputs[2226] = (inputs[707]) ^ (inputs[360]);
    assign layer0_outputs[2227] = ~(inputs[301]) | (inputs[526]);
    assign layer0_outputs[2228] = (inputs[301]) ^ (inputs[166]);
    assign layer0_outputs[2229] = (inputs[658]) | (inputs[688]);
    assign layer0_outputs[2230] = inputs[591];
    assign layer0_outputs[2231] = inputs[862];
    assign layer0_outputs[2232] = inputs[880];
    assign layer0_outputs[2233] = (inputs[877]) ^ (inputs[133]);
    assign layer0_outputs[2234] = inputs[848];
    assign layer0_outputs[2235] = inputs[233];
    assign layer0_outputs[2236] = ~(inputs[697]) | (inputs[609]);
    assign layer0_outputs[2237] = (inputs[816]) & ~(inputs[300]);
    assign layer0_outputs[2238] = ~(inputs[487]) | (inputs[616]);
    assign layer0_outputs[2239] = (inputs[475]) ^ (inputs[432]);
    assign layer0_outputs[2240] = 1'b0;
    assign layer0_outputs[2241] = inputs[168];
    assign layer0_outputs[2242] = inputs[689];
    assign layer0_outputs[2243] = (inputs[128]) | (inputs[633]);
    assign layer0_outputs[2244] = (inputs[307]) & (inputs[254]);
    assign layer0_outputs[2245] = ~(inputs[6]);
    assign layer0_outputs[2246] = inputs[814];
    assign layer0_outputs[2247] = ~(inputs[528]);
    assign layer0_outputs[2248] = ~(inputs[455]);
    assign layer0_outputs[2249] = ~((inputs[71]) & (inputs[68]));
    assign layer0_outputs[2250] = ~((inputs[365]) ^ (inputs[470]));
    assign layer0_outputs[2251] = ~((inputs[800]) & (inputs[884]));
    assign layer0_outputs[2252] = ~(inputs[791]) | (inputs[205]);
    assign layer0_outputs[2253] = ~(inputs[852]) | (inputs[62]);
    assign layer0_outputs[2254] = ~((inputs[673]) & (inputs[892]));
    assign layer0_outputs[2255] = ~(inputs[677]);
    assign layer0_outputs[2256] = ~((inputs[54]) ^ (inputs[20]));
    assign layer0_outputs[2257] = ~(inputs[305]) | (inputs[153]);
    assign layer0_outputs[2258] = 1'b1;
    assign layer0_outputs[2259] = 1'b1;
    assign layer0_outputs[2260] = (inputs[959]) & ~(inputs[836]);
    assign layer0_outputs[2261] = ~(inputs[458]) | (inputs[964]);
    assign layer0_outputs[2262] = ~((inputs[425]) | (inputs[876]));
    assign layer0_outputs[2263] = ~(inputs[700]);
    assign layer0_outputs[2264] = (inputs[997]) & ~(inputs[905]);
    assign layer0_outputs[2265] = 1'b0;
    assign layer0_outputs[2266] = ~((inputs[615]) ^ (inputs[452]));
    assign layer0_outputs[2267] = 1'b1;
    assign layer0_outputs[2268] = inputs[487];
    assign layer0_outputs[2269] = (inputs[309]) | (inputs[808]);
    assign layer0_outputs[2270] = ~(inputs[361]);
    assign layer0_outputs[2271] = (inputs[972]) & ~(inputs[672]);
    assign layer0_outputs[2272] = (inputs[635]) & ~(inputs[888]);
    assign layer0_outputs[2273] = ~((inputs[329]) ^ (inputs[524]));
    assign layer0_outputs[2274] = (inputs[30]) & (inputs[56]);
    assign layer0_outputs[2275] = (inputs[136]) | (inputs[155]);
    assign layer0_outputs[2276] = inputs[585];
    assign layer0_outputs[2277] = ~(inputs[411]) | (inputs[735]);
    assign layer0_outputs[2278] = ~((inputs[832]) ^ (inputs[872]));
    assign layer0_outputs[2279] = inputs[302];
    assign layer0_outputs[2280] = ~((inputs[561]) | (inputs[239]));
    assign layer0_outputs[2281] = (inputs[294]) | (inputs[228]);
    assign layer0_outputs[2282] = ~(inputs[819]) | (inputs[217]);
    assign layer0_outputs[2283] = ~(inputs[193]) | (inputs[290]);
    assign layer0_outputs[2284] = (inputs[488]) & ~(inputs[53]);
    assign layer0_outputs[2285] = (inputs[594]) & ~(inputs[149]);
    assign layer0_outputs[2286] = inputs[340];
    assign layer0_outputs[2287] = (inputs[828]) | (inputs[285]);
    assign layer0_outputs[2288] = (inputs[178]) & ~(inputs[979]);
    assign layer0_outputs[2289] = inputs[361];
    assign layer0_outputs[2290] = (inputs[904]) & ~(inputs[161]);
    assign layer0_outputs[2291] = ~(inputs[762]);
    assign layer0_outputs[2292] = (inputs[600]) & ~(inputs[358]);
    assign layer0_outputs[2293] = (inputs[964]) & (inputs[542]);
    assign layer0_outputs[2294] = ~(inputs[716]) | (inputs[318]);
    assign layer0_outputs[2295] = 1'b1;
    assign layer0_outputs[2296] = ~(inputs[890]) | (inputs[1004]);
    assign layer0_outputs[2297] = ~(inputs[617]) | (inputs[153]);
    assign layer0_outputs[2298] = (inputs[720]) & ~(inputs[767]);
    assign layer0_outputs[2299] = ~(inputs[433]);
    assign layer0_outputs[2300] = ~(inputs[775]);
    assign layer0_outputs[2301] = (inputs[489]) ^ (inputs[265]);
    assign layer0_outputs[2302] = ~((inputs[115]) & (inputs[995]));
    assign layer0_outputs[2303] = (inputs[304]) & (inputs[863]);
    assign layer0_outputs[2304] = inputs[684];
    assign layer0_outputs[2305] = ~((inputs[278]) | (inputs[681]));
    assign layer0_outputs[2306] = ~((inputs[210]) | (inputs[673]));
    assign layer0_outputs[2307] = inputs[25];
    assign layer0_outputs[2308] = (inputs[211]) & ~(inputs[992]);
    assign layer0_outputs[2309] = (inputs[905]) & ~(inputs[736]);
    assign layer0_outputs[2310] = (inputs[760]) & ~(inputs[150]);
    assign layer0_outputs[2311] = ~((inputs[191]) | (inputs[59]));
    assign layer0_outputs[2312] = ~((inputs[946]) | (inputs[638]));
    assign layer0_outputs[2313] = inputs[875];
    assign layer0_outputs[2314] = ~((inputs[825]) | (inputs[734]));
    assign layer0_outputs[2315] = ~(inputs[252]);
    assign layer0_outputs[2316] = (inputs[203]) & ~(inputs[862]);
    assign layer0_outputs[2317] = 1'b0;
    assign layer0_outputs[2318] = inputs[872];
    assign layer0_outputs[2319] = (inputs[597]) ^ (inputs[506]);
    assign layer0_outputs[2320] = ~(inputs[875]);
    assign layer0_outputs[2321] = (inputs[282]) ^ (inputs[990]);
    assign layer0_outputs[2322] = 1'b1;
    assign layer0_outputs[2323] = ~(inputs[927]) | (inputs[508]);
    assign layer0_outputs[2324] = ~((inputs[915]) ^ (inputs[283]));
    assign layer0_outputs[2325] = ~((inputs[797]) ^ (inputs[858]));
    assign layer0_outputs[2326] = ~((inputs[359]) ^ (inputs[361]));
    assign layer0_outputs[2327] = (inputs[668]) & ~(inputs[483]);
    assign layer0_outputs[2328] = ~((inputs[853]) ^ (inputs[574]));
    assign layer0_outputs[2329] = ~((inputs[516]) & (inputs[150]));
    assign layer0_outputs[2330] = ~(inputs[333]);
    assign layer0_outputs[2331] = (inputs[348]) | (inputs[619]);
    assign layer0_outputs[2332] = ~((inputs[875]) ^ (inputs[310]));
    assign layer0_outputs[2333] = ~((inputs[360]) ^ (inputs[612]));
    assign layer0_outputs[2334] = ~(inputs[764]) | (inputs[194]);
    assign layer0_outputs[2335] = inputs[682];
    assign layer0_outputs[2336] = (inputs[242]) | (inputs[925]);
    assign layer0_outputs[2337] = ~((inputs[757]) | (inputs[113]));
    assign layer0_outputs[2338] = ~(inputs[458]);
    assign layer0_outputs[2339] = (inputs[136]) ^ (inputs[120]);
    assign layer0_outputs[2340] = (inputs[438]) & ~(inputs[113]);
    assign layer0_outputs[2341] = ~(inputs[464]) | (inputs[1014]);
    assign layer0_outputs[2342] = (inputs[281]) | (inputs[991]);
    assign layer0_outputs[2343] = ~((inputs[482]) | (inputs[996]));
    assign layer0_outputs[2344] = 1'b0;
    assign layer0_outputs[2345] = ~((inputs[929]) ^ (inputs[891]));
    assign layer0_outputs[2346] = (inputs[639]) ^ (inputs[1020]);
    assign layer0_outputs[2347] = (inputs[872]) | (inputs[475]);
    assign layer0_outputs[2348] = inputs[592];
    assign layer0_outputs[2349] = (inputs[366]) ^ (inputs[349]);
    assign layer0_outputs[2350] = (inputs[293]) & ~(inputs[737]);
    assign layer0_outputs[2351] = (inputs[436]) & ~(inputs[539]);
    assign layer0_outputs[2352] = (inputs[37]) ^ (inputs[1023]);
    assign layer0_outputs[2353] = (inputs[704]) ^ (inputs[847]);
    assign layer0_outputs[2354] = inputs[658];
    assign layer0_outputs[2355] = ~(inputs[426]) | (inputs[108]);
    assign layer0_outputs[2356] = inputs[932];
    assign layer0_outputs[2357] = 1'b0;
    assign layer0_outputs[2358] = inputs[809];
    assign layer0_outputs[2359] = ~(inputs[818]);
    assign layer0_outputs[2360] = inputs[754];
    assign layer0_outputs[2361] = ~((inputs[467]) | (inputs[101]));
    assign layer0_outputs[2362] = ~(inputs[471]) | (inputs[436]);
    assign layer0_outputs[2363] = (inputs[268]) & ~(inputs[763]);
    assign layer0_outputs[2364] = inputs[426];
    assign layer0_outputs[2365] = (inputs[184]) & ~(inputs[961]);
    assign layer0_outputs[2366] = ~((inputs[668]) | (inputs[557]));
    assign layer0_outputs[2367] = ~(inputs[720]);
    assign layer0_outputs[2368] = ~(inputs[496]);
    assign layer0_outputs[2369] = ~(inputs[362]);
    assign layer0_outputs[2370] = ~((inputs[646]) | (inputs[305]));
    assign layer0_outputs[2371] = (inputs[174]) & ~(inputs[907]);
    assign layer0_outputs[2372] = (inputs[984]) ^ (inputs[228]);
    assign layer0_outputs[2373] = ~(inputs[556]);
    assign layer0_outputs[2374] = (inputs[737]) ^ (inputs[800]);
    assign layer0_outputs[2375] = inputs[175];
    assign layer0_outputs[2376] = (inputs[972]) & ~(inputs[126]);
    assign layer0_outputs[2377] = (inputs[680]) & ~(inputs[2]);
    assign layer0_outputs[2378] = ~(inputs[534]);
    assign layer0_outputs[2379] = ~(inputs[817]) | (inputs[545]);
    assign layer0_outputs[2380] = inputs[327];
    assign layer0_outputs[2381] = (inputs[604]) ^ (inputs[536]);
    assign layer0_outputs[2382] = ~((inputs[432]) | (inputs[963]));
    assign layer0_outputs[2383] = inputs[773];
    assign layer0_outputs[2384] = (inputs[112]) ^ (inputs[278]);
    assign layer0_outputs[2385] = (inputs[972]) ^ (inputs[206]);
    assign layer0_outputs[2386] = ~((inputs[265]) | (inputs[642]));
    assign layer0_outputs[2387] = (inputs[844]) & ~(inputs[442]);
    assign layer0_outputs[2388] = ~(inputs[262]) | (inputs[99]);
    assign layer0_outputs[2389] = (inputs[803]) ^ (inputs[809]);
    assign layer0_outputs[2390] = (inputs[605]) & ~(inputs[2]);
    assign layer0_outputs[2391] = ~(inputs[939]);
    assign layer0_outputs[2392] = (inputs[234]) | (inputs[728]);
    assign layer0_outputs[2393] = ~(inputs[547]) | (inputs[15]);
    assign layer0_outputs[2394] = inputs[460];
    assign layer0_outputs[2395] = ~(inputs[775]) | (inputs[799]);
    assign layer0_outputs[2396] = (inputs[852]) | (inputs[709]);
    assign layer0_outputs[2397] = ~((inputs[695]) | (inputs[150]));
    assign layer0_outputs[2398] = (inputs[312]) & ~(inputs[582]);
    assign layer0_outputs[2399] = ~((inputs[59]) ^ (inputs[522]));
    assign layer0_outputs[2400] = ~((inputs[387]) & (inputs[761]));
    assign layer0_outputs[2401] = ~(inputs[871]) | (inputs[549]);
    assign layer0_outputs[2402] = 1'b1;
    assign layer0_outputs[2403] = ~((inputs[391]) ^ (inputs[891]));
    assign layer0_outputs[2404] = 1'b0;
    assign layer0_outputs[2405] = (inputs[207]) & ~(inputs[406]);
    assign layer0_outputs[2406] = 1'b0;
    assign layer0_outputs[2407] = ~((inputs[600]) | (inputs[806]));
    assign layer0_outputs[2408] = ~(inputs[599]);
    assign layer0_outputs[2409] = ~(inputs[271]);
    assign layer0_outputs[2410] = ~(inputs[609]) | (inputs[220]);
    assign layer0_outputs[2411] = (inputs[336]) ^ (inputs[810]);
    assign layer0_outputs[2412] = (inputs[179]) | (inputs[801]);
    assign layer0_outputs[2413] = (inputs[456]) & ~(inputs[281]);
    assign layer0_outputs[2414] = ~(inputs[71]) | (inputs[547]);
    assign layer0_outputs[2415] = (inputs[260]) ^ (inputs[739]);
    assign layer0_outputs[2416] = ~(inputs[232]);
    assign layer0_outputs[2417] = (inputs[812]) ^ (inputs[345]);
    assign layer0_outputs[2418] = ~((inputs[386]) & (inputs[595]));
    assign layer0_outputs[2419] = 1'b1;
    assign layer0_outputs[2420] = (inputs[1015]) & ~(inputs[318]);
    assign layer0_outputs[2421] = ~((inputs[250]) ^ (inputs[861]));
    assign layer0_outputs[2422] = ~(inputs[51]) | (inputs[142]);
    assign layer0_outputs[2423] = ~(inputs[505]) | (inputs[866]);
    assign layer0_outputs[2424] = ~(inputs[313]);
    assign layer0_outputs[2425] = 1'b1;
    assign layer0_outputs[2426] = 1'b0;
    assign layer0_outputs[2427] = 1'b0;
    assign layer0_outputs[2428] = ~(inputs[690]);
    assign layer0_outputs[2429] = (inputs[510]) ^ (inputs[536]);
    assign layer0_outputs[2430] = (inputs[477]) ^ (inputs[789]);
    assign layer0_outputs[2431] = inputs[306];
    assign layer0_outputs[2432] = ~(inputs[640]) | (inputs[423]);
    assign layer0_outputs[2433] = ~(inputs[342]) | (inputs[537]);
    assign layer0_outputs[2434] = (inputs[307]) | (inputs[392]);
    assign layer0_outputs[2435] = ~(inputs[532]);
    assign layer0_outputs[2436] = (inputs[523]) & ~(inputs[375]);
    assign layer0_outputs[2437] = (inputs[912]) ^ (inputs[915]);
    assign layer0_outputs[2438] = ~(inputs[532]);
    assign layer0_outputs[2439] = (inputs[148]) ^ (inputs[145]);
    assign layer0_outputs[2440] = inputs[760];
    assign layer0_outputs[2441] = ~((inputs[934]) ^ (inputs[183]));
    assign layer0_outputs[2442] = (inputs[378]) | (inputs[789]);
    assign layer0_outputs[2443] = inputs[954];
    assign layer0_outputs[2444] = ~((inputs[508]) ^ (inputs[679]));
    assign layer0_outputs[2445] = ~(inputs[918]);
    assign layer0_outputs[2446] = inputs[340];
    assign layer0_outputs[2447] = ~(inputs[523]) | (inputs[792]);
    assign layer0_outputs[2448] = (inputs[279]) ^ (inputs[227]);
    assign layer0_outputs[2449] = ~(inputs[249]) | (inputs[295]);
    assign layer0_outputs[2450] = ~((inputs[991]) | (inputs[37]));
    assign layer0_outputs[2451] = ~(inputs[245]);
    assign layer0_outputs[2452] = inputs[400];
    assign layer0_outputs[2453] = ~(inputs[83]);
    assign layer0_outputs[2454] = (inputs[630]) & ~(inputs[644]);
    assign layer0_outputs[2455] = ~(inputs[551]) | (inputs[288]);
    assign layer0_outputs[2456] = inputs[284];
    assign layer0_outputs[2457] = inputs[646];
    assign layer0_outputs[2458] = ~((inputs[326]) ^ (inputs[178]));
    assign layer0_outputs[2459] = ~(inputs[442]) | (inputs[983]);
    assign layer0_outputs[2460] = ~(inputs[780]) | (inputs[374]);
    assign layer0_outputs[2461] = (inputs[214]) ^ (inputs[239]);
    assign layer0_outputs[2462] = ~(inputs[952]) | (inputs[184]);
    assign layer0_outputs[2463] = ~(inputs[397]) | (inputs[1012]);
    assign layer0_outputs[2464] = (inputs[303]) & ~(inputs[772]);
    assign layer0_outputs[2465] = ~(inputs[635]) | (inputs[543]);
    assign layer0_outputs[2466] = ~(inputs[334]) | (inputs[552]);
    assign layer0_outputs[2467] = (inputs[577]) | (inputs[293]);
    assign layer0_outputs[2468] = ~((inputs[64]) | (inputs[499]));
    assign layer0_outputs[2469] = ~(inputs[522]) | (inputs[421]);
    assign layer0_outputs[2470] = ~(inputs[674]);
    assign layer0_outputs[2471] = (inputs[214]) ^ (inputs[339]);
    assign layer0_outputs[2472] = inputs[559];
    assign layer0_outputs[2473] = ~(inputs[32]);
    assign layer0_outputs[2474] = ~(inputs[877]) | (inputs[711]);
    assign layer0_outputs[2475] = (inputs[310]) | (inputs[345]);
    assign layer0_outputs[2476] = ~((inputs[630]) ^ (inputs[173]));
    assign layer0_outputs[2477] = ~(inputs[786]);
    assign layer0_outputs[2478] = ~(inputs[32]) | (inputs[74]);
    assign layer0_outputs[2479] = ~(inputs[875]);
    assign layer0_outputs[2480] = inputs[550];
    assign layer0_outputs[2481] = ~(inputs[418]) | (inputs[1015]);
    assign layer0_outputs[2482] = (inputs[322]) ^ (inputs[777]);
    assign layer0_outputs[2483] = inputs[467];
    assign layer0_outputs[2484] = ~(inputs[193]);
    assign layer0_outputs[2485] = (inputs[876]) | (inputs[856]);
    assign layer0_outputs[2486] = ~((inputs[433]) ^ (inputs[172]));
    assign layer0_outputs[2487] = (inputs[958]) ^ (inputs[746]);
    assign layer0_outputs[2488] = ~((inputs[941]) & (inputs[59]));
    assign layer0_outputs[2489] = inputs[716];
    assign layer0_outputs[2490] = (inputs[88]) & (inputs[355]);
    assign layer0_outputs[2491] = ~((inputs[780]) | (inputs[211]));
    assign layer0_outputs[2492] = (inputs[1006]) | (inputs[214]);
    assign layer0_outputs[2493] = inputs[139];
    assign layer0_outputs[2494] = inputs[931];
    assign layer0_outputs[2495] = (inputs[811]) ^ (inputs[670]);
    assign layer0_outputs[2496] = ~(inputs[770]);
    assign layer0_outputs[2497] = (inputs[163]) | (inputs[879]);
    assign layer0_outputs[2498] = (inputs[220]) & (inputs[929]);
    assign layer0_outputs[2499] = ~((inputs[275]) & (inputs[430]));
    assign layer0_outputs[2500] = ~(inputs[159]) | (inputs[730]);
    assign layer0_outputs[2501] = ~(inputs[530]);
    assign layer0_outputs[2502] = ~((inputs[239]) ^ (inputs[174]));
    assign layer0_outputs[2503] = (inputs[240]) ^ (inputs[44]);
    assign layer0_outputs[2504] = ~(inputs[474]) | (inputs[324]);
    assign layer0_outputs[2505] = ~(inputs[541]) | (inputs[873]);
    assign layer0_outputs[2506] = ~((inputs[330]) & (inputs[328]));
    assign layer0_outputs[2507] = (inputs[658]) | (inputs[159]);
    assign layer0_outputs[2508] = inputs[613];
    assign layer0_outputs[2509] = ~(inputs[380]);
    assign layer0_outputs[2510] = (inputs[508]) & ~(inputs[827]);
    assign layer0_outputs[2511] = (inputs[174]) ^ (inputs[696]);
    assign layer0_outputs[2512] = ~((inputs[597]) | (inputs[441]));
    assign layer0_outputs[2513] = ~(inputs[278]) | (inputs[144]);
    assign layer0_outputs[2514] = inputs[402];
    assign layer0_outputs[2515] = (inputs[528]) | (inputs[642]);
    assign layer0_outputs[2516] = ~((inputs[898]) ^ (inputs[372]));
    assign layer0_outputs[2517] = 1'b0;
    assign layer0_outputs[2518] = 1'b0;
    assign layer0_outputs[2519] = (inputs[271]) | (inputs[489]);
    assign layer0_outputs[2520] = (inputs[341]) & ~(inputs[47]);
    assign layer0_outputs[2521] = ~((inputs[258]) | (inputs[610]));
    assign layer0_outputs[2522] = ~(inputs[660]);
    assign layer0_outputs[2523] = (inputs[609]) | (inputs[888]);
    assign layer0_outputs[2524] = (inputs[310]) & ~(inputs[657]);
    assign layer0_outputs[2525] = (inputs[414]) & (inputs[167]);
    assign layer0_outputs[2526] = ~(inputs[283]) | (inputs[159]);
    assign layer0_outputs[2527] = ~((inputs[100]) | (inputs[829]));
    assign layer0_outputs[2528] = ~((inputs[772]) | (inputs[797]));
    assign layer0_outputs[2529] = inputs[130];
    assign layer0_outputs[2530] = ~(inputs[487]);
    assign layer0_outputs[2531] = (inputs[864]) ^ (inputs[380]);
    assign layer0_outputs[2532] = (inputs[843]) | (inputs[267]);
    assign layer0_outputs[2533] = ~((inputs[25]) | (inputs[856]));
    assign layer0_outputs[2534] = 1'b1;
    assign layer0_outputs[2535] = (inputs[149]) & ~(inputs[516]);
    assign layer0_outputs[2536] = ~((inputs[603]) | (inputs[416]));
    assign layer0_outputs[2537] = (inputs[568]) & ~(inputs[708]);
    assign layer0_outputs[2538] = (inputs[213]) & ~(inputs[463]);
    assign layer0_outputs[2539] = (inputs[841]) & ~(inputs[198]);
    assign layer0_outputs[2540] = (inputs[1023]) & ~(inputs[36]);
    assign layer0_outputs[2541] = ~(inputs[858]) | (inputs[1018]);
    assign layer0_outputs[2542] = ~((inputs[994]) & (inputs[375]));
    assign layer0_outputs[2543] = ~(inputs[523]);
    assign layer0_outputs[2544] = (inputs[980]) ^ (inputs[381]);
    assign layer0_outputs[2545] = inputs[941];
    assign layer0_outputs[2546] = ~(inputs[348]);
    assign layer0_outputs[2547] = ~(inputs[540]) | (inputs[481]);
    assign layer0_outputs[2548] = ~((inputs[253]) | (inputs[61]));
    assign layer0_outputs[2549] = inputs[666];
    assign layer0_outputs[2550] = (inputs[445]) ^ (inputs[347]);
    assign layer0_outputs[2551] = inputs[861];
    assign layer0_outputs[2552] = (inputs[16]) ^ (inputs[89]);
    assign layer0_outputs[2553] = (inputs[939]) | (inputs[738]);
    assign layer0_outputs[2554] = ~(inputs[271]) | (inputs[943]);
    assign layer0_outputs[2555] = (inputs[486]) | (inputs[915]);
    assign layer0_outputs[2556] = (inputs[247]) ^ (inputs[119]);
    assign layer0_outputs[2557] = (inputs[639]) & ~(inputs[390]);
    assign layer0_outputs[2558] = ~(inputs[400]);
    assign layer0_outputs[2559] = ~((inputs[62]) & (inputs[4]));
    assign layer0_outputs[2560] = inputs[611];
    assign layer0_outputs[2561] = (inputs[60]) & (inputs[646]);
    assign layer0_outputs[2562] = (inputs[384]) & ~(inputs[66]);
    assign layer0_outputs[2563] = ~((inputs[464]) | (inputs[723]));
    assign layer0_outputs[2564] = (inputs[96]) & ~(inputs[287]);
    assign layer0_outputs[2565] = ~(inputs[216]) | (inputs[751]);
    assign layer0_outputs[2566] = (inputs[911]) | (inputs[1019]);
    assign layer0_outputs[2567] = 1'b1;
    assign layer0_outputs[2568] = ~((inputs[526]) | (inputs[627]));
    assign layer0_outputs[2569] = (inputs[9]) & (inputs[162]);
    assign layer0_outputs[2570] = ~((inputs[1014]) | (inputs[16]));
    assign layer0_outputs[2571] = inputs[537];
    assign layer0_outputs[2572] = (inputs[487]) & ~(inputs[230]);
    assign layer0_outputs[2573] = (inputs[194]) & ~(inputs[815]);
    assign layer0_outputs[2574] = ~(inputs[7]);
    assign layer0_outputs[2575] = ~(inputs[299]);
    assign layer0_outputs[2576] = ~(inputs[938]);
    assign layer0_outputs[2577] = ~((inputs[284]) ^ (inputs[368]));
    assign layer0_outputs[2578] = (inputs[344]) | (inputs[232]);
    assign layer0_outputs[2579] = (inputs[627]) & ~(inputs[391]);
    assign layer0_outputs[2580] = (inputs[796]) & ~(inputs[27]);
    assign layer0_outputs[2581] = inputs[10];
    assign layer0_outputs[2582] = (inputs[989]) & ~(inputs[501]);
    assign layer0_outputs[2583] = inputs[987];
    assign layer0_outputs[2584] = (inputs[634]) ^ (inputs[124]);
    assign layer0_outputs[2585] = (inputs[619]) ^ (inputs[29]);
    assign layer0_outputs[2586] = (inputs[92]) | (inputs[245]);
    assign layer0_outputs[2587] = (inputs[379]) | (inputs[490]);
    assign layer0_outputs[2588] = ~((inputs[56]) & (inputs[354]));
    assign layer0_outputs[2589] = (inputs[598]) ^ (inputs[463]);
    assign layer0_outputs[2590] = inputs[449];
    assign layer0_outputs[2591] = ~(inputs[921]);
    assign layer0_outputs[2592] = ~((inputs[980]) & (inputs[1012]));
    assign layer0_outputs[2593] = ~((inputs[1017]) & (inputs[66]));
    assign layer0_outputs[2594] = ~(inputs[975]) | (inputs[135]);
    assign layer0_outputs[2595] = (inputs[114]) & ~(inputs[229]);
    assign layer0_outputs[2596] = (inputs[807]) | (inputs[267]);
    assign layer0_outputs[2597] = ~((inputs[557]) | (inputs[203]));
    assign layer0_outputs[2598] = ~(inputs[457]) | (inputs[806]);
    assign layer0_outputs[2599] = (inputs[774]) & ~(inputs[421]);
    assign layer0_outputs[2600] = ~(inputs[853]) | (inputs[446]);
    assign layer0_outputs[2601] = ~((inputs[247]) ^ (inputs[380]));
    assign layer0_outputs[2602] = ~((inputs[300]) & (inputs[1018]));
    assign layer0_outputs[2603] = ~(inputs[450]) | (inputs[51]);
    assign layer0_outputs[2604] = (inputs[1012]) & ~(inputs[301]);
    assign layer0_outputs[2605] = ~(inputs[683]);
    assign layer0_outputs[2606] = inputs[264];
    assign layer0_outputs[2607] = (inputs[799]) ^ (inputs[166]);
    assign layer0_outputs[2608] = inputs[274];
    assign layer0_outputs[2609] = (inputs[237]) ^ (inputs[398]);
    assign layer0_outputs[2610] = (inputs[418]) & (inputs[802]);
    assign layer0_outputs[2611] = ~(inputs[474]) | (inputs[822]);
    assign layer0_outputs[2612] = ~(inputs[554]) | (inputs[144]);
    assign layer0_outputs[2613] = (inputs[789]) & (inputs[476]);
    assign layer0_outputs[2614] = (inputs[340]) & ~(inputs[167]);
    assign layer0_outputs[2615] = ~(inputs[834]) | (inputs[721]);
    assign layer0_outputs[2616] = ~(inputs[272]);
    assign layer0_outputs[2617] = 1'b0;
    assign layer0_outputs[2618] = 1'b0;
    assign layer0_outputs[2619] = ~((inputs[82]) | (inputs[741]));
    assign layer0_outputs[2620] = (inputs[931]) ^ (inputs[685]);
    assign layer0_outputs[2621] = ~(inputs[790]);
    assign layer0_outputs[2622] = (inputs[783]) & ~(inputs[167]);
    assign layer0_outputs[2623] = ~((inputs[849]) | (inputs[205]));
    assign layer0_outputs[2624] = ~(inputs[250]);
    assign layer0_outputs[2625] = ~((inputs[728]) | (inputs[208]));
    assign layer0_outputs[2626] = ~(inputs[88]) | (inputs[228]);
    assign layer0_outputs[2627] = (inputs[522]) & ~(inputs[939]);
    assign layer0_outputs[2628] = ~(inputs[546]);
    assign layer0_outputs[2629] = ~((inputs[792]) ^ (inputs[509]));
    assign layer0_outputs[2630] = (inputs[469]) | (inputs[147]);
    assign layer0_outputs[2631] = (inputs[86]) & ~(inputs[285]);
    assign layer0_outputs[2632] = (inputs[550]) & ~(inputs[386]);
    assign layer0_outputs[2633] = ~((inputs[415]) | (inputs[273]));
    assign layer0_outputs[2634] = (inputs[374]) & ~(inputs[498]);
    assign layer0_outputs[2635] = inputs[588];
    assign layer0_outputs[2636] = ~((inputs[302]) | (inputs[129]));
    assign layer0_outputs[2637] = (inputs[253]) | (inputs[696]);
    assign layer0_outputs[2638] = ~(inputs[55]);
    assign layer0_outputs[2639] = (inputs[663]) | (inputs[75]);
    assign layer0_outputs[2640] = (inputs[259]) ^ (inputs[923]);
    assign layer0_outputs[2641] = ~(inputs[672]) | (inputs[80]);
    assign layer0_outputs[2642] = (inputs[972]) & ~(inputs[138]);
    assign layer0_outputs[2643] = ~((inputs[586]) | (inputs[698]));
    assign layer0_outputs[2644] = 1'b0;
    assign layer0_outputs[2645] = ~(inputs[650]) | (inputs[825]);
    assign layer0_outputs[2646] = ~((inputs[29]) & (inputs[1008]));
    assign layer0_outputs[2647] = (inputs[429]) | (inputs[120]);
    assign layer0_outputs[2648] = (inputs[753]) | (inputs[947]);
    assign layer0_outputs[2649] = ~(inputs[775]) | (inputs[551]);
    assign layer0_outputs[2650] = ~((inputs[831]) ^ (inputs[443]));
    assign layer0_outputs[2651] = (inputs[502]) & ~(inputs[70]);
    assign layer0_outputs[2652] = inputs[759];
    assign layer0_outputs[2653] = ~(inputs[237]) | (inputs[1020]);
    assign layer0_outputs[2654] = (inputs[69]) | (inputs[837]);
    assign layer0_outputs[2655] = (inputs[688]) | (inputs[108]);
    assign layer0_outputs[2656] = ~((inputs[548]) | (inputs[944]));
    assign layer0_outputs[2657] = ~((inputs[87]) | (inputs[1000]));
    assign layer0_outputs[2658] = (inputs[649]) & ~(inputs[518]);
    assign layer0_outputs[2659] = 1'b1;
    assign layer0_outputs[2660] = inputs[107];
    assign layer0_outputs[2661] = inputs[945];
    assign layer0_outputs[2662] = ~((inputs[116]) | (inputs[944]));
    assign layer0_outputs[2663] = inputs[203];
    assign layer0_outputs[2664] = ~(inputs[398]);
    assign layer0_outputs[2665] = (inputs[514]) & (inputs[703]);
    assign layer0_outputs[2666] = (inputs[830]) | (inputs[261]);
    assign layer0_outputs[2667] = 1'b0;
    assign layer0_outputs[2668] = (inputs[444]) & (inputs[978]);
    assign layer0_outputs[2669] = inputs[904];
    assign layer0_outputs[2670] = (inputs[474]) & ~(inputs[3]);
    assign layer0_outputs[2671] = ~(inputs[751]) | (inputs[856]);
    assign layer0_outputs[2672] = ~((inputs[63]) ^ (inputs[704]));
    assign layer0_outputs[2673] = (inputs[917]) ^ (inputs[624]);
    assign layer0_outputs[2674] = inputs[646];
    assign layer0_outputs[2675] = ~(inputs[591]);
    assign layer0_outputs[2676] = ~(inputs[399]);
    assign layer0_outputs[2677] = ~(inputs[937]);
    assign layer0_outputs[2678] = ~((inputs[631]) | (inputs[442]));
    assign layer0_outputs[2679] = ~((inputs[783]) | (inputs[55]));
    assign layer0_outputs[2680] = ~(inputs[204]);
    assign layer0_outputs[2681] = (inputs[607]) & ~(inputs[150]);
    assign layer0_outputs[2682] = ~(inputs[186]) | (inputs[671]);
    assign layer0_outputs[2683] = inputs[653];
    assign layer0_outputs[2684] = inputs[694];
    assign layer0_outputs[2685] = ~(inputs[877]) | (inputs[356]);
    assign layer0_outputs[2686] = ~((inputs[34]) | (inputs[340]));
    assign layer0_outputs[2687] = ~((inputs[253]) | (inputs[605]));
    assign layer0_outputs[2688] = ~((inputs[411]) | (inputs[259]));
    assign layer0_outputs[2689] = ~(inputs[528]);
    assign layer0_outputs[2690] = inputs[906];
    assign layer0_outputs[2691] = ~((inputs[822]) | (inputs[319]));
    assign layer0_outputs[2692] = ~(inputs[172]);
    assign layer0_outputs[2693] = ~(inputs[674]);
    assign layer0_outputs[2694] = ~(inputs[356]);
    assign layer0_outputs[2695] = ~(inputs[46]);
    assign layer0_outputs[2696] = ~((inputs[279]) ^ (inputs[613]));
    assign layer0_outputs[2697] = ~((inputs[134]) | (inputs[945]));
    assign layer0_outputs[2698] = ~((inputs[565]) | (inputs[386]));
    assign layer0_outputs[2699] = (inputs[113]) & (inputs[443]);
    assign layer0_outputs[2700] = (inputs[101]) ^ (inputs[746]);
    assign layer0_outputs[2701] = inputs[811];
    assign layer0_outputs[2702] = (inputs[349]) & ~(inputs[967]);
    assign layer0_outputs[2703] = ~(inputs[401]) | (inputs[383]);
    assign layer0_outputs[2704] = ~((inputs[240]) & (inputs[274]));
    assign layer0_outputs[2705] = (inputs[367]) ^ (inputs[129]);
    assign layer0_outputs[2706] = ~(inputs[387]);
    assign layer0_outputs[2707] = (inputs[262]) ^ (inputs[927]);
    assign layer0_outputs[2708] = ~((inputs[976]) ^ (inputs[637]));
    assign layer0_outputs[2709] = (inputs[223]) & (inputs[62]);
    assign layer0_outputs[2710] = ~(inputs[679]);
    assign layer0_outputs[2711] = ~(inputs[528]) | (inputs[245]);
    assign layer0_outputs[2712] = (inputs[179]) | (inputs[834]);
    assign layer0_outputs[2713] = (inputs[517]) & ~(inputs[548]);
    assign layer0_outputs[2714] = ~((inputs[414]) ^ (inputs[455]));
    assign layer0_outputs[2715] = ~((inputs[537]) ^ (inputs[1005]));
    assign layer0_outputs[2716] = ~(inputs[188]) | (inputs[123]);
    assign layer0_outputs[2717] = ~((inputs[355]) ^ (inputs[70]));
    assign layer0_outputs[2718] = ~(inputs[588]) | (inputs[111]);
    assign layer0_outputs[2719] = inputs[826];
    assign layer0_outputs[2720] = ~((inputs[261]) | (inputs[568]));
    assign layer0_outputs[2721] = ~(inputs[569]);
    assign layer0_outputs[2722] = 1'b1;
    assign layer0_outputs[2723] = ~(inputs[650]);
    assign layer0_outputs[2724] = (inputs[839]) ^ (inputs[861]);
    assign layer0_outputs[2725] = ~(inputs[380]);
    assign layer0_outputs[2726] = (inputs[394]) ^ (inputs[918]);
    assign layer0_outputs[2727] = 1'b0;
    assign layer0_outputs[2728] = 1'b1;
    assign layer0_outputs[2729] = ~((inputs[366]) | (inputs[503]));
    assign layer0_outputs[2730] = inputs[171];
    assign layer0_outputs[2731] = ~(inputs[883]) | (inputs[10]);
    assign layer0_outputs[2732] = ~(inputs[492]) | (inputs[697]);
    assign layer0_outputs[2733] = 1'b1;
    assign layer0_outputs[2734] = ~(inputs[490]) | (inputs[612]);
    assign layer0_outputs[2735] = ~((inputs[247]) | (inputs[863]));
    assign layer0_outputs[2736] = (inputs[35]) & (inputs[98]);
    assign layer0_outputs[2737] = ~((inputs[655]) | (inputs[510]));
    assign layer0_outputs[2738] = (inputs[426]) & ~(inputs[1017]);
    assign layer0_outputs[2739] = ~(inputs[187]) | (inputs[418]);
    assign layer0_outputs[2740] = ~((inputs[231]) | (inputs[222]));
    assign layer0_outputs[2741] = (inputs[864]) ^ (inputs[399]);
    assign layer0_outputs[2742] = inputs[658];
    assign layer0_outputs[2743] = ~((inputs[478]) ^ (inputs[736]));
    assign layer0_outputs[2744] = ~((inputs[100]) | (inputs[831]));
    assign layer0_outputs[2745] = (inputs[33]) | (inputs[13]);
    assign layer0_outputs[2746] = inputs[77];
    assign layer0_outputs[2747] = ~(inputs[491]) | (inputs[89]);
    assign layer0_outputs[2748] = (inputs[538]) | (inputs[900]);
    assign layer0_outputs[2749] = ~(inputs[678]);
    assign layer0_outputs[2750] = 1'b0;
    assign layer0_outputs[2751] = inputs[3];
    assign layer0_outputs[2752] = (inputs[614]) & ~(inputs[415]);
    assign layer0_outputs[2753] = 1'b1;
    assign layer0_outputs[2754] = inputs[386];
    assign layer0_outputs[2755] = 1'b0;
    assign layer0_outputs[2756] = (inputs[904]) & ~(inputs[34]);
    assign layer0_outputs[2757] = (inputs[618]) | (inputs[205]);
    assign layer0_outputs[2758] = ~(inputs[364]) | (inputs[926]);
    assign layer0_outputs[2759] = ~(inputs[317]);
    assign layer0_outputs[2760] = ~((inputs[932]) | (inputs[216]));
    assign layer0_outputs[2761] = (inputs[755]) ^ (inputs[1005]);
    assign layer0_outputs[2762] = 1'b1;
    assign layer0_outputs[2763] = inputs[418];
    assign layer0_outputs[2764] = (inputs[433]) ^ (inputs[543]);
    assign layer0_outputs[2765] = inputs[262];
    assign layer0_outputs[2766] = ~(inputs[890]);
    assign layer0_outputs[2767] = inputs[685];
    assign layer0_outputs[2768] = 1'b1;
    assign layer0_outputs[2769] = ~(inputs[593]);
    assign layer0_outputs[2770] = 1'b1;
    assign layer0_outputs[2771] = ~((inputs[544]) | (inputs[488]));
    assign layer0_outputs[2772] = (inputs[5]) ^ (inputs[258]);
    assign layer0_outputs[2773] = (inputs[461]) ^ (inputs[537]);
    assign layer0_outputs[2774] = inputs[218];
    assign layer0_outputs[2775] = (inputs[712]) | (inputs[629]);
    assign layer0_outputs[2776] = inputs[430];
    assign layer0_outputs[2777] = inputs[276];
    assign layer0_outputs[2778] = (inputs[132]) & ~(inputs[762]);
    assign layer0_outputs[2779] = (inputs[77]) ^ (inputs[84]);
    assign layer0_outputs[2780] = (inputs[379]) | (inputs[762]);
    assign layer0_outputs[2781] = ~(inputs[486]);
    assign layer0_outputs[2782] = ~(inputs[367]) | (inputs[385]);
    assign layer0_outputs[2783] = inputs[237];
    assign layer0_outputs[2784] = ~(inputs[975]) | (inputs[317]);
    assign layer0_outputs[2785] = (inputs[107]) | (inputs[570]);
    assign layer0_outputs[2786] = inputs[213];
    assign layer0_outputs[2787] = ~(inputs[45]) | (inputs[1021]);
    assign layer0_outputs[2788] = (inputs[411]) ^ (inputs[118]);
    assign layer0_outputs[2789] = ~(inputs[935]);
    assign layer0_outputs[2790] = (inputs[888]) & (inputs[200]);
    assign layer0_outputs[2791] = (inputs[1004]) & ~(inputs[65]);
    assign layer0_outputs[2792] = ~(inputs[386]) | (inputs[823]);
    assign layer0_outputs[2793] = ~((inputs[434]) ^ (inputs[543]));
    assign layer0_outputs[2794] = ~(inputs[967]);
    assign layer0_outputs[2795] = ~((inputs[315]) | (inputs[533]));
    assign layer0_outputs[2796] = ~(inputs[637]);
    assign layer0_outputs[2797] = ~((inputs[328]) ^ (inputs[173]));
    assign layer0_outputs[2798] = (inputs[965]) | (inputs[397]);
    assign layer0_outputs[2799] = ~((inputs[143]) | (inputs[821]));
    assign layer0_outputs[2800] = ~((inputs[25]) | (inputs[153]));
    assign layer0_outputs[2801] = ~(inputs[207]);
    assign layer0_outputs[2802] = ~((inputs[225]) | (inputs[440]));
    assign layer0_outputs[2803] = (inputs[96]) ^ (inputs[295]);
    assign layer0_outputs[2804] = (inputs[772]) | (inputs[732]);
    assign layer0_outputs[2805] = ~((inputs[692]) | (inputs[106]));
    assign layer0_outputs[2806] = ~((inputs[662]) & (inputs[534]));
    assign layer0_outputs[2807] = ~(inputs[591]);
    assign layer0_outputs[2808] = ~((inputs[996]) | (inputs[651]));
    assign layer0_outputs[2809] = ~((inputs[196]) | (inputs[236]));
    assign layer0_outputs[2810] = ~(inputs[365]) | (inputs[88]);
    assign layer0_outputs[2811] = ~(inputs[638]);
    assign layer0_outputs[2812] = (inputs[957]) | (inputs[317]);
    assign layer0_outputs[2813] = ~(inputs[273]);
    assign layer0_outputs[2814] = ~((inputs[195]) & (inputs[321]));
    assign layer0_outputs[2815] = ~(inputs[432]);
    assign layer0_outputs[2816] = ~(inputs[787]);
    assign layer0_outputs[2817] = ~(inputs[942]) | (inputs[950]);
    assign layer0_outputs[2818] = ~(inputs[639]) | (inputs[83]);
    assign layer0_outputs[2819] = inputs[1014];
    assign layer0_outputs[2820] = inputs[11];
    assign layer0_outputs[2821] = ~((inputs[248]) | (inputs[428]));
    assign layer0_outputs[2822] = inputs[205];
    assign layer0_outputs[2823] = (inputs[163]) | (inputs[504]);
    assign layer0_outputs[2824] = ~((inputs[412]) ^ (inputs[304]));
    assign layer0_outputs[2825] = ~((inputs[975]) & (inputs[88]));
    assign layer0_outputs[2826] = (inputs[649]) | (inputs[815]);
    assign layer0_outputs[2827] = (inputs[271]) | (inputs[743]);
    assign layer0_outputs[2828] = ~(inputs[446]) | (inputs[72]);
    assign layer0_outputs[2829] = ~(inputs[657]);
    assign layer0_outputs[2830] = inputs[467];
    assign layer0_outputs[2831] = (inputs[758]) & ~(inputs[103]);
    assign layer0_outputs[2832] = ~(inputs[472]);
    assign layer0_outputs[2833] = (inputs[77]) & (inputs[198]);
    assign layer0_outputs[2834] = ~((inputs[210]) ^ (inputs[840]));
    assign layer0_outputs[2835] = inputs[534];
    assign layer0_outputs[2836] = ~((inputs[623]) | (inputs[628]));
    assign layer0_outputs[2837] = inputs[838];
    assign layer0_outputs[2838] = ~(inputs[961]) | (inputs[452]);
    assign layer0_outputs[2839] = inputs[306];
    assign layer0_outputs[2840] = ~((inputs[441]) | (inputs[860]));
    assign layer0_outputs[2841] = ~((inputs[194]) | (inputs[573]));
    assign layer0_outputs[2842] = (inputs[1002]) & ~(inputs[561]);
    assign layer0_outputs[2843] = (inputs[787]) & ~(inputs[513]);
    assign layer0_outputs[2844] = (inputs[259]) & (inputs[676]);
    assign layer0_outputs[2845] = ~(inputs[552]);
    assign layer0_outputs[2846] = inputs[806];
    assign layer0_outputs[2847] = ~((inputs[75]) | (inputs[696]));
    assign layer0_outputs[2848] = ~((inputs[213]) ^ (inputs[885]));
    assign layer0_outputs[2849] = inputs[817];
    assign layer0_outputs[2850] = (inputs[605]) | (inputs[367]);
    assign layer0_outputs[2851] = ~(inputs[774]) | (inputs[165]);
    assign layer0_outputs[2852] = (inputs[201]) | (inputs[167]);
    assign layer0_outputs[2853] = inputs[908];
    assign layer0_outputs[2854] = ~(inputs[614]) | (inputs[79]);
    assign layer0_outputs[2855] = ~((inputs[864]) | (inputs[902]));
    assign layer0_outputs[2856] = ~(inputs[89]) | (inputs[966]);
    assign layer0_outputs[2857] = ~(inputs[461]) | (inputs[579]);
    assign layer0_outputs[2858] = inputs[689];
    assign layer0_outputs[2859] = ~(inputs[64]);
    assign layer0_outputs[2860] = ~(inputs[529]) | (inputs[827]);
    assign layer0_outputs[2861] = (inputs[171]) | (inputs[721]);
    assign layer0_outputs[2862] = ~(inputs[302]);
    assign layer0_outputs[2863] = ~(inputs[404]) | (inputs[963]);
    assign layer0_outputs[2864] = 1'b0;
    assign layer0_outputs[2865] = (inputs[396]) & ~(inputs[212]);
    assign layer0_outputs[2866] = (inputs[414]) ^ (inputs[315]);
    assign layer0_outputs[2867] = inputs[593];
    assign layer0_outputs[2868] = ~((inputs[945]) ^ (inputs[928]));
    assign layer0_outputs[2869] = ~((inputs[252]) ^ (inputs[20]));
    assign layer0_outputs[2870] = ~((inputs[713]) | (inputs[691]));
    assign layer0_outputs[2871] = 1'b0;
    assign layer0_outputs[2872] = ~(inputs[252]) | (inputs[547]);
    assign layer0_outputs[2873] = ~((inputs[740]) | (inputs[79]));
    assign layer0_outputs[2874] = ~(inputs[273]) | (inputs[249]);
    assign layer0_outputs[2875] = inputs[32];
    assign layer0_outputs[2876] = (inputs[533]) & ~(inputs[390]);
    assign layer0_outputs[2877] = (inputs[170]) ^ (inputs[903]);
    assign layer0_outputs[2878] = 1'b1;
    assign layer0_outputs[2879] = ~(inputs[587]);
    assign layer0_outputs[2880] = (inputs[814]) & ~(inputs[804]);
    assign layer0_outputs[2881] = ~((inputs[579]) ^ (inputs[557]));
    assign layer0_outputs[2882] = ~(inputs[814]) | (inputs[544]);
    assign layer0_outputs[2883] = (inputs[323]) | (inputs[967]);
    assign layer0_outputs[2884] = ~((inputs[982]) | (inputs[51]));
    assign layer0_outputs[2885] = ~(inputs[615]);
    assign layer0_outputs[2886] = (inputs[146]) & ~(inputs[284]);
    assign layer0_outputs[2887] = (inputs[919]) & (inputs[18]);
    assign layer0_outputs[2888] = (inputs[98]) & (inputs[756]);
    assign layer0_outputs[2889] = ~(inputs[48]);
    assign layer0_outputs[2890] = (inputs[596]) & ~(inputs[940]);
    assign layer0_outputs[2891] = ~(inputs[463]);
    assign layer0_outputs[2892] = ~((inputs[632]) ^ (inputs[960]));
    assign layer0_outputs[2893] = ~((inputs[758]) ^ (inputs[56]));
    assign layer0_outputs[2894] = ~(inputs[740]);
    assign layer0_outputs[2895] = ~(inputs[368]);
    assign layer0_outputs[2896] = ~((inputs[704]) & (inputs[447]));
    assign layer0_outputs[2897] = ~((inputs[829]) | (inputs[907]));
    assign layer0_outputs[2898] = (inputs[943]) & (inputs[738]);
    assign layer0_outputs[2899] = 1'b1;
    assign layer0_outputs[2900] = inputs[862];
    assign layer0_outputs[2901] = ~(inputs[675]);
    assign layer0_outputs[2902] = ~((inputs[792]) | (inputs[316]));
    assign layer0_outputs[2903] = ~(inputs[822]);
    assign layer0_outputs[2904] = (inputs[411]) | (inputs[1012]);
    assign layer0_outputs[2905] = ~(inputs[295]);
    assign layer0_outputs[2906] = ~(inputs[882]);
    assign layer0_outputs[2907] = (inputs[844]) | (inputs[288]);
    assign layer0_outputs[2908] = ~((inputs[844]) ^ (inputs[378]));
    assign layer0_outputs[2909] = ~(inputs[216]) | (inputs[1003]);
    assign layer0_outputs[2910] = ~(inputs[363]) | (inputs[55]);
    assign layer0_outputs[2911] = inputs[847];
    assign layer0_outputs[2912] = (inputs[1018]) & ~(inputs[594]);
    assign layer0_outputs[2913] = ~((inputs[116]) ^ (inputs[294]));
    assign layer0_outputs[2914] = ~(inputs[972]) | (inputs[905]);
    assign layer0_outputs[2915] = ~(inputs[586]);
    assign layer0_outputs[2916] = ~(inputs[920]);
    assign layer0_outputs[2917] = (inputs[458]) | (inputs[831]);
    assign layer0_outputs[2918] = ~(inputs[809]) | (inputs[392]);
    assign layer0_outputs[2919] = inputs[523];
    assign layer0_outputs[2920] = ~((inputs[159]) | (inputs[679]));
    assign layer0_outputs[2921] = ~((inputs[205]) | (inputs[777]));
    assign layer0_outputs[2922] = ~(inputs[592]);
    assign layer0_outputs[2923] = ~(inputs[641]);
    assign layer0_outputs[2924] = (inputs[885]) & (inputs[905]);
    assign layer0_outputs[2925] = ~((inputs[700]) | (inputs[643]));
    assign layer0_outputs[2926] = (inputs[383]) ^ (inputs[798]);
    assign layer0_outputs[2927] = (inputs[381]) | (inputs[80]);
    assign layer0_outputs[2928] = ~(inputs[504]);
    assign layer0_outputs[2929] = (inputs[579]) & ~(inputs[124]);
    assign layer0_outputs[2930] = inputs[671];
    assign layer0_outputs[2931] = (inputs[973]) & ~(inputs[141]);
    assign layer0_outputs[2932] = (inputs[543]) & ~(inputs[13]);
    assign layer0_outputs[2933] = ~(inputs[49]);
    assign layer0_outputs[2934] = (inputs[965]) ^ (inputs[870]);
    assign layer0_outputs[2935] = (inputs[511]) ^ (inputs[981]);
    assign layer0_outputs[2936] = (inputs[159]) ^ (inputs[994]);
    assign layer0_outputs[2937] = (inputs[246]) ^ (inputs[727]);
    assign layer0_outputs[2938] = ~(inputs[141]);
    assign layer0_outputs[2939] = (inputs[347]) | (inputs[189]);
    assign layer0_outputs[2940] = (inputs[89]) & (inputs[950]);
    assign layer0_outputs[2941] = ~(inputs[502]);
    assign layer0_outputs[2942] = inputs[385];
    assign layer0_outputs[2943] = (inputs[81]) & (inputs[874]);
    assign layer0_outputs[2944] = ~((inputs[943]) | (inputs[107]));
    assign layer0_outputs[2945] = (inputs[516]) | (inputs[917]);
    assign layer0_outputs[2946] = ~((inputs[451]) | (inputs[684]));
    assign layer0_outputs[2947] = ~(inputs[405]);
    assign layer0_outputs[2948] = ~(inputs[407]);
    assign layer0_outputs[2949] = ~((inputs[1011]) | (inputs[568]));
    assign layer0_outputs[2950] = 1'b0;
    assign layer0_outputs[2951] = ~((inputs[917]) ^ (inputs[532]));
    assign layer0_outputs[2952] = inputs[400];
    assign layer0_outputs[2953] = ~((inputs[811]) ^ (inputs[749]));
    assign layer0_outputs[2954] = ~(inputs[50]) | (inputs[346]);
    assign layer0_outputs[2955] = (inputs[372]) ^ (inputs[893]);
    assign layer0_outputs[2956] = (inputs[878]) | (inputs[975]);
    assign layer0_outputs[2957] = (inputs[52]) | (inputs[251]);
    assign layer0_outputs[2958] = ~(inputs[582]);
    assign layer0_outputs[2959] = (inputs[406]) | (inputs[519]);
    assign layer0_outputs[2960] = ~(inputs[841]) | (inputs[999]);
    assign layer0_outputs[2961] = (inputs[518]) & ~(inputs[734]);
    assign layer0_outputs[2962] = (inputs[716]) & ~(inputs[316]);
    assign layer0_outputs[2963] = (inputs[792]) | (inputs[17]);
    assign layer0_outputs[2964] = inputs[313];
    assign layer0_outputs[2965] = (inputs[723]) ^ (inputs[235]);
    assign layer0_outputs[2966] = ~(inputs[332]) | (inputs[628]);
    assign layer0_outputs[2967] = ~((inputs[156]) | (inputs[603]));
    assign layer0_outputs[2968] = ~(inputs[816]) | (inputs[212]);
    assign layer0_outputs[2969] = ~(inputs[647]);
    assign layer0_outputs[2970] = (inputs[510]) ^ (inputs[997]);
    assign layer0_outputs[2971] = inputs[797];
    assign layer0_outputs[2972] = ~((inputs[843]) ^ (inputs[371]));
    assign layer0_outputs[2973] = inputs[277];
    assign layer0_outputs[2974] = ~((inputs[116]) ^ (inputs[338]));
    assign layer0_outputs[2975] = inputs[283];
    assign layer0_outputs[2976] = ~(inputs[152]);
    assign layer0_outputs[2977] = ~((inputs[68]) ^ (inputs[782]));
    assign layer0_outputs[2978] = (inputs[274]) & ~(inputs[997]);
    assign layer0_outputs[2979] = ~((inputs[700]) | (inputs[482]));
    assign layer0_outputs[2980] = inputs[625];
    assign layer0_outputs[2981] = (inputs[624]) ^ (inputs[47]);
    assign layer0_outputs[2982] = (inputs[632]) & ~(inputs[998]);
    assign layer0_outputs[2983] = inputs[438];
    assign layer0_outputs[2984] = ~((inputs[741]) | (inputs[924]));
    assign layer0_outputs[2985] = 1'b0;
    assign layer0_outputs[2986] = (inputs[312]) ^ (inputs[954]);
    assign layer0_outputs[2987] = ~(inputs[7]) | (inputs[99]);
    assign layer0_outputs[2988] = (inputs[678]) ^ (inputs[664]);
    assign layer0_outputs[2989] = ~((inputs[808]) | (inputs[669]));
    assign layer0_outputs[2990] = (inputs[837]) | (inputs[301]);
    assign layer0_outputs[2991] = ~((inputs[135]) ^ (inputs[883]));
    assign layer0_outputs[2992] = ~(inputs[204]);
    assign layer0_outputs[2993] = ~(inputs[282]);
    assign layer0_outputs[2994] = ~(inputs[120]);
    assign layer0_outputs[2995] = ~(inputs[938]) | (inputs[46]);
    assign layer0_outputs[2996] = ~((inputs[485]) ^ (inputs[98]));
    assign layer0_outputs[2997] = inputs[652];
    assign layer0_outputs[2998] = (inputs[1008]) | (inputs[89]);
    assign layer0_outputs[2999] = (inputs[431]) & (inputs[550]);
    assign layer0_outputs[3000] = 1'b0;
    assign layer0_outputs[3001] = ~(inputs[12]);
    assign layer0_outputs[3002] = ~((inputs[309]) | (inputs[379]));
    assign layer0_outputs[3003] = (inputs[280]) & ~(inputs[383]);
    assign layer0_outputs[3004] = ~(inputs[504]);
    assign layer0_outputs[3005] = (inputs[1]) | (inputs[473]);
    assign layer0_outputs[3006] = ~((inputs[873]) ^ (inputs[104]));
    assign layer0_outputs[3007] = inputs[97];
    assign layer0_outputs[3008] = (inputs[36]) ^ (inputs[788]);
    assign layer0_outputs[3009] = ~((inputs[952]) | (inputs[7]));
    assign layer0_outputs[3010] = (inputs[113]) & ~(inputs[105]);
    assign layer0_outputs[3011] = ~(inputs[790]) | (inputs[571]);
    assign layer0_outputs[3012] = (inputs[1005]) ^ (inputs[533]);
    assign layer0_outputs[3013] = ~(inputs[845]);
    assign layer0_outputs[3014] = (inputs[305]) & ~(inputs[769]);
    assign layer0_outputs[3015] = inputs[840];
    assign layer0_outputs[3016] = inputs[845];
    assign layer0_outputs[3017] = (inputs[869]) | (inputs[202]);
    assign layer0_outputs[3018] = ~(inputs[717]) | (inputs[363]);
    assign layer0_outputs[3019] = inputs[778];
    assign layer0_outputs[3020] = 1'b1;
    assign layer0_outputs[3021] = ~(inputs[717]);
    assign layer0_outputs[3022] = inputs[553];
    assign layer0_outputs[3023] = ~(inputs[239]) | (inputs[732]);
    assign layer0_outputs[3024] = ~((inputs[686]) ^ (inputs[766]));
    assign layer0_outputs[3025] = ~((inputs[411]) | (inputs[378]));
    assign layer0_outputs[3026] = inputs[368];
    assign layer0_outputs[3027] = inputs[971];
    assign layer0_outputs[3028] = (inputs[776]) | (inputs[134]);
    assign layer0_outputs[3029] = ~((inputs[118]) & (inputs[445]));
    assign layer0_outputs[3030] = ~(inputs[266]) | (inputs[921]);
    assign layer0_outputs[3031] = ~(inputs[802]) | (inputs[21]);
    assign layer0_outputs[3032] = ~(inputs[158]);
    assign layer0_outputs[3033] = (inputs[332]) | (inputs[996]);
    assign layer0_outputs[3034] = ~((inputs[454]) | (inputs[935]));
    assign layer0_outputs[3035] = inputs[78];
    assign layer0_outputs[3036] = ~((inputs[231]) & (inputs[919]));
    assign layer0_outputs[3037] = ~((inputs[266]) ^ (inputs[67]));
    assign layer0_outputs[3038] = (inputs[988]) ^ (inputs[417]);
    assign layer0_outputs[3039] = (inputs[459]) & ~(inputs[630]);
    assign layer0_outputs[3040] = inputs[845];
    assign layer0_outputs[3041] = (inputs[307]) | (inputs[958]);
    assign layer0_outputs[3042] = ~(inputs[942]);
    assign layer0_outputs[3043] = (inputs[952]) ^ (inputs[433]);
    assign layer0_outputs[3044] = (inputs[3]) ^ (inputs[572]);
    assign layer0_outputs[3045] = inputs[821];
    assign layer0_outputs[3046] = (inputs[903]) | (inputs[870]);
    assign layer0_outputs[3047] = (inputs[421]) | (inputs[681]);
    assign layer0_outputs[3048] = (inputs[964]) ^ (inputs[773]);
    assign layer0_outputs[3049] = ~((inputs[266]) | (inputs[251]));
    assign layer0_outputs[3050] = inputs[496];
    assign layer0_outputs[3051] = inputs[749];
    assign layer0_outputs[3052] = (inputs[707]) & (inputs[955]);
    assign layer0_outputs[3053] = 1'b1;
    assign layer0_outputs[3054] = inputs[223];
    assign layer0_outputs[3055] = (inputs[251]) & ~(inputs[987]);
    assign layer0_outputs[3056] = (inputs[184]) | (inputs[689]);
    assign layer0_outputs[3057] = inputs[466];
    assign layer0_outputs[3058] = (inputs[298]) ^ (inputs[189]);
    assign layer0_outputs[3059] = ~((inputs[56]) | (inputs[401]));
    assign layer0_outputs[3060] = ~((inputs[169]) | (inputs[475]));
    assign layer0_outputs[3061] = (inputs[768]) ^ (inputs[445]);
    assign layer0_outputs[3062] = 1'b1;
    assign layer0_outputs[3063] = (inputs[610]) ^ (inputs[554]);
    assign layer0_outputs[3064] = ~((inputs[654]) ^ (inputs[618]));
    assign layer0_outputs[3065] = (inputs[164]) & ~(inputs[972]);
    assign layer0_outputs[3066] = (inputs[427]) & (inputs[919]);
    assign layer0_outputs[3067] = inputs[495];
    assign layer0_outputs[3068] = ~(inputs[812]) | (inputs[486]);
    assign layer0_outputs[3069] = ~(inputs[441]);
    assign layer0_outputs[3070] = ~(inputs[430]);
    assign layer0_outputs[3071] = (inputs[889]) & ~(inputs[249]);
    assign layer0_outputs[3072] = ~((inputs[232]) ^ (inputs[19]));
    assign layer0_outputs[3073] = (inputs[394]) & ~(inputs[183]);
    assign layer0_outputs[3074] = inputs[164];
    assign layer0_outputs[3075] = ~(inputs[80]) | (inputs[887]);
    assign layer0_outputs[3076] = ~((inputs[50]) | (inputs[202]));
    assign layer0_outputs[3077] = (inputs[377]) & (inputs[699]);
    assign layer0_outputs[3078] = ~(inputs[311]) | (inputs[898]);
    assign layer0_outputs[3079] = inputs[715];
    assign layer0_outputs[3080] = ~(inputs[696]) | (inputs[904]);
    assign layer0_outputs[3081] = ~(inputs[977]);
    assign layer0_outputs[3082] = ~((inputs[732]) | (inputs[950]));
    assign layer0_outputs[3083] = ~((inputs[161]) | (inputs[65]));
    assign layer0_outputs[3084] = (inputs[673]) & ~(inputs[480]);
    assign layer0_outputs[3085] = (inputs[501]) | (inputs[1002]);
    assign layer0_outputs[3086] = 1'b1;
    assign layer0_outputs[3087] = (inputs[23]) | (inputs[123]);
    assign layer0_outputs[3088] = ~(inputs[669]);
    assign layer0_outputs[3089] = inputs[346];
    assign layer0_outputs[3090] = inputs[652];
    assign layer0_outputs[3091] = ~(inputs[680]);
    assign layer0_outputs[3092] = ~((inputs[474]) | (inputs[684]));
    assign layer0_outputs[3093] = ~(inputs[924]) | (inputs[698]);
    assign layer0_outputs[3094] = ~(inputs[595]);
    assign layer0_outputs[3095] = ~(inputs[887]) | (inputs[641]);
    assign layer0_outputs[3096] = (inputs[80]) ^ (inputs[221]);
    assign layer0_outputs[3097] = 1'b1;
    assign layer0_outputs[3098] = inputs[728];
    assign layer0_outputs[3099] = ~((inputs[780]) | (inputs[988]));
    assign layer0_outputs[3100] = (inputs[834]) & ~(inputs[735]);
    assign layer0_outputs[3101] = inputs[704];
    assign layer0_outputs[3102] = (inputs[879]) | (inputs[360]);
    assign layer0_outputs[3103] = ~(inputs[973]);
    assign layer0_outputs[3104] = 1'b0;
    assign layer0_outputs[3105] = (inputs[443]) & ~(inputs[320]);
    assign layer0_outputs[3106] = ~(inputs[994]) | (inputs[316]);
    assign layer0_outputs[3107] = ~((inputs[993]) | (inputs[813]));
    assign layer0_outputs[3108] = (inputs[183]) | (inputs[753]);
    assign layer0_outputs[3109] = (inputs[667]) & (inputs[350]);
    assign layer0_outputs[3110] = ~(inputs[156]) | (inputs[941]);
    assign layer0_outputs[3111] = (inputs[882]) | (inputs[986]);
    assign layer0_outputs[3112] = (inputs[607]) | (inputs[270]);
    assign layer0_outputs[3113] = ~(inputs[845]);
    assign layer0_outputs[3114] = ~((inputs[413]) | (inputs[848]));
    assign layer0_outputs[3115] = (inputs[436]) & ~(inputs[392]);
    assign layer0_outputs[3116] = ~(inputs[775]) | (inputs[926]);
    assign layer0_outputs[3117] = ~(inputs[489]);
    assign layer0_outputs[3118] = 1'b1;
    assign layer0_outputs[3119] = ~(inputs[635]);
    assign layer0_outputs[3120] = ~(inputs[335]) | (inputs[836]);
    assign layer0_outputs[3121] = (inputs[58]) & (inputs[222]);
    assign layer0_outputs[3122] = ~(inputs[280]);
    assign layer0_outputs[3123] = (inputs[515]) & (inputs[769]);
    assign layer0_outputs[3124] = (inputs[90]) | (inputs[858]);
    assign layer0_outputs[3125] = (inputs[964]) & ~(inputs[735]);
    assign layer0_outputs[3126] = ~((inputs[792]) | (inputs[268]));
    assign layer0_outputs[3127] = (inputs[152]) & ~(inputs[290]);
    assign layer0_outputs[3128] = inputs[495];
    assign layer0_outputs[3129] = (inputs[624]) & ~(inputs[268]);
    assign layer0_outputs[3130] = ~((inputs[327]) | (inputs[689]));
    assign layer0_outputs[3131] = (inputs[375]) & ~(inputs[58]);
    assign layer0_outputs[3132] = ~(inputs[821]) | (inputs[770]);
    assign layer0_outputs[3133] = (inputs[295]) & (inputs[448]);
    assign layer0_outputs[3134] = (inputs[388]) & ~(inputs[305]);
    assign layer0_outputs[3135] = ~(inputs[411]);
    assign layer0_outputs[3136] = inputs[331];
    assign layer0_outputs[3137] = inputs[18];
    assign layer0_outputs[3138] = ~(inputs[216]) | (inputs[1001]);
    assign layer0_outputs[3139] = ~(inputs[168]);
    assign layer0_outputs[3140] = ~((inputs[52]) ^ (inputs[690]));
    assign layer0_outputs[3141] = (inputs[299]) & ~(inputs[256]);
    assign layer0_outputs[3142] = ~(inputs[463]);
    assign layer0_outputs[3143] = ~((inputs[181]) | (inputs[128]));
    assign layer0_outputs[3144] = ~((inputs[719]) ^ (inputs[780]));
    assign layer0_outputs[3145] = (inputs[937]) & ~(inputs[90]);
    assign layer0_outputs[3146] = ~((inputs[52]) & (inputs[329]));
    assign layer0_outputs[3147] = inputs[540];
    assign layer0_outputs[3148] = ~(inputs[819]);
    assign layer0_outputs[3149] = ~((inputs[96]) | (inputs[941]));
    assign layer0_outputs[3150] = ~(inputs[993]) | (inputs[774]);
    assign layer0_outputs[3151] = ~((inputs[539]) ^ (inputs[735]));
    assign layer0_outputs[3152] = inputs[67];
    assign layer0_outputs[3153] = ~(inputs[884]) | (inputs[607]);
    assign layer0_outputs[3154] = inputs[786];
    assign layer0_outputs[3155] = 1'b1;
    assign layer0_outputs[3156] = (inputs[633]) ^ (inputs[176]);
    assign layer0_outputs[3157] = ~((inputs[557]) | (inputs[362]));
    assign layer0_outputs[3158] = ~(inputs[845]);
    assign layer0_outputs[3159] = ~(inputs[596]);
    assign layer0_outputs[3160] = ~((inputs[718]) ^ (inputs[1003]));
    assign layer0_outputs[3161] = (inputs[354]) & ~(inputs[639]);
    assign layer0_outputs[3162] = 1'b0;
    assign layer0_outputs[3163] = ~((inputs[347]) | (inputs[370]));
    assign layer0_outputs[3164] = (inputs[731]) & ~(inputs[960]);
    assign layer0_outputs[3165] = (inputs[1010]) | (inputs[8]);
    assign layer0_outputs[3166] = (inputs[846]) | (inputs[18]);
    assign layer0_outputs[3167] = ~(inputs[645]) | (inputs[747]);
    assign layer0_outputs[3168] = ~((inputs[630]) | (inputs[628]));
    assign layer0_outputs[3169] = inputs[169];
    assign layer0_outputs[3170] = ~(inputs[922]) | (inputs[369]);
    assign layer0_outputs[3171] = ~(inputs[345]);
    assign layer0_outputs[3172] = ~(inputs[161]);
    assign layer0_outputs[3173] = ~((inputs[714]) ^ (inputs[427]));
    assign layer0_outputs[3174] = (inputs[476]) | (inputs[571]);
    assign layer0_outputs[3175] = (inputs[330]) ^ (inputs[775]);
    assign layer0_outputs[3176] = ~(inputs[540]) | (inputs[143]);
    assign layer0_outputs[3177] = ~(inputs[541]);
    assign layer0_outputs[3178] = (inputs[154]) | (inputs[430]);
    assign layer0_outputs[3179] = (inputs[678]) & (inputs[856]);
    assign layer0_outputs[3180] = (inputs[699]) | (inputs[742]);
    assign layer0_outputs[3181] = ~((inputs[697]) ^ (inputs[78]));
    assign layer0_outputs[3182] = (inputs[164]) | (inputs[545]);
    assign layer0_outputs[3183] = (inputs[602]) ^ (inputs[55]);
    assign layer0_outputs[3184] = inputs[580];
    assign layer0_outputs[3185] = ~((inputs[1001]) | (inputs[304]));
    assign layer0_outputs[3186] = (inputs[71]) ^ (inputs[278]);
    assign layer0_outputs[3187] = ~((inputs[629]) | (inputs[283]));
    assign layer0_outputs[3188] = ~(inputs[426]) | (inputs[479]);
    assign layer0_outputs[3189] = ~(inputs[986]) | (inputs[113]);
    assign layer0_outputs[3190] = (inputs[698]) & ~(inputs[158]);
    assign layer0_outputs[3191] = ~((inputs[444]) | (inputs[654]));
    assign layer0_outputs[3192] = inputs[339];
    assign layer0_outputs[3193] = ~((inputs[69]) ^ (inputs[265]));
    assign layer0_outputs[3194] = inputs[590];
    assign layer0_outputs[3195] = (inputs[985]) ^ (inputs[999]);
    assign layer0_outputs[3196] = ~(inputs[551]);
    assign layer0_outputs[3197] = ~((inputs[840]) & (inputs[478]));
    assign layer0_outputs[3198] = ~(inputs[653]) | (inputs[179]);
    assign layer0_outputs[3199] = ~((inputs[1011]) ^ (inputs[576]));
    assign layer0_outputs[3200] = (inputs[565]) & ~(inputs[45]);
    assign layer0_outputs[3201] = inputs[782];
    assign layer0_outputs[3202] = ~(inputs[1022]) | (inputs[191]);
    assign layer0_outputs[3203] = inputs[751];
    assign layer0_outputs[3204] = inputs[79];
    assign layer0_outputs[3205] = ~((inputs[795]) | (inputs[835]));
    assign layer0_outputs[3206] = inputs[506];
    assign layer0_outputs[3207] = ~((inputs[528]) ^ (inputs[937]));
    assign layer0_outputs[3208] = (inputs[888]) ^ (inputs[3]);
    assign layer0_outputs[3209] = inputs[752];
    assign layer0_outputs[3210] = ~((inputs[978]) | (inputs[751]));
    assign layer0_outputs[3211] = (inputs[749]) & ~(inputs[162]);
    assign layer0_outputs[3212] = inputs[956];
    assign layer0_outputs[3213] = ~((inputs[807]) | (inputs[162]));
    assign layer0_outputs[3214] = (inputs[281]) | (inputs[727]);
    assign layer0_outputs[3215] = ~((inputs[395]) ^ (inputs[26]));
    assign layer0_outputs[3216] = (inputs[540]) & (inputs[355]);
    assign layer0_outputs[3217] = ~((inputs[270]) | (inputs[105]));
    assign layer0_outputs[3218] = (inputs[725]) & ~(inputs[443]);
    assign layer0_outputs[3219] = ~((inputs[577]) | (inputs[191]));
    assign layer0_outputs[3220] = ~(inputs[786]);
    assign layer0_outputs[3221] = (inputs[552]) & ~(inputs[998]);
    assign layer0_outputs[3222] = ~((inputs[673]) ^ (inputs[777]));
    assign layer0_outputs[3223] = ~(inputs[396]);
    assign layer0_outputs[3224] = ~((inputs[146]) ^ (inputs[962]));
    assign layer0_outputs[3225] = ~(inputs[923]);
    assign layer0_outputs[3226] = ~(inputs[454]) | (inputs[807]);
    assign layer0_outputs[3227] = (inputs[868]) & ~(inputs[57]);
    assign layer0_outputs[3228] = ~(inputs[935]) | (inputs[836]);
    assign layer0_outputs[3229] = (inputs[784]) & ~(inputs[403]);
    assign layer0_outputs[3230] = (inputs[530]) & ~(inputs[403]);
    assign layer0_outputs[3231] = (inputs[786]) | (inputs[714]);
    assign layer0_outputs[3232] = (inputs[861]) | (inputs[148]);
    assign layer0_outputs[3233] = ~(inputs[397]);
    assign layer0_outputs[3234] = (inputs[858]) & ~(inputs[290]);
    assign layer0_outputs[3235] = ~(inputs[747]) | (inputs[950]);
    assign layer0_outputs[3236] = (inputs[529]) & ~(inputs[731]);
    assign layer0_outputs[3237] = (inputs[121]) | (inputs[331]);
    assign layer0_outputs[3238] = ~((inputs[135]) & (inputs[146]));
    assign layer0_outputs[3239] = 1'b1;
    assign layer0_outputs[3240] = inputs[368];
    assign layer0_outputs[3241] = (inputs[39]) ^ (inputs[573]);
    assign layer0_outputs[3242] = (inputs[757]) & (inputs[848]);
    assign layer0_outputs[3243] = (inputs[344]) & ~(inputs[79]);
    assign layer0_outputs[3244] = ~((inputs[573]) | (inputs[172]));
    assign layer0_outputs[3245] = 1'b0;
    assign layer0_outputs[3246] = ~(inputs[116]) | (inputs[574]);
    assign layer0_outputs[3247] = (inputs[903]) & (inputs[994]);
    assign layer0_outputs[3248] = (inputs[680]) | (inputs[804]);
    assign layer0_outputs[3249] = inputs[1000];
    assign layer0_outputs[3250] = (inputs[36]) & ~(inputs[317]);
    assign layer0_outputs[3251] = ~((inputs[324]) | (inputs[482]));
    assign layer0_outputs[3252] = (inputs[763]) ^ (inputs[866]);
    assign layer0_outputs[3253] = ~((inputs[295]) ^ (inputs[564]));
    assign layer0_outputs[3254] = ~((inputs[213]) & (inputs[102]));
    assign layer0_outputs[3255] = ~(inputs[342]);
    assign layer0_outputs[3256] = ~(inputs[518]);
    assign layer0_outputs[3257] = (inputs[750]) & ~(inputs[486]);
    assign layer0_outputs[3258] = ~(inputs[437]);
    assign layer0_outputs[3259] = (inputs[353]) & ~(inputs[866]);
    assign layer0_outputs[3260] = (inputs[918]) & (inputs[989]);
    assign layer0_outputs[3261] = inputs[375];
    assign layer0_outputs[3262] = (inputs[777]) ^ (inputs[862]);
    assign layer0_outputs[3263] = ~(inputs[145]);
    assign layer0_outputs[3264] = inputs[695];
    assign layer0_outputs[3265] = ~((inputs[369]) | (inputs[1007]));
    assign layer0_outputs[3266] = ~((inputs[37]) ^ (inputs[13]));
    assign layer0_outputs[3267] = inputs[300];
    assign layer0_outputs[3268] = ~((inputs[501]) ^ (inputs[830]));
    assign layer0_outputs[3269] = (inputs[726]) & ~(inputs[823]);
    assign layer0_outputs[3270] = (inputs[425]) | (inputs[956]);
    assign layer0_outputs[3271] = (inputs[524]) | (inputs[494]);
    assign layer0_outputs[3272] = (inputs[261]) | (inputs[439]);
    assign layer0_outputs[3273] = (inputs[717]) & ~(inputs[379]);
    assign layer0_outputs[3274] = (inputs[641]) & (inputs[50]);
    assign layer0_outputs[3275] = (inputs[342]) & ~(inputs[996]);
    assign layer0_outputs[3276] = 1'b0;
    assign layer0_outputs[3277] = (inputs[969]) ^ (inputs[517]);
    assign layer0_outputs[3278] = ~(inputs[52]);
    assign layer0_outputs[3279] = (inputs[456]) & ~(inputs[874]);
    assign layer0_outputs[3280] = (inputs[266]) & (inputs[864]);
    assign layer0_outputs[3281] = (inputs[996]) & (inputs[982]);
    assign layer0_outputs[3282] = 1'b0;
    assign layer0_outputs[3283] = ~(inputs[241]);
    assign layer0_outputs[3284] = (inputs[611]) ^ (inputs[985]);
    assign layer0_outputs[3285] = ~((inputs[554]) ^ (inputs[897]));
    assign layer0_outputs[3286] = (inputs[1016]) | (inputs[336]);
    assign layer0_outputs[3287] = (inputs[760]) ^ (inputs[906]);
    assign layer0_outputs[3288] = (inputs[158]) & ~(inputs[143]);
    assign layer0_outputs[3289] = ~(inputs[416]) | (inputs[870]);
    assign layer0_outputs[3290] = ~(inputs[16]) | (inputs[121]);
    assign layer0_outputs[3291] = ~(inputs[167]);
    assign layer0_outputs[3292] = ~(inputs[60]);
    assign layer0_outputs[3293] = ~((inputs[857]) ^ (inputs[910]));
    assign layer0_outputs[3294] = (inputs[267]) & (inputs[768]);
    assign layer0_outputs[3295] = ~(inputs[366]) | (inputs[681]);
    assign layer0_outputs[3296] = ~((inputs[994]) | (inputs[808]));
    assign layer0_outputs[3297] = (inputs[584]) & ~(inputs[607]);
    assign layer0_outputs[3298] = (inputs[973]) | (inputs[301]);
    assign layer0_outputs[3299] = inputs[130];
    assign layer0_outputs[3300] = 1'b0;
    assign layer0_outputs[3301] = (inputs[887]) ^ (inputs[213]);
    assign layer0_outputs[3302] = inputs[623];
    assign layer0_outputs[3303] = ~((inputs[836]) & (inputs[276]));
    assign layer0_outputs[3304] = ~(inputs[23]);
    assign layer0_outputs[3305] = (inputs[959]) & (inputs[109]);
    assign layer0_outputs[3306] = ~(inputs[664]);
    assign layer0_outputs[3307] = ~((inputs[784]) | (inputs[329]));
    assign layer0_outputs[3308] = ~((inputs[838]) & (inputs[93]));
    assign layer0_outputs[3309] = ~((inputs[1003]) & (inputs[855]));
    assign layer0_outputs[3310] = ~(inputs[85]) | (inputs[914]);
    assign layer0_outputs[3311] = ~((inputs[231]) | (inputs[752]));
    assign layer0_outputs[3312] = 1'b0;
    assign layer0_outputs[3313] = ~((inputs[148]) ^ (inputs[593]));
    assign layer0_outputs[3314] = ~((inputs[661]) ^ (inputs[859]));
    assign layer0_outputs[3315] = (inputs[662]) | (inputs[243]);
    assign layer0_outputs[3316] = inputs[724];
    assign layer0_outputs[3317] = ~(inputs[674]) | (inputs[86]);
    assign layer0_outputs[3318] = (inputs[644]) ^ (inputs[481]);
    assign layer0_outputs[3319] = ~(inputs[159]);
    assign layer0_outputs[3320] = (inputs[756]) ^ (inputs[580]);
    assign layer0_outputs[3321] = 1'b0;
    assign layer0_outputs[3322] = ~((inputs[935]) | (inputs[724]));
    assign layer0_outputs[3323] = ~((inputs[815]) ^ (inputs[403]));
    assign layer0_outputs[3324] = ~(inputs[979]) | (inputs[293]);
    assign layer0_outputs[3325] = (inputs[542]) ^ (inputs[172]);
    assign layer0_outputs[3326] = (inputs[547]) | (inputs[612]);
    assign layer0_outputs[3327] = ~(inputs[293]) | (inputs[83]);
    assign layer0_outputs[3328] = ~((inputs[765]) | (inputs[918]));
    assign layer0_outputs[3329] = (inputs[619]) ^ (inputs[802]);
    assign layer0_outputs[3330] = (inputs[250]) & (inputs[760]);
    assign layer0_outputs[3331] = (inputs[133]) | (inputs[337]);
    assign layer0_outputs[3332] = ~(inputs[987]);
    assign layer0_outputs[3333] = ~(inputs[110]);
    assign layer0_outputs[3334] = ~((inputs[421]) | (inputs[703]));
    assign layer0_outputs[3335] = ~((inputs[893]) | (inputs[788]));
    assign layer0_outputs[3336] = ~(inputs[97]);
    assign layer0_outputs[3337] = (inputs[797]) & ~(inputs[326]);
    assign layer0_outputs[3338] = inputs[713];
    assign layer0_outputs[3339] = ~(inputs[54]);
    assign layer0_outputs[3340] = (inputs[365]) ^ (inputs[571]);
    assign layer0_outputs[3341] = ~(inputs[213]) | (inputs[187]);
    assign layer0_outputs[3342] = ~(inputs[376]);
    assign layer0_outputs[3343] = (inputs[536]) & ~(inputs[916]);
    assign layer0_outputs[3344] = (inputs[609]) | (inputs[344]);
    assign layer0_outputs[3345] = ~(inputs[359]) | (inputs[1002]);
    assign layer0_outputs[3346] = (inputs[131]) ^ (inputs[600]);
    assign layer0_outputs[3347] = ~((inputs[876]) | (inputs[49]));
    assign layer0_outputs[3348] = ~((inputs[666]) | (inputs[695]));
    assign layer0_outputs[3349] = (inputs[989]) ^ (inputs[614]);
    assign layer0_outputs[3350] = ~(inputs[655]);
    assign layer0_outputs[3351] = ~(inputs[141]);
    assign layer0_outputs[3352] = (inputs[397]) ^ (inputs[681]);
    assign layer0_outputs[3353] = ~(inputs[812]);
    assign layer0_outputs[3354] = (inputs[123]) & (inputs[100]);
    assign layer0_outputs[3355] = 1'b1;
    assign layer0_outputs[3356] = ~((inputs[726]) ^ (inputs[1005]));
    assign layer0_outputs[3357] = ~(inputs[391]);
    assign layer0_outputs[3358] = ~(inputs[810]) | (inputs[612]);
    assign layer0_outputs[3359] = ~((inputs[234]) ^ (inputs[988]));
    assign layer0_outputs[3360] = (inputs[323]) ^ (inputs[609]);
    assign layer0_outputs[3361] = (inputs[85]) ^ (inputs[840]);
    assign layer0_outputs[3362] = ~((inputs[481]) | (inputs[565]));
    assign layer0_outputs[3363] = inputs[719];
    assign layer0_outputs[3364] = (inputs[847]) ^ (inputs[222]);
    assign layer0_outputs[3365] = ~((inputs[355]) | (inputs[502]));
    assign layer0_outputs[3366] = (inputs[362]) ^ (inputs[477]);
    assign layer0_outputs[3367] = ~((inputs[704]) | (inputs[218]));
    assign layer0_outputs[3368] = ~(inputs[402]) | (inputs[313]);
    assign layer0_outputs[3369] = (inputs[950]) & ~(inputs[1016]);
    assign layer0_outputs[3370] = inputs[284];
    assign layer0_outputs[3371] = 1'b0;
    assign layer0_outputs[3372] = (inputs[859]) | (inputs[502]);
    assign layer0_outputs[3373] = ~((inputs[542]) | (inputs[871]));
    assign layer0_outputs[3374] = (inputs[304]) & ~(inputs[281]);
    assign layer0_outputs[3375] = ~(inputs[320]) | (inputs[263]);
    assign layer0_outputs[3376] = (inputs[620]) ^ (inputs[216]);
    assign layer0_outputs[3377] = inputs[22];
    assign layer0_outputs[3378] = (inputs[238]) | (inputs[364]);
    assign layer0_outputs[3379] = (inputs[932]) | (inputs[76]);
    assign layer0_outputs[3380] = ~((inputs[573]) ^ (inputs[167]));
    assign layer0_outputs[3381] = (inputs[888]) | (inputs[211]);
    assign layer0_outputs[3382] = (inputs[853]) & ~(inputs[73]);
    assign layer0_outputs[3383] = ~((inputs[845]) ^ (inputs[749]));
    assign layer0_outputs[3384] = ~(inputs[490]);
    assign layer0_outputs[3385] = ~(inputs[199]);
    assign layer0_outputs[3386] = ~(inputs[463]);
    assign layer0_outputs[3387] = inputs[867];
    assign layer0_outputs[3388] = inputs[599];
    assign layer0_outputs[3389] = ~((inputs[960]) | (inputs[572]));
    assign layer0_outputs[3390] = ~(inputs[15]);
    assign layer0_outputs[3391] = ~((inputs[760]) ^ (inputs[768]));
    assign layer0_outputs[3392] = (inputs[288]) & ~(inputs[442]);
    assign layer0_outputs[3393] = inputs[707];
    assign layer0_outputs[3394] = (inputs[812]) & ~(inputs[829]);
    assign layer0_outputs[3395] = ~(inputs[241]);
    assign layer0_outputs[3396] = ~((inputs[702]) | (inputs[979]));
    assign layer0_outputs[3397] = ~(inputs[741]);
    assign layer0_outputs[3398] = (inputs[466]) & ~(inputs[349]);
    assign layer0_outputs[3399] = (inputs[231]) | (inputs[563]);
    assign layer0_outputs[3400] = (inputs[591]) | (inputs[452]);
    assign layer0_outputs[3401] = (inputs[94]) & (inputs[958]);
    assign layer0_outputs[3402] = ~((inputs[123]) ^ (inputs[879]));
    assign layer0_outputs[3403] = 1'b0;
    assign layer0_outputs[3404] = ~(inputs[527]);
    assign layer0_outputs[3405] = (inputs[211]) & ~(inputs[387]);
    assign layer0_outputs[3406] = (inputs[287]) & (inputs[65]);
    assign layer0_outputs[3407] = (inputs[152]) ^ (inputs[79]);
    assign layer0_outputs[3408] = (inputs[220]) & ~(inputs[907]);
    assign layer0_outputs[3409] = inputs[983];
    assign layer0_outputs[3410] = (inputs[185]) & ~(inputs[641]);
    assign layer0_outputs[3411] = ~((inputs[377]) | (inputs[717]));
    assign layer0_outputs[3412] = ~(inputs[438]) | (inputs[907]);
    assign layer0_outputs[3413] = (inputs[474]) | (inputs[329]);
    assign layer0_outputs[3414] = ~(inputs[265]);
    assign layer0_outputs[3415] = (inputs[1000]) ^ (inputs[612]);
    assign layer0_outputs[3416] = (inputs[594]) & ~(inputs[143]);
    assign layer0_outputs[3417] = 1'b0;
    assign layer0_outputs[3418] = (inputs[661]) ^ (inputs[263]);
    assign layer0_outputs[3419] = (inputs[431]) ^ (inputs[797]);
    assign layer0_outputs[3420] = ~((inputs[631]) ^ (inputs[642]));
    assign layer0_outputs[3421] = (inputs[938]) | (inputs[405]);
    assign layer0_outputs[3422] = (inputs[128]) & ~(inputs[611]);
    assign layer0_outputs[3423] = ~((inputs[278]) ^ (inputs[57]));
    assign layer0_outputs[3424] = ~((inputs[438]) | (inputs[121]));
    assign layer0_outputs[3425] = (inputs[631]) ^ (inputs[793]);
    assign layer0_outputs[3426] = 1'b0;
    assign layer0_outputs[3427] = ~(inputs[73]);
    assign layer0_outputs[3428] = (inputs[102]) ^ (inputs[739]);
    assign layer0_outputs[3429] = ~((inputs[87]) | (inputs[750]));
    assign layer0_outputs[3430] = ~((inputs[810]) | (inputs[388]));
    assign layer0_outputs[3431] = ~((inputs[990]) | (inputs[363]));
    assign layer0_outputs[3432] = ~((inputs[115]) | (inputs[565]));
    assign layer0_outputs[3433] = (inputs[525]) ^ (inputs[634]);
    assign layer0_outputs[3434] = ~((inputs[411]) | (inputs[143]));
    assign layer0_outputs[3435] = inputs[202];
    assign layer0_outputs[3436] = (inputs[722]) & ~(inputs[998]);
    assign layer0_outputs[3437] = ~((inputs[490]) ^ (inputs[68]));
    assign layer0_outputs[3438] = ~((inputs[595]) | (inputs[308]));
    assign layer0_outputs[3439] = (inputs[600]) & ~(inputs[936]);
    assign layer0_outputs[3440] = (inputs[300]) | (inputs[727]);
    assign layer0_outputs[3441] = ~((inputs[25]) | (inputs[20]));
    assign layer0_outputs[3442] = (inputs[535]) | (inputs[189]);
    assign layer0_outputs[3443] = (inputs[309]) & ~(inputs[124]);
    assign layer0_outputs[3444] = inputs[269];
    assign layer0_outputs[3445] = (inputs[828]) ^ (inputs[364]);
    assign layer0_outputs[3446] = ~(inputs[496]) | (inputs[1003]);
    assign layer0_outputs[3447] = ~((inputs[820]) | (inputs[898]));
    assign layer0_outputs[3448] = (inputs[177]) | (inputs[742]);
    assign layer0_outputs[3449] = inputs[724];
    assign layer0_outputs[3450] = (inputs[169]) & ~(inputs[381]);
    assign layer0_outputs[3451] = (inputs[592]) & ~(inputs[556]);
    assign layer0_outputs[3452] = 1'b1;
    assign layer0_outputs[3453] = ~(inputs[740]);
    assign layer0_outputs[3454] = ~(inputs[403]);
    assign layer0_outputs[3455] = ~((inputs[780]) | (inputs[680]));
    assign layer0_outputs[3456] = inputs[632];
    assign layer0_outputs[3457] = (inputs[880]) | (inputs[963]);
    assign layer0_outputs[3458] = ~((inputs[974]) | (inputs[966]));
    assign layer0_outputs[3459] = inputs[903];
    assign layer0_outputs[3460] = ~((inputs[835]) & (inputs[44]));
    assign layer0_outputs[3461] = (inputs[657]) & ~(inputs[965]);
    assign layer0_outputs[3462] = (inputs[891]) | (inputs[716]);
    assign layer0_outputs[3463] = ~(inputs[333]);
    assign layer0_outputs[3464] = ~(inputs[5]) | (inputs[783]);
    assign layer0_outputs[3465] = inputs[456];
    assign layer0_outputs[3466] = ~(inputs[402]);
    assign layer0_outputs[3467] = (inputs[52]) | (inputs[755]);
    assign layer0_outputs[3468] = inputs[523];
    assign layer0_outputs[3469] = (inputs[312]) | (inputs[634]);
    assign layer0_outputs[3470] = ~(inputs[774]) | (inputs[451]);
    assign layer0_outputs[3471] = 1'b0;
    assign layer0_outputs[3472] = (inputs[256]) ^ (inputs[199]);
    assign layer0_outputs[3473] = (inputs[701]) & (inputs[260]);
    assign layer0_outputs[3474] = ~((inputs[132]) ^ (inputs[366]));
    assign layer0_outputs[3475] = (inputs[669]) & ~(inputs[826]);
    assign layer0_outputs[3476] = ~(inputs[814]) | (inputs[147]);
    assign layer0_outputs[3477] = ~(inputs[786]) | (inputs[328]);
    assign layer0_outputs[3478] = ~(inputs[934]);
    assign layer0_outputs[3479] = ~(inputs[713]);
    assign layer0_outputs[3480] = ~((inputs[808]) ^ (inputs[970]));
    assign layer0_outputs[3481] = (inputs[991]) & ~(inputs[348]);
    assign layer0_outputs[3482] = (inputs[585]) ^ (inputs[460]);
    assign layer0_outputs[3483] = (inputs[1007]) & (inputs[899]);
    assign layer0_outputs[3484] = (inputs[922]) & ~(inputs[1011]);
    assign layer0_outputs[3485] = (inputs[968]) ^ (inputs[1008]);
    assign layer0_outputs[3486] = (inputs[22]) ^ (inputs[946]);
    assign layer0_outputs[3487] = ~((inputs[962]) ^ (inputs[607]));
    assign layer0_outputs[3488] = ~(inputs[790]) | (inputs[865]);
    assign layer0_outputs[3489] = inputs[372];
    assign layer0_outputs[3490] = ~((inputs[744]) | (inputs[270]));
    assign layer0_outputs[3491] = 1'b1;
    assign layer0_outputs[3492] = (inputs[206]) ^ (inputs[867]);
    assign layer0_outputs[3493] = (inputs[586]) | (inputs[54]);
    assign layer0_outputs[3494] = (inputs[331]) ^ (inputs[41]);
    assign layer0_outputs[3495] = (inputs[360]) & ~(inputs[447]);
    assign layer0_outputs[3496] = (inputs[35]) | (inputs[852]);
    assign layer0_outputs[3497] = inputs[393];
    assign layer0_outputs[3498] = (inputs[681]) & ~(inputs[230]);
    assign layer0_outputs[3499] = inputs[563];
    assign layer0_outputs[3500] = (inputs[615]) & (inputs[974]);
    assign layer0_outputs[3501] = (inputs[471]) & ~(inputs[857]);
    assign layer0_outputs[3502] = (inputs[187]) | (inputs[247]);
    assign layer0_outputs[3503] = (inputs[686]) & (inputs[656]);
    assign layer0_outputs[3504] = ~(inputs[589]) | (inputs[164]);
    assign layer0_outputs[3505] = (inputs[600]) & (inputs[728]);
    assign layer0_outputs[3506] = ~(inputs[612]);
    assign layer0_outputs[3507] = (inputs[846]) & ~(inputs[19]);
    assign layer0_outputs[3508] = ~((inputs[490]) ^ (inputs[63]));
    assign layer0_outputs[3509] = ~((inputs[741]) | (inputs[431]));
    assign layer0_outputs[3510] = ~(inputs[753]) | (inputs[452]);
    assign layer0_outputs[3511] = (inputs[893]) & (inputs[865]);
    assign layer0_outputs[3512] = inputs[87];
    assign layer0_outputs[3513] = ~(inputs[967]);
    assign layer0_outputs[3514] = inputs[565];
    assign layer0_outputs[3515] = ~(inputs[956]) | (inputs[709]);
    assign layer0_outputs[3516] = inputs[912];
    assign layer0_outputs[3517] = (inputs[48]) | (inputs[353]);
    assign layer0_outputs[3518] = (inputs[409]) & (inputs[441]);
    assign layer0_outputs[3519] = (inputs[282]) & ~(inputs[123]);
    assign layer0_outputs[3520] = ~(inputs[312]) | (inputs[83]);
    assign layer0_outputs[3521] = (inputs[530]) ^ (inputs[257]);
    assign layer0_outputs[3522] = ~(inputs[541]);
    assign layer0_outputs[3523] = ~(inputs[64]);
    assign layer0_outputs[3524] = 1'b1;
    assign layer0_outputs[3525] = ~((inputs[405]) ^ (inputs[355]));
    assign layer0_outputs[3526] = ~(inputs[265]);
    assign layer0_outputs[3527] = inputs[275];
    assign layer0_outputs[3528] = 1'b1;
    assign layer0_outputs[3529] = inputs[24];
    assign layer0_outputs[3530] = (inputs[37]) ^ (inputs[783]);
    assign layer0_outputs[3531] = ~(inputs[957]) | (inputs[328]);
    assign layer0_outputs[3532] = ~((inputs[750]) ^ (inputs[813]));
    assign layer0_outputs[3533] = inputs[242];
    assign layer0_outputs[3534] = 1'b0;
    assign layer0_outputs[3535] = 1'b0;
    assign layer0_outputs[3536] = inputs[631];
    assign layer0_outputs[3537] = ~(inputs[503]) | (inputs[131]);
    assign layer0_outputs[3538] = ~((inputs[824]) | (inputs[1023]));
    assign layer0_outputs[3539] = ~((inputs[130]) | (inputs[503]));
    assign layer0_outputs[3540] = ~(inputs[276]) | (inputs[256]);
    assign layer0_outputs[3541] = ~((inputs[927]) ^ (inputs[477]));
    assign layer0_outputs[3542] = ~((inputs[379]) | (inputs[496]));
    assign layer0_outputs[3543] = (inputs[337]) & ~(inputs[779]);
    assign layer0_outputs[3544] = inputs[437];
    assign layer0_outputs[3545] = 1'b0;
    assign layer0_outputs[3546] = ~(inputs[130]);
    assign layer0_outputs[3547] = inputs[41];
    assign layer0_outputs[3548] = ~(inputs[108]) | (inputs[736]);
    assign layer0_outputs[3549] = ~((inputs[851]) | (inputs[58]));
    assign layer0_outputs[3550] = (inputs[959]) & ~(inputs[352]);
    assign layer0_outputs[3551] = (inputs[235]) | (inputs[296]);
    assign layer0_outputs[3552] = inputs[815];
    assign layer0_outputs[3553] = (inputs[485]) ^ (inputs[934]);
    assign layer0_outputs[3554] = ~((inputs[860]) | (inputs[912]));
    assign layer0_outputs[3555] = ~((inputs[97]) ^ (inputs[95]));
    assign layer0_outputs[3556] = ~(inputs[728]);
    assign layer0_outputs[3557] = (inputs[711]) & ~(inputs[4]);
    assign layer0_outputs[3558] = ~(inputs[149]) | (inputs[70]);
    assign layer0_outputs[3559] = (inputs[597]) | (inputs[494]);
    assign layer0_outputs[3560] = (inputs[860]) | (inputs[902]);
    assign layer0_outputs[3561] = ~((inputs[294]) ^ (inputs[78]));
    assign layer0_outputs[3562] = inputs[395];
    assign layer0_outputs[3563] = inputs[597];
    assign layer0_outputs[3564] = inputs[532];
    assign layer0_outputs[3565] = ~(inputs[651]) | (inputs[132]);
    assign layer0_outputs[3566] = (inputs[210]) | (inputs[952]);
    assign layer0_outputs[3567] = ~((inputs[1002]) ^ (inputs[781]));
    assign layer0_outputs[3568] = ~(inputs[247]) | (inputs[643]);
    assign layer0_outputs[3569] = ~(inputs[623]);
    assign layer0_outputs[3570] = (inputs[962]) ^ (inputs[610]);
    assign layer0_outputs[3571] = ~((inputs[156]) | (inputs[906]));
    assign layer0_outputs[3572] = inputs[810];
    assign layer0_outputs[3573] = (inputs[418]) & ~(inputs[549]);
    assign layer0_outputs[3574] = ~((inputs[519]) ^ (inputs[921]));
    assign layer0_outputs[3575] = ~((inputs[178]) ^ (inputs[977]));
    assign layer0_outputs[3576] = inputs[313];
    assign layer0_outputs[3577] = ~((inputs[57]) & (inputs[610]));
    assign layer0_outputs[3578] = ~((inputs[797]) & (inputs[41]));
    assign layer0_outputs[3579] = ~(inputs[827]);
    assign layer0_outputs[3580] = (inputs[438]) & ~(inputs[282]);
    assign layer0_outputs[3581] = ~((inputs[461]) | (inputs[26]));
    assign layer0_outputs[3582] = ~((inputs[407]) ^ (inputs[510]));
    assign layer0_outputs[3583] = inputs[92];
    assign layer0_outputs[3584] = inputs[41];
    assign layer0_outputs[3585] = ~(inputs[424]);
    assign layer0_outputs[3586] = (inputs[585]) & ~(inputs[71]);
    assign layer0_outputs[3587] = (inputs[730]) & ~(inputs[489]);
    assign layer0_outputs[3588] = (inputs[493]) & ~(inputs[769]);
    assign layer0_outputs[3589] = ~((inputs[4]) & (inputs[1007]));
    assign layer0_outputs[3590] = (inputs[40]) & ~(inputs[269]);
    assign layer0_outputs[3591] = ~(inputs[784]);
    assign layer0_outputs[3592] = ~((inputs[117]) & (inputs[166]));
    assign layer0_outputs[3593] = (inputs[469]) | (inputs[909]);
    assign layer0_outputs[3594] = (inputs[915]) | (inputs[27]);
    assign layer0_outputs[3595] = inputs[842];
    assign layer0_outputs[3596] = ~(inputs[128]) | (inputs[136]);
    assign layer0_outputs[3597] = (inputs[697]) & ~(inputs[486]);
    assign layer0_outputs[3598] = (inputs[404]) ^ (inputs[981]);
    assign layer0_outputs[3599] = (inputs[433]) ^ (inputs[404]);
    assign layer0_outputs[3600] = ~(inputs[663]);
    assign layer0_outputs[3601] = ~(inputs[488]);
    assign layer0_outputs[3602] = ~((inputs[194]) & (inputs[601]));
    assign layer0_outputs[3603] = inputs[378];
    assign layer0_outputs[3604] = (inputs[172]) | (inputs[854]);
    assign layer0_outputs[3605] = ~(inputs[103]);
    assign layer0_outputs[3606] = ~(inputs[782]) | (inputs[892]);
    assign layer0_outputs[3607] = ~(inputs[376]);
    assign layer0_outputs[3608] = ~(inputs[756]);
    assign layer0_outputs[3609] = (inputs[366]) | (inputs[226]);
    assign layer0_outputs[3610] = (inputs[928]) ^ (inputs[568]);
    assign layer0_outputs[3611] = ~(inputs[33]) | (inputs[945]);
    assign layer0_outputs[3612] = ~(inputs[672]) | (inputs[706]);
    assign layer0_outputs[3613] = (inputs[960]) & (inputs[916]);
    assign layer0_outputs[3614] = (inputs[416]) | (inputs[676]);
    assign layer0_outputs[3615] = 1'b1;
    assign layer0_outputs[3616] = ~((inputs[742]) | (inputs[423]));
    assign layer0_outputs[3617] = inputs[583];
    assign layer0_outputs[3618] = ~(inputs[924]) | (inputs[23]);
    assign layer0_outputs[3619] = (inputs[512]) | (inputs[301]);
    assign layer0_outputs[3620] = 1'b1;
    assign layer0_outputs[3621] = ~((inputs[278]) | (inputs[793]));
    assign layer0_outputs[3622] = ~(inputs[163]);
    assign layer0_outputs[3623] = ~(inputs[322]) | (inputs[509]);
    assign layer0_outputs[3624] = ~((inputs[419]) & (inputs[193]));
    assign layer0_outputs[3625] = inputs[956];
    assign layer0_outputs[3626] = 1'b0;
    assign layer0_outputs[3627] = 1'b1;
    assign layer0_outputs[3628] = ~((inputs[616]) | (inputs[637]));
    assign layer0_outputs[3629] = (inputs[962]) & ~(inputs[50]);
    assign layer0_outputs[3630] = ~((inputs[19]) | (inputs[528]));
    assign layer0_outputs[3631] = inputs[217];
    assign layer0_outputs[3632] = inputs[520];
    assign layer0_outputs[3633] = 1'b1;
    assign layer0_outputs[3634] = ~((inputs[629]) | (inputs[375]));
    assign layer0_outputs[3635] = inputs[800];
    assign layer0_outputs[3636] = ~((inputs[1003]) | (inputs[599]));
    assign layer0_outputs[3637] = (inputs[467]) ^ (inputs[615]);
    assign layer0_outputs[3638] = ~(inputs[173]);
    assign layer0_outputs[3639] = inputs[343];
    assign layer0_outputs[3640] = (inputs[968]) & ~(inputs[787]);
    assign layer0_outputs[3641] = ~((inputs[966]) | (inputs[687]));
    assign layer0_outputs[3642] = (inputs[421]) ^ (inputs[489]);
    assign layer0_outputs[3643] = ~(inputs[360]);
    assign layer0_outputs[3644] = ~((inputs[948]) ^ (inputs[117]));
    assign layer0_outputs[3645] = (inputs[664]) | (inputs[616]);
    assign layer0_outputs[3646] = ~((inputs[380]) ^ (inputs[884]));
    assign layer0_outputs[3647] = (inputs[825]) & (inputs[781]);
    assign layer0_outputs[3648] = ~((inputs[275]) | (inputs[708]));
    assign layer0_outputs[3649] = (inputs[16]) & ~(inputs[270]);
    assign layer0_outputs[3650] = ~((inputs[54]) | (inputs[161]));
    assign layer0_outputs[3651] = ~((inputs[778]) ^ (inputs[448]));
    assign layer0_outputs[3652] = inputs[593];
    assign layer0_outputs[3653] = ~(inputs[339]);
    assign layer0_outputs[3654] = ~(inputs[958]);
    assign layer0_outputs[3655] = ~(inputs[259]);
    assign layer0_outputs[3656] = (inputs[179]) ^ (inputs[291]);
    assign layer0_outputs[3657] = (inputs[287]) & (inputs[670]);
    assign layer0_outputs[3658] = 1'b1;
    assign layer0_outputs[3659] = ~(inputs[432]);
    assign layer0_outputs[3660] = (inputs[176]) ^ (inputs[263]);
    assign layer0_outputs[3661] = inputs[827];
    assign layer0_outputs[3662] = ~(inputs[615]);
    assign layer0_outputs[3663] = inputs[440];
    assign layer0_outputs[3664] = (inputs[617]) | (inputs[763]);
    assign layer0_outputs[3665] = (inputs[1023]) | (inputs[200]);
    assign layer0_outputs[3666] = inputs[145];
    assign layer0_outputs[3667] = ~(inputs[77]) | (inputs[23]);
    assign layer0_outputs[3668] = ~(inputs[618]) | (inputs[259]);
    assign layer0_outputs[3669] = (inputs[652]) & ~(inputs[152]);
    assign layer0_outputs[3670] = (inputs[551]) & ~(inputs[140]);
    assign layer0_outputs[3671] = ~(inputs[526]) | (inputs[863]);
    assign layer0_outputs[3672] = ~(inputs[439]) | (inputs[232]);
    assign layer0_outputs[3673] = ~((inputs[110]) ^ (inputs[575]));
    assign layer0_outputs[3674] = inputs[984];
    assign layer0_outputs[3675] = ~(inputs[301]) | (inputs[649]);
    assign layer0_outputs[3676] = (inputs[658]) | (inputs[836]);
    assign layer0_outputs[3677] = (inputs[526]) | (inputs[133]);
    assign layer0_outputs[3678] = ~((inputs[809]) | (inputs[11]));
    assign layer0_outputs[3679] = ~(inputs[791]) | (inputs[47]);
    assign layer0_outputs[3680] = 1'b0;
    assign layer0_outputs[3681] = inputs[74];
    assign layer0_outputs[3682] = (inputs[523]) & ~(inputs[835]);
    assign layer0_outputs[3683] = ~((inputs[570]) ^ (inputs[830]));
    assign layer0_outputs[3684] = (inputs[639]) | (inputs[472]);
    assign layer0_outputs[3685] = ~(inputs[764]) | (inputs[641]);
    assign layer0_outputs[3686] = ~((inputs[389]) ^ (inputs[874]));
    assign layer0_outputs[3687] = (inputs[882]) & ~(inputs[871]);
    assign layer0_outputs[3688] = (inputs[540]) ^ (inputs[905]);
    assign layer0_outputs[3689] = inputs[930];
    assign layer0_outputs[3690] = (inputs[757]) ^ (inputs[85]);
    assign layer0_outputs[3691] = ~((inputs[702]) & (inputs[834]));
    assign layer0_outputs[3692] = inputs[435];
    assign layer0_outputs[3693] = ~(inputs[345]) | (inputs[121]);
    assign layer0_outputs[3694] = inputs[608];
    assign layer0_outputs[3695] = (inputs[191]) | (inputs[146]);
    assign layer0_outputs[3696] = ~((inputs[815]) | (inputs[391]));
    assign layer0_outputs[3697] = ~((inputs[556]) | (inputs[605]));
    assign layer0_outputs[3698] = 1'b1;
    assign layer0_outputs[3699] = (inputs[661]) | (inputs[582]);
    assign layer0_outputs[3700] = 1'b1;
    assign layer0_outputs[3701] = (inputs[1019]) & ~(inputs[985]);
    assign layer0_outputs[3702] = (inputs[904]) | (inputs[845]);
    assign layer0_outputs[3703] = (inputs[517]) | (inputs[633]);
    assign layer0_outputs[3704] = (inputs[406]) & ~(inputs[297]);
    assign layer0_outputs[3705] = (inputs[343]) | (inputs[864]);
    assign layer0_outputs[3706] = ~((inputs[580]) | (inputs[705]));
    assign layer0_outputs[3707] = ~((inputs[252]) & (inputs[1017]));
    assign layer0_outputs[3708] = (inputs[692]) | (inputs[352]);
    assign layer0_outputs[3709] = ~((inputs[364]) ^ (inputs[529]));
    assign layer0_outputs[3710] = ~(inputs[516]) | (inputs[480]);
    assign layer0_outputs[3711] = (inputs[177]) & ~(inputs[372]);
    assign layer0_outputs[3712] = ~((inputs[906]) & (inputs[130]));
    assign layer0_outputs[3713] = (inputs[308]) & ~(inputs[590]);
    assign layer0_outputs[3714] = ~(inputs[332]) | (inputs[438]);
    assign layer0_outputs[3715] = (inputs[667]) & (inputs[352]);
    assign layer0_outputs[3716] = (inputs[244]) & ~(inputs[977]);
    assign layer0_outputs[3717] = (inputs[615]) & ~(inputs[341]);
    assign layer0_outputs[3718] = (inputs[781]) | (inputs[6]);
    assign layer0_outputs[3719] = inputs[954];
    assign layer0_outputs[3720] = (inputs[552]) & ~(inputs[980]);
    assign layer0_outputs[3721] = (inputs[932]) | (inputs[963]);
    assign layer0_outputs[3722] = ~(inputs[116]);
    assign layer0_outputs[3723] = (inputs[721]) & ~(inputs[380]);
    assign layer0_outputs[3724] = ~(inputs[369]);
    assign layer0_outputs[3725] = (inputs[201]) | (inputs[795]);
    assign layer0_outputs[3726] = ~((inputs[469]) | (inputs[910]));
    assign layer0_outputs[3727] = inputs[1021];
    assign layer0_outputs[3728] = ~(inputs[265]);
    assign layer0_outputs[3729] = ~(inputs[62]) | (inputs[898]);
    assign layer0_outputs[3730] = ~((inputs[714]) | (inputs[184]));
    assign layer0_outputs[3731] = (inputs[585]) ^ (inputs[869]);
    assign layer0_outputs[3732] = ~(inputs[648]) | (inputs[138]);
    assign layer0_outputs[3733] = ~((inputs[147]) | (inputs[778]));
    assign layer0_outputs[3734] = (inputs[458]) ^ (inputs[430]);
    assign layer0_outputs[3735] = 1'b0;
    assign layer0_outputs[3736] = ~((inputs[298]) | (inputs[621]));
    assign layer0_outputs[3737] = ~(inputs[436]);
    assign layer0_outputs[3738] = ~((inputs[321]) ^ (inputs[597]));
    assign layer0_outputs[3739] = ~(inputs[716]);
    assign layer0_outputs[3740] = ~((inputs[886]) | (inputs[394]));
    assign layer0_outputs[3741] = (inputs[919]) ^ (inputs[698]);
    assign layer0_outputs[3742] = (inputs[418]) | (inputs[155]);
    assign layer0_outputs[3743] = (inputs[268]) | (inputs[697]);
    assign layer0_outputs[3744] = (inputs[241]) & (inputs[714]);
    assign layer0_outputs[3745] = inputs[206];
    assign layer0_outputs[3746] = ~((inputs[596]) ^ (inputs[532]));
    assign layer0_outputs[3747] = ~(inputs[455]) | (inputs[976]);
    assign layer0_outputs[3748] = ~(inputs[339]) | (inputs[80]);
    assign layer0_outputs[3749] = 1'b1;
    assign layer0_outputs[3750] = ~(inputs[978]) | (inputs[455]);
    assign layer0_outputs[3751] = (inputs[381]) & ~(inputs[605]);
    assign layer0_outputs[3752] = ~((inputs[704]) & (inputs[605]));
    assign layer0_outputs[3753] = inputs[906];
    assign layer0_outputs[3754] = inputs[782];
    assign layer0_outputs[3755] = (inputs[91]) ^ (inputs[489]);
    assign layer0_outputs[3756] = (inputs[563]) ^ (inputs[973]);
    assign layer0_outputs[3757] = ~((inputs[640]) ^ (inputs[472]));
    assign layer0_outputs[3758] = inputs[765];
    assign layer0_outputs[3759] = (inputs[653]) & ~(inputs[385]);
    assign layer0_outputs[3760] = 1'b0;
    assign layer0_outputs[3761] = ~((inputs[606]) | (inputs[706]));
    assign layer0_outputs[3762] = ~(inputs[760]);
    assign layer0_outputs[3763] = ~((inputs[289]) ^ (inputs[9]));
    assign layer0_outputs[3764] = ~(inputs[811]);
    assign layer0_outputs[3765] = (inputs[264]) & ~(inputs[648]);
    assign layer0_outputs[3766] = ~(inputs[621]) | (inputs[397]);
    assign layer0_outputs[3767] = ~((inputs[885]) | (inputs[878]));
    assign layer0_outputs[3768] = ~(inputs[914]) | (inputs[114]);
    assign layer0_outputs[3769] = (inputs[287]) | (inputs[314]);
    assign layer0_outputs[3770] = ~((inputs[872]) ^ (inputs[544]));
    assign layer0_outputs[3771] = (inputs[864]) | (inputs[971]);
    assign layer0_outputs[3772] = ~((inputs[571]) & (inputs[779]));
    assign layer0_outputs[3773] = ~((inputs[781]) | (inputs[925]));
    assign layer0_outputs[3774] = (inputs[181]) ^ (inputs[717]);
    assign layer0_outputs[3775] = ~(inputs[5]) | (inputs[478]);
    assign layer0_outputs[3776] = inputs[104];
    assign layer0_outputs[3777] = ~(inputs[373]);
    assign layer0_outputs[3778] = 1'b1;
    assign layer0_outputs[3779] = (inputs[79]) ^ (inputs[996]);
    assign layer0_outputs[3780] = (inputs[635]) & ~(inputs[483]);
    assign layer0_outputs[3781] = ~(inputs[527]);
    assign layer0_outputs[3782] = (inputs[814]) & ~(inputs[838]);
    assign layer0_outputs[3783] = (inputs[610]) | (inputs[206]);
    assign layer0_outputs[3784] = ~((inputs[431]) | (inputs[668]));
    assign layer0_outputs[3785] = ~(inputs[634]) | (inputs[955]);
    assign layer0_outputs[3786] = inputs[163];
    assign layer0_outputs[3787] = ~(inputs[887]);
    assign layer0_outputs[3788] = (inputs[556]) ^ (inputs[764]);
    assign layer0_outputs[3789] = ~(inputs[457]) | (inputs[847]);
    assign layer0_outputs[3790] = (inputs[505]) & ~(inputs[68]);
    assign layer0_outputs[3791] = (inputs[785]) ^ (inputs[253]);
    assign layer0_outputs[3792] = (inputs[510]) & (inputs[439]);
    assign layer0_outputs[3793] = ~((inputs[949]) & (inputs[1020]));
    assign layer0_outputs[3794] = ~((inputs[287]) ^ (inputs[811]));
    assign layer0_outputs[3795] = (inputs[212]) & ~(inputs[825]);
    assign layer0_outputs[3796] = (inputs[986]) & ~(inputs[990]);
    assign layer0_outputs[3797] = (inputs[324]) & (inputs[154]);
    assign layer0_outputs[3798] = (inputs[665]) ^ (inputs[779]);
    assign layer0_outputs[3799] = ~(inputs[847]);
    assign layer0_outputs[3800] = ~(inputs[53]) | (inputs[838]);
    assign layer0_outputs[3801] = (inputs[764]) | (inputs[325]);
    assign layer0_outputs[3802] = inputs[246];
    assign layer0_outputs[3803] = ~((inputs[765]) | (inputs[909]));
    assign layer0_outputs[3804] = ~(inputs[889]);
    assign layer0_outputs[3805] = (inputs[589]) & (inputs[440]);
    assign layer0_outputs[3806] = ~((inputs[554]) | (inputs[119]));
    assign layer0_outputs[3807] = (inputs[254]) & ~(inputs[906]);
    assign layer0_outputs[3808] = ~((inputs[627]) ^ (inputs[233]));
    assign layer0_outputs[3809] = ~((inputs[741]) | (inputs[194]));
    assign layer0_outputs[3810] = (inputs[614]) | (inputs[683]);
    assign layer0_outputs[3811] = (inputs[604]) & ~(inputs[642]);
    assign layer0_outputs[3812] = (inputs[822]) | (inputs[702]);
    assign layer0_outputs[3813] = (inputs[588]) | (inputs[317]);
    assign layer0_outputs[3814] = (inputs[239]) & ~(inputs[53]);
    assign layer0_outputs[3815] = (inputs[109]) & ~(inputs[740]);
    assign layer0_outputs[3816] = ~(inputs[58]);
    assign layer0_outputs[3817] = inputs[493];
    assign layer0_outputs[3818] = ~((inputs[378]) | (inputs[327]));
    assign layer0_outputs[3819] = inputs[244];
    assign layer0_outputs[3820] = (inputs[738]) | (inputs[157]);
    assign layer0_outputs[3821] = (inputs[664]) | (inputs[687]);
    assign layer0_outputs[3822] = (inputs[525]) | (inputs[1004]);
    assign layer0_outputs[3823] = 1'b1;
    assign layer0_outputs[3824] = inputs[655];
    assign layer0_outputs[3825] = ~(inputs[663]);
    assign layer0_outputs[3826] = (inputs[984]) | (inputs[461]);
    assign layer0_outputs[3827] = ~((inputs[513]) | (inputs[938]));
    assign layer0_outputs[3828] = ~(inputs[1023]);
    assign layer0_outputs[3829] = ~((inputs[233]) ^ (inputs[44]));
    assign layer0_outputs[3830] = ~((inputs[997]) ^ (inputs[610]));
    assign layer0_outputs[3831] = (inputs[803]) & (inputs[954]);
    assign layer0_outputs[3832] = ~(inputs[242]);
    assign layer0_outputs[3833] = 1'b0;
    assign layer0_outputs[3834] = ~(inputs[663]) | (inputs[218]);
    assign layer0_outputs[3835] = ~(inputs[250]) | (inputs[286]);
    assign layer0_outputs[3836] = (inputs[625]) & ~(inputs[991]);
    assign layer0_outputs[3837] = ~(inputs[778]) | (inputs[960]);
    assign layer0_outputs[3838] = ~(inputs[631]);
    assign layer0_outputs[3839] = ~((inputs[655]) | (inputs[675]));
    assign layer0_outputs[3840] = (inputs[188]) ^ (inputs[871]);
    assign layer0_outputs[3841] = (inputs[649]) | (inputs[556]);
    assign layer0_outputs[3842] = ~(inputs[616]);
    assign layer0_outputs[3843] = ~(inputs[700]);
    assign layer0_outputs[3844] = ~((inputs[559]) | (inputs[825]));
    assign layer0_outputs[3845] = ~(inputs[136]);
    assign layer0_outputs[3846] = ~(inputs[394]);
    assign layer0_outputs[3847] = ~(inputs[500]);
    assign layer0_outputs[3848] = inputs[229];
    assign layer0_outputs[3849] = (inputs[1021]) & ~(inputs[895]);
    assign layer0_outputs[3850] = 1'b1;
    assign layer0_outputs[3851] = ~(inputs[429]);
    assign layer0_outputs[3852] = (inputs[651]) & ~(inputs[770]);
    assign layer0_outputs[3853] = (inputs[303]) & ~(inputs[900]);
    assign layer0_outputs[3854] = ~(inputs[1009]);
    assign layer0_outputs[3855] = (inputs[592]) & ~(inputs[103]);
    assign layer0_outputs[3856] = (inputs[284]) & ~(inputs[669]);
    assign layer0_outputs[3857] = ~((inputs[690]) & (inputs[416]));
    assign layer0_outputs[3858] = ~(inputs[838]) | (inputs[911]);
    assign layer0_outputs[3859] = (inputs[424]) & (inputs[908]);
    assign layer0_outputs[3860] = ~((inputs[860]) | (inputs[364]));
    assign layer0_outputs[3861] = inputs[712];
    assign layer0_outputs[3862] = ~(inputs[825]);
    assign layer0_outputs[3863] = 1'b1;
    assign layer0_outputs[3864] = inputs[613];
    assign layer0_outputs[3865] = ~((inputs[815]) ^ (inputs[791]));
    assign layer0_outputs[3866] = ~(inputs[629]) | (inputs[796]);
    assign layer0_outputs[3867] = 1'b0;
    assign layer0_outputs[3868] = (inputs[447]) & (inputs[13]);
    assign layer0_outputs[3869] = (inputs[1021]) | (inputs[695]);
    assign layer0_outputs[3870] = (inputs[151]) & ~(inputs[987]);
    assign layer0_outputs[3871] = (inputs[472]) | (inputs[556]);
    assign layer0_outputs[3872] = ~((inputs[323]) ^ (inputs[874]));
    assign layer0_outputs[3873] = (inputs[318]) ^ (inputs[151]);
    assign layer0_outputs[3874] = 1'b1;
    assign layer0_outputs[3875] = (inputs[595]) & ~(inputs[336]);
    assign layer0_outputs[3876] = inputs[875];
    assign layer0_outputs[3877] = ~((inputs[25]) ^ (inputs[110]));
    assign layer0_outputs[3878] = (inputs[919]) | (inputs[957]);
    assign layer0_outputs[3879] = ~(inputs[926]);
    assign layer0_outputs[3880] = ~((inputs[586]) | (inputs[941]));
    assign layer0_outputs[3881] = inputs[228];
    assign layer0_outputs[3882] = ~((inputs[197]) | (inputs[219]));
    assign layer0_outputs[3883] = inputs[429];
    assign layer0_outputs[3884] = ~((inputs[82]) ^ (inputs[174]));
    assign layer0_outputs[3885] = inputs[727];
    assign layer0_outputs[3886] = (inputs[631]) & ~(inputs[363]);
    assign layer0_outputs[3887] = inputs[165];
    assign layer0_outputs[3888] = inputs[130];
    assign layer0_outputs[3889] = inputs[61];
    assign layer0_outputs[3890] = (inputs[759]) & ~(inputs[224]);
    assign layer0_outputs[3891] = inputs[376];
    assign layer0_outputs[3892] = inputs[340];
    assign layer0_outputs[3893] = ~((inputs[108]) ^ (inputs[43]));
    assign layer0_outputs[3894] = ~(inputs[522]) | (inputs[94]);
    assign layer0_outputs[3895] = ~((inputs[682]) | (inputs[692]));
    assign layer0_outputs[3896] = ~(inputs[405]);
    assign layer0_outputs[3897] = ~(inputs[1003]);
    assign layer0_outputs[3898] = ~((inputs[440]) | (inputs[951]));
    assign layer0_outputs[3899] = (inputs[25]) ^ (inputs[181]);
    assign layer0_outputs[3900] = ~(inputs[784]) | (inputs[243]);
    assign layer0_outputs[3901] = ~(inputs[466]) | (inputs[762]);
    assign layer0_outputs[3902] = ~((inputs[799]) ^ (inputs[616]));
    assign layer0_outputs[3903] = inputs[286];
    assign layer0_outputs[3904] = (inputs[691]) ^ (inputs[388]);
    assign layer0_outputs[3905] = ~(inputs[539]);
    assign layer0_outputs[3906] = (inputs[59]) & ~(inputs[998]);
    assign layer0_outputs[3907] = ~((inputs[908]) ^ (inputs[350]));
    assign layer0_outputs[3908] = (inputs[365]) & ~(inputs[322]);
    assign layer0_outputs[3909] = ~(inputs[134]);
    assign layer0_outputs[3910] = ~((inputs[610]) ^ (inputs[608]));
    assign layer0_outputs[3911] = ~((inputs[493]) & (inputs[330]));
    assign layer0_outputs[3912] = ~(inputs[90]) | (inputs[353]);
    assign layer0_outputs[3913] = ~(inputs[243]) | (inputs[1021]);
    assign layer0_outputs[3914] = (inputs[145]) | (inputs[706]);
    assign layer0_outputs[3915] = (inputs[560]) | (inputs[384]);
    assign layer0_outputs[3916] = ~(inputs[455]) | (inputs[606]);
    assign layer0_outputs[3917] = inputs[546];
    assign layer0_outputs[3918] = ~((inputs[412]) | (inputs[203]));
    assign layer0_outputs[3919] = (inputs[288]) | (inputs[781]);
    assign layer0_outputs[3920] = (inputs[794]) | (inputs[273]);
    assign layer0_outputs[3921] = (inputs[559]) & ~(inputs[767]);
    assign layer0_outputs[3922] = (inputs[324]) | (inputs[504]);
    assign layer0_outputs[3923] = ~(inputs[554]);
    assign layer0_outputs[3924] = ~(inputs[353]);
    assign layer0_outputs[3925] = ~(inputs[306]);
    assign layer0_outputs[3926] = ~((inputs[263]) & (inputs[419]));
    assign layer0_outputs[3927] = (inputs[368]) ^ (inputs[988]);
    assign layer0_outputs[3928] = (inputs[148]) | (inputs[724]);
    assign layer0_outputs[3929] = ~((inputs[1001]) ^ (inputs[355]));
    assign layer0_outputs[3930] = (inputs[747]) & ~(inputs[842]);
    assign layer0_outputs[3931] = ~((inputs[601]) & (inputs[102]));
    assign layer0_outputs[3932] = ~((inputs[621]) | (inputs[520]));
    assign layer0_outputs[3933] = ~(inputs[591]);
    assign layer0_outputs[3934] = inputs[333];
    assign layer0_outputs[3935] = inputs[227];
    assign layer0_outputs[3936] = ~((inputs[520]) ^ (inputs[288]));
    assign layer0_outputs[3937] = ~(inputs[193]);
    assign layer0_outputs[3938] = ~(inputs[866]) | (inputs[472]);
    assign layer0_outputs[3939] = (inputs[274]) & ~(inputs[421]);
    assign layer0_outputs[3940] = (inputs[413]) & (inputs[472]);
    assign layer0_outputs[3941] = ~(inputs[463]);
    assign layer0_outputs[3942] = inputs[596];
    assign layer0_outputs[3943] = (inputs[16]) | (inputs[816]);
    assign layer0_outputs[3944] = ~(inputs[176]) | (inputs[128]);
    assign layer0_outputs[3945] = (inputs[524]) & ~(inputs[960]);
    assign layer0_outputs[3946] = ~(inputs[497]) | (inputs[136]);
    assign layer0_outputs[3947] = (inputs[657]) & ~(inputs[749]);
    assign layer0_outputs[3948] = 1'b0;
    assign layer0_outputs[3949] = ~((inputs[747]) | (inputs[477]));
    assign layer0_outputs[3950] = (inputs[365]) & ~(inputs[167]);
    assign layer0_outputs[3951] = ~(inputs[360]) | (inputs[651]);
    assign layer0_outputs[3952] = ~((inputs[670]) | (inputs[697]));
    assign layer0_outputs[3953] = ~(inputs[246]) | (inputs[19]);
    assign layer0_outputs[3954] = (inputs[974]) & (inputs[605]);
    assign layer0_outputs[3955] = inputs[146];
    assign layer0_outputs[3956] = (inputs[104]) | (inputs[943]);
    assign layer0_outputs[3957] = (inputs[203]) & ~(inputs[86]);
    assign layer0_outputs[3958] = (inputs[729]) ^ (inputs[113]);
    assign layer0_outputs[3959] = (inputs[675]) | (inputs[494]);
    assign layer0_outputs[3960] = ~(inputs[663]);
    assign layer0_outputs[3961] = (inputs[733]) ^ (inputs[764]);
    assign layer0_outputs[3962] = ~(inputs[455]);
    assign layer0_outputs[3963] = 1'b0;
    assign layer0_outputs[3964] = 1'b0;
    assign layer0_outputs[3965] = ~(inputs[877]);
    assign layer0_outputs[3966] = (inputs[330]) & ~(inputs[985]);
    assign layer0_outputs[3967] = (inputs[385]) | (inputs[314]);
    assign layer0_outputs[3968] = ~((inputs[85]) ^ (inputs[121]));
    assign layer0_outputs[3969] = (inputs[476]) ^ (inputs[803]);
    assign layer0_outputs[3970] = ~(inputs[347]) | (inputs[295]);
    assign layer0_outputs[3971] = ~((inputs[654]) & (inputs[880]));
    assign layer0_outputs[3972] = ~(inputs[932]) | (inputs[473]);
    assign layer0_outputs[3973] = (inputs[731]) ^ (inputs[823]);
    assign layer0_outputs[3974] = ~(inputs[34]) | (inputs[681]);
    assign layer0_outputs[3975] = (inputs[34]) ^ (inputs[9]);
    assign layer0_outputs[3976] = ~(inputs[487]) | (inputs[940]);
    assign layer0_outputs[3977] = (inputs[520]) & ~(inputs[69]);
    assign layer0_outputs[3978] = inputs[725];
    assign layer0_outputs[3979] = ~(inputs[794]);
    assign layer0_outputs[3980] = (inputs[158]) ^ (inputs[578]);
    assign layer0_outputs[3981] = ~(inputs[59]) | (inputs[515]);
    assign layer0_outputs[3982] = ~((inputs[214]) | (inputs[678]));
    assign layer0_outputs[3983] = ~(inputs[469]) | (inputs[117]);
    assign layer0_outputs[3984] = 1'b1;
    assign layer0_outputs[3985] = ~((inputs[574]) & (inputs[942]));
    assign layer0_outputs[3986] = ~(inputs[627]);
    assign layer0_outputs[3987] = ~((inputs[529]) ^ (inputs[632]));
    assign layer0_outputs[3988] = (inputs[845]) & ~(inputs[70]);
    assign layer0_outputs[3989] = inputs[759];
    assign layer0_outputs[3990] = ~(inputs[521]) | (inputs[80]);
    assign layer0_outputs[3991] = (inputs[437]) & ~(inputs[20]);
    assign layer0_outputs[3992] = ~(inputs[947]) | (inputs[438]);
    assign layer0_outputs[3993] = ~(inputs[10]) | (inputs[985]);
    assign layer0_outputs[3994] = (inputs[627]) | (inputs[409]);
    assign layer0_outputs[3995] = ~((inputs[286]) | (inputs[44]));
    assign layer0_outputs[3996] = (inputs[143]) ^ (inputs[337]);
    assign layer0_outputs[3997] = (inputs[863]) | (inputs[186]);
    assign layer0_outputs[3998] = (inputs[713]) & ~(inputs[771]);
    assign layer0_outputs[3999] = inputs[818];
    assign layer0_outputs[4000] = ~((inputs[665]) | (inputs[597]));
    assign layer0_outputs[4001] = (inputs[914]) & (inputs[253]);
    assign layer0_outputs[4002] = ~(inputs[401]) | (inputs[485]);
    assign layer0_outputs[4003] = ~(inputs[434]) | (inputs[808]);
    assign layer0_outputs[4004] = ~((inputs[933]) ^ (inputs[851]));
    assign layer0_outputs[4005] = (inputs[946]) ^ (inputs[881]);
    assign layer0_outputs[4006] = inputs[723];
    assign layer0_outputs[4007] = ~(inputs[504]) | (inputs[544]);
    assign layer0_outputs[4008] = ~(inputs[733]) | (inputs[391]);
    assign layer0_outputs[4009] = inputs[280];
    assign layer0_outputs[4010] = (inputs[770]) | (inputs[753]);
    assign layer0_outputs[4011] = ~(inputs[806]);
    assign layer0_outputs[4012] = (inputs[366]) & ~(inputs[282]);
    assign layer0_outputs[4013] = ~(inputs[717]) | (inputs[702]);
    assign layer0_outputs[4014] = ~((inputs[984]) | (inputs[301]));
    assign layer0_outputs[4015] = ~((inputs[773]) | (inputs[568]));
    assign layer0_outputs[4016] = (inputs[151]) | (inputs[736]);
    assign layer0_outputs[4017] = inputs[544];
    assign layer0_outputs[4018] = (inputs[913]) ^ (inputs[503]);
    assign layer0_outputs[4019] = (inputs[719]) ^ (inputs[814]);
    assign layer0_outputs[4020] = (inputs[316]) | (inputs[618]);
    assign layer0_outputs[4021] = ~((inputs[226]) & (inputs[803]));
    assign layer0_outputs[4022] = ~(inputs[144]) | (inputs[581]);
    assign layer0_outputs[4023] = (inputs[408]) | (inputs[148]);
    assign layer0_outputs[4024] = ~((inputs[316]) ^ (inputs[953]));
    assign layer0_outputs[4025] = 1'b1;
    assign layer0_outputs[4026] = (inputs[421]) ^ (inputs[49]);
    assign layer0_outputs[4027] = (inputs[335]) & ~(inputs[140]);
    assign layer0_outputs[4028] = ~((inputs[403]) ^ (inputs[841]));
    assign layer0_outputs[4029] = ~(inputs[907]);
    assign layer0_outputs[4030] = (inputs[399]) ^ (inputs[317]);
    assign layer0_outputs[4031] = inputs[712];
    assign layer0_outputs[4032] = (inputs[162]) | (inputs[543]);
    assign layer0_outputs[4033] = ~(inputs[429]);
    assign layer0_outputs[4034] = ~(inputs[595]) | (inputs[154]);
    assign layer0_outputs[4035] = (inputs[617]) & ~(inputs[381]);
    assign layer0_outputs[4036] = ~(inputs[539]) | (inputs[960]);
    assign layer0_outputs[4037] = ~(inputs[517]);
    assign layer0_outputs[4038] = ~((inputs[629]) ^ (inputs[138]));
    assign layer0_outputs[4039] = (inputs[702]) ^ (inputs[973]);
    assign layer0_outputs[4040] = 1'b1;
    assign layer0_outputs[4041] = (inputs[794]) | (inputs[712]);
    assign layer0_outputs[4042] = inputs[935];
    assign layer0_outputs[4043] = ~(inputs[373]) | (inputs[381]);
    assign layer0_outputs[4044] = inputs[585];
    assign layer0_outputs[4045] = inputs[99];
    assign layer0_outputs[4046] = (inputs[451]) | (inputs[5]);
    assign layer0_outputs[4047] = (inputs[657]) | (inputs[76]);
    assign layer0_outputs[4048] = ~(inputs[295]) | (inputs[3]);
    assign layer0_outputs[4049] = ~((inputs[880]) | (inputs[651]));
    assign layer0_outputs[4050] = inputs[454];
    assign layer0_outputs[4051] = ~((inputs[678]) | (inputs[679]));
    assign layer0_outputs[4052] = inputs[658];
    assign layer0_outputs[4053] = ~(inputs[447]);
    assign layer0_outputs[4054] = ~(inputs[283]) | (inputs[995]);
    assign layer0_outputs[4055] = ~(inputs[185]);
    assign layer0_outputs[4056] = (inputs[623]) & ~(inputs[891]);
    assign layer0_outputs[4057] = (inputs[937]) | (inputs[332]);
    assign layer0_outputs[4058] = ~(inputs[461]) | (inputs[347]);
    assign layer0_outputs[4059] = inputs[535];
    assign layer0_outputs[4060] = ~(inputs[381]) | (inputs[804]);
    assign layer0_outputs[4061] = ~(inputs[329]);
    assign layer0_outputs[4062] = (inputs[520]) & (inputs[679]);
    assign layer0_outputs[4063] = ~((inputs[665]) | (inputs[655]));
    assign layer0_outputs[4064] = ~((inputs[267]) ^ (inputs[963]));
    assign layer0_outputs[4065] = inputs[404];
    assign layer0_outputs[4066] = ~((inputs[939]) | (inputs[868]));
    assign layer0_outputs[4067] = ~((inputs[209]) | (inputs[474]));
    assign layer0_outputs[4068] = ~((inputs[687]) ^ (inputs[866]));
    assign layer0_outputs[4069] = ~(inputs[351]) | (inputs[797]);
    assign layer0_outputs[4070] = ~((inputs[728]) | (inputs[295]));
    assign layer0_outputs[4071] = (inputs[125]) & ~(inputs[229]);
    assign layer0_outputs[4072] = ~(inputs[637]) | (inputs[872]);
    assign layer0_outputs[4073] = inputs[789];
    assign layer0_outputs[4074] = ~((inputs[801]) ^ (inputs[421]));
    assign layer0_outputs[4075] = ~(inputs[207]);
    assign layer0_outputs[4076] = 1'b0;
    assign layer0_outputs[4077] = ~((inputs[1002]) ^ (inputs[471]));
    assign layer0_outputs[4078] = ~(inputs[585]);
    assign layer0_outputs[4079] = ~(inputs[616]) | (inputs[6]);
    assign layer0_outputs[4080] = (inputs[123]) | (inputs[207]);
    assign layer0_outputs[4081] = ~((inputs[231]) | (inputs[774]));
    assign layer0_outputs[4082] = inputs[233];
    assign layer0_outputs[4083] = inputs[57];
    assign layer0_outputs[4084] = ~((inputs[380]) | (inputs[863]));
    assign layer0_outputs[4085] = (inputs[235]) | (inputs[939]);
    assign layer0_outputs[4086] = inputs[637];
    assign layer0_outputs[4087] = ~(inputs[878]) | (inputs[707]);
    assign layer0_outputs[4088] = ~(inputs[796]);
    assign layer0_outputs[4089] = (inputs[76]) | (inputs[781]);
    assign layer0_outputs[4090] = 1'b0;
    assign layer0_outputs[4091] = ~(inputs[959]) | (inputs[607]);
    assign layer0_outputs[4092] = ~((inputs[466]) | (inputs[475]));
    assign layer0_outputs[4093] = (inputs[488]) ^ (inputs[256]);
    assign layer0_outputs[4094] = ~((inputs[646]) ^ (inputs[684]));
    assign layer0_outputs[4095] = (inputs[418]) | (inputs[724]);
    assign layer0_outputs[4096] = ~(inputs[989]);
    assign layer0_outputs[4097] = ~(inputs[913]);
    assign layer0_outputs[4098] = ~(inputs[528]);
    assign layer0_outputs[4099] = (inputs[807]) & ~(inputs[752]);
    assign layer0_outputs[4100] = 1'b0;
    assign layer0_outputs[4101] = inputs[123];
    assign layer0_outputs[4102] = (inputs[782]) ^ (inputs[388]);
    assign layer0_outputs[4103] = ~(inputs[810]) | (inputs[513]);
    assign layer0_outputs[4104] = (inputs[309]) ^ (inputs[118]);
    assign layer0_outputs[4105] = inputs[308];
    assign layer0_outputs[4106] = (inputs[254]) | (inputs[583]);
    assign layer0_outputs[4107] = (inputs[396]) | (inputs[241]);
    assign layer0_outputs[4108] = ~((inputs[87]) | (inputs[496]));
    assign layer0_outputs[4109] = ~(inputs[759]);
    assign layer0_outputs[4110] = inputs[248];
    assign layer0_outputs[4111] = inputs[3];
    assign layer0_outputs[4112] = (inputs[886]) | (inputs[276]);
    assign layer0_outputs[4113] = ~(inputs[229]) | (inputs[44]);
    assign layer0_outputs[4114] = ~((inputs[205]) ^ (inputs[18]));
    assign layer0_outputs[4115] = (inputs[713]) & ~(inputs[950]);
    assign layer0_outputs[4116] = (inputs[133]) & ~(inputs[237]);
    assign layer0_outputs[4117] = ~(inputs[190]) | (inputs[387]);
    assign layer0_outputs[4118] = (inputs[592]) ^ (inputs[955]);
    assign layer0_outputs[4119] = ~((inputs[601]) | (inputs[918]));
    assign layer0_outputs[4120] = inputs[815];
    assign layer0_outputs[4121] = inputs[881];
    assign layer0_outputs[4122] = (inputs[136]) ^ (inputs[319]);
    assign layer0_outputs[4123] = (inputs[839]) & ~(inputs[642]);
    assign layer0_outputs[4124] = (inputs[429]) ^ (inputs[523]);
    assign layer0_outputs[4125] = ~(inputs[152]);
    assign layer0_outputs[4126] = ~(inputs[470]) | (inputs[233]);
    assign layer0_outputs[4127] = (inputs[871]) & (inputs[69]);
    assign layer0_outputs[4128] = ~((inputs[985]) ^ (inputs[169]));
    assign layer0_outputs[4129] = (inputs[560]) & ~(inputs[607]);
    assign layer0_outputs[4130] = (inputs[247]) & ~(inputs[728]);
    assign layer0_outputs[4131] = ~(inputs[217]);
    assign layer0_outputs[4132] = inputs[930];
    assign layer0_outputs[4133] = ~(inputs[569]) | (inputs[135]);
    assign layer0_outputs[4134] = ~((inputs[248]) ^ (inputs[378]));
    assign layer0_outputs[4135] = (inputs[593]) & (inputs[1007]);
    assign layer0_outputs[4136] = inputs[385];
    assign layer0_outputs[4137] = ~((inputs[714]) ^ (inputs[1004]));
    assign layer0_outputs[4138] = ~((inputs[561]) | (inputs[132]));
    assign layer0_outputs[4139] = (inputs[261]) & ~(inputs[158]);
    assign layer0_outputs[4140] = (inputs[880]) & ~(inputs[978]);
    assign layer0_outputs[4141] = ~((inputs[996]) | (inputs[872]));
    assign layer0_outputs[4142] = (inputs[907]) & ~(inputs[322]);
    assign layer0_outputs[4143] = inputs[396];
    assign layer0_outputs[4144] = ~((inputs[107]) | (inputs[854]));
    assign layer0_outputs[4145] = ~((inputs[435]) ^ (inputs[69]));
    assign layer0_outputs[4146] = inputs[430];
    assign layer0_outputs[4147] = ~(inputs[993]) | (inputs[611]);
    assign layer0_outputs[4148] = (inputs[545]) & ~(inputs[481]);
    assign layer0_outputs[4149] = inputs[338];
    assign layer0_outputs[4150] = ~(inputs[88]) | (inputs[102]);
    assign layer0_outputs[4151] = ~(inputs[908]);
    assign layer0_outputs[4152] = (inputs[538]) | (inputs[645]);
    assign layer0_outputs[4153] = ~(inputs[655]) | (inputs[259]);
    assign layer0_outputs[4154] = ~((inputs[494]) | (inputs[349]));
    assign layer0_outputs[4155] = ~((inputs[662]) ^ (inputs[519]));
    assign layer0_outputs[4156] = (inputs[938]) & (inputs[377]);
    assign layer0_outputs[4157] = ~((inputs[156]) ^ (inputs[815]));
    assign layer0_outputs[4158] = ~((inputs[776]) | (inputs[981]));
    assign layer0_outputs[4159] = inputs[21];
    assign layer0_outputs[4160] = inputs[391];
    assign layer0_outputs[4161] = (inputs[735]) & ~(inputs[261]);
    assign layer0_outputs[4162] = (inputs[747]) & ~(inputs[275]);
    assign layer0_outputs[4163] = (inputs[345]) ^ (inputs[975]);
    assign layer0_outputs[4164] = ~((inputs[38]) | (inputs[209]));
    assign layer0_outputs[4165] = ~(inputs[925]);
    assign layer0_outputs[4166] = (inputs[481]) & ~(inputs[822]);
    assign layer0_outputs[4167] = ~((inputs[452]) ^ (inputs[909]));
    assign layer0_outputs[4168] = ~((inputs[322]) ^ (inputs[666]));
    assign layer0_outputs[4169] = ~(inputs[321]);
    assign layer0_outputs[4170] = ~(inputs[505]);
    assign layer0_outputs[4171] = ~((inputs[881]) ^ (inputs[704]));
    assign layer0_outputs[4172] = inputs[40];
    assign layer0_outputs[4173] = ~(inputs[402]) | (inputs[359]);
    assign layer0_outputs[4174] = (inputs[293]) & ~(inputs[91]);
    assign layer0_outputs[4175] = (inputs[85]) ^ (inputs[728]);
    assign layer0_outputs[4176] = 1'b0;
    assign layer0_outputs[4177] = (inputs[623]) & ~(inputs[324]);
    assign layer0_outputs[4178] = ~((inputs[770]) ^ (inputs[393]));
    assign layer0_outputs[4179] = inputs[862];
    assign layer0_outputs[4180] = (inputs[594]) & ~(inputs[70]);
    assign layer0_outputs[4181] = inputs[127];
    assign layer0_outputs[4182] = ~(inputs[336]);
    assign layer0_outputs[4183] = (inputs[752]) | (inputs[953]);
    assign layer0_outputs[4184] = ~(inputs[210]) | (inputs[968]);
    assign layer0_outputs[4185] = inputs[1019];
    assign layer0_outputs[4186] = ~(inputs[632]);
    assign layer0_outputs[4187] = ~(inputs[615]);
    assign layer0_outputs[4188] = (inputs[617]) | (inputs[1020]);
    assign layer0_outputs[4189] = (inputs[875]) & ~(inputs[88]);
    assign layer0_outputs[4190] = inputs[82];
    assign layer0_outputs[4191] = ~(inputs[377]);
    assign layer0_outputs[4192] = (inputs[659]) | (inputs[1000]);
    assign layer0_outputs[4193] = inputs[66];
    assign layer0_outputs[4194] = ~(inputs[247]) | (inputs[244]);
    assign layer0_outputs[4195] = (inputs[666]) | (inputs[807]);
    assign layer0_outputs[4196] = ~((inputs[791]) | (inputs[202]));
    assign layer0_outputs[4197] = ~(inputs[970]) | (inputs[262]);
    assign layer0_outputs[4198] = inputs[842];
    assign layer0_outputs[4199] = (inputs[744]) ^ (inputs[940]);
    assign layer0_outputs[4200] = ~((inputs[531]) | (inputs[484]));
    assign layer0_outputs[4201] = 1'b1;
    assign layer0_outputs[4202] = (inputs[970]) & ~(inputs[320]);
    assign layer0_outputs[4203] = ~((inputs[415]) ^ (inputs[695]));
    assign layer0_outputs[4204] = ~(inputs[839]) | (inputs[1014]);
    assign layer0_outputs[4205] = ~(inputs[173]);
    assign layer0_outputs[4206] = (inputs[649]) & ~(inputs[902]);
    assign layer0_outputs[4207] = ~((inputs[292]) | (inputs[367]));
    assign layer0_outputs[4208] = (inputs[483]) & ~(inputs[142]);
    assign layer0_outputs[4209] = ~(inputs[181]);
    assign layer0_outputs[4210] = ~((inputs[496]) & (inputs[562]));
    assign layer0_outputs[4211] = ~(inputs[773]) | (inputs[596]);
    assign layer0_outputs[4212] = ~((inputs[985]) | (inputs[238]));
    assign layer0_outputs[4213] = ~(inputs[235]) | (inputs[22]);
    assign layer0_outputs[4214] = (inputs[57]) & (inputs[15]);
    assign layer0_outputs[4215] = inputs[849];
    assign layer0_outputs[4216] = (inputs[239]) & ~(inputs[186]);
    assign layer0_outputs[4217] = ~((inputs[243]) ^ (inputs[468]));
    assign layer0_outputs[4218] = (inputs[789]) & ~(inputs[964]);
    assign layer0_outputs[4219] = ~((inputs[579]) ^ (inputs[459]));
    assign layer0_outputs[4220] = inputs[756];
    assign layer0_outputs[4221] = (inputs[1022]) ^ (inputs[856]);
    assign layer0_outputs[4222] = ~((inputs[931]) & (inputs[801]));
    assign layer0_outputs[4223] = ~((inputs[147]) & (inputs[22]));
    assign layer0_outputs[4224] = ~((inputs[897]) & (inputs[1004]));
    assign layer0_outputs[4225] = ~((inputs[39]) ^ (inputs[813]));
    assign layer0_outputs[4226] = (inputs[741]) ^ (inputs[585]);
    assign layer0_outputs[4227] = (inputs[809]) ^ (inputs[579]);
    assign layer0_outputs[4228] = ~((inputs[577]) ^ (inputs[144]));
    assign layer0_outputs[4229] = inputs[312];
    assign layer0_outputs[4230] = (inputs[573]) ^ (inputs[367]);
    assign layer0_outputs[4231] = ~((inputs[924]) ^ (inputs[789]));
    assign layer0_outputs[4232] = inputs[391];
    assign layer0_outputs[4233] = (inputs[216]) | (inputs[256]);
    assign layer0_outputs[4234] = (inputs[330]) | (inputs[131]);
    assign layer0_outputs[4235] = (inputs[249]) & ~(inputs[861]);
    assign layer0_outputs[4236] = 1'b0;
    assign layer0_outputs[4237] = (inputs[643]) | (inputs[376]);
    assign layer0_outputs[4238] = (inputs[197]) | (inputs[696]);
    assign layer0_outputs[4239] = ~(inputs[538]) | (inputs[990]);
    assign layer0_outputs[4240] = ~((inputs[321]) ^ (inputs[474]));
    assign layer0_outputs[4241] = (inputs[567]) | (inputs[897]);
    assign layer0_outputs[4242] = ~((inputs[154]) ^ (inputs[521]));
    assign layer0_outputs[4243] = ~((inputs[639]) ^ (inputs[482]));
    assign layer0_outputs[4244] = (inputs[919]) & ~(inputs[27]);
    assign layer0_outputs[4245] = ~(inputs[748]) | (inputs[38]);
    assign layer0_outputs[4246] = ~((inputs[220]) ^ (inputs[448]));
    assign layer0_outputs[4247] = inputs[918];
    assign layer0_outputs[4248] = ~(inputs[849]);
    assign layer0_outputs[4249] = ~(inputs[682]) | (inputs[323]);
    assign layer0_outputs[4250] = ~(inputs[348]);
    assign layer0_outputs[4251] = ~(inputs[861]);
    assign layer0_outputs[4252] = (inputs[19]) & (inputs[62]);
    assign layer0_outputs[4253] = ~((inputs[428]) | (inputs[21]));
    assign layer0_outputs[4254] = (inputs[702]) & ~(inputs[227]);
    assign layer0_outputs[4255] = ~((inputs[193]) | (inputs[693]));
    assign layer0_outputs[4256] = (inputs[688]) ^ (inputs[956]);
    assign layer0_outputs[4257] = ~(inputs[245]) | (inputs[588]);
    assign layer0_outputs[4258] = inputs[780];
    assign layer0_outputs[4259] = ~(inputs[342]) | (inputs[893]);
    assign layer0_outputs[4260] = (inputs[229]) ^ (inputs[1023]);
    assign layer0_outputs[4261] = ~(inputs[431]) | (inputs[389]);
    assign layer0_outputs[4262] = (inputs[450]) | (inputs[883]);
    assign layer0_outputs[4263] = (inputs[254]) | (inputs[656]);
    assign layer0_outputs[4264] = inputs[470];
    assign layer0_outputs[4265] = ~(inputs[517]) | (inputs[1016]);
    assign layer0_outputs[4266] = ~((inputs[149]) ^ (inputs[1018]));
    assign layer0_outputs[4267] = (inputs[712]) ^ (inputs[570]);
    assign layer0_outputs[4268] = ~((inputs[603]) ^ (inputs[975]));
    assign layer0_outputs[4269] = inputs[239];
    assign layer0_outputs[4270] = ~(inputs[753]) | (inputs[279]);
    assign layer0_outputs[4271] = ~((inputs[976]) & (inputs[168]));
    assign layer0_outputs[4272] = (inputs[429]) & ~(inputs[575]);
    assign layer0_outputs[4273] = ~((inputs[2]) ^ (inputs[400]));
    assign layer0_outputs[4274] = (inputs[307]) & ~(inputs[233]);
    assign layer0_outputs[4275] = inputs[249];
    assign layer0_outputs[4276] = ~(inputs[730]);
    assign layer0_outputs[4277] = inputs[489];
    assign layer0_outputs[4278] = (inputs[273]) ^ (inputs[789]);
    assign layer0_outputs[4279] = ~(inputs[212]) | (inputs[515]);
    assign layer0_outputs[4280] = ~(inputs[675]) | (inputs[64]);
    assign layer0_outputs[4281] = (inputs[428]) | (inputs[876]);
    assign layer0_outputs[4282] = ~(inputs[332]) | (inputs[190]);
    assign layer0_outputs[4283] = (inputs[912]) ^ (inputs[720]);
    assign layer0_outputs[4284] = (inputs[181]) | (inputs[420]);
    assign layer0_outputs[4285] = (inputs[1003]) | (inputs[1021]);
    assign layer0_outputs[4286] = ~(inputs[355]) | (inputs[477]);
    assign layer0_outputs[4287] = (inputs[796]) & ~(inputs[48]);
    assign layer0_outputs[4288] = (inputs[710]) & ~(inputs[72]);
    assign layer0_outputs[4289] = inputs[211];
    assign layer0_outputs[4290] = (inputs[589]) & ~(inputs[55]);
    assign layer0_outputs[4291] = ~(inputs[854]) | (inputs[451]);
    assign layer0_outputs[4292] = (inputs[899]) & ~(inputs[738]);
    assign layer0_outputs[4293] = (inputs[793]) | (inputs[225]);
    assign layer0_outputs[4294] = (inputs[689]) & ~(inputs[804]);
    assign layer0_outputs[4295] = ~(inputs[235]);
    assign layer0_outputs[4296] = ~(inputs[372]);
    assign layer0_outputs[4297] = ~(inputs[525]);
    assign layer0_outputs[4298] = (inputs[465]) ^ (inputs[85]);
    assign layer0_outputs[4299] = ~((inputs[774]) ^ (inputs[951]));
    assign layer0_outputs[4300] = ~((inputs[777]) ^ (inputs[786]));
    assign layer0_outputs[4301] = ~(inputs[726]) | (inputs[573]);
    assign layer0_outputs[4302] = ~(inputs[676]);
    assign layer0_outputs[4303] = ~((inputs[189]) & (inputs[787]));
    assign layer0_outputs[4304] = inputs[380];
    assign layer0_outputs[4305] = (inputs[690]) ^ (inputs[693]);
    assign layer0_outputs[4306] = ~(inputs[329]);
    assign layer0_outputs[4307] = ~(inputs[980]);
    assign layer0_outputs[4308] = ~((inputs[3]) | (inputs[704]));
    assign layer0_outputs[4309] = ~(inputs[778]) | (inputs[316]);
    assign layer0_outputs[4310] = (inputs[738]) | (inputs[489]);
    assign layer0_outputs[4311] = (inputs[123]) & ~(inputs[1009]);
    assign layer0_outputs[4312] = inputs[846];
    assign layer0_outputs[4313] = ~((inputs[848]) | (inputs[670]));
    assign layer0_outputs[4314] = (inputs[862]) ^ (inputs[790]);
    assign layer0_outputs[4315] = (inputs[570]) & ~(inputs[832]);
    assign layer0_outputs[4316] = inputs[778];
    assign layer0_outputs[4317] = ~((inputs[793]) | (inputs[740]));
    assign layer0_outputs[4318] = (inputs[87]) | (inputs[154]);
    assign layer0_outputs[4319] = (inputs[812]) ^ (inputs[749]);
    assign layer0_outputs[4320] = ~((inputs[294]) | (inputs[433]));
    assign layer0_outputs[4321] = (inputs[344]) ^ (inputs[645]);
    assign layer0_outputs[4322] = (inputs[941]) & ~(inputs[940]);
    assign layer0_outputs[4323] = ~(inputs[60]) | (inputs[1020]);
    assign layer0_outputs[4324] = ~((inputs[415]) | (inputs[749]));
    assign layer0_outputs[4325] = (inputs[408]) | (inputs[878]);
    assign layer0_outputs[4326] = ~((inputs[914]) ^ (inputs[855]));
    assign layer0_outputs[4327] = inputs[493];
    assign layer0_outputs[4328] = (inputs[167]) & ~(inputs[849]);
    assign layer0_outputs[4329] = inputs[686];
    assign layer0_outputs[4330] = (inputs[752]) & ~(inputs[789]);
    assign layer0_outputs[4331] = ~((inputs[238]) ^ (inputs[533]));
    assign layer0_outputs[4332] = (inputs[49]) | (inputs[756]);
    assign layer0_outputs[4333] = (inputs[331]) & ~(inputs[641]);
    assign layer0_outputs[4334] = ~(inputs[986]) | (inputs[556]);
    assign layer0_outputs[4335] = ~(inputs[343]);
    assign layer0_outputs[4336] = (inputs[916]) ^ (inputs[150]);
    assign layer0_outputs[4337] = inputs[948];
    assign layer0_outputs[4338] = inputs[561];
    assign layer0_outputs[4339] = ~(inputs[733]);
    assign layer0_outputs[4340] = (inputs[390]) ^ (inputs[873]);
    assign layer0_outputs[4341] = ~(inputs[868]);
    assign layer0_outputs[4342] = (inputs[76]) ^ (inputs[404]);
    assign layer0_outputs[4343] = 1'b1;
    assign layer0_outputs[4344] = 1'b1;
    assign layer0_outputs[4345] = ~((inputs[1005]) ^ (inputs[237]));
    assign layer0_outputs[4346] = ~((inputs[392]) ^ (inputs[695]));
    assign layer0_outputs[4347] = (inputs[873]) | (inputs[97]);
    assign layer0_outputs[4348] = ~(inputs[1021]);
    assign layer0_outputs[4349] = ~((inputs[639]) ^ (inputs[260]));
    assign layer0_outputs[4350] = (inputs[557]) ^ (inputs[93]);
    assign layer0_outputs[4351] = 1'b1;
    assign layer0_outputs[4352] = ~(inputs[309]);
    assign layer0_outputs[4353] = ~(inputs[823]) | (inputs[570]);
    assign layer0_outputs[4354] = (inputs[832]) & ~(inputs[234]);
    assign layer0_outputs[4355] = ~((inputs[557]) ^ (inputs[515]));
    assign layer0_outputs[4356] = ~((inputs[887]) ^ (inputs[639]));
    assign layer0_outputs[4357] = (inputs[940]) & ~(inputs[170]);
    assign layer0_outputs[4358] = (inputs[389]) ^ (inputs[60]);
    assign layer0_outputs[4359] = (inputs[528]) & ~(inputs[838]);
    assign layer0_outputs[4360] = (inputs[505]) & ~(inputs[609]);
    assign layer0_outputs[4361] = ~(inputs[591]) | (inputs[285]);
    assign layer0_outputs[4362] = (inputs[105]) | (inputs[863]);
    assign layer0_outputs[4363] = (inputs[714]) & ~(inputs[548]);
    assign layer0_outputs[4364] = ~(inputs[279]) | (inputs[55]);
    assign layer0_outputs[4365] = (inputs[536]) | (inputs[216]);
    assign layer0_outputs[4366] = (inputs[626]) ^ (inputs[778]);
    assign layer0_outputs[4367] = ~(inputs[933]);
    assign layer0_outputs[4368] = ~((inputs[150]) ^ (inputs[710]));
    assign layer0_outputs[4369] = 1'b1;
    assign layer0_outputs[4370] = ~(inputs[305]);
    assign layer0_outputs[4371] = inputs[481];
    assign layer0_outputs[4372] = ~((inputs[748]) | (inputs[98]));
    assign layer0_outputs[4373] = (inputs[719]) | (inputs[702]);
    assign layer0_outputs[4374] = ~(inputs[877]);
    assign layer0_outputs[4375] = ~((inputs[586]) | (inputs[137]));
    assign layer0_outputs[4376] = ~((inputs[791]) | (inputs[907]));
    assign layer0_outputs[4377] = (inputs[103]) | (inputs[566]);
    assign layer0_outputs[4378] = inputs[62];
    assign layer0_outputs[4379] = ~((inputs[273]) | (inputs[741]));
    assign layer0_outputs[4380] = ~(inputs[510]);
    assign layer0_outputs[4381] = ~(inputs[243]);
    assign layer0_outputs[4382] = ~(inputs[910]);
    assign layer0_outputs[4383] = ~(inputs[467]) | (inputs[816]);
    assign layer0_outputs[4384] = (inputs[689]) ^ (inputs[630]);
    assign layer0_outputs[4385] = (inputs[750]) & ~(inputs[347]);
    assign layer0_outputs[4386] = ~((inputs[125]) & (inputs[479]));
    assign layer0_outputs[4387] = ~((inputs[869]) ^ (inputs[792]));
    assign layer0_outputs[4388] = (inputs[929]) & ~(inputs[439]);
    assign layer0_outputs[4389] = ~(inputs[279]) | (inputs[94]);
    assign layer0_outputs[4390] = ~(inputs[596]);
    assign layer0_outputs[4391] = ~(inputs[106]) | (inputs[350]);
    assign layer0_outputs[4392] = (inputs[366]) & ~(inputs[187]);
    assign layer0_outputs[4393] = (inputs[138]) | (inputs[320]);
    assign layer0_outputs[4394] = ~((inputs[208]) & (inputs[407]));
    assign layer0_outputs[4395] = inputs[432];
    assign layer0_outputs[4396] = inputs[384];
    assign layer0_outputs[4397] = ~(inputs[683]);
    assign layer0_outputs[4398] = ~((inputs[169]) ^ (inputs[667]));
    assign layer0_outputs[4399] = inputs[459];
    assign layer0_outputs[4400] = ~(inputs[300]) | (inputs[846]);
    assign layer0_outputs[4401] = ~((inputs[329]) ^ (inputs[992]));
    assign layer0_outputs[4402] = ~(inputs[342]) | (inputs[1019]);
    assign layer0_outputs[4403] = inputs[655];
    assign layer0_outputs[4404] = inputs[857];
    assign layer0_outputs[4405] = inputs[1017];
    assign layer0_outputs[4406] = inputs[152];
    assign layer0_outputs[4407] = ~(inputs[359]) | (inputs[256]);
    assign layer0_outputs[4408] = (inputs[645]) & ~(inputs[358]);
    assign layer0_outputs[4409] = inputs[339];
    assign layer0_outputs[4410] = inputs[1001];
    assign layer0_outputs[4411] = ~(inputs[755]) | (inputs[442]);
    assign layer0_outputs[4412] = (inputs[12]) | (inputs[648]);
    assign layer0_outputs[4413] = (inputs[569]) ^ (inputs[124]);
    assign layer0_outputs[4414] = ~(inputs[777]);
    assign layer0_outputs[4415] = ~((inputs[13]) ^ (inputs[305]));
    assign layer0_outputs[4416] = 1'b1;
    assign layer0_outputs[4417] = (inputs[979]) | (inputs[926]);
    assign layer0_outputs[4418] = ~(inputs[359]) | (inputs[952]);
    assign layer0_outputs[4419] = (inputs[235]) | (inputs[179]);
    assign layer0_outputs[4420] = (inputs[823]) ^ (inputs[913]);
    assign layer0_outputs[4421] = ~((inputs[964]) | (inputs[984]));
    assign layer0_outputs[4422] = (inputs[897]) ^ (inputs[386]);
    assign layer0_outputs[4423] = ~(inputs[846]) | (inputs[37]);
    assign layer0_outputs[4424] = ~((inputs[513]) & (inputs[139]));
    assign layer0_outputs[4425] = inputs[457];
    assign layer0_outputs[4426] = (inputs[622]) ^ (inputs[945]);
    assign layer0_outputs[4427] = ~((inputs[995]) ^ (inputs[200]));
    assign layer0_outputs[4428] = ~((inputs[199]) | (inputs[80]));
    assign layer0_outputs[4429] = (inputs[72]) & ~(inputs[158]);
    assign layer0_outputs[4430] = (inputs[294]) & ~(inputs[700]);
    assign layer0_outputs[4431] = ~(inputs[370]);
    assign layer0_outputs[4432] = (inputs[301]) ^ (inputs[237]);
    assign layer0_outputs[4433] = (inputs[396]) & ~(inputs[643]);
    assign layer0_outputs[4434] = (inputs[649]) & ~(inputs[14]);
    assign layer0_outputs[4435] = ~((inputs[937]) ^ (inputs[218]));
    assign layer0_outputs[4436] = inputs[469];
    assign layer0_outputs[4437] = ~((inputs[23]) | (inputs[612]));
    assign layer0_outputs[4438] = ~(inputs[930]) | (inputs[414]);
    assign layer0_outputs[4439] = (inputs[533]) ^ (inputs[35]);
    assign layer0_outputs[4440] = ~(inputs[621]);
    assign layer0_outputs[4441] = (inputs[733]) ^ (inputs[407]);
    assign layer0_outputs[4442] = inputs[651];
    assign layer0_outputs[4443] = ~((inputs[48]) | (inputs[891]));
    assign layer0_outputs[4444] = inputs[195];
    assign layer0_outputs[4445] = (inputs[457]) | (inputs[617]);
    assign layer0_outputs[4446] = (inputs[425]) & ~(inputs[106]);
    assign layer0_outputs[4447] = ~((inputs[867]) | (inputs[552]));
    assign layer0_outputs[4448] = (inputs[920]) & (inputs[952]);
    assign layer0_outputs[4449] = inputs[532];
    assign layer0_outputs[4450] = ~((inputs[234]) | (inputs[148]));
    assign layer0_outputs[4451] = (inputs[41]) & ~(inputs[471]);
    assign layer0_outputs[4452] = ~((inputs[45]) ^ (inputs[757]));
    assign layer0_outputs[4453] = (inputs[869]) ^ (inputs[397]);
    assign layer0_outputs[4454] = inputs[825];
    assign layer0_outputs[4455] = (inputs[836]) ^ (inputs[547]);
    assign layer0_outputs[4456] = ~((inputs[629]) | (inputs[618]));
    assign layer0_outputs[4457] = ~(inputs[560]);
    assign layer0_outputs[4458] = ~((inputs[460]) | (inputs[256]));
    assign layer0_outputs[4459] = (inputs[406]) ^ (inputs[341]);
    assign layer0_outputs[4460] = ~((inputs[913]) | (inputs[566]));
    assign layer0_outputs[4461] = ~((inputs[708]) ^ (inputs[419]));
    assign layer0_outputs[4462] = inputs[463];
    assign layer0_outputs[4463] = ~(inputs[622]);
    assign layer0_outputs[4464] = ~(inputs[881]) | (inputs[1006]);
    assign layer0_outputs[4465] = ~((inputs[953]) ^ (inputs[974]));
    assign layer0_outputs[4466] = ~(inputs[647]);
    assign layer0_outputs[4467] = (inputs[128]) | (inputs[281]);
    assign layer0_outputs[4468] = ~((inputs[682]) ^ (inputs[591]));
    assign layer0_outputs[4469] = 1'b1;
    assign layer0_outputs[4470] = (inputs[364]) ^ (inputs[998]);
    assign layer0_outputs[4471] = ~((inputs[196]) | (inputs[708]));
    assign layer0_outputs[4472] = (inputs[389]) & ~(inputs[327]);
    assign layer0_outputs[4473] = ~((inputs[38]) | (inputs[32]));
    assign layer0_outputs[4474] = (inputs[595]) & ~(inputs[876]);
    assign layer0_outputs[4475] = ~((inputs[851]) ^ (inputs[361]));
    assign layer0_outputs[4476] = ~(inputs[821]) | (inputs[977]);
    assign layer0_outputs[4477] = inputs[589];
    assign layer0_outputs[4478] = ~((inputs[147]) | (inputs[15]));
    assign layer0_outputs[4479] = ~(inputs[78]) | (inputs[23]);
    assign layer0_outputs[4480] = ~((inputs[405]) ^ (inputs[215]));
    assign layer0_outputs[4481] = ~((inputs[768]) & (inputs[547]));
    assign layer0_outputs[4482] = ~((inputs[84]) ^ (inputs[97]));
    assign layer0_outputs[4483] = 1'b1;
    assign layer0_outputs[4484] = (inputs[114]) | (inputs[138]);
    assign layer0_outputs[4485] = ~(inputs[505]);
    assign layer0_outputs[4486] = inputs[394];
    assign layer0_outputs[4487] = ~((inputs[448]) | (inputs[916]));
    assign layer0_outputs[4488] = inputs[491];
    assign layer0_outputs[4489] = ~((inputs[469]) | (inputs[824]));
    assign layer0_outputs[4490] = (inputs[871]) | (inputs[669]);
    assign layer0_outputs[4491] = ~(inputs[455]) | (inputs[28]);
    assign layer0_outputs[4492] = ~((inputs[443]) | (inputs[476]));
    assign layer0_outputs[4493] = ~((inputs[264]) ^ (inputs[770]));
    assign layer0_outputs[4494] = inputs[683];
    assign layer0_outputs[4495] = 1'b1;
    assign layer0_outputs[4496] = inputs[535];
    assign layer0_outputs[4497] = ~((inputs[796]) ^ (inputs[747]));
    assign layer0_outputs[4498] = (inputs[36]) | (inputs[655]);
    assign layer0_outputs[4499] = (inputs[660]) | (inputs[441]);
    assign layer0_outputs[4500] = (inputs[234]) | (inputs[251]);
    assign layer0_outputs[4501] = (inputs[489]) | (inputs[409]);
    assign layer0_outputs[4502] = (inputs[896]) | (inputs[684]);
    assign layer0_outputs[4503] = (inputs[953]) | (inputs[530]);
    assign layer0_outputs[4504] = (inputs[752]) & ~(inputs[72]);
    assign layer0_outputs[4505] = (inputs[821]) & ~(inputs[950]);
    assign layer0_outputs[4506] = ~(inputs[146]);
    assign layer0_outputs[4507] = ~(inputs[1006]);
    assign layer0_outputs[4508] = (inputs[385]) ^ (inputs[57]);
    assign layer0_outputs[4509] = ~(inputs[794]);
    assign layer0_outputs[4510] = 1'b1;
    assign layer0_outputs[4511] = (inputs[708]) & ~(inputs[550]);
    assign layer0_outputs[4512] = ~((inputs[268]) | (inputs[530]));
    assign layer0_outputs[4513] = (inputs[442]) & ~(inputs[640]);
    assign layer0_outputs[4514] = (inputs[460]) & ~(inputs[1010]);
    assign layer0_outputs[4515] = (inputs[685]) ^ (inputs[681]);
    assign layer0_outputs[4516] = inputs[142];
    assign layer0_outputs[4517] = (inputs[823]) | (inputs[1017]);
    assign layer0_outputs[4518] = ~(inputs[71]) | (inputs[61]);
    assign layer0_outputs[4519] = ~(inputs[234]);
    assign layer0_outputs[4520] = ~(inputs[783]) | (inputs[743]);
    assign layer0_outputs[4521] = (inputs[353]) & ~(inputs[985]);
    assign layer0_outputs[4522] = ~(inputs[527]) | (inputs[456]);
    assign layer0_outputs[4523] = inputs[706];
    assign layer0_outputs[4524] = 1'b0;
    assign layer0_outputs[4525] = ~(inputs[528]);
    assign layer0_outputs[4526] = ~(inputs[524]);
    assign layer0_outputs[4527] = inputs[483];
    assign layer0_outputs[4528] = ~(inputs[61]);
    assign layer0_outputs[4529] = ~(inputs[716]);
    assign layer0_outputs[4530] = ~(inputs[493]);
    assign layer0_outputs[4531] = (inputs[658]) & ~(inputs[922]);
    assign layer0_outputs[4532] = ~((inputs[166]) | (inputs[557]));
    assign layer0_outputs[4533] = ~((inputs[926]) | (inputs[826]));
    assign layer0_outputs[4534] = ~(inputs[737]) | (inputs[449]);
    assign layer0_outputs[4535] = (inputs[710]) | (inputs[549]);
    assign layer0_outputs[4536] = (inputs[254]) ^ (inputs[465]);
    assign layer0_outputs[4537] = ~((inputs[883]) ^ (inputs[174]));
    assign layer0_outputs[4538] = ~(inputs[987]) | (inputs[732]);
    assign layer0_outputs[4539] = inputs[456];
    assign layer0_outputs[4540] = ~(inputs[42]) | (inputs[22]);
    assign layer0_outputs[4541] = ~(inputs[907]) | (inputs[549]);
    assign layer0_outputs[4542] = ~(inputs[956]);
    assign layer0_outputs[4543] = (inputs[5]) & ~(inputs[794]);
    assign layer0_outputs[4544] = inputs[112];
    assign layer0_outputs[4545] = (inputs[478]) ^ (inputs[483]);
    assign layer0_outputs[4546] = (inputs[272]) & ~(inputs[7]);
    assign layer0_outputs[4547] = (inputs[437]) ^ (inputs[718]);
    assign layer0_outputs[4548] = (inputs[142]) ^ (inputs[587]);
    assign layer0_outputs[4549] = ~((inputs[564]) | (inputs[501]));
    assign layer0_outputs[4550] = ~((inputs[522]) | (inputs[579]));
    assign layer0_outputs[4551] = ~(inputs[339]) | (inputs[177]);
    assign layer0_outputs[4552] = ~((inputs[20]) | (inputs[244]));
    assign layer0_outputs[4553] = (inputs[754]) ^ (inputs[226]);
    assign layer0_outputs[4554] = ~(inputs[382]) | (inputs[518]);
    assign layer0_outputs[4555] = ~((inputs[356]) & (inputs[93]));
    assign layer0_outputs[4556] = ~((inputs[565]) ^ (inputs[511]));
    assign layer0_outputs[4557] = 1'b0;
    assign layer0_outputs[4558] = (inputs[259]) ^ (inputs[482]);
    assign layer0_outputs[4559] = inputs[241];
    assign layer0_outputs[4560] = ~((inputs[893]) ^ (inputs[47]));
    assign layer0_outputs[4561] = inputs[120];
    assign layer0_outputs[4562] = (inputs[102]) | (inputs[837]);
    assign layer0_outputs[4563] = inputs[277];
    assign layer0_outputs[4564] = ~(inputs[738]) | (inputs[558]);
    assign layer0_outputs[4565] = ~((inputs[269]) ^ (inputs[387]));
    assign layer0_outputs[4566] = 1'b0;
    assign layer0_outputs[4567] = (inputs[461]) ^ (inputs[487]);
    assign layer0_outputs[4568] = (inputs[977]) ^ (inputs[243]);
    assign layer0_outputs[4569] = ~((inputs[340]) ^ (inputs[341]));
    assign layer0_outputs[4570] = (inputs[422]) | (inputs[411]);
    assign layer0_outputs[4571] = (inputs[238]) | (inputs[30]);
    assign layer0_outputs[4572] = (inputs[614]) ^ (inputs[312]);
    assign layer0_outputs[4573] = ~(inputs[363]);
    assign layer0_outputs[4574] = (inputs[234]) & ~(inputs[900]);
    assign layer0_outputs[4575] = ~(inputs[361]) | (inputs[805]);
    assign layer0_outputs[4576] = inputs[244];
    assign layer0_outputs[4577] = (inputs[11]) & ~(inputs[998]);
    assign layer0_outputs[4578] = (inputs[185]) & ~(inputs[769]);
    assign layer0_outputs[4579] = inputs[345];
    assign layer0_outputs[4580] = (inputs[295]) | (inputs[764]);
    assign layer0_outputs[4581] = (inputs[346]) | (inputs[129]);
    assign layer0_outputs[4582] = ~((inputs[27]) & (inputs[55]));
    assign layer0_outputs[4583] = (inputs[957]) ^ (inputs[265]);
    assign layer0_outputs[4584] = (inputs[195]) ^ (inputs[241]);
    assign layer0_outputs[4585] = inputs[681];
    assign layer0_outputs[4586] = ~((inputs[942]) ^ (inputs[994]));
    assign layer0_outputs[4587] = (inputs[113]) | (inputs[267]);
    assign layer0_outputs[4588] = (inputs[357]) | (inputs[406]);
    assign layer0_outputs[4589] = (inputs[57]) ^ (inputs[132]);
    assign layer0_outputs[4590] = (inputs[335]) | (inputs[10]);
    assign layer0_outputs[4591] = (inputs[911]) & ~(inputs[60]);
    assign layer0_outputs[4592] = ~((inputs[636]) | (inputs[743]));
    assign layer0_outputs[4593] = 1'b0;
    assign layer0_outputs[4594] = 1'b1;
    assign layer0_outputs[4595] = ~((inputs[540]) | (inputs[923]));
    assign layer0_outputs[4596] = ~((inputs[236]) | (inputs[609]));
    assign layer0_outputs[4597] = ~((inputs[714]) | (inputs[779]));
    assign layer0_outputs[4598] = ~(inputs[363]);
    assign layer0_outputs[4599] = (inputs[56]) & ~(inputs[552]);
    assign layer0_outputs[4600] = (inputs[405]) & ~(inputs[223]);
    assign layer0_outputs[4601] = ~((inputs[795]) ^ (inputs[615]));
    assign layer0_outputs[4602] = inputs[675];
    assign layer0_outputs[4603] = ~((inputs[603]) ^ (inputs[692]));
    assign layer0_outputs[4604] = (inputs[834]) | (inputs[202]);
    assign layer0_outputs[4605] = ~(inputs[457]) | (inputs[981]);
    assign layer0_outputs[4606] = ~(inputs[777]) | (inputs[537]);
    assign layer0_outputs[4607] = ~(inputs[1001]) | (inputs[425]);
    assign layer0_outputs[4608] = (inputs[956]) | (inputs[690]);
    assign layer0_outputs[4609] = inputs[533];
    assign layer0_outputs[4610] = ~((inputs[445]) ^ (inputs[581]));
    assign layer0_outputs[4611] = ~(inputs[15]);
    assign layer0_outputs[4612] = ~((inputs[93]) | (inputs[363]));
    assign layer0_outputs[4613] = inputs[952];
    assign layer0_outputs[4614] = ~(inputs[302]) | (inputs[643]);
    assign layer0_outputs[4615] = ~(inputs[592]) | (inputs[139]);
    assign layer0_outputs[4616] = (inputs[464]) ^ (inputs[25]);
    assign layer0_outputs[4617] = inputs[366];
    assign layer0_outputs[4618] = (inputs[816]) & ~(inputs[477]);
    assign layer0_outputs[4619] = inputs[297];
    assign layer0_outputs[4620] = ~(inputs[832]);
    assign layer0_outputs[4621] = (inputs[135]) ^ (inputs[719]);
    assign layer0_outputs[4622] = inputs[651];
    assign layer0_outputs[4623] = (inputs[799]) | (inputs[7]);
    assign layer0_outputs[4624] = ~((inputs[178]) | (inputs[922]));
    assign layer0_outputs[4625] = ~(inputs[975]) | (inputs[701]);
    assign layer0_outputs[4626] = ~(inputs[241]);
    assign layer0_outputs[4627] = (inputs[351]) | (inputs[344]);
    assign layer0_outputs[4628] = ~((inputs[700]) | (inputs[495]));
    assign layer0_outputs[4629] = (inputs[281]) | (inputs[406]);
    assign layer0_outputs[4630] = (inputs[1017]) | (inputs[736]);
    assign layer0_outputs[4631] = ~(inputs[685]);
    assign layer0_outputs[4632] = inputs[544];
    assign layer0_outputs[4633] = (inputs[388]) | (inputs[395]);
    assign layer0_outputs[4634] = (inputs[983]) | (inputs[517]);
    assign layer0_outputs[4635] = (inputs[664]) | (inputs[144]);
    assign layer0_outputs[4636] = ~((inputs[321]) & (inputs[959]));
    assign layer0_outputs[4637] = (inputs[304]) ^ (inputs[58]);
    assign layer0_outputs[4638] = (inputs[109]) | (inputs[204]);
    assign layer0_outputs[4639] = (inputs[756]) ^ (inputs[93]);
    assign layer0_outputs[4640] = inputs[836];
    assign layer0_outputs[4641] = ~((inputs[280]) ^ (inputs[368]));
    assign layer0_outputs[4642] = 1'b0;
    assign layer0_outputs[4643] = 1'b1;
    assign layer0_outputs[4644] = ~(inputs[483]) | (inputs[1022]);
    assign layer0_outputs[4645] = (inputs[636]) | (inputs[92]);
    assign layer0_outputs[4646] = ~(inputs[141]);
    assign layer0_outputs[4647] = (inputs[251]) ^ (inputs[312]);
    assign layer0_outputs[4648] = ~((inputs[805]) | (inputs[304]));
    assign layer0_outputs[4649] = ~(inputs[199]);
    assign layer0_outputs[4650] = (inputs[371]) ^ (inputs[829]);
    assign layer0_outputs[4651] = ~((inputs[411]) ^ (inputs[360]));
    assign layer0_outputs[4652] = ~((inputs[766]) | (inputs[604]));
    assign layer0_outputs[4653] = ~(inputs[178]);
    assign layer0_outputs[4654] = ~(inputs[578]);
    assign layer0_outputs[4655] = ~((inputs[45]) | (inputs[320]));
    assign layer0_outputs[4656] = inputs[319];
    assign layer0_outputs[4657] = inputs[600];
    assign layer0_outputs[4658] = (inputs[901]) ^ (inputs[83]);
    assign layer0_outputs[4659] = (inputs[654]) & ~(inputs[119]);
    assign layer0_outputs[4660] = (inputs[761]) | (inputs[124]);
    assign layer0_outputs[4661] = (inputs[686]) | (inputs[319]);
    assign layer0_outputs[4662] = (inputs[178]) | (inputs[253]);
    assign layer0_outputs[4663] = ~((inputs[392]) | (inputs[1008]));
    assign layer0_outputs[4664] = (inputs[358]) | (inputs[310]);
    assign layer0_outputs[4665] = (inputs[831]) ^ (inputs[408]);
    assign layer0_outputs[4666] = (inputs[43]) & ~(inputs[418]);
    assign layer0_outputs[4667] = (inputs[641]) | (inputs[227]);
    assign layer0_outputs[4668] = ~(inputs[789]) | (inputs[995]);
    assign layer0_outputs[4669] = ~(inputs[755]) | (inputs[881]);
    assign layer0_outputs[4670] = ~((inputs[1002]) | (inputs[215]));
    assign layer0_outputs[4671] = ~((inputs[294]) | (inputs[371]));
    assign layer0_outputs[4672] = (inputs[732]) & ~(inputs[360]);
    assign layer0_outputs[4673] = (inputs[175]) & ~(inputs[376]);
    assign layer0_outputs[4674] = inputs[847];
    assign layer0_outputs[4675] = (inputs[654]) | (inputs[91]);
    assign layer0_outputs[4676] = ~(inputs[600]) | (inputs[453]);
    assign layer0_outputs[4677] = (inputs[825]) | (inputs[395]);
    assign layer0_outputs[4678] = inputs[473];
    assign layer0_outputs[4679] = 1'b0;
    assign layer0_outputs[4680] = inputs[831];
    assign layer0_outputs[4681] = (inputs[399]) | (inputs[694]);
    assign layer0_outputs[4682] = ~((inputs[416]) ^ (inputs[168]));
    assign layer0_outputs[4683] = ~(inputs[365]);
    assign layer0_outputs[4684] = (inputs[583]) ^ (inputs[626]);
    assign layer0_outputs[4685] = (inputs[93]) & (inputs[280]);
    assign layer0_outputs[4686] = 1'b0;
    assign layer0_outputs[4687] = ~(inputs[242]);
    assign layer0_outputs[4688] = (inputs[86]) | (inputs[267]);
    assign layer0_outputs[4689] = (inputs[416]) & ~(inputs[614]);
    assign layer0_outputs[4690] = ~(inputs[397]);
    assign layer0_outputs[4691] = ~((inputs[787]) | (inputs[540]));
    assign layer0_outputs[4692] = inputs[330];
    assign layer0_outputs[4693] = ~(inputs[556]);
    assign layer0_outputs[4694] = (inputs[1015]) | (inputs[679]);
    assign layer0_outputs[4695] = (inputs[934]) & (inputs[450]);
    assign layer0_outputs[4696] = ~(inputs[372]) | (inputs[606]);
    assign layer0_outputs[4697] = ~((inputs[369]) | (inputs[696]));
    assign layer0_outputs[4698] = inputs[933];
    assign layer0_outputs[4699] = inputs[780];
    assign layer0_outputs[4700] = ~((inputs[99]) & (inputs[291]));
    assign layer0_outputs[4701] = ~(inputs[141]) | (inputs[229]);
    assign layer0_outputs[4702] = ~(inputs[886]);
    assign layer0_outputs[4703] = inputs[371];
    assign layer0_outputs[4704] = ~(inputs[477]) | (inputs[522]);
    assign layer0_outputs[4705] = ~((inputs[303]) | (inputs[165]));
    assign layer0_outputs[4706] = (inputs[153]) | (inputs[724]);
    assign layer0_outputs[4707] = 1'b0;
    assign layer0_outputs[4708] = ~((inputs[177]) ^ (inputs[751]));
    assign layer0_outputs[4709] = (inputs[74]) & ~(inputs[174]);
    assign layer0_outputs[4710] = ~(inputs[948]) | (inputs[862]);
    assign layer0_outputs[4711] = (inputs[84]) ^ (inputs[127]);
    assign layer0_outputs[4712] = (inputs[585]) & ~(inputs[127]);
    assign layer0_outputs[4713] = ~(inputs[558]) | (inputs[122]);
    assign layer0_outputs[4714] = inputs[464];
    assign layer0_outputs[4715] = ~(inputs[136]) | (inputs[275]);
    assign layer0_outputs[4716] = ~(inputs[361]);
    assign layer0_outputs[4717] = ~((inputs[184]) ^ (inputs[58]));
    assign layer0_outputs[4718] = ~((inputs[748]) | (inputs[53]));
    assign layer0_outputs[4719] = ~((inputs[119]) | (inputs[491]));
    assign layer0_outputs[4720] = (inputs[657]) & ~(inputs[905]);
    assign layer0_outputs[4721] = ~((inputs[799]) ^ (inputs[749]));
    assign layer0_outputs[4722] = ~((inputs[503]) | (inputs[217]));
    assign layer0_outputs[4723] = ~(inputs[651]);
    assign layer0_outputs[4724] = (inputs[227]) & (inputs[349]);
    assign layer0_outputs[4725] = ~(inputs[153]) | (inputs[12]);
    assign layer0_outputs[4726] = ~((inputs[423]) | (inputs[183]));
    assign layer0_outputs[4727] = ~(inputs[818]);
    assign layer0_outputs[4728] = (inputs[979]) & ~(inputs[149]);
    assign layer0_outputs[4729] = ~((inputs[101]) & (inputs[62]));
    assign layer0_outputs[4730] = (inputs[773]) & ~(inputs[452]);
    assign layer0_outputs[4731] = 1'b1;
    assign layer0_outputs[4732] = 1'b1;
    assign layer0_outputs[4733] = (inputs[483]) ^ (inputs[865]);
    assign layer0_outputs[4734] = ~(inputs[619]);
    assign layer0_outputs[4735] = ~((inputs[21]) ^ (inputs[59]));
    assign layer0_outputs[4736] = inputs[971];
    assign layer0_outputs[4737] = inputs[208];
    assign layer0_outputs[4738] = ~(inputs[844]);
    assign layer0_outputs[4739] = ~((inputs[337]) ^ (inputs[255]));
    assign layer0_outputs[4740] = (inputs[109]) ^ (inputs[948]);
    assign layer0_outputs[4741] = ~(inputs[292]);
    assign layer0_outputs[4742] = ~(inputs[748]);
    assign layer0_outputs[4743] = 1'b0;
    assign layer0_outputs[4744] = (inputs[727]) ^ (inputs[636]);
    assign layer0_outputs[4745] = ~((inputs[240]) | (inputs[768]));
    assign layer0_outputs[4746] = ~((inputs[112]) | (inputs[95]));
    assign layer0_outputs[4747] = inputs[624];
    assign layer0_outputs[4748] = ~((inputs[659]) | (inputs[579]));
    assign layer0_outputs[4749] = (inputs[450]) & ~(inputs[788]);
    assign layer0_outputs[4750] = ~(inputs[43]);
    assign layer0_outputs[4751] = (inputs[457]) | (inputs[855]);
    assign layer0_outputs[4752] = ~((inputs[283]) ^ (inputs[452]));
    assign layer0_outputs[4753] = ~((inputs[717]) ^ (inputs[578]));
    assign layer0_outputs[4754] = 1'b0;
    assign layer0_outputs[4755] = ~((inputs[660]) | (inputs[126]));
    assign layer0_outputs[4756] = ~(inputs[496]);
    assign layer0_outputs[4757] = (inputs[741]) ^ (inputs[871]);
    assign layer0_outputs[4758] = (inputs[249]) & ~(inputs[710]);
    assign layer0_outputs[4759] = (inputs[325]) | (inputs[371]);
    assign layer0_outputs[4760] = ~(inputs[616]);
    assign layer0_outputs[4761] = inputs[521];
    assign layer0_outputs[4762] = (inputs[473]) | (inputs[452]);
    assign layer0_outputs[4763] = ~(inputs[152]) | (inputs[957]);
    assign layer0_outputs[4764] = ~((inputs[353]) | (inputs[277]));
    assign layer0_outputs[4765] = (inputs[367]) & ~(inputs[683]);
    assign layer0_outputs[4766] = (inputs[840]) ^ (inputs[276]);
    assign layer0_outputs[4767] = ~((inputs[355]) ^ (inputs[948]));
    assign layer0_outputs[4768] = ~((inputs[450]) | (inputs[340]));
    assign layer0_outputs[4769] = ~(inputs[442]) | (inputs[434]);
    assign layer0_outputs[4770] = ~((inputs[30]) | (inputs[888]));
    assign layer0_outputs[4771] = 1'b1;
    assign layer0_outputs[4772] = (inputs[983]) ^ (inputs[665]);
    assign layer0_outputs[4773] = 1'b0;
    assign layer0_outputs[4774] = (inputs[165]) ^ (inputs[425]);
    assign layer0_outputs[4775] = (inputs[400]) & (inputs[892]);
    assign layer0_outputs[4776] = ~(inputs[899]);
    assign layer0_outputs[4777] = ~(inputs[637]);
    assign layer0_outputs[4778] = (inputs[188]) ^ (inputs[685]);
    assign layer0_outputs[4779] = (inputs[183]) | (inputs[268]);
    assign layer0_outputs[4780] = ~((inputs[775]) & (inputs[626]));
    assign layer0_outputs[4781] = ~(inputs[605]);
    assign layer0_outputs[4782] = ~((inputs[282]) | (inputs[779]));
    assign layer0_outputs[4783] = ~(inputs[618]);
    assign layer0_outputs[4784] = 1'b1;
    assign layer0_outputs[4785] = (inputs[434]) ^ (inputs[990]);
    assign layer0_outputs[4786] = ~((inputs[911]) & (inputs[232]));
    assign layer0_outputs[4787] = (inputs[776]) | (inputs[880]);
    assign layer0_outputs[4788] = (inputs[167]) | (inputs[207]);
    assign layer0_outputs[4789] = ~((inputs[709]) ^ (inputs[167]));
    assign layer0_outputs[4790] = (inputs[433]) ^ (inputs[479]);
    assign layer0_outputs[4791] = ~(inputs[543]);
    assign layer0_outputs[4792] = 1'b1;
    assign layer0_outputs[4793] = inputs[409];
    assign layer0_outputs[4794] = 1'b1;
    assign layer0_outputs[4795] = ~(inputs[528]);
    assign layer0_outputs[4796] = ~((inputs[330]) ^ (inputs[843]));
    assign layer0_outputs[4797] = ~(inputs[335]) | (inputs[969]);
    assign layer0_outputs[4798] = ~(inputs[806]);
    assign layer0_outputs[4799] = ~((inputs[417]) | (inputs[1006]));
    assign layer0_outputs[4800] = ~((inputs[796]) & (inputs[28]));
    assign layer0_outputs[4801] = 1'b1;
    assign layer0_outputs[4802] = ~((inputs[701]) | (inputs[207]));
    assign layer0_outputs[4803] = (inputs[964]) | (inputs[468]);
    assign layer0_outputs[4804] = (inputs[555]) & ~(inputs[914]);
    assign layer0_outputs[4805] = inputs[274];
    assign layer0_outputs[4806] = (inputs[712]) | (inputs[947]);
    assign layer0_outputs[4807] = ~(inputs[410]);
    assign layer0_outputs[4808] = ~(inputs[597]) | (inputs[223]);
    assign layer0_outputs[4809] = ~(inputs[361]);
    assign layer0_outputs[4810] = (inputs[1004]) | (inputs[420]);
    assign layer0_outputs[4811] = ~(inputs[283]);
    assign layer0_outputs[4812] = ~((inputs[172]) ^ (inputs[217]));
    assign layer0_outputs[4813] = (inputs[892]) | (inputs[459]);
    assign layer0_outputs[4814] = (inputs[439]) & (inputs[407]);
    assign layer0_outputs[4815] = (inputs[978]) | (inputs[404]);
    assign layer0_outputs[4816] = ~(inputs[406]) | (inputs[221]);
    assign layer0_outputs[4817] = (inputs[225]) | (inputs[784]);
    assign layer0_outputs[4818] = ~((inputs[880]) | (inputs[745]));
    assign layer0_outputs[4819] = (inputs[459]) ^ (inputs[506]);
    assign layer0_outputs[4820] = (inputs[268]) | (inputs[444]);
    assign layer0_outputs[4821] = 1'b1;
    assign layer0_outputs[4822] = ~((inputs[231]) ^ (inputs[470]));
    assign layer0_outputs[4823] = ~(inputs[456]);
    assign layer0_outputs[4824] = ~(inputs[333]);
    assign layer0_outputs[4825] = ~((inputs[17]) | (inputs[294]));
    assign layer0_outputs[4826] = (inputs[744]) & ~(inputs[433]);
    assign layer0_outputs[4827] = ~((inputs[893]) & (inputs[895]));
    assign layer0_outputs[4828] = (inputs[458]) & ~(inputs[655]);
    assign layer0_outputs[4829] = ~(inputs[1020]) | (inputs[511]);
    assign layer0_outputs[4830] = (inputs[640]) | (inputs[415]);
    assign layer0_outputs[4831] = (inputs[283]) & (inputs[383]);
    assign layer0_outputs[4832] = (inputs[847]) & ~(inputs[579]);
    assign layer0_outputs[4833] = ~(inputs[745]) | (inputs[324]);
    assign layer0_outputs[4834] = inputs[260];
    assign layer0_outputs[4835] = inputs[506];
    assign layer0_outputs[4836] = ~(inputs[141]) | (inputs[949]);
    assign layer0_outputs[4837] = ~((inputs[1005]) ^ (inputs[172]));
    assign layer0_outputs[4838] = (inputs[173]) ^ (inputs[739]);
    assign layer0_outputs[4839] = (inputs[897]) | (inputs[855]);
    assign layer0_outputs[4840] = 1'b0;
    assign layer0_outputs[4841] = 1'b0;
    assign layer0_outputs[4842] = (inputs[171]) ^ (inputs[898]);
    assign layer0_outputs[4843] = ~((inputs[157]) ^ (inputs[296]));
    assign layer0_outputs[4844] = 1'b1;
    assign layer0_outputs[4845] = (inputs[77]) & (inputs[679]);
    assign layer0_outputs[4846] = ~((inputs[186]) ^ (inputs[986]));
    assign layer0_outputs[4847] = ~(inputs[651]);
    assign layer0_outputs[4848] = inputs[249];
    assign layer0_outputs[4849] = (inputs[510]) ^ (inputs[1011]);
    assign layer0_outputs[4850] = (inputs[518]) & ~(inputs[82]);
    assign layer0_outputs[4851] = (inputs[738]) ^ (inputs[647]);
    assign layer0_outputs[4852] = ~((inputs[751]) ^ (inputs[511]));
    assign layer0_outputs[4853] = (inputs[155]) ^ (inputs[89]);
    assign layer0_outputs[4854] = inputs[400];
    assign layer0_outputs[4855] = ~((inputs[723]) | (inputs[1009]));
    assign layer0_outputs[4856] = ~((inputs[309]) | (inputs[445]));
    assign layer0_outputs[4857] = (inputs[552]) & ~(inputs[997]);
    assign layer0_outputs[4858] = (inputs[813]) & ~(inputs[482]);
    assign layer0_outputs[4859] = ~((inputs[889]) | (inputs[741]));
    assign layer0_outputs[4860] = (inputs[450]) ^ (inputs[991]);
    assign layer0_outputs[4861] = (inputs[581]) ^ (inputs[709]);
    assign layer0_outputs[4862] = ~((inputs[825]) | (inputs[944]));
    assign layer0_outputs[4863] = ~(inputs[293]);
    assign layer0_outputs[4864] = (inputs[775]) & ~(inputs[885]);
    assign layer0_outputs[4865] = ~((inputs[735]) | (inputs[299]));
    assign layer0_outputs[4866] = (inputs[598]) | (inputs[438]);
    assign layer0_outputs[4867] = ~(inputs[233]) | (inputs[213]);
    assign layer0_outputs[4868] = (inputs[409]) | (inputs[682]);
    assign layer0_outputs[4869] = 1'b1;
    assign layer0_outputs[4870] = (inputs[161]) ^ (inputs[606]);
    assign layer0_outputs[4871] = (inputs[373]) & ~(inputs[587]);
    assign layer0_outputs[4872] = (inputs[667]) | (inputs[210]);
    assign layer0_outputs[4873] = inputs[272];
    assign layer0_outputs[4874] = (inputs[365]) ^ (inputs[448]);
    assign layer0_outputs[4875] = (inputs[608]) & (inputs[56]);
    assign layer0_outputs[4876] = ~(inputs[336]);
    assign layer0_outputs[4877] = (inputs[103]) ^ (inputs[357]);
    assign layer0_outputs[4878] = ~(inputs[196]);
    assign layer0_outputs[4879] = (inputs[445]) ^ (inputs[172]);
    assign layer0_outputs[4880] = ~(inputs[682]);
    assign layer0_outputs[4881] = inputs[836];
    assign layer0_outputs[4882] = ~(inputs[332]);
    assign layer0_outputs[4883] = ~(inputs[876]);
    assign layer0_outputs[4884] = ~((inputs[721]) | (inputs[672]));
    assign layer0_outputs[4885] = ~(inputs[160]) | (inputs[246]);
    assign layer0_outputs[4886] = (inputs[182]) & ~(inputs[873]);
    assign layer0_outputs[4887] = inputs[922];
    assign layer0_outputs[4888] = inputs[668];
    assign layer0_outputs[4889] = inputs[223];
    assign layer0_outputs[4890] = (inputs[767]) ^ (inputs[244]);
    assign layer0_outputs[4891] = (inputs[813]) & ~(inputs[475]);
    assign layer0_outputs[4892] = (inputs[990]) & ~(inputs[952]);
    assign layer0_outputs[4893] = (inputs[142]) | (inputs[757]);
    assign layer0_outputs[4894] = ~(inputs[566]) | (inputs[837]);
    assign layer0_outputs[4895] = ~(inputs[585]) | (inputs[195]);
    assign layer0_outputs[4896] = ~((inputs[272]) ^ (inputs[363]));
    assign layer0_outputs[4897] = ~(inputs[339]) | (inputs[150]);
    assign layer0_outputs[4898] = (inputs[72]) ^ (inputs[312]);
    assign layer0_outputs[4899] = ~(inputs[256]);
    assign layer0_outputs[4900] = ~((inputs[945]) & (inputs[424]));
    assign layer0_outputs[4901] = inputs[273];
    assign layer0_outputs[4902] = ~((inputs[8]) | (inputs[551]));
    assign layer0_outputs[4903] = inputs[865];
    assign layer0_outputs[4904] = ~((inputs[476]) | (inputs[586]));
    assign layer0_outputs[4905] = 1'b1;
    assign layer0_outputs[4906] = 1'b0;
    assign layer0_outputs[4907] = (inputs[240]) ^ (inputs[352]);
    assign layer0_outputs[4908] = ~((inputs[912]) | (inputs[594]));
    assign layer0_outputs[4909] = (inputs[298]) ^ (inputs[706]);
    assign layer0_outputs[4910] = 1'b0;
    assign layer0_outputs[4911] = ~((inputs[828]) & (inputs[7]));
    assign layer0_outputs[4912] = ~(inputs[81]) | (inputs[576]);
    assign layer0_outputs[4913] = inputs[762];
    assign layer0_outputs[4914] = ~((inputs[184]) ^ (inputs[470]));
    assign layer0_outputs[4915] = inputs[231];
    assign layer0_outputs[4916] = ~((inputs[578]) | (inputs[464]));
    assign layer0_outputs[4917] = ~((inputs[476]) ^ (inputs[85]));
    assign layer0_outputs[4918] = ~(inputs[513]);
    assign layer0_outputs[4919] = (inputs[783]) & ~(inputs[348]);
    assign layer0_outputs[4920] = ~((inputs[112]) ^ (inputs[606]));
    assign layer0_outputs[4921] = ~(inputs[597]) | (inputs[604]);
    assign layer0_outputs[4922] = (inputs[651]) ^ (inputs[496]);
    assign layer0_outputs[4923] = inputs[529];
    assign layer0_outputs[4924] = ~(inputs[287]) | (inputs[443]);
    assign layer0_outputs[4925] = ~(inputs[777]);
    assign layer0_outputs[4926] = ~(inputs[497]);
    assign layer0_outputs[4927] = (inputs[164]) | (inputs[648]);
    assign layer0_outputs[4928] = ~((inputs[909]) | (inputs[462]));
    assign layer0_outputs[4929] = ~((inputs[386]) & (inputs[160]));
    assign layer0_outputs[4930] = (inputs[347]) & ~(inputs[17]);
    assign layer0_outputs[4931] = ~(inputs[881]) | (inputs[736]);
    assign layer0_outputs[4932] = (inputs[940]) ^ (inputs[572]);
    assign layer0_outputs[4933] = ~(inputs[498]);
    assign layer0_outputs[4934] = (inputs[428]) & ~(inputs[1015]);
    assign layer0_outputs[4935] = (inputs[740]) | (inputs[19]);
    assign layer0_outputs[4936] = ~(inputs[533]);
    assign layer0_outputs[4937] = ~(inputs[67]) | (inputs[688]);
    assign layer0_outputs[4938] = (inputs[908]) ^ (inputs[75]);
    assign layer0_outputs[4939] = ~((inputs[325]) | (inputs[512]));
    assign layer0_outputs[4940] = ~((inputs[182]) | (inputs[969]));
    assign layer0_outputs[4941] = ~((inputs[1003]) ^ (inputs[471]));
    assign layer0_outputs[4942] = 1'b0;
    assign layer0_outputs[4943] = ~(inputs[961]);
    assign layer0_outputs[4944] = ~((inputs[663]) | (inputs[208]));
    assign layer0_outputs[4945] = (inputs[45]) | (inputs[636]);
    assign layer0_outputs[4946] = (inputs[324]) & ~(inputs[86]);
    assign layer0_outputs[4947] = ~((inputs[362]) | (inputs[376]));
    assign layer0_outputs[4948] = inputs[297];
    assign layer0_outputs[4949] = ~(inputs[254]);
    assign layer0_outputs[4950] = ~(inputs[268]);
    assign layer0_outputs[4951] = ~((inputs[295]) | (inputs[871]));
    assign layer0_outputs[4952] = (inputs[634]) & ~(inputs[544]);
    assign layer0_outputs[4953] = ~(inputs[657]);
    assign layer0_outputs[4954] = ~(inputs[486]) | (inputs[315]);
    assign layer0_outputs[4955] = (inputs[494]) & ~(inputs[27]);
    assign layer0_outputs[4956] = ~((inputs[909]) | (inputs[630]));
    assign layer0_outputs[4957] = inputs[181];
    assign layer0_outputs[4958] = inputs[518];
    assign layer0_outputs[4959] = (inputs[124]) & ~(inputs[990]);
    assign layer0_outputs[4960] = ~((inputs[482]) ^ (inputs[726]));
    assign layer0_outputs[4961] = inputs[884];
    assign layer0_outputs[4962] = (inputs[331]) | (inputs[552]);
    assign layer0_outputs[4963] = ~(inputs[532]);
    assign layer0_outputs[4964] = inputs[914];
    assign layer0_outputs[4965] = ~((inputs[364]) & (inputs[921]));
    assign layer0_outputs[4966] = (inputs[83]) ^ (inputs[208]);
    assign layer0_outputs[4967] = 1'b0;
    assign layer0_outputs[4968] = ~((inputs[289]) | (inputs[40]));
    assign layer0_outputs[4969] = (inputs[702]) & ~(inputs[792]);
    assign layer0_outputs[4970] = ~((inputs[592]) ^ (inputs[1003]));
    assign layer0_outputs[4971] = ~((inputs[313]) | (inputs[484]));
    assign layer0_outputs[4972] = ~(inputs[160]);
    assign layer0_outputs[4973] = (inputs[817]) & ~(inputs[971]);
    assign layer0_outputs[4974] = (inputs[398]) & (inputs[775]);
    assign layer0_outputs[4975] = (inputs[370]) & ~(inputs[1014]);
    assign layer0_outputs[4976] = ~((inputs[891]) & (inputs[601]));
    assign layer0_outputs[4977] = ~(inputs[244]);
    assign layer0_outputs[4978] = (inputs[504]) | (inputs[599]);
    assign layer0_outputs[4979] = (inputs[378]) | (inputs[87]);
    assign layer0_outputs[4980] = inputs[231];
    assign layer0_outputs[4981] = (inputs[41]) | (inputs[336]);
    assign layer0_outputs[4982] = ~(inputs[149]) | (inputs[575]);
    assign layer0_outputs[4983] = inputs[764];
    assign layer0_outputs[4984] = ~((inputs[218]) | (inputs[587]));
    assign layer0_outputs[4985] = inputs[494];
    assign layer0_outputs[4986] = ~((inputs[692]) ^ (inputs[699]));
    assign layer0_outputs[4987] = ~(inputs[685]);
    assign layer0_outputs[4988] = (inputs[434]) & ~(inputs[503]);
    assign layer0_outputs[4989] = (inputs[531]) & (inputs[442]);
    assign layer0_outputs[4990] = ~((inputs[776]) | (inputs[49]));
    assign layer0_outputs[4991] = (inputs[561]) ^ (inputs[1000]);
    assign layer0_outputs[4992] = ~(inputs[142]);
    assign layer0_outputs[4993] = (inputs[41]) | (inputs[350]);
    assign layer0_outputs[4994] = (inputs[492]) | (inputs[349]);
    assign layer0_outputs[4995] = (inputs[906]) & (inputs[353]);
    assign layer0_outputs[4996] = ~((inputs[101]) ^ (inputs[101]));
    assign layer0_outputs[4997] = ~(inputs[435]) | (inputs[731]);
    assign layer0_outputs[4998] = ~(inputs[887]) | (inputs[382]);
    assign layer0_outputs[4999] = (inputs[853]) | (inputs[360]);
    assign layer0_outputs[5000] = (inputs[309]) ^ (inputs[629]);
    assign layer0_outputs[5001] = ~(inputs[299]) | (inputs[1011]);
    assign layer0_outputs[5002] = inputs[465];
    assign layer0_outputs[5003] = ~((inputs[53]) & (inputs[73]));
    assign layer0_outputs[5004] = (inputs[11]) | (inputs[917]);
    assign layer0_outputs[5005] = ~((inputs[132]) & (inputs[60]));
    assign layer0_outputs[5006] = inputs[616];
    assign layer0_outputs[5007] = ~((inputs[615]) ^ (inputs[286]));
    assign layer0_outputs[5008] = ~((inputs[891]) | (inputs[782]));
    assign layer0_outputs[5009] = (inputs[113]) ^ (inputs[151]);
    assign layer0_outputs[5010] = ~(inputs[510]) | (inputs[129]);
    assign layer0_outputs[5011] = inputs[652];
    assign layer0_outputs[5012] = (inputs[931]) & (inputs[548]);
    assign layer0_outputs[5013] = inputs[156];
    assign layer0_outputs[5014] = (inputs[387]) | (inputs[513]);
    assign layer0_outputs[5015] = ~(inputs[1020]);
    assign layer0_outputs[5016] = ~(inputs[824]);
    assign layer0_outputs[5017] = (inputs[927]) ^ (inputs[27]);
    assign layer0_outputs[5018] = ~(inputs[905]);
    assign layer0_outputs[5019] = ~(inputs[754]);
    assign layer0_outputs[5020] = ~((inputs[972]) ^ (inputs[256]));
    assign layer0_outputs[5021] = inputs[923];
    assign layer0_outputs[5022] = ~(inputs[808]);
    assign layer0_outputs[5023] = ~((inputs[74]) ^ (inputs[471]));
    assign layer0_outputs[5024] = ~(inputs[794]) | (inputs[882]);
    assign layer0_outputs[5025] = ~((inputs[996]) ^ (inputs[40]));
    assign layer0_outputs[5026] = (inputs[795]) | (inputs[821]);
    assign layer0_outputs[5027] = inputs[843];
    assign layer0_outputs[5028] = (inputs[410]) | (inputs[582]);
    assign layer0_outputs[5029] = ~((inputs[990]) ^ (inputs[371]));
    assign layer0_outputs[5030] = inputs[534];
    assign layer0_outputs[5031] = inputs[387];
    assign layer0_outputs[5032] = ~((inputs[34]) | (inputs[985]));
    assign layer0_outputs[5033] = (inputs[686]) & ~(inputs[933]);
    assign layer0_outputs[5034] = ~((inputs[816]) | (inputs[166]));
    assign layer0_outputs[5035] = ~((inputs[1006]) | (inputs[428]));
    assign layer0_outputs[5036] = (inputs[939]) & (inputs[66]);
    assign layer0_outputs[5037] = (inputs[345]) & ~(inputs[166]);
    assign layer0_outputs[5038] = (inputs[838]) & (inputs[838]);
    assign layer0_outputs[5039] = inputs[823];
    assign layer0_outputs[5040] = ~((inputs[468]) | (inputs[253]));
    assign layer0_outputs[5041] = (inputs[650]) & ~(inputs[264]);
    assign layer0_outputs[5042] = ~(inputs[105]) | (inputs[262]);
    assign layer0_outputs[5043] = ~(inputs[167]) | (inputs[126]);
    assign layer0_outputs[5044] = ~(inputs[118]);
    assign layer0_outputs[5045] = (inputs[1016]) | (inputs[840]);
    assign layer0_outputs[5046] = (inputs[519]) & ~(inputs[1008]);
    assign layer0_outputs[5047] = ~((inputs[101]) | (inputs[652]));
    assign layer0_outputs[5048] = ~((inputs[109]) | (inputs[652]));
    assign layer0_outputs[5049] = ~(inputs[777]);
    assign layer0_outputs[5050] = inputs[557];
    assign layer0_outputs[5051] = ~((inputs[826]) | (inputs[458]));
    assign layer0_outputs[5052] = (inputs[993]) | (inputs[624]);
    assign layer0_outputs[5053] = (inputs[178]) | (inputs[865]);
    assign layer0_outputs[5054] = ~((inputs[386]) | (inputs[549]));
    assign layer0_outputs[5055] = ~((inputs[261]) | (inputs[548]));
    assign layer0_outputs[5056] = inputs[749];
    assign layer0_outputs[5057] = ~(inputs[659]) | (inputs[354]);
    assign layer0_outputs[5058] = (inputs[618]) & ~(inputs[910]);
    assign layer0_outputs[5059] = inputs[238];
    assign layer0_outputs[5060] = 1'b1;
    assign layer0_outputs[5061] = (inputs[938]) | (inputs[785]);
    assign layer0_outputs[5062] = ~((inputs[774]) ^ (inputs[165]));
    assign layer0_outputs[5063] = ~(inputs[189]) | (inputs[669]);
    assign layer0_outputs[5064] = ~(inputs[636]) | (inputs[7]);
    assign layer0_outputs[5065] = inputs[348];
    assign layer0_outputs[5066] = inputs[273];
    assign layer0_outputs[5067] = inputs[995];
    assign layer0_outputs[5068] = inputs[722];
    assign layer0_outputs[5069] = (inputs[497]) & ~(inputs[297]);
    assign layer0_outputs[5070] = ~(inputs[442]);
    assign layer0_outputs[5071] = ~(inputs[302]) | (inputs[1019]);
    assign layer0_outputs[5072] = ~((inputs[837]) ^ (inputs[60]));
    assign layer0_outputs[5073] = inputs[788];
    assign layer0_outputs[5074] = ~(inputs[464]) | (inputs[21]);
    assign layer0_outputs[5075] = ~((inputs[723]) | (inputs[772]));
    assign layer0_outputs[5076] = ~((inputs[56]) ^ (inputs[767]));
    assign layer0_outputs[5077] = ~(inputs[833]) | (inputs[389]);
    assign layer0_outputs[5078] = ~((inputs[418]) | (inputs[375]));
    assign layer0_outputs[5079] = ~((inputs[127]) | (inputs[321]));
    assign layer0_outputs[5080] = ~(inputs[709]);
    assign layer0_outputs[5081] = (inputs[262]) | (inputs[769]);
    assign layer0_outputs[5082] = (inputs[328]) & (inputs[373]);
    assign layer0_outputs[5083] = 1'b1;
    assign layer0_outputs[5084] = ~((inputs[196]) | (inputs[548]));
    assign layer0_outputs[5085] = ~((inputs[874]) ^ (inputs[996]));
    assign layer0_outputs[5086] = (inputs[304]) & ~(inputs[216]);
    assign layer0_outputs[5087] = (inputs[597]) ^ (inputs[786]);
    assign layer0_outputs[5088] = (inputs[292]) ^ (inputs[22]);
    assign layer0_outputs[5089] = ~(inputs[725]) | (inputs[189]);
    assign layer0_outputs[5090] = (inputs[721]) ^ (inputs[234]);
    assign layer0_outputs[5091] = (inputs[195]) | (inputs[858]);
    assign layer0_outputs[5092] = (inputs[867]) & ~(inputs[318]);
    assign layer0_outputs[5093] = ~((inputs[117]) ^ (inputs[532]));
    assign layer0_outputs[5094] = ~(inputs[948]);
    assign layer0_outputs[5095] = ~(inputs[243]) | (inputs[927]);
    assign layer0_outputs[5096] = ~(inputs[622]) | (inputs[772]);
    assign layer0_outputs[5097] = ~((inputs[14]) & (inputs[927]));
    assign layer0_outputs[5098] = (inputs[304]) & ~(inputs[30]);
    assign layer0_outputs[5099] = (inputs[275]) & ~(inputs[281]);
    assign layer0_outputs[5100] = ~(inputs[688]) | (inputs[608]);
    assign layer0_outputs[5101] = inputs[374];
    assign layer0_outputs[5102] = ~(inputs[259]);
    assign layer0_outputs[5103] = ~(inputs[961]);
    assign layer0_outputs[5104] = ~(inputs[505]);
    assign layer0_outputs[5105] = ~((inputs[316]) ^ (inputs[918]));
    assign layer0_outputs[5106] = ~(inputs[866]);
    assign layer0_outputs[5107] = (inputs[4]) ^ (inputs[790]);
    assign layer0_outputs[5108] = inputs[949];
    assign layer0_outputs[5109] = ~((inputs[991]) & (inputs[1019]));
    assign layer0_outputs[5110] = inputs[772];
    assign layer0_outputs[5111] = (inputs[12]) & ~(inputs[415]);
    assign layer0_outputs[5112] = ~(inputs[991]) | (inputs[228]);
    assign layer0_outputs[5113] = (inputs[765]) ^ (inputs[418]);
    assign layer0_outputs[5114] = ~(inputs[358]) | (inputs[761]);
    assign layer0_outputs[5115] = (inputs[915]) ^ (inputs[711]);
    assign layer0_outputs[5116] = ~((inputs[215]) ^ (inputs[453]));
    assign layer0_outputs[5117] = inputs[231];
    assign layer0_outputs[5118] = (inputs[430]) ^ (inputs[358]);
    assign layer0_outputs[5119] = inputs[99];
    assign layer0_outputs[5120] = ~(inputs[465]) | (inputs[585]);
    assign layer0_outputs[5121] = ~(inputs[372]);
    assign layer0_outputs[5122] = (inputs[207]) ^ (inputs[222]);
    assign layer0_outputs[5123] = inputs[876];
    assign layer0_outputs[5124] = 1'b0;
    assign layer0_outputs[5125] = ~(inputs[459]);
    assign layer0_outputs[5126] = (inputs[513]) & ~(inputs[321]);
    assign layer0_outputs[5127] = (inputs[17]) ^ (inputs[46]);
    assign layer0_outputs[5128] = ~(inputs[136]) | (inputs[260]);
    assign layer0_outputs[5129] = (inputs[366]) & ~(inputs[921]);
    assign layer0_outputs[5130] = (inputs[393]) & ~(inputs[587]);
    assign layer0_outputs[5131] = inputs[76];
    assign layer0_outputs[5132] = ~(inputs[539]) | (inputs[64]);
    assign layer0_outputs[5133] = inputs[432];
    assign layer0_outputs[5134] = ~((inputs[455]) | (inputs[820]));
    assign layer0_outputs[5135] = ~((inputs[317]) | (inputs[744]));
    assign layer0_outputs[5136] = inputs[224];
    assign layer0_outputs[5137] = ~(inputs[87]);
    assign layer0_outputs[5138] = ~((inputs[380]) ^ (inputs[748]));
    assign layer0_outputs[5139] = ~((inputs[725]) | (inputs[108]));
    assign layer0_outputs[5140] = ~((inputs[691]) ^ (inputs[51]));
    assign layer0_outputs[5141] = (inputs[760]) | (inputs[696]);
    assign layer0_outputs[5142] = ~(inputs[831]) | (inputs[1001]);
    assign layer0_outputs[5143] = 1'b1;
    assign layer0_outputs[5144] = ~((inputs[779]) | (inputs[726]));
    assign layer0_outputs[5145] = 1'b0;
    assign layer0_outputs[5146] = ~((inputs[644]) | (inputs[148]));
    assign layer0_outputs[5147] = ~((inputs[812]) | (inputs[145]));
    assign layer0_outputs[5148] = ~((inputs[903]) | (inputs[578]));
    assign layer0_outputs[5149] = ~(inputs[684]);
    assign layer0_outputs[5150] = ~(inputs[90]) | (inputs[459]);
    assign layer0_outputs[5151] = ~(inputs[180]);
    assign layer0_outputs[5152] = ~((inputs[233]) | (inputs[110]));
    assign layer0_outputs[5153] = (inputs[438]) | (inputs[639]);
    assign layer0_outputs[5154] = (inputs[290]) ^ (inputs[994]);
    assign layer0_outputs[5155] = inputs[170];
    assign layer0_outputs[5156] = (inputs[961]) & ~(inputs[136]);
    assign layer0_outputs[5157] = ~((inputs[861]) ^ (inputs[777]));
    assign layer0_outputs[5158] = ~(inputs[525]) | (inputs[144]);
    assign layer0_outputs[5159] = ~((inputs[455]) & (inputs[161]));
    assign layer0_outputs[5160] = (inputs[316]) & ~(inputs[290]);
    assign layer0_outputs[5161] = (inputs[619]) | (inputs[760]);
    assign layer0_outputs[5162] = ~(inputs[64]);
    assign layer0_outputs[5163] = (inputs[1018]) & ~(inputs[493]);
    assign layer0_outputs[5164] = ~(inputs[406]);
    assign layer0_outputs[5165] = inputs[553];
    assign layer0_outputs[5166] = ~((inputs[281]) ^ (inputs[41]));
    assign layer0_outputs[5167] = ~(inputs[467]);
    assign layer0_outputs[5168] = ~((inputs[134]) | (inputs[381]));
    assign layer0_outputs[5169] = (inputs[11]) | (inputs[876]);
    assign layer0_outputs[5170] = (inputs[504]) | (inputs[144]);
    assign layer0_outputs[5171] = ~(inputs[554]) | (inputs[709]);
    assign layer0_outputs[5172] = (inputs[727]) | (inputs[888]);
    assign layer0_outputs[5173] = ~((inputs[783]) & (inputs[811]));
    assign layer0_outputs[5174] = (inputs[154]) & ~(inputs[265]);
    assign layer0_outputs[5175] = ~(inputs[945]) | (inputs[854]);
    assign layer0_outputs[5176] = ~((inputs[872]) | (inputs[601]));
    assign layer0_outputs[5177] = 1'b0;
    assign layer0_outputs[5178] = ~((inputs[407]) | (inputs[832]));
    assign layer0_outputs[5179] = ~((inputs[277]) ^ (inputs[599]));
    assign layer0_outputs[5180] = inputs[191];
    assign layer0_outputs[5181] = ~(inputs[598]) | (inputs[27]);
    assign layer0_outputs[5182] = ~((inputs[460]) | (inputs[639]));
    assign layer0_outputs[5183] = ~((inputs[216]) | (inputs[785]));
    assign layer0_outputs[5184] = ~(inputs[248]);
    assign layer0_outputs[5185] = (inputs[873]) & (inputs[76]);
    assign layer0_outputs[5186] = inputs[428];
    assign layer0_outputs[5187] = ~((inputs[276]) | (inputs[833]));
    assign layer0_outputs[5188] = (inputs[314]) | (inputs[588]);
    assign layer0_outputs[5189] = ~(inputs[246]) | (inputs[153]);
    assign layer0_outputs[5190] = (inputs[513]) ^ (inputs[237]);
    assign layer0_outputs[5191] = 1'b0;
    assign layer0_outputs[5192] = ~((inputs[533]) | (inputs[182]));
    assign layer0_outputs[5193] = ~((inputs[134]) & (inputs[105]));
    assign layer0_outputs[5194] = ~(inputs[837]);
    assign layer0_outputs[5195] = ~(inputs[436]) | (inputs[130]);
    assign layer0_outputs[5196] = inputs[553];
    assign layer0_outputs[5197] = (inputs[679]) & (inputs[588]);
    assign layer0_outputs[5198] = ~((inputs[322]) | (inputs[213]));
    assign layer0_outputs[5199] = (inputs[310]) ^ (inputs[1019]);
    assign layer0_outputs[5200] = ~((inputs[674]) | (inputs[471]));
    assign layer0_outputs[5201] = ~((inputs[1017]) | (inputs[803]));
    assign layer0_outputs[5202] = inputs[258];
    assign layer0_outputs[5203] = inputs[508];
    assign layer0_outputs[5204] = ~(inputs[115]);
    assign layer0_outputs[5205] = inputs[720];
    assign layer0_outputs[5206] = (inputs[282]) ^ (inputs[451]);
    assign layer0_outputs[5207] = (inputs[529]) & ~(inputs[230]);
    assign layer0_outputs[5208] = (inputs[890]) | (inputs[948]);
    assign layer0_outputs[5209] = (inputs[310]) & ~(inputs[190]);
    assign layer0_outputs[5210] = ~(inputs[790]) | (inputs[666]);
    assign layer0_outputs[5211] = inputs[809];
    assign layer0_outputs[5212] = ~((inputs[331]) | (inputs[650]));
    assign layer0_outputs[5213] = (inputs[171]) & (inputs[224]);
    assign layer0_outputs[5214] = inputs[111];
    assign layer0_outputs[5215] = ~(inputs[492]);
    assign layer0_outputs[5216] = ~(inputs[257]);
    assign layer0_outputs[5217] = ~((inputs[986]) | (inputs[812]));
    assign layer0_outputs[5218] = (inputs[88]) | (inputs[1014]);
    assign layer0_outputs[5219] = (inputs[927]) & ~(inputs[416]);
    assign layer0_outputs[5220] = 1'b0;
    assign layer0_outputs[5221] = (inputs[983]) ^ (inputs[529]);
    assign layer0_outputs[5222] = ~((inputs[208]) ^ (inputs[121]));
    assign layer0_outputs[5223] = ~(inputs[622]);
    assign layer0_outputs[5224] = (inputs[715]) | (inputs[681]);
    assign layer0_outputs[5225] = inputs[682];
    assign layer0_outputs[5226] = inputs[334];
    assign layer0_outputs[5227] = ~((inputs[199]) | (inputs[598]));
    assign layer0_outputs[5228] = inputs[810];
    assign layer0_outputs[5229] = ~((inputs[439]) ^ (inputs[856]));
    assign layer0_outputs[5230] = ~(inputs[866]);
    assign layer0_outputs[5231] = ~(inputs[260]);
    assign layer0_outputs[5232] = ~(inputs[791]) | (inputs[572]);
    assign layer0_outputs[5233] = (inputs[175]) | (inputs[417]);
    assign layer0_outputs[5234] = ~(inputs[562]) | (inputs[246]);
    assign layer0_outputs[5235] = ~((inputs[899]) & (inputs[27]));
    assign layer0_outputs[5236] = (inputs[420]) ^ (inputs[684]);
    assign layer0_outputs[5237] = ~(inputs[621]) | (inputs[1020]);
    assign layer0_outputs[5238] = inputs[846];
    assign layer0_outputs[5239] = ~(inputs[567]);
    assign layer0_outputs[5240] = (inputs[1022]) & ~(inputs[808]);
    assign layer0_outputs[5241] = (inputs[399]) | (inputs[129]);
    assign layer0_outputs[5242] = (inputs[236]) & ~(inputs[472]);
    assign layer0_outputs[5243] = ~((inputs[945]) | (inputs[157]));
    assign layer0_outputs[5244] = ~(inputs[42]) | (inputs[128]);
    assign layer0_outputs[5245] = ~(inputs[310]) | (inputs[862]);
    assign layer0_outputs[5246] = (inputs[874]) | (inputs[390]);
    assign layer0_outputs[5247] = ~(inputs[623]);
    assign layer0_outputs[5248] = ~(inputs[416]);
    assign layer0_outputs[5249] = (inputs[759]) & ~(inputs[911]);
    assign layer0_outputs[5250] = (inputs[750]) & ~(inputs[873]);
    assign layer0_outputs[5251] = ~((inputs[644]) | (inputs[369]));
    assign layer0_outputs[5252] = inputs[803];
    assign layer0_outputs[5253] = ~((inputs[931]) | (inputs[662]));
    assign layer0_outputs[5254] = (inputs[1004]) & ~(inputs[326]);
    assign layer0_outputs[5255] = ~(inputs[29]);
    assign layer0_outputs[5256] = (inputs[394]) & ~(inputs[215]);
    assign layer0_outputs[5257] = ~(inputs[276]);
    assign layer0_outputs[5258] = inputs[1];
    assign layer0_outputs[5259] = ~((inputs[371]) ^ (inputs[77]));
    assign layer0_outputs[5260] = ~(inputs[964]);
    assign layer0_outputs[5261] = (inputs[526]) & ~(inputs[731]);
    assign layer0_outputs[5262] = (inputs[246]) ^ (inputs[819]);
    assign layer0_outputs[5263] = inputs[240];
    assign layer0_outputs[5264] = (inputs[947]) ^ (inputs[602]);
    assign layer0_outputs[5265] = (inputs[509]) ^ (inputs[249]);
    assign layer0_outputs[5266] = inputs[308];
    assign layer0_outputs[5267] = ~(inputs[284]) | (inputs[447]);
    assign layer0_outputs[5268] = (inputs[799]) & (inputs[604]);
    assign layer0_outputs[5269] = (inputs[381]) ^ (inputs[55]);
    assign layer0_outputs[5270] = (inputs[808]) & ~(inputs[799]);
    assign layer0_outputs[5271] = ~((inputs[546]) ^ (inputs[520]));
    assign layer0_outputs[5272] = (inputs[804]) & ~(inputs[354]);
    assign layer0_outputs[5273] = inputs[589];
    assign layer0_outputs[5274] = ~(inputs[499]);
    assign layer0_outputs[5275] = ~(inputs[457]);
    assign layer0_outputs[5276] = (inputs[477]) | (inputs[872]);
    assign layer0_outputs[5277] = inputs[404];
    assign layer0_outputs[5278] = ~((inputs[458]) & (inputs[663]));
    assign layer0_outputs[5279] = 1'b0;
    assign layer0_outputs[5280] = ~(inputs[413]);
    assign layer0_outputs[5281] = ~((inputs[856]) | (inputs[791]));
    assign layer0_outputs[5282] = ~((inputs[886]) | (inputs[801]));
    assign layer0_outputs[5283] = ~(inputs[970]) | (inputs[297]);
    assign layer0_outputs[5284] = (inputs[46]) ^ (inputs[480]);
    assign layer0_outputs[5285] = ~(inputs[40]) | (inputs[594]);
    assign layer0_outputs[5286] = (inputs[215]) ^ (inputs[180]);
    assign layer0_outputs[5287] = ~(inputs[558]);
    assign layer0_outputs[5288] = ~(inputs[365]);
    assign layer0_outputs[5289] = inputs[171];
    assign layer0_outputs[5290] = 1'b1;
    assign layer0_outputs[5291] = ~((inputs[183]) | (inputs[346]));
    assign layer0_outputs[5292] = (inputs[672]) & ~(inputs[772]);
    assign layer0_outputs[5293] = ~((inputs[647]) ^ (inputs[964]));
    assign layer0_outputs[5294] = (inputs[555]) | (inputs[289]);
    assign layer0_outputs[5295] = ~(inputs[32]);
    assign layer0_outputs[5296] = ~(inputs[742]) | (inputs[353]);
    assign layer0_outputs[5297] = ~(inputs[889]) | (inputs[287]);
    assign layer0_outputs[5298] = (inputs[647]) | (inputs[859]);
    assign layer0_outputs[5299] = (inputs[950]) | (inputs[227]);
    assign layer0_outputs[5300] = ~((inputs[402]) | (inputs[1007]));
    assign layer0_outputs[5301] = ~(inputs[596]) | (inputs[110]);
    assign layer0_outputs[5302] = ~(inputs[582]) | (inputs[598]);
    assign layer0_outputs[5303] = ~(inputs[810]) | (inputs[801]);
    assign layer0_outputs[5304] = (inputs[522]) | (inputs[421]);
    assign layer0_outputs[5305] = inputs[269];
    assign layer0_outputs[5306] = inputs[202];
    assign layer0_outputs[5307] = (inputs[92]) ^ (inputs[460]);
    assign layer0_outputs[5308] = ~((inputs[801]) ^ (inputs[608]));
    assign layer0_outputs[5309] = (inputs[474]) | (inputs[291]);
    assign layer0_outputs[5310] = ~((inputs[997]) & (inputs[225]));
    assign layer0_outputs[5311] = (inputs[737]) ^ (inputs[369]);
    assign layer0_outputs[5312] = ~((inputs[581]) | (inputs[196]));
    assign layer0_outputs[5313] = (inputs[276]) ^ (inputs[196]);
    assign layer0_outputs[5314] = (inputs[58]) | (inputs[277]);
    assign layer0_outputs[5315] = ~(inputs[566]);
    assign layer0_outputs[5316] = (inputs[303]) | (inputs[879]);
    assign layer0_outputs[5317] = (inputs[107]) & (inputs[161]);
    assign layer0_outputs[5318] = ~(inputs[337]);
    assign layer0_outputs[5319] = 1'b1;
    assign layer0_outputs[5320] = (inputs[637]) & (inputs[157]);
    assign layer0_outputs[5321] = ~((inputs[156]) ^ (inputs[438]));
    assign layer0_outputs[5322] = ~(inputs[22]);
    assign layer0_outputs[5323] = (inputs[356]) & ~(inputs[130]);
    assign layer0_outputs[5324] = ~((inputs[636]) | (inputs[12]));
    assign layer0_outputs[5325] = 1'b1;
    assign layer0_outputs[5326] = (inputs[481]) ^ (inputs[273]);
    assign layer0_outputs[5327] = ~(inputs[644]) | (inputs[761]);
    assign layer0_outputs[5328] = (inputs[946]) | (inputs[971]);
    assign layer0_outputs[5329] = ~(inputs[81]);
    assign layer0_outputs[5330] = (inputs[624]) | (inputs[167]);
    assign layer0_outputs[5331] = inputs[241];
    assign layer0_outputs[5332] = inputs[146];
    assign layer0_outputs[5333] = ~(inputs[619]);
    assign layer0_outputs[5334] = ~(inputs[93]);
    assign layer0_outputs[5335] = (inputs[748]) | (inputs[365]);
    assign layer0_outputs[5336] = (inputs[277]) & ~(inputs[732]);
    assign layer0_outputs[5337] = ~(inputs[424]) | (inputs[1014]);
    assign layer0_outputs[5338] = (inputs[846]) & ~(inputs[953]);
    assign layer0_outputs[5339] = inputs[780];
    assign layer0_outputs[5340] = (inputs[282]) & ~(inputs[60]);
    assign layer0_outputs[5341] = ~((inputs[477]) | (inputs[177]));
    assign layer0_outputs[5342] = ~((inputs[103]) ^ (inputs[781]));
    assign layer0_outputs[5343] = (inputs[409]) & ~(inputs[224]);
    assign layer0_outputs[5344] = (inputs[215]) & ~(inputs[978]);
    assign layer0_outputs[5345] = inputs[649];
    assign layer0_outputs[5346] = ~(inputs[504]) | (inputs[44]);
    assign layer0_outputs[5347] = ~(inputs[966]);
    assign layer0_outputs[5348] = (inputs[631]) | (inputs[679]);
    assign layer0_outputs[5349] = (inputs[68]) | (inputs[460]);
    assign layer0_outputs[5350] = (inputs[689]) & ~(inputs[913]);
    assign layer0_outputs[5351] = 1'b1;
    assign layer0_outputs[5352] = ~((inputs[779]) | (inputs[632]));
    assign layer0_outputs[5353] = (inputs[405]) & ~(inputs[710]);
    assign layer0_outputs[5354] = (inputs[822]) & ~(inputs[350]);
    assign layer0_outputs[5355] = ~((inputs[541]) & (inputs[481]));
    assign layer0_outputs[5356] = ~(inputs[687]);
    assign layer0_outputs[5357] = (inputs[838]) | (inputs[387]);
    assign layer0_outputs[5358] = ~(inputs[622]) | (inputs[772]);
    assign layer0_outputs[5359] = ~(inputs[806]) | (inputs[257]);
    assign layer0_outputs[5360] = (inputs[673]) | (inputs[363]);
    assign layer0_outputs[5361] = ~((inputs[321]) | (inputs[179]));
    assign layer0_outputs[5362] = ~(inputs[112]);
    assign layer0_outputs[5363] = (inputs[782]) & ~(inputs[33]);
    assign layer0_outputs[5364] = (inputs[317]) ^ (inputs[474]);
    assign layer0_outputs[5365] = inputs[698];
    assign layer0_outputs[5366] = (inputs[101]) ^ (inputs[810]);
    assign layer0_outputs[5367] = inputs[587];
    assign layer0_outputs[5368] = 1'b0;
    assign layer0_outputs[5369] = (inputs[331]) | (inputs[350]);
    assign layer0_outputs[5370] = (inputs[579]) | (inputs[834]);
    assign layer0_outputs[5371] = inputs[637];
    assign layer0_outputs[5372] = ~((inputs[1009]) | (inputs[723]));
    assign layer0_outputs[5373] = 1'b1;
    assign layer0_outputs[5374] = inputs[44];
    assign layer0_outputs[5375] = ~(inputs[835]);
    assign layer0_outputs[5376] = ~(inputs[420]);
    assign layer0_outputs[5377] = ~(inputs[435]);
    assign layer0_outputs[5378] = 1'b0;
    assign layer0_outputs[5379] = ~(inputs[427]) | (inputs[805]);
    assign layer0_outputs[5380] = ~((inputs[794]) ^ (inputs[182]));
    assign layer0_outputs[5381] = inputs[319];
    assign layer0_outputs[5382] = ~((inputs[849]) | (inputs[19]));
    assign layer0_outputs[5383] = (inputs[784]) & ~(inputs[905]);
    assign layer0_outputs[5384] = ~((inputs[760]) ^ (inputs[809]));
    assign layer0_outputs[5385] = ~(inputs[402]);
    assign layer0_outputs[5386] = inputs[487];
    assign layer0_outputs[5387] = ~((inputs[675]) ^ (inputs[631]));
    assign layer0_outputs[5388] = ~((inputs[8]) ^ (inputs[106]));
    assign layer0_outputs[5389] = (inputs[898]) ^ (inputs[519]);
    assign layer0_outputs[5390] = (inputs[949]) & (inputs[271]);
    assign layer0_outputs[5391] = (inputs[227]) & (inputs[93]);
    assign layer0_outputs[5392] = (inputs[155]) & ~(inputs[227]);
    assign layer0_outputs[5393] = (inputs[132]) ^ (inputs[479]);
    assign layer0_outputs[5394] = ~(inputs[179]) | (inputs[984]);
    assign layer0_outputs[5395] = 1'b1;
    assign layer0_outputs[5396] = ~(inputs[703]) | (inputs[39]);
    assign layer0_outputs[5397] = (inputs[183]) | (inputs[600]);
    assign layer0_outputs[5398] = (inputs[811]) & ~(inputs[655]);
    assign layer0_outputs[5399] = ~(inputs[916]);
    assign layer0_outputs[5400] = inputs[123];
    assign layer0_outputs[5401] = ~((inputs[142]) ^ (inputs[676]));
    assign layer0_outputs[5402] = ~(inputs[518]);
    assign layer0_outputs[5403] = (inputs[599]) ^ (inputs[850]);
    assign layer0_outputs[5404] = ~(inputs[728]);
    assign layer0_outputs[5405] = ~((inputs[528]) ^ (inputs[633]));
    assign layer0_outputs[5406] = (inputs[42]) | (inputs[490]);
    assign layer0_outputs[5407] = (inputs[955]) & ~(inputs[350]);
    assign layer0_outputs[5408] = (inputs[443]) ^ (inputs[31]);
    assign layer0_outputs[5409] = ~((inputs[269]) | (inputs[125]));
    assign layer0_outputs[5410] = ~((inputs[559]) ^ (inputs[5]));
    assign layer0_outputs[5411] = (inputs[684]) ^ (inputs[744]);
    assign layer0_outputs[5412] = ~((inputs[297]) ^ (inputs[828]));
    assign layer0_outputs[5413] = ~((inputs[238]) | (inputs[910]));
    assign layer0_outputs[5414] = (inputs[691]) & ~(inputs[735]);
    assign layer0_outputs[5415] = (inputs[669]) ^ (inputs[649]);
    assign layer0_outputs[5416] = ~((inputs[980]) | (inputs[656]));
    assign layer0_outputs[5417] = ~((inputs[10]) ^ (inputs[661]));
    assign layer0_outputs[5418] = ~(inputs[427]);
    assign layer0_outputs[5419] = ~((inputs[605]) ^ (inputs[826]));
    assign layer0_outputs[5420] = (inputs[809]) | (inputs[417]);
    assign layer0_outputs[5421] = ~((inputs[798]) | (inputs[87]));
    assign layer0_outputs[5422] = (inputs[628]) ^ (inputs[999]);
    assign layer0_outputs[5423] = (inputs[421]) & ~(inputs[209]);
    assign layer0_outputs[5424] = ~((inputs[999]) | (inputs[275]));
    assign layer0_outputs[5425] = (inputs[1002]) & ~(inputs[28]);
    assign layer0_outputs[5426] = (inputs[578]) & ~(inputs[167]);
    assign layer0_outputs[5427] = ~(inputs[182]);
    assign layer0_outputs[5428] = ~((inputs[48]) ^ (inputs[582]));
    assign layer0_outputs[5429] = ~((inputs[939]) | (inputs[21]));
    assign layer0_outputs[5430] = ~(inputs[384]);
    assign layer0_outputs[5431] = (inputs[844]) | (inputs[68]);
    assign layer0_outputs[5432] = ~((inputs[133]) ^ (inputs[308]));
    assign layer0_outputs[5433] = ~((inputs[169]) | (inputs[269]));
    assign layer0_outputs[5434] = ~(inputs[466]);
    assign layer0_outputs[5435] = ~(inputs[550]);
    assign layer0_outputs[5436] = ~(inputs[424]) | (inputs[114]);
    assign layer0_outputs[5437] = ~(inputs[527]) | (inputs[428]);
    assign layer0_outputs[5438] = ~(inputs[399]) | (inputs[528]);
    assign layer0_outputs[5439] = ~(inputs[440]);
    assign layer0_outputs[5440] = (inputs[366]) | (inputs[904]);
    assign layer0_outputs[5441] = (inputs[1014]) | (inputs[589]);
    assign layer0_outputs[5442] = (inputs[357]) | (inputs[469]);
    assign layer0_outputs[5443] = ~(inputs[433]) | (inputs[64]);
    assign layer0_outputs[5444] = (inputs[336]) | (inputs[948]);
    assign layer0_outputs[5445] = ~((inputs[147]) | (inputs[632]));
    assign layer0_outputs[5446] = (inputs[508]) | (inputs[730]);
    assign layer0_outputs[5447] = inputs[228];
    assign layer0_outputs[5448] = inputs[424];
    assign layer0_outputs[5449] = ~((inputs[668]) | (inputs[937]));
    assign layer0_outputs[5450] = (inputs[427]) & (inputs[531]);
    assign layer0_outputs[5451] = ~(inputs[49]);
    assign layer0_outputs[5452] = (inputs[860]) & ~(inputs[707]);
    assign layer0_outputs[5453] = (inputs[143]) & ~(inputs[800]);
    assign layer0_outputs[5454] = (inputs[889]) | (inputs[512]);
    assign layer0_outputs[5455] = ~(inputs[501]) | (inputs[736]);
    assign layer0_outputs[5456] = inputs[179];
    assign layer0_outputs[5457] = 1'b0;
    assign layer0_outputs[5458] = (inputs[441]) & ~(inputs[130]);
    assign layer0_outputs[5459] = (inputs[160]) ^ (inputs[242]);
    assign layer0_outputs[5460] = inputs[637];
    assign layer0_outputs[5461] = ~((inputs[976]) | (inputs[96]));
    assign layer0_outputs[5462] = inputs[413];
    assign layer0_outputs[5463] = inputs[809];
    assign layer0_outputs[5464] = ~(inputs[511]);
    assign layer0_outputs[5465] = ~((inputs[1014]) ^ (inputs[797]));
    assign layer0_outputs[5466] = 1'b0;
    assign layer0_outputs[5467] = ~(inputs[402]);
    assign layer0_outputs[5468] = (inputs[105]) ^ (inputs[594]);
    assign layer0_outputs[5469] = ~((inputs[875]) | (inputs[310]));
    assign layer0_outputs[5470] = ~(inputs[918]) | (inputs[71]);
    assign layer0_outputs[5471] = ~((inputs[631]) ^ (inputs[350]));
    assign layer0_outputs[5472] = ~(inputs[851]) | (inputs[42]);
    assign layer0_outputs[5473] = (inputs[212]) | (inputs[458]);
    assign layer0_outputs[5474] = inputs[334];
    assign layer0_outputs[5475] = inputs[85];
    assign layer0_outputs[5476] = (inputs[128]) ^ (inputs[942]);
    assign layer0_outputs[5477] = ~((inputs[929]) & (inputs[924]));
    assign layer0_outputs[5478] = ~((inputs[994]) ^ (inputs[877]));
    assign layer0_outputs[5479] = ~(inputs[588]);
    assign layer0_outputs[5480] = ~(inputs[406]);
    assign layer0_outputs[5481] = ~((inputs[545]) ^ (inputs[13]));
    assign layer0_outputs[5482] = inputs[546];
    assign layer0_outputs[5483] = inputs[434];
    assign layer0_outputs[5484] = ~((inputs[894]) | (inputs[481]));
    assign layer0_outputs[5485] = (inputs[183]) | (inputs[593]);
    assign layer0_outputs[5486] = ~(inputs[600]);
    assign layer0_outputs[5487] = ~((inputs[352]) ^ (inputs[263]));
    assign layer0_outputs[5488] = ~(inputs[432]) | (inputs[140]);
    assign layer0_outputs[5489] = inputs[296];
    assign layer0_outputs[5490] = (inputs[856]) | (inputs[413]);
    assign layer0_outputs[5491] = (inputs[541]) & ~(inputs[133]);
    assign layer0_outputs[5492] = ~((inputs[597]) ^ (inputs[456]));
    assign layer0_outputs[5493] = 1'b0;
    assign layer0_outputs[5494] = ~(inputs[189]) | (inputs[43]);
    assign layer0_outputs[5495] = 1'b0;
    assign layer0_outputs[5496] = ~(inputs[510]);
    assign layer0_outputs[5497] = (inputs[870]) ^ (inputs[326]);
    assign layer0_outputs[5498] = 1'b1;
    assign layer0_outputs[5499] = 1'b1;
    assign layer0_outputs[5500] = ~((inputs[939]) | (inputs[307]));
    assign layer0_outputs[5501] = ~(inputs[398]);
    assign layer0_outputs[5502] = ~(inputs[616]) | (inputs[881]);
    assign layer0_outputs[5503] = (inputs[273]) & ~(inputs[91]);
    assign layer0_outputs[5504] = inputs[817];
    assign layer0_outputs[5505] = ~((inputs[810]) & (inputs[592]));
    assign layer0_outputs[5506] = (inputs[90]) ^ (inputs[783]);
    assign layer0_outputs[5507] = ~(inputs[412]);
    assign layer0_outputs[5508] = (inputs[977]) ^ (inputs[953]);
    assign layer0_outputs[5509] = inputs[748];
    assign layer0_outputs[5510] = ~((inputs[866]) & (inputs[37]));
    assign layer0_outputs[5511] = (inputs[454]) & ~(inputs[84]);
    assign layer0_outputs[5512] = (inputs[903]) | (inputs[120]);
    assign layer0_outputs[5513] = ~(inputs[290]);
    assign layer0_outputs[5514] = ~(inputs[747]) | (inputs[919]);
    assign layer0_outputs[5515] = ~((inputs[307]) | (inputs[660]));
    assign layer0_outputs[5516] = (inputs[75]) & ~(inputs[15]);
    assign layer0_outputs[5517] = inputs[13];
    assign layer0_outputs[5518] = (inputs[338]) & ~(inputs[916]);
    assign layer0_outputs[5519] = ~(inputs[493]);
    assign layer0_outputs[5520] = ~((inputs[706]) | (inputs[521]));
    assign layer0_outputs[5521] = (inputs[835]) & ~(inputs[121]);
    assign layer0_outputs[5522] = ~(inputs[265]);
    assign layer0_outputs[5523] = ~(inputs[607]) | (inputs[24]);
    assign layer0_outputs[5524] = inputs[432];
    assign layer0_outputs[5525] = inputs[553];
    assign layer0_outputs[5526] = inputs[129];
    assign layer0_outputs[5527] = inputs[20];
    assign layer0_outputs[5528] = ~((inputs[188]) ^ (inputs[154]));
    assign layer0_outputs[5529] = ~((inputs[885]) | (inputs[249]));
    assign layer0_outputs[5530] = inputs[107];
    assign layer0_outputs[5531] = (inputs[574]) ^ (inputs[655]);
    assign layer0_outputs[5532] = (inputs[585]) | (inputs[827]);
    assign layer0_outputs[5533] = inputs[217];
    assign layer0_outputs[5534] = (inputs[127]) ^ (inputs[493]);
    assign layer0_outputs[5535] = (inputs[713]) ^ (inputs[917]);
    assign layer0_outputs[5536] = (inputs[790]) | (inputs[223]);
    assign layer0_outputs[5537] = ~((inputs[261]) ^ (inputs[636]));
    assign layer0_outputs[5538] = ~(inputs[519]);
    assign layer0_outputs[5539] = 1'b0;
    assign layer0_outputs[5540] = ~((inputs[248]) | (inputs[124]));
    assign layer0_outputs[5541] = ~((inputs[713]) & (inputs[562]));
    assign layer0_outputs[5542] = ~((inputs[946]) | (inputs[584]));
    assign layer0_outputs[5543] = inputs[534];
    assign layer0_outputs[5544] = inputs[620];
    assign layer0_outputs[5545] = 1'b0;
    assign layer0_outputs[5546] = ~(inputs[650]);
    assign layer0_outputs[5547] = inputs[528];
    assign layer0_outputs[5548] = inputs[713];
    assign layer0_outputs[5549] = (inputs[196]) & ~(inputs[474]);
    assign layer0_outputs[5550] = 1'b0;
    assign layer0_outputs[5551] = ~((inputs[229]) ^ (inputs[279]));
    assign layer0_outputs[5552] = (inputs[100]) | (inputs[490]);
    assign layer0_outputs[5553] = (inputs[683]) | (inputs[931]);
    assign layer0_outputs[5554] = ~((inputs[950]) | (inputs[665]));
    assign layer0_outputs[5555] = ~((inputs[539]) | (inputs[473]));
    assign layer0_outputs[5556] = (inputs[786]) & ~(inputs[39]);
    assign layer0_outputs[5557] = ~(inputs[125]) | (inputs[179]);
    assign layer0_outputs[5558] = ~((inputs[564]) ^ (inputs[334]));
    assign layer0_outputs[5559] = (inputs[754]) ^ (inputs[156]);
    assign layer0_outputs[5560] = ~(inputs[941]);
    assign layer0_outputs[5561] = ~((inputs[472]) ^ (inputs[769]));
    assign layer0_outputs[5562] = (inputs[241]) & ~(inputs[4]);
    assign layer0_outputs[5563] = (inputs[816]) | (inputs[690]);
    assign layer0_outputs[5564] = (inputs[462]) | (inputs[315]);
    assign layer0_outputs[5565] = ~(inputs[65]);
    assign layer0_outputs[5566] = ~((inputs[580]) ^ (inputs[305]));
    assign layer0_outputs[5567] = ~((inputs[22]) ^ (inputs[521]));
    assign layer0_outputs[5568] = inputs[197];
    assign layer0_outputs[5569] = inputs[159];
    assign layer0_outputs[5570] = ~(inputs[614]);
    assign layer0_outputs[5571] = inputs[537];
    assign layer0_outputs[5572] = ~((inputs[305]) | (inputs[635]));
    assign layer0_outputs[5573] = (inputs[649]) ^ (inputs[327]);
    assign layer0_outputs[5574] = (inputs[840]) & (inputs[535]);
    assign layer0_outputs[5575] = (inputs[884]) & ~(inputs[841]);
    assign layer0_outputs[5576] = 1'b0;
    assign layer0_outputs[5577] = (inputs[473]) ^ (inputs[30]);
    assign layer0_outputs[5578] = inputs[685];
    assign layer0_outputs[5579] = ~((inputs[271]) | (inputs[346]));
    assign layer0_outputs[5580] = ~((inputs[389]) ^ (inputs[84]));
    assign layer0_outputs[5581] = ~((inputs[91]) | (inputs[13]));
    assign layer0_outputs[5582] = (inputs[1000]) ^ (inputs[270]);
    assign layer0_outputs[5583] = inputs[555];
    assign layer0_outputs[5584] = (inputs[314]) & ~(inputs[383]);
    assign layer0_outputs[5585] = inputs[379];
    assign layer0_outputs[5586] = ~(inputs[949]);
    assign layer0_outputs[5587] = (inputs[659]) & ~(inputs[866]);
    assign layer0_outputs[5588] = (inputs[889]) ^ (inputs[74]);
    assign layer0_outputs[5589] = ~((inputs[667]) | (inputs[722]));
    assign layer0_outputs[5590] = inputs[721];
    assign layer0_outputs[5591] = inputs[585];
    assign layer0_outputs[5592] = (inputs[620]) & ~(inputs[100]);
    assign layer0_outputs[5593] = (inputs[176]) & ~(inputs[186]);
    assign layer0_outputs[5594] = (inputs[976]) | (inputs[812]);
    assign layer0_outputs[5595] = ~((inputs[462]) | (inputs[363]));
    assign layer0_outputs[5596] = ~((inputs[710]) | (inputs[179]));
    assign layer0_outputs[5597] = ~(inputs[561]) | (inputs[255]);
    assign layer0_outputs[5598] = ~(inputs[713]);
    assign layer0_outputs[5599] = ~(inputs[662]) | (inputs[201]);
    assign layer0_outputs[5600] = ~(inputs[457]);
    assign layer0_outputs[5601] = inputs[596];
    assign layer0_outputs[5602] = ~(inputs[347]);
    assign layer0_outputs[5603] = ~(inputs[634]) | (inputs[85]);
    assign layer0_outputs[5604] = ~(inputs[159]);
    assign layer0_outputs[5605] = ~((inputs[81]) | (inputs[520]));
    assign layer0_outputs[5606] = 1'b0;
    assign layer0_outputs[5607] = inputs[69];
    assign layer0_outputs[5608] = inputs[582];
    assign layer0_outputs[5609] = inputs[182];
    assign layer0_outputs[5610] = inputs[558];
    assign layer0_outputs[5611] = (inputs[88]) | (inputs[750]);
    assign layer0_outputs[5612] = 1'b1;
    assign layer0_outputs[5613] = 1'b1;
    assign layer0_outputs[5614] = 1'b0;
    assign layer0_outputs[5615] = inputs[849];
    assign layer0_outputs[5616] = ~((inputs[1012]) ^ (inputs[58]));
    assign layer0_outputs[5617] = ~((inputs[189]) ^ (inputs[168]));
    assign layer0_outputs[5618] = inputs[67];
    assign layer0_outputs[5619] = ~((inputs[399]) | (inputs[712]));
    assign layer0_outputs[5620] = ~((inputs[784]) | (inputs[700]));
    assign layer0_outputs[5621] = inputs[953];
    assign layer0_outputs[5622] = 1'b1;
    assign layer0_outputs[5623] = 1'b0;
    assign layer0_outputs[5624] = ~(inputs[675]);
    assign layer0_outputs[5625] = ~((inputs[1008]) | (inputs[478]));
    assign layer0_outputs[5626] = (inputs[152]) & ~(inputs[100]);
    assign layer0_outputs[5627] = ~((inputs[801]) | (inputs[422]));
    assign layer0_outputs[5628] = ~((inputs[6]) ^ (inputs[883]));
    assign layer0_outputs[5629] = (inputs[393]) ^ (inputs[9]);
    assign layer0_outputs[5630] = ~((inputs[667]) | (inputs[847]));
    assign layer0_outputs[5631] = ~(inputs[146]) | (inputs[995]);
    assign layer0_outputs[5632] = (inputs[610]) | (inputs[997]);
    assign layer0_outputs[5633] = (inputs[574]) & (inputs[31]);
    assign layer0_outputs[5634] = ~(inputs[934]) | (inputs[800]);
    assign layer0_outputs[5635] = ~((inputs[767]) | (inputs[584]));
    assign layer0_outputs[5636] = (inputs[748]) | (inputs[538]);
    assign layer0_outputs[5637] = ~((inputs[980]) | (inputs[707]));
    assign layer0_outputs[5638] = ~(inputs[508]) | (inputs[190]);
    assign layer0_outputs[5639] = ~(inputs[689]);
    assign layer0_outputs[5640] = (inputs[508]) | (inputs[371]);
    assign layer0_outputs[5641] = ~(inputs[505]) | (inputs[417]);
    assign layer0_outputs[5642] = 1'b0;
    assign layer0_outputs[5643] = ~((inputs[198]) | (inputs[182]));
    assign layer0_outputs[5644] = (inputs[949]) | (inputs[483]);
    assign layer0_outputs[5645] = (inputs[330]) & ~(inputs[104]);
    assign layer0_outputs[5646] = ~((inputs[851]) | (inputs[901]));
    assign layer0_outputs[5647] = inputs[964];
    assign layer0_outputs[5648] = ~(inputs[824]);
    assign layer0_outputs[5649] = (inputs[214]) & ~(inputs[891]);
    assign layer0_outputs[5650] = (inputs[1014]) & ~(inputs[181]);
    assign layer0_outputs[5651] = 1'b1;
    assign layer0_outputs[5652] = ~((inputs[897]) | (inputs[534]));
    assign layer0_outputs[5653] = ~((inputs[731]) | (inputs[158]));
    assign layer0_outputs[5654] = 1'b0;
    assign layer0_outputs[5655] = 1'b0;
    assign layer0_outputs[5656] = (inputs[784]) | (inputs[27]);
    assign layer0_outputs[5657] = ~((inputs[758]) & (inputs[908]));
    assign layer0_outputs[5658] = (inputs[820]) & ~(inputs[288]);
    assign layer0_outputs[5659] = ~(inputs[374]) | (inputs[105]);
    assign layer0_outputs[5660] = ~(inputs[837]);
    assign layer0_outputs[5661] = ~(inputs[880]) | (inputs[514]);
    assign layer0_outputs[5662] = ~((inputs[887]) ^ (inputs[856]));
    assign layer0_outputs[5663] = ~(inputs[770]) | (inputs[640]);
    assign layer0_outputs[5664] = (inputs[439]) | (inputs[624]);
    assign layer0_outputs[5665] = (inputs[98]) | (inputs[904]);
    assign layer0_outputs[5666] = ~((inputs[94]) & (inputs[954]));
    assign layer0_outputs[5667] = (inputs[111]) ^ (inputs[805]);
    assign layer0_outputs[5668] = (inputs[719]) | (inputs[676]);
    assign layer0_outputs[5669] = inputs[590];
    assign layer0_outputs[5670] = ~(inputs[564]);
    assign layer0_outputs[5671] = inputs[335];
    assign layer0_outputs[5672] = ~(inputs[786]);
    assign layer0_outputs[5673] = ~(inputs[585]);
    assign layer0_outputs[5674] = ~((inputs[332]) ^ (inputs[193]));
    assign layer0_outputs[5675] = ~((inputs[863]) | (inputs[777]));
    assign layer0_outputs[5676] = ~(inputs[586]) | (inputs[868]);
    assign layer0_outputs[5677] = (inputs[122]) ^ (inputs[1018]);
    assign layer0_outputs[5678] = (inputs[20]) ^ (inputs[147]);
    assign layer0_outputs[5679] = ~(inputs[743]) | (inputs[127]);
    assign layer0_outputs[5680] = (inputs[553]) ^ (inputs[930]);
    assign layer0_outputs[5681] = (inputs[911]) | (inputs[825]);
    assign layer0_outputs[5682] = inputs[671];
    assign layer0_outputs[5683] = ~((inputs[66]) ^ (inputs[786]));
    assign layer0_outputs[5684] = ~(inputs[120]);
    assign layer0_outputs[5685] = ~((inputs[933]) ^ (inputs[224]));
    assign layer0_outputs[5686] = (inputs[233]) | (inputs[904]);
    assign layer0_outputs[5687] = ~(inputs[229]);
    assign layer0_outputs[5688] = ~(inputs[907]);
    assign layer0_outputs[5689] = (inputs[55]) | (inputs[786]);
    assign layer0_outputs[5690] = ~(inputs[625]);
    assign layer0_outputs[5691] = (inputs[131]) & (inputs[1017]);
    assign layer0_outputs[5692] = inputs[59];
    assign layer0_outputs[5693] = ~(inputs[250]);
    assign layer0_outputs[5694] = ~((inputs[746]) | (inputs[711]));
    assign layer0_outputs[5695] = (inputs[1015]) | (inputs[232]);
    assign layer0_outputs[5696] = ~(inputs[167]) | (inputs[1017]);
    assign layer0_outputs[5697] = ~(inputs[151]);
    assign layer0_outputs[5698] = (inputs[813]) | (inputs[282]);
    assign layer0_outputs[5699] = ~(inputs[775]);
    assign layer0_outputs[5700] = (inputs[100]) & (inputs[959]);
    assign layer0_outputs[5701] = (inputs[76]) & ~(inputs[34]);
    assign layer0_outputs[5702] = ~(inputs[622]);
    assign layer0_outputs[5703] = ~(inputs[274]) | (inputs[97]);
    assign layer0_outputs[5704] = (inputs[987]) | (inputs[444]);
    assign layer0_outputs[5705] = ~((inputs[937]) | (inputs[609]));
    assign layer0_outputs[5706] = (inputs[346]) | (inputs[781]);
    assign layer0_outputs[5707] = ~(inputs[618]);
    assign layer0_outputs[5708] = inputs[567];
    assign layer0_outputs[5709] = inputs[127];
    assign layer0_outputs[5710] = inputs[552];
    assign layer0_outputs[5711] = ~((inputs[305]) | (inputs[251]));
    assign layer0_outputs[5712] = (inputs[816]) ^ (inputs[990]);
    assign layer0_outputs[5713] = (inputs[210]) & ~(inputs[3]);
    assign layer0_outputs[5714] = ~((inputs[56]) ^ (inputs[717]));
    assign layer0_outputs[5715] = inputs[714];
    assign layer0_outputs[5716] = (inputs[243]) & ~(inputs[815]);
    assign layer0_outputs[5717] = ~((inputs[416]) & (inputs[93]));
    assign layer0_outputs[5718] = (inputs[176]) | (inputs[85]);
    assign layer0_outputs[5719] = ~((inputs[31]) ^ (inputs[678]));
    assign layer0_outputs[5720] = (inputs[686]) & ~(inputs[437]);
    assign layer0_outputs[5721] = ~((inputs[356]) | (inputs[801]));
    assign layer0_outputs[5722] = inputs[245];
    assign layer0_outputs[5723] = (inputs[906]) & ~(inputs[859]);
    assign layer0_outputs[5724] = ~(inputs[758]) | (inputs[473]);
    assign layer0_outputs[5725] = ~((inputs[375]) | (inputs[221]));
    assign layer0_outputs[5726] = inputs[727];
    assign layer0_outputs[5727] = (inputs[729]) & (inputs[681]);
    assign layer0_outputs[5728] = (inputs[329]) & ~(inputs[131]);
    assign layer0_outputs[5729] = ~((inputs[943]) | (inputs[806]));
    assign layer0_outputs[5730] = ~((inputs[286]) | (inputs[591]));
    assign layer0_outputs[5731] = inputs[832];
    assign layer0_outputs[5732] = ~(inputs[501]) | (inputs[710]);
    assign layer0_outputs[5733] = (inputs[727]) & ~(inputs[789]);
    assign layer0_outputs[5734] = (inputs[759]) | (inputs[662]);
    assign layer0_outputs[5735] = ~((inputs[521]) | (inputs[120]));
    assign layer0_outputs[5736] = ~(inputs[742]) | (inputs[118]);
    assign layer0_outputs[5737] = ~(inputs[674]) | (inputs[644]);
    assign layer0_outputs[5738] = ~((inputs[939]) ^ (inputs[860]));
    assign layer0_outputs[5739] = ~((inputs[609]) ^ (inputs[907]));
    assign layer0_outputs[5740] = ~((inputs[500]) ^ (inputs[451]));
    assign layer0_outputs[5741] = (inputs[196]) & ~(inputs[165]);
    assign layer0_outputs[5742] = (inputs[302]) ^ (inputs[410]);
    assign layer0_outputs[5743] = (inputs[607]) | (inputs[1004]);
    assign layer0_outputs[5744] = (inputs[665]) & ~(inputs[89]);
    assign layer0_outputs[5745] = ~((inputs[468]) ^ (inputs[454]));
    assign layer0_outputs[5746] = ~(inputs[781]);
    assign layer0_outputs[5747] = (inputs[899]) & ~(inputs[129]);
    assign layer0_outputs[5748] = (inputs[538]) | (inputs[980]);
    assign layer0_outputs[5749] = inputs[145];
    assign layer0_outputs[5750] = ~((inputs[151]) ^ (inputs[209]));
    assign layer0_outputs[5751] = ~((inputs[177]) | (inputs[190]));
    assign layer0_outputs[5752] = ~(inputs[596]) | (inputs[74]);
    assign layer0_outputs[5753] = ~(inputs[461]) | (inputs[515]);
    assign layer0_outputs[5754] = ~((inputs[857]) ^ (inputs[146]));
    assign layer0_outputs[5755] = ~((inputs[757]) | (inputs[203]));
    assign layer0_outputs[5756] = (inputs[374]) & ~(inputs[725]);
    assign layer0_outputs[5757] = ~(inputs[978]);
    assign layer0_outputs[5758] = (inputs[436]) & ~(inputs[997]);
    assign layer0_outputs[5759] = ~(inputs[669]);
    assign layer0_outputs[5760] = (inputs[147]) & ~(inputs[314]);
    assign layer0_outputs[5761] = ~(inputs[683]);
    assign layer0_outputs[5762] = ~(inputs[656]);
    assign layer0_outputs[5763] = (inputs[818]) ^ (inputs[83]);
    assign layer0_outputs[5764] = ~((inputs[170]) ^ (inputs[111]));
    assign layer0_outputs[5765] = ~(inputs[333]);
    assign layer0_outputs[5766] = ~(inputs[561]) | (inputs[971]);
    assign layer0_outputs[5767] = (inputs[389]) | (inputs[152]);
    assign layer0_outputs[5768] = inputs[635];
    assign layer0_outputs[5769] = inputs[28];
    assign layer0_outputs[5770] = ~(inputs[303]);
    assign layer0_outputs[5771] = ~((inputs[539]) | (inputs[895]));
    assign layer0_outputs[5772] = (inputs[148]) | (inputs[452]);
    assign layer0_outputs[5773] = ~((inputs[820]) | (inputs[711]));
    assign layer0_outputs[5774] = (inputs[397]) & ~(inputs[980]);
    assign layer0_outputs[5775] = ~(inputs[339]) | (inputs[42]);
    assign layer0_outputs[5776] = (inputs[230]) ^ (inputs[455]);
    assign layer0_outputs[5777] = ~((inputs[704]) | (inputs[986]));
    assign layer0_outputs[5778] = ~((inputs[760]) | (inputs[745]));
    assign layer0_outputs[5779] = ~((inputs[306]) | (inputs[43]));
    assign layer0_outputs[5780] = ~((inputs[413]) | (inputs[816]));
    assign layer0_outputs[5781] = (inputs[390]) & ~(inputs[989]);
    assign layer0_outputs[5782] = inputs[563];
    assign layer0_outputs[5783] = ~(inputs[480]);
    assign layer0_outputs[5784] = (inputs[761]) ^ (inputs[742]);
    assign layer0_outputs[5785] = ~(inputs[393]) | (inputs[106]);
    assign layer0_outputs[5786] = ~((inputs[186]) ^ (inputs[879]));
    assign layer0_outputs[5787] = ~((inputs[560]) ^ (inputs[605]));
    assign layer0_outputs[5788] = ~((inputs[362]) ^ (inputs[701]));
    assign layer0_outputs[5789] = (inputs[685]) ^ (inputs[552]);
    assign layer0_outputs[5790] = ~(inputs[475]);
    assign layer0_outputs[5791] = (inputs[499]) & ~(inputs[683]);
    assign layer0_outputs[5792] = (inputs[381]) | (inputs[754]);
    assign layer0_outputs[5793] = ~(inputs[840]) | (inputs[6]);
    assign layer0_outputs[5794] = ~(inputs[144]) | (inputs[468]);
    assign layer0_outputs[5795] = 1'b0;
    assign layer0_outputs[5796] = (inputs[257]) | (inputs[336]);
    assign layer0_outputs[5797] = (inputs[223]) & ~(inputs[792]);
    assign layer0_outputs[5798] = (inputs[453]) & ~(inputs[737]);
    assign layer0_outputs[5799] = ~(inputs[731]) | (inputs[951]);
    assign layer0_outputs[5800] = ~((inputs[738]) ^ (inputs[895]));
    assign layer0_outputs[5801] = inputs[11];
    assign layer0_outputs[5802] = (inputs[221]) & ~(inputs[341]);
    assign layer0_outputs[5803] = ~((inputs[230]) ^ (inputs[86]));
    assign layer0_outputs[5804] = inputs[32];
    assign layer0_outputs[5805] = (inputs[268]) & ~(inputs[50]);
    assign layer0_outputs[5806] = inputs[695];
    assign layer0_outputs[5807] = ~(inputs[108]);
    assign layer0_outputs[5808] = (inputs[516]) & ~(inputs[519]);
    assign layer0_outputs[5809] = 1'b1;
    assign layer0_outputs[5810] = (inputs[542]) & (inputs[599]);
    assign layer0_outputs[5811] = ~(inputs[31]) | (inputs[229]);
    assign layer0_outputs[5812] = ~((inputs[525]) | (inputs[587]));
    assign layer0_outputs[5813] = 1'b0;
    assign layer0_outputs[5814] = (inputs[252]) ^ (inputs[867]);
    assign layer0_outputs[5815] = inputs[716];
    assign layer0_outputs[5816] = ~(inputs[614]);
    assign layer0_outputs[5817] = ~(inputs[855]) | (inputs[390]);
    assign layer0_outputs[5818] = (inputs[768]) ^ (inputs[894]);
    assign layer0_outputs[5819] = ~(inputs[941]);
    assign layer0_outputs[5820] = ~((inputs[799]) | (inputs[436]));
    assign layer0_outputs[5821] = (inputs[443]) & (inputs[255]);
    assign layer0_outputs[5822] = ~((inputs[466]) ^ (inputs[382]));
    assign layer0_outputs[5823] = ~(inputs[272]);
    assign layer0_outputs[5824] = ~((inputs[704]) & (inputs[225]));
    assign layer0_outputs[5825] = inputs[58];
    assign layer0_outputs[5826] = (inputs[786]) & ~(inputs[159]);
    assign layer0_outputs[5827] = ~((inputs[806]) ^ (inputs[797]));
    assign layer0_outputs[5828] = ~(inputs[779]) | (inputs[126]);
    assign layer0_outputs[5829] = (inputs[204]) ^ (inputs[190]);
    assign layer0_outputs[5830] = (inputs[84]) | (inputs[513]);
    assign layer0_outputs[5831] = (inputs[404]) | (inputs[932]);
    assign layer0_outputs[5832] = inputs[312];
    assign layer0_outputs[5833] = ~(inputs[56]) | (inputs[859]);
    assign layer0_outputs[5834] = ~(inputs[519]);
    assign layer0_outputs[5835] = ~(inputs[590]);
    assign layer0_outputs[5836] = ~(inputs[238]) | (inputs[568]);
    assign layer0_outputs[5837] = ~(inputs[262]);
    assign layer0_outputs[5838] = ~((inputs[1017]) ^ (inputs[513]));
    assign layer0_outputs[5839] = ~((inputs[876]) ^ (inputs[657]));
    assign layer0_outputs[5840] = (inputs[879]) ^ (inputs[21]);
    assign layer0_outputs[5841] = ~(inputs[111]) | (inputs[796]);
    assign layer0_outputs[5842] = ~((inputs[384]) | (inputs[568]));
    assign layer0_outputs[5843] = ~(inputs[419]) | (inputs[3]);
    assign layer0_outputs[5844] = ~((inputs[106]) ^ (inputs[258]));
    assign layer0_outputs[5845] = ~((inputs[651]) ^ (inputs[605]));
    assign layer0_outputs[5846] = (inputs[64]) & ~(inputs[480]);
    assign layer0_outputs[5847] = ~(inputs[297]);
    assign layer0_outputs[5848] = inputs[522];
    assign layer0_outputs[5849] = (inputs[432]) | (inputs[470]);
    assign layer0_outputs[5850] = (inputs[589]) & ~(inputs[962]);
    assign layer0_outputs[5851] = ~((inputs[37]) | (inputs[222]));
    assign layer0_outputs[5852] = (inputs[593]) | (inputs[342]);
    assign layer0_outputs[5853] = ~(inputs[13]) | (inputs[89]);
    assign layer0_outputs[5854] = (inputs[919]) ^ (inputs[218]);
    assign layer0_outputs[5855] = inputs[1023];
    assign layer0_outputs[5856] = (inputs[907]) & ~(inputs[737]);
    assign layer0_outputs[5857] = 1'b1;
    assign layer0_outputs[5858] = (inputs[309]) ^ (inputs[216]);
    assign layer0_outputs[5859] = ~((inputs[141]) | (inputs[48]));
    assign layer0_outputs[5860] = (inputs[434]) & ~(inputs[459]);
    assign layer0_outputs[5861] = ~((inputs[546]) ^ (inputs[17]));
    assign layer0_outputs[5862] = 1'b1;
    assign layer0_outputs[5863] = (inputs[147]) ^ (inputs[283]);
    assign layer0_outputs[5864] = (inputs[625]) & ~(inputs[286]);
    assign layer0_outputs[5865] = ~(inputs[148]) | (inputs[733]);
    assign layer0_outputs[5866] = ~(inputs[367]);
    assign layer0_outputs[5867] = ~((inputs[564]) ^ (inputs[119]));
    assign layer0_outputs[5868] = inputs[254];
    assign layer0_outputs[5869] = (inputs[359]) ^ (inputs[483]);
    assign layer0_outputs[5870] = inputs[297];
    assign layer0_outputs[5871] = (inputs[212]) & ~(inputs[232]);
    assign layer0_outputs[5872] = 1'b0;
    assign layer0_outputs[5873] = (inputs[80]) & ~(inputs[835]);
    assign layer0_outputs[5874] = ~(inputs[710]) | (inputs[283]);
    assign layer0_outputs[5875] = (inputs[645]) | (inputs[311]);
    assign layer0_outputs[5876] = ~(inputs[300]);
    assign layer0_outputs[5877] = ~((inputs[132]) ^ (inputs[773]));
    assign layer0_outputs[5878] = (inputs[13]) | (inputs[870]);
    assign layer0_outputs[5879] = (inputs[980]) | (inputs[910]);
    assign layer0_outputs[5880] = ~((inputs[411]) | (inputs[240]));
    assign layer0_outputs[5881] = 1'b0;
    assign layer0_outputs[5882] = (inputs[602]) | (inputs[53]);
    assign layer0_outputs[5883] = ~((inputs[178]) ^ (inputs[958]));
    assign layer0_outputs[5884] = (inputs[581]) ^ (inputs[524]);
    assign layer0_outputs[5885] = inputs[82];
    assign layer0_outputs[5886] = ~(inputs[305]);
    assign layer0_outputs[5887] = (inputs[6]) & ~(inputs[17]);
    assign layer0_outputs[5888] = ~(inputs[391]);
    assign layer0_outputs[5889] = ~((inputs[627]) ^ (inputs[740]));
    assign layer0_outputs[5890] = 1'b1;
    assign layer0_outputs[5891] = inputs[271];
    assign layer0_outputs[5892] = (inputs[678]) | (inputs[815]);
    assign layer0_outputs[5893] = (inputs[522]) | (inputs[619]);
    assign layer0_outputs[5894] = ~((inputs[523]) ^ (inputs[933]));
    assign layer0_outputs[5895] = ~(inputs[243]) | (inputs[594]);
    assign layer0_outputs[5896] = (inputs[576]) ^ (inputs[723]);
    assign layer0_outputs[5897] = ~((inputs[404]) & (inputs[301]));
    assign layer0_outputs[5898] = ~((inputs[31]) ^ (inputs[123]));
    assign layer0_outputs[5899] = ~((inputs[990]) ^ (inputs[705]));
    assign layer0_outputs[5900] = inputs[837];
    assign layer0_outputs[5901] = ~(inputs[271]);
    assign layer0_outputs[5902] = ~((inputs[946]) ^ (inputs[730]));
    assign layer0_outputs[5903] = ~(inputs[652]);
    assign layer0_outputs[5904] = ~(inputs[604]) | (inputs[351]);
    assign layer0_outputs[5905] = ~(inputs[626]) | (inputs[435]);
    assign layer0_outputs[5906] = 1'b0;
    assign layer0_outputs[5907] = 1'b1;
    assign layer0_outputs[5908] = inputs[295];
    assign layer0_outputs[5909] = inputs[774];
    assign layer0_outputs[5910] = ~(inputs[834]) | (inputs[380]);
    assign layer0_outputs[5911] = ~(inputs[751]);
    assign layer0_outputs[5912] = (inputs[869]) ^ (inputs[643]);
    assign layer0_outputs[5913] = ~((inputs[567]) & (inputs[535]));
    assign layer0_outputs[5914] = (inputs[618]) & ~(inputs[950]);
    assign layer0_outputs[5915] = ~((inputs[143]) | (inputs[659]));
    assign layer0_outputs[5916] = inputs[594];
    assign layer0_outputs[5917] = ~((inputs[608]) | (inputs[545]));
    assign layer0_outputs[5918] = ~(inputs[738]);
    assign layer0_outputs[5919] = (inputs[357]) ^ (inputs[12]);
    assign layer0_outputs[5920] = 1'b0;
    assign layer0_outputs[5921] = ~((inputs[314]) | (inputs[788]));
    assign layer0_outputs[5922] = (inputs[925]) & ~(inputs[288]);
    assign layer0_outputs[5923] = (inputs[565]) & ~(inputs[64]);
    assign layer0_outputs[5924] = ~((inputs[341]) ^ (inputs[639]));
    assign layer0_outputs[5925] = (inputs[493]) | (inputs[645]);
    assign layer0_outputs[5926] = ~(inputs[495]) | (inputs[220]);
    assign layer0_outputs[5927] = inputs[2];
    assign layer0_outputs[5928] = ~(inputs[636]);
    assign layer0_outputs[5929] = (inputs[78]) ^ (inputs[726]);
    assign layer0_outputs[5930] = (inputs[834]) | (inputs[142]);
    assign layer0_outputs[5931] = ~((inputs[436]) | (inputs[954]));
    assign layer0_outputs[5932] = ~(inputs[574]) | (inputs[120]);
    assign layer0_outputs[5933] = inputs[210];
    assign layer0_outputs[5934] = ~(inputs[799]) | (inputs[928]);
    assign layer0_outputs[5935] = 1'b0;
    assign layer0_outputs[5936] = ~(inputs[272]);
    assign layer0_outputs[5937] = 1'b0;
    assign layer0_outputs[5938] = ~((inputs[668]) ^ (inputs[135]));
    assign layer0_outputs[5939] = ~(inputs[467]);
    assign layer0_outputs[5940] = ~(inputs[877]);
    assign layer0_outputs[5941] = inputs[40];
    assign layer0_outputs[5942] = ~(inputs[149]) | (inputs[858]);
    assign layer0_outputs[5943] = inputs[493];
    assign layer0_outputs[5944] = inputs[277];
    assign layer0_outputs[5945] = ~((inputs[507]) ^ (inputs[94]));
    assign layer0_outputs[5946] = ~(inputs[101]) | (inputs[324]);
    assign layer0_outputs[5947] = 1'b0;
    assign layer0_outputs[5948] = (inputs[447]) & (inputs[12]);
    assign layer0_outputs[5949] = ~((inputs[890]) & (inputs[962]));
    assign layer0_outputs[5950] = (inputs[490]) & ~(inputs[1006]);
    assign layer0_outputs[5951] = ~(inputs[760]) | (inputs[767]);
    assign layer0_outputs[5952] = inputs[193];
    assign layer0_outputs[5953] = (inputs[475]) | (inputs[236]);
    assign layer0_outputs[5954] = ~((inputs[457]) ^ (inputs[931]));
    assign layer0_outputs[5955] = ~((inputs[339]) ^ (inputs[728]));
    assign layer0_outputs[5956] = (inputs[751]) & ~(inputs[839]);
    assign layer0_outputs[5957] = inputs[217];
    assign layer0_outputs[5958] = ~(inputs[912]) | (inputs[1021]);
    assign layer0_outputs[5959] = (inputs[133]) & (inputs[921]);
    assign layer0_outputs[5960] = (inputs[467]) ^ (inputs[298]);
    assign layer0_outputs[5961] = ~(inputs[21]);
    assign layer0_outputs[5962] = ~(inputs[747]) | (inputs[644]);
    assign layer0_outputs[5963] = 1'b0;
    assign layer0_outputs[5964] = ~((inputs[640]) | (inputs[78]));
    assign layer0_outputs[5965] = (inputs[653]) & ~(inputs[710]);
    assign layer0_outputs[5966] = inputs[131];
    assign layer0_outputs[5967] = ~(inputs[854]) | (inputs[319]);
    assign layer0_outputs[5968] = ~((inputs[372]) | (inputs[417]));
    assign layer0_outputs[5969] = (inputs[970]) | (inputs[81]);
    assign layer0_outputs[5970] = ~(inputs[499]) | (inputs[68]);
    assign layer0_outputs[5971] = 1'b1;
    assign layer0_outputs[5972] = ~((inputs[640]) ^ (inputs[478]));
    assign layer0_outputs[5973] = (inputs[646]) & ~(inputs[444]);
    assign layer0_outputs[5974] = inputs[102];
    assign layer0_outputs[5975] = inputs[577];
    assign layer0_outputs[5976] = inputs[454];
    assign layer0_outputs[5977] = ~((inputs[880]) ^ (inputs[561]));
    assign layer0_outputs[5978] = ~(inputs[936]) | (inputs[850]);
    assign layer0_outputs[5979] = (inputs[707]) | (inputs[746]);
    assign layer0_outputs[5980] = ~((inputs[201]) | (inputs[665]));
    assign layer0_outputs[5981] = ~(inputs[658]) | (inputs[993]);
    assign layer0_outputs[5982] = ~((inputs[724]) ^ (inputs[450]));
    assign layer0_outputs[5983] = (inputs[807]) & ~(inputs[1003]);
    assign layer0_outputs[5984] = (inputs[151]) | (inputs[673]);
    assign layer0_outputs[5985] = ~((inputs[3]) | (inputs[872]));
    assign layer0_outputs[5986] = (inputs[558]) | (inputs[445]);
    assign layer0_outputs[5987] = ~(inputs[498]) | (inputs[772]);
    assign layer0_outputs[5988] = (inputs[149]) ^ (inputs[258]);
    assign layer0_outputs[5989] = ~(inputs[519]) | (inputs[487]);
    assign layer0_outputs[5990] = ~((inputs[778]) | (inputs[52]));
    assign layer0_outputs[5991] = ~((inputs[231]) ^ (inputs[662]));
    assign layer0_outputs[5992] = ~(inputs[968]);
    assign layer0_outputs[5993] = (inputs[624]) ^ (inputs[1011]);
    assign layer0_outputs[5994] = inputs[596];
    assign layer0_outputs[5995] = inputs[629];
    assign layer0_outputs[5996] = ~(inputs[543]);
    assign layer0_outputs[5997] = ~((inputs[951]) ^ (inputs[732]));
    assign layer0_outputs[5998] = (inputs[775]) & (inputs[834]);
    assign layer0_outputs[5999] = inputs[613];
    assign layer0_outputs[6000] = 1'b1;
    assign layer0_outputs[6001] = (inputs[943]) & ~(inputs[431]);
    assign layer0_outputs[6002] = ~((inputs[68]) & (inputs[165]));
    assign layer0_outputs[6003] = ~(inputs[298]) | (inputs[473]);
    assign layer0_outputs[6004] = ~(inputs[710]) | (inputs[415]);
    assign layer0_outputs[6005] = ~(inputs[343]) | (inputs[969]);
    assign layer0_outputs[6006] = ~(inputs[824]);
    assign layer0_outputs[6007] = ~(inputs[506]);
    assign layer0_outputs[6008] = inputs[846];
    assign layer0_outputs[6009] = ~(inputs[533]) | (inputs[451]);
    assign layer0_outputs[6010] = ~((inputs[470]) & (inputs[864]));
    assign layer0_outputs[6011] = ~(inputs[654]);
    assign layer0_outputs[6012] = ~((inputs[882]) | (inputs[424]));
    assign layer0_outputs[6013] = (inputs[468]) | (inputs[857]);
    assign layer0_outputs[6014] = (inputs[185]) | (inputs[491]);
    assign layer0_outputs[6015] = inputs[571];
    assign layer0_outputs[6016] = ~(inputs[905]) | (inputs[18]);
    assign layer0_outputs[6017] = ~(inputs[530]) | (inputs[65]);
    assign layer0_outputs[6018] = inputs[544];
    assign layer0_outputs[6019] = ~(inputs[246]);
    assign layer0_outputs[6020] = 1'b0;
    assign layer0_outputs[6021] = (inputs[970]) | (inputs[475]);
    assign layer0_outputs[6022] = ~((inputs[869]) | (inputs[1014]));
    assign layer0_outputs[6023] = (inputs[194]) & (inputs[384]);
    assign layer0_outputs[6024] = (inputs[208]) | (inputs[936]);
    assign layer0_outputs[6025] = (inputs[521]) | (inputs[764]);
    assign layer0_outputs[6026] = (inputs[538]) | (inputs[684]);
    assign layer0_outputs[6027] = ~((inputs[794]) ^ (inputs[466]));
    assign layer0_outputs[6028] = inputs[278];
    assign layer0_outputs[6029] = ~(inputs[236]) | (inputs[46]);
    assign layer0_outputs[6030] = (inputs[825]) ^ (inputs[332]);
    assign layer0_outputs[6031] = (inputs[511]) ^ (inputs[901]);
    assign layer0_outputs[6032] = (inputs[456]) & ~(inputs[698]);
    assign layer0_outputs[6033] = ~(inputs[461]) | (inputs[838]);
    assign layer0_outputs[6034] = ~(inputs[652]) | (inputs[906]);
    assign layer0_outputs[6035] = (inputs[746]) | (inputs[354]);
    assign layer0_outputs[6036] = (inputs[630]) & ~(inputs[435]);
    assign layer0_outputs[6037] = 1'b0;
    assign layer0_outputs[6038] = ~(inputs[757]);
    assign layer0_outputs[6039] = (inputs[163]) | (inputs[975]);
    assign layer0_outputs[6040] = ~((inputs[590]) | (inputs[13]));
    assign layer0_outputs[6041] = (inputs[796]) | (inputs[817]);
    assign layer0_outputs[6042] = inputs[495];
    assign layer0_outputs[6043] = ~(inputs[591]) | (inputs[257]);
    assign layer0_outputs[6044] = inputs[116];
    assign layer0_outputs[6045] = ~(inputs[505]);
    assign layer0_outputs[6046] = ~((inputs[120]) | (inputs[610]));
    assign layer0_outputs[6047] = 1'b0;
    assign layer0_outputs[6048] = 1'b0;
    assign layer0_outputs[6049] = ~(inputs[715]);
    assign layer0_outputs[6050] = ~(inputs[1000]) | (inputs[844]);
    assign layer0_outputs[6051] = (inputs[68]) | (inputs[839]);
    assign layer0_outputs[6052] = (inputs[277]) ^ (inputs[730]);
    assign layer0_outputs[6053] = (inputs[899]) | (inputs[488]);
    assign layer0_outputs[6054] = inputs[323];
    assign layer0_outputs[6055] = ~(inputs[242]);
    assign layer0_outputs[6056] = ~((inputs[717]) | (inputs[853]));
    assign layer0_outputs[6057] = (inputs[851]) & (inputs[552]);
    assign layer0_outputs[6058] = ~((inputs[1015]) | (inputs[64]));
    assign layer0_outputs[6059] = ~(inputs[789]);
    assign layer0_outputs[6060] = ~(inputs[362]);
    assign layer0_outputs[6061] = ~((inputs[266]) ^ (inputs[146]));
    assign layer0_outputs[6062] = (inputs[127]) | (inputs[949]);
    assign layer0_outputs[6063] = (inputs[951]) & ~(inputs[580]);
    assign layer0_outputs[6064] = inputs[271];
    assign layer0_outputs[6065] = ~((inputs[382]) ^ (inputs[1012]));
    assign layer0_outputs[6066] = ~((inputs[539]) | (inputs[594]));
    assign layer0_outputs[6067] = 1'b1;
    assign layer0_outputs[6068] = ~((inputs[309]) ^ (inputs[387]));
    assign layer0_outputs[6069] = (inputs[619]) & ~(inputs[49]);
    assign layer0_outputs[6070] = (inputs[99]) | (inputs[451]);
    assign layer0_outputs[6071] = ~((inputs[263]) | (inputs[804]));
    assign layer0_outputs[6072] = ~(inputs[569]);
    assign layer0_outputs[6073] = ~((inputs[910]) ^ (inputs[450]));
    assign layer0_outputs[6074] = (inputs[556]) ^ (inputs[797]);
    assign layer0_outputs[6075] = (inputs[921]) ^ (inputs[972]);
    assign layer0_outputs[6076] = ~(inputs[470]);
    assign layer0_outputs[6077] = 1'b0;
    assign layer0_outputs[6078] = (inputs[805]) | (inputs[706]);
    assign layer0_outputs[6079] = ~(inputs[841]);
    assign layer0_outputs[6080] = ~(inputs[942]);
    assign layer0_outputs[6081] = ~((inputs[991]) | (inputs[440]));
    assign layer0_outputs[6082] = (inputs[944]) ^ (inputs[76]);
    assign layer0_outputs[6083] = ~((inputs[693]) & (inputs[997]));
    assign layer0_outputs[6084] = (inputs[465]) & ~(inputs[508]);
    assign layer0_outputs[6085] = (inputs[294]) | (inputs[811]);
    assign layer0_outputs[6086] = ~((inputs[702]) | (inputs[721]));
    assign layer0_outputs[6087] = ~(inputs[1012]);
    assign layer0_outputs[6088] = ~(inputs[370]) | (inputs[947]);
    assign layer0_outputs[6089] = (inputs[180]) ^ (inputs[876]);
    assign layer0_outputs[6090] = ~((inputs[909]) ^ (inputs[45]));
    assign layer0_outputs[6091] = ~(inputs[522]);
    assign layer0_outputs[6092] = ~((inputs[509]) ^ (inputs[299]));
    assign layer0_outputs[6093] = (inputs[378]) | (inputs[943]);
    assign layer0_outputs[6094] = (inputs[856]) ^ (inputs[1011]);
    assign layer0_outputs[6095] = ~(inputs[719]);
    assign layer0_outputs[6096] = (inputs[976]) & ~(inputs[95]);
    assign layer0_outputs[6097] = ~(inputs[210]);
    assign layer0_outputs[6098] = ~(inputs[867]) | (inputs[192]);
    assign layer0_outputs[6099] = (inputs[347]) | (inputs[430]);
    assign layer0_outputs[6100] = ~(inputs[417]) | (inputs[50]);
    assign layer0_outputs[6101] = ~(inputs[941]);
    assign layer0_outputs[6102] = inputs[957];
    assign layer0_outputs[6103] = ~((inputs[444]) | (inputs[150]));
    assign layer0_outputs[6104] = (inputs[692]) | (inputs[249]);
    assign layer0_outputs[6105] = ~((inputs[937]) ^ (inputs[940]));
    assign layer0_outputs[6106] = (inputs[40]) & ~(inputs[1005]);
    assign layer0_outputs[6107] = ~(inputs[492]);
    assign layer0_outputs[6108] = (inputs[694]) | (inputs[205]);
    assign layer0_outputs[6109] = ~(inputs[911]) | (inputs[550]);
    assign layer0_outputs[6110] = ~((inputs[675]) | (inputs[798]));
    assign layer0_outputs[6111] = inputs[488];
    assign layer0_outputs[6112] = ~(inputs[506]);
    assign layer0_outputs[6113] = (inputs[588]) | (inputs[734]);
    assign layer0_outputs[6114] = (inputs[389]) | (inputs[621]);
    assign layer0_outputs[6115] = ~(inputs[308]);
    assign layer0_outputs[6116] = ~(inputs[688]) | (inputs[1008]);
    assign layer0_outputs[6117] = ~(inputs[396]);
    assign layer0_outputs[6118] = inputs[176];
    assign layer0_outputs[6119] = ~(inputs[361]) | (inputs[164]);
    assign layer0_outputs[6120] = (inputs[569]) & ~(inputs[888]);
    assign layer0_outputs[6121] = ~(inputs[552]) | (inputs[737]);
    assign layer0_outputs[6122] = inputs[201];
    assign layer0_outputs[6123] = ~(inputs[327]);
    assign layer0_outputs[6124] = ~((inputs[375]) ^ (inputs[543]));
    assign layer0_outputs[6125] = 1'b0;
    assign layer0_outputs[6126] = ~((inputs[383]) ^ (inputs[719]));
    assign layer0_outputs[6127] = ~((inputs[47]) ^ (inputs[761]));
    assign layer0_outputs[6128] = ~(inputs[556]) | (inputs[583]);
    assign layer0_outputs[6129] = inputs[151];
    assign layer0_outputs[6130] = inputs[654];
    assign layer0_outputs[6131] = ~(inputs[884]) | (inputs[169]);
    assign layer0_outputs[6132] = (inputs[393]) & ~(inputs[939]);
    assign layer0_outputs[6133] = (inputs[92]) & ~(inputs[509]);
    assign layer0_outputs[6134] = ~((inputs[815]) | (inputs[178]));
    assign layer0_outputs[6135] = ~((inputs[471]) | (inputs[467]));
    assign layer0_outputs[6136] = ~((inputs[971]) | (inputs[302]));
    assign layer0_outputs[6137] = 1'b1;
    assign layer0_outputs[6138] = ~(inputs[492]);
    assign layer0_outputs[6139] = (inputs[337]) & ~(inputs[994]);
    assign layer0_outputs[6140] = (inputs[433]) | (inputs[773]);
    assign layer0_outputs[6141] = ~((inputs[1023]) | (inputs[433]));
    assign layer0_outputs[6142] = ~(inputs[370]);
    assign layer0_outputs[6143] = (inputs[570]) ^ (inputs[928]);
    assign layer0_outputs[6144] = (inputs[544]) ^ (inputs[763]);
    assign layer0_outputs[6145] = ~((inputs[936]) | (inputs[674]));
    assign layer0_outputs[6146] = ~((inputs[808]) ^ (inputs[736]));
    assign layer0_outputs[6147] = (inputs[315]) & ~(inputs[806]);
    assign layer0_outputs[6148] = ~((inputs[177]) & (inputs[766]));
    assign layer0_outputs[6149] = ~(inputs[621]);
    assign layer0_outputs[6150] = (inputs[311]) | (inputs[909]);
    assign layer0_outputs[6151] = (inputs[978]) | (inputs[881]);
    assign layer0_outputs[6152] = ~(inputs[326]);
    assign layer0_outputs[6153] = ~(inputs[531]);
    assign layer0_outputs[6154] = ~((inputs[755]) ^ (inputs[382]));
    assign layer0_outputs[6155] = (inputs[969]) ^ (inputs[645]);
    assign layer0_outputs[6156] = (inputs[548]) & ~(inputs[114]);
    assign layer0_outputs[6157] = ~(inputs[429]) | (inputs[671]);
    assign layer0_outputs[6158] = (inputs[539]) & ~(inputs[524]);
    assign layer0_outputs[6159] = ~(inputs[693]) | (inputs[289]);
    assign layer0_outputs[6160] = ~((inputs[778]) | (inputs[698]));
    assign layer0_outputs[6161] = ~((inputs[555]) ^ (inputs[834]));
    assign layer0_outputs[6162] = ~((inputs[816]) | (inputs[391]));
    assign layer0_outputs[6163] = (inputs[662]) & ~(inputs[226]);
    assign layer0_outputs[6164] = (inputs[476]) | (inputs[40]);
    assign layer0_outputs[6165] = 1'b0;
    assign layer0_outputs[6166] = inputs[963];
    assign layer0_outputs[6167] = (inputs[423]) | (inputs[688]);
    assign layer0_outputs[6168] = ~(inputs[14]) | (inputs[1019]);
    assign layer0_outputs[6169] = (inputs[207]) & ~(inputs[72]);
    assign layer0_outputs[6170] = ~((inputs[575]) | (inputs[817]));
    assign layer0_outputs[6171] = ~(inputs[949]) | (inputs[1018]);
    assign layer0_outputs[6172] = inputs[83];
    assign layer0_outputs[6173] = ~((inputs[285]) | (inputs[10]));
    assign layer0_outputs[6174] = ~(inputs[881]) | (inputs[729]);
    assign layer0_outputs[6175] = ~(inputs[712]);
    assign layer0_outputs[6176] = (inputs[951]) | (inputs[1022]);
    assign layer0_outputs[6177] = ~(inputs[531]);
    assign layer0_outputs[6178] = ~((inputs[22]) | (inputs[744]));
    assign layer0_outputs[6179] = 1'b0;
    assign layer0_outputs[6180] = ~(inputs[177]) | (inputs[123]);
    assign layer0_outputs[6181] = ~(inputs[479]);
    assign layer0_outputs[6182] = (inputs[674]) ^ (inputs[941]);
    assign layer0_outputs[6183] = (inputs[654]) ^ (inputs[524]);
    assign layer0_outputs[6184] = (inputs[769]) & ~(inputs[377]);
    assign layer0_outputs[6185] = (inputs[574]) ^ (inputs[140]);
    assign layer0_outputs[6186] = ~(inputs[63]) | (inputs[322]);
    assign layer0_outputs[6187] = ~((inputs[439]) | (inputs[819]));
    assign layer0_outputs[6188] = (inputs[776]) & ~(inputs[830]);
    assign layer0_outputs[6189] = 1'b0;
    assign layer0_outputs[6190] = (inputs[38]) ^ (inputs[286]);
    assign layer0_outputs[6191] = inputs[438];
    assign layer0_outputs[6192] = (inputs[114]) ^ (inputs[662]);
    assign layer0_outputs[6193] = inputs[768];
    assign layer0_outputs[6194] = ~((inputs[546]) & (inputs[481]));
    assign layer0_outputs[6195] = (inputs[437]) & ~(inputs[81]);
    assign layer0_outputs[6196] = (inputs[807]) | (inputs[239]);
    assign layer0_outputs[6197] = inputs[416];
    assign layer0_outputs[6198] = 1'b0;
    assign layer0_outputs[6199] = (inputs[182]) ^ (inputs[752]);
    assign layer0_outputs[6200] = ~((inputs[638]) | (inputs[887]));
    assign layer0_outputs[6201] = ~((inputs[388]) & (inputs[639]));
    assign layer0_outputs[6202] = ~((inputs[915]) ^ (inputs[301]));
    assign layer0_outputs[6203] = (inputs[125]) ^ (inputs[313]);
    assign layer0_outputs[6204] = (inputs[157]) | (inputs[972]);
    assign layer0_outputs[6205] = ~((inputs[543]) & (inputs[602]));
    assign layer0_outputs[6206] = ~((inputs[811]) ^ (inputs[648]));
    assign layer0_outputs[6207] = ~((inputs[349]) & (inputs[475]));
    assign layer0_outputs[6208] = (inputs[416]) ^ (inputs[61]);
    assign layer0_outputs[6209] = 1'b1;
    assign layer0_outputs[6210] = (inputs[793]) ^ (inputs[58]);
    assign layer0_outputs[6211] = (inputs[245]) & ~(inputs[972]);
    assign layer0_outputs[6212] = ~((inputs[799]) | (inputs[426]));
    assign layer0_outputs[6213] = (inputs[691]) ^ (inputs[982]);
    assign layer0_outputs[6214] = 1'b1;
    assign layer0_outputs[6215] = ~(inputs[494]);
    assign layer0_outputs[6216] = ~(inputs[672]);
    assign layer0_outputs[6217] = ~((inputs[1005]) | (inputs[197]));
    assign layer0_outputs[6218] = ~(inputs[686]);
    assign layer0_outputs[6219] = ~(inputs[2]);
    assign layer0_outputs[6220] = ~(inputs[24]) | (inputs[219]);
    assign layer0_outputs[6221] = ~((inputs[124]) | (inputs[456]));
    assign layer0_outputs[6222] = ~(inputs[498]);
    assign layer0_outputs[6223] = ~((inputs[620]) | (inputs[695]));
    assign layer0_outputs[6224] = (inputs[372]) & ~(inputs[918]);
    assign layer0_outputs[6225] = ~(inputs[633]);
    assign layer0_outputs[6226] = ~((inputs[788]) | (inputs[192]));
    assign layer0_outputs[6227] = ~(inputs[590]);
    assign layer0_outputs[6228] = (inputs[269]) | (inputs[476]);
    assign layer0_outputs[6229] = ~((inputs[381]) & (inputs[918]));
    assign layer0_outputs[6230] = ~(inputs[232]);
    assign layer0_outputs[6231] = (inputs[367]) & ~(inputs[807]);
    assign layer0_outputs[6232] = ~(inputs[55]);
    assign layer0_outputs[6233] = (inputs[427]) & ~(inputs[185]);
    assign layer0_outputs[6234] = inputs[843];
    assign layer0_outputs[6235] = ~((inputs[673]) ^ (inputs[919]));
    assign layer0_outputs[6236] = inputs[613];
    assign layer0_outputs[6237] = (inputs[238]) & (inputs[725]);
    assign layer0_outputs[6238] = ~((inputs[69]) | (inputs[857]));
    assign layer0_outputs[6239] = ~(inputs[518]) | (inputs[891]);
    assign layer0_outputs[6240] = ~(inputs[869]) | (inputs[335]);
    assign layer0_outputs[6241] = (inputs[385]) ^ (inputs[232]);
    assign layer0_outputs[6242] = inputs[41];
    assign layer0_outputs[6243] = ~(inputs[281]) | (inputs[192]);
    assign layer0_outputs[6244] = (inputs[6]) ^ (inputs[460]);
    assign layer0_outputs[6245] = ~((inputs[47]) ^ (inputs[717]));
    assign layer0_outputs[6246] = (inputs[182]) & ~(inputs[874]);
    assign layer0_outputs[6247] = ~((inputs[703]) ^ (inputs[336]));
    assign layer0_outputs[6248] = ~(inputs[202]) | (inputs[89]);
    assign layer0_outputs[6249] = (inputs[977]) | (inputs[361]);
    assign layer0_outputs[6250] = (inputs[525]) ^ (inputs[81]);
    assign layer0_outputs[6251] = (inputs[412]) & (inputs[196]);
    assign layer0_outputs[6252] = ~(inputs[514]);
    assign layer0_outputs[6253] = inputs[569];
    assign layer0_outputs[6254] = inputs[584];
    assign layer0_outputs[6255] = (inputs[334]) ^ (inputs[830]);
    assign layer0_outputs[6256] = ~((inputs[33]) | (inputs[147]));
    assign layer0_outputs[6257] = ~((inputs[925]) | (inputs[199]));
    assign layer0_outputs[6258] = ~(inputs[223]);
    assign layer0_outputs[6259] = ~((inputs[259]) ^ (inputs[338]));
    assign layer0_outputs[6260] = ~((inputs[363]) | (inputs[954]));
    assign layer0_outputs[6261] = (inputs[453]) ^ (inputs[68]);
    assign layer0_outputs[6262] = (inputs[365]) ^ (inputs[326]);
    assign layer0_outputs[6263] = ~(inputs[325]);
    assign layer0_outputs[6264] = inputs[429];
    assign layer0_outputs[6265] = (inputs[911]) | (inputs[938]);
    assign layer0_outputs[6266] = inputs[105];
    assign layer0_outputs[6267] = ~((inputs[599]) | (inputs[360]));
    assign layer0_outputs[6268] = ~((inputs[602]) | (inputs[501]));
    assign layer0_outputs[6269] = ~((inputs[501]) ^ (inputs[481]));
    assign layer0_outputs[6270] = ~((inputs[1003]) ^ (inputs[237]));
    assign layer0_outputs[6271] = inputs[584];
    assign layer0_outputs[6272] = (inputs[220]) | (inputs[672]);
    assign layer0_outputs[6273] = inputs[495];
    assign layer0_outputs[6274] = (inputs[743]) | (inputs[760]);
    assign layer0_outputs[6275] = ~(inputs[376]);
    assign layer0_outputs[6276] = ~((inputs[664]) ^ (inputs[531]));
    assign layer0_outputs[6277] = ~(inputs[230]);
    assign layer0_outputs[6278] = inputs[683];
    assign layer0_outputs[6279] = ~((inputs[737]) ^ (inputs[127]));
    assign layer0_outputs[6280] = ~(inputs[584]);
    assign layer0_outputs[6281] = (inputs[727]) & ~(inputs[923]);
    assign layer0_outputs[6282] = (inputs[531]) | (inputs[8]);
    assign layer0_outputs[6283] = inputs[477];
    assign layer0_outputs[6284] = ~((inputs[750]) | (inputs[224]));
    assign layer0_outputs[6285] = (inputs[562]) | (inputs[886]);
    assign layer0_outputs[6286] = (inputs[573]) | (inputs[362]);
    assign layer0_outputs[6287] = ~(inputs[716]) | (inputs[604]);
    assign layer0_outputs[6288] = ~((inputs[24]) | (inputs[979]));
    assign layer0_outputs[6289] = ~(inputs[151]);
    assign layer0_outputs[6290] = inputs[721];
    assign layer0_outputs[6291] = (inputs[942]) & ~(inputs[1011]);
    assign layer0_outputs[6292] = ~(inputs[233]);
    assign layer0_outputs[6293] = inputs[467];
    assign layer0_outputs[6294] = ~(inputs[656]);
    assign layer0_outputs[6295] = ~((inputs[687]) | (inputs[442]));
    assign layer0_outputs[6296] = (inputs[4]) | (inputs[428]);
    assign layer0_outputs[6297] = (inputs[376]) & ~(inputs[64]);
    assign layer0_outputs[6298] = (inputs[681]) & ~(inputs[53]);
    assign layer0_outputs[6299] = ~(inputs[458]);
    assign layer0_outputs[6300] = ~(inputs[402]);
    assign layer0_outputs[6301] = ~((inputs[894]) & (inputs[766]));
    assign layer0_outputs[6302] = ~((inputs[551]) | (inputs[810]));
    assign layer0_outputs[6303] = ~(inputs[460]) | (inputs[741]);
    assign layer0_outputs[6304] = inputs[369];
    assign layer0_outputs[6305] = ~(inputs[622]);
    assign layer0_outputs[6306] = ~((inputs[974]) & (inputs[515]));
    assign layer0_outputs[6307] = (inputs[383]) & ~(inputs[1005]);
    assign layer0_outputs[6308] = ~(inputs[537]) | (inputs[886]);
    assign layer0_outputs[6309] = inputs[428];
    assign layer0_outputs[6310] = inputs[776];
    assign layer0_outputs[6311] = ~(inputs[63]) | (inputs[262]);
    assign layer0_outputs[6312] = ~((inputs[204]) ^ (inputs[629]));
    assign layer0_outputs[6313] = ~((inputs[379]) ^ (inputs[397]));
    assign layer0_outputs[6314] = ~(inputs[91]) | (inputs[63]);
    assign layer0_outputs[6315] = ~(inputs[588]);
    assign layer0_outputs[6316] = ~(inputs[114]) | (inputs[479]);
    assign layer0_outputs[6317] = (inputs[61]) & (inputs[607]);
    assign layer0_outputs[6318] = ~((inputs[714]) | (inputs[173]));
    assign layer0_outputs[6319] = (inputs[906]) | (inputs[306]);
    assign layer0_outputs[6320] = inputs[93];
    assign layer0_outputs[6321] = ~((inputs[882]) ^ (inputs[78]));
    assign layer0_outputs[6322] = ~((inputs[37]) & (inputs[61]));
    assign layer0_outputs[6323] = ~(inputs[948]) | (inputs[88]);
    assign layer0_outputs[6324] = ~(inputs[68]) | (inputs[735]);
    assign layer0_outputs[6325] = ~(inputs[724]);
    assign layer0_outputs[6326] = (inputs[53]) & ~(inputs[947]);
    assign layer0_outputs[6327] = (inputs[840]) & ~(inputs[21]);
    assign layer0_outputs[6328] = ~(inputs[235]) | (inputs[758]);
    assign layer0_outputs[6329] = inputs[132];
    assign layer0_outputs[6330] = ~((inputs[752]) ^ (inputs[800]));
    assign layer0_outputs[6331] = (inputs[599]) | (inputs[131]);
    assign layer0_outputs[6332] = (inputs[773]) | (inputs[196]);
    assign layer0_outputs[6333] = inputs[11];
    assign layer0_outputs[6334] = inputs[582];
    assign layer0_outputs[6335] = inputs[953];
    assign layer0_outputs[6336] = ~((inputs[634]) ^ (inputs[448]));
    assign layer0_outputs[6337] = ~(inputs[476]) | (inputs[471]);
    assign layer0_outputs[6338] = ~(inputs[917]);
    assign layer0_outputs[6339] = (inputs[227]) | (inputs[257]);
    assign layer0_outputs[6340] = ~(inputs[832]);
    assign layer0_outputs[6341] = ~((inputs[311]) ^ (inputs[631]));
    assign layer0_outputs[6342] = ~(inputs[443]);
    assign layer0_outputs[6343] = 1'b0;
    assign layer0_outputs[6344] = ~((inputs[207]) | (inputs[862]));
    assign layer0_outputs[6345] = ~((inputs[239]) | (inputs[443]));
    assign layer0_outputs[6346] = (inputs[427]) | (inputs[155]);
    assign layer0_outputs[6347] = (inputs[945]) & ~(inputs[147]);
    assign layer0_outputs[6348] = (inputs[829]) & ~(inputs[42]);
    assign layer0_outputs[6349] = inputs[467];
    assign layer0_outputs[6350] = ~((inputs[526]) ^ (inputs[95]));
    assign layer0_outputs[6351] = inputs[694];
    assign layer0_outputs[6352] = ~(inputs[642]) | (inputs[824]);
    assign layer0_outputs[6353] = ~(inputs[725]);
    assign layer0_outputs[6354] = (inputs[6]) ^ (inputs[88]);
    assign layer0_outputs[6355] = inputs[146];
    assign layer0_outputs[6356] = ~(inputs[696]);
    assign layer0_outputs[6357] = (inputs[420]) | (inputs[943]);
    assign layer0_outputs[6358] = (inputs[394]) | (inputs[249]);
    assign layer0_outputs[6359] = ~(inputs[900]);
    assign layer0_outputs[6360] = (inputs[902]) ^ (inputs[771]);
    assign layer0_outputs[6361] = ~((inputs[238]) ^ (inputs[219]));
    assign layer0_outputs[6362] = (inputs[244]) & ~(inputs[466]);
    assign layer0_outputs[6363] = (inputs[573]) | (inputs[407]);
    assign layer0_outputs[6364] = ~(inputs[377]) | (inputs[61]);
    assign layer0_outputs[6365] = (inputs[591]) | (inputs[421]);
    assign layer0_outputs[6366] = inputs[877];
    assign layer0_outputs[6367] = (inputs[291]) | (inputs[729]);
    assign layer0_outputs[6368] = ~((inputs[359]) ^ (inputs[741]));
    assign layer0_outputs[6369] = ~((inputs[408]) ^ (inputs[723]));
    assign layer0_outputs[6370] = ~(inputs[314]);
    assign layer0_outputs[6371] = (inputs[409]) & (inputs[516]);
    assign layer0_outputs[6372] = ~((inputs[437]) & (inputs[248]));
    assign layer0_outputs[6373] = 1'b0;
    assign layer0_outputs[6374] = ~((inputs[855]) | (inputs[875]));
    assign layer0_outputs[6375] = ~((inputs[758]) ^ (inputs[490]));
    assign layer0_outputs[6376] = ~(inputs[168]);
    assign layer0_outputs[6377] = ~(inputs[382]) | (inputs[790]);
    assign layer0_outputs[6378] = ~(inputs[220]);
    assign layer0_outputs[6379] = (inputs[569]) ^ (inputs[336]);
    assign layer0_outputs[6380] = (inputs[151]) ^ (inputs[523]);
    assign layer0_outputs[6381] = inputs[944];
    assign layer0_outputs[6382] = (inputs[699]) & ~(inputs[903]);
    assign layer0_outputs[6383] = ~((inputs[790]) ^ (inputs[210]));
    assign layer0_outputs[6384] = inputs[431];
    assign layer0_outputs[6385] = ~(inputs[725]) | (inputs[349]);
    assign layer0_outputs[6386] = inputs[740];
    assign layer0_outputs[6387] = ~((inputs[607]) | (inputs[501]));
    assign layer0_outputs[6388] = inputs[913];
    assign layer0_outputs[6389] = (inputs[470]) & ~(inputs[539]);
    assign layer0_outputs[6390] = inputs[457];
    assign layer0_outputs[6391] = (inputs[965]) & ~(inputs[13]);
    assign layer0_outputs[6392] = ~((inputs[665]) & (inputs[542]));
    assign layer0_outputs[6393] = ~(inputs[305]);
    assign layer0_outputs[6394] = (inputs[964]) & ~(inputs[1000]);
    assign layer0_outputs[6395] = 1'b0;
    assign layer0_outputs[6396] = inputs[555];
    assign layer0_outputs[6397] = (inputs[990]) | (inputs[475]);
    assign layer0_outputs[6398] = ~(inputs[658]);
    assign layer0_outputs[6399] = ~((inputs[989]) & (inputs[567]));
    assign layer0_outputs[6400] = (inputs[218]) ^ (inputs[608]);
    assign layer0_outputs[6401] = (inputs[248]) | (inputs[894]);
    assign layer0_outputs[6402] = (inputs[38]) ^ (inputs[285]);
    assign layer0_outputs[6403] = ~((inputs[992]) ^ (inputs[331]));
    assign layer0_outputs[6404] = (inputs[26]) & (inputs[298]);
    assign layer0_outputs[6405] = ~(inputs[995]) | (inputs[961]);
    assign layer0_outputs[6406] = (inputs[409]) | (inputs[884]);
    assign layer0_outputs[6407] = (inputs[210]) | (inputs[1011]);
    assign layer0_outputs[6408] = ~(inputs[422]) | (inputs[612]);
    assign layer0_outputs[6409] = ~(inputs[290]) | (inputs[556]);
    assign layer0_outputs[6410] = inputs[866];
    assign layer0_outputs[6411] = inputs[646];
    assign layer0_outputs[6412] = 1'b1;
    assign layer0_outputs[6413] = 1'b1;
    assign layer0_outputs[6414] = inputs[907];
    assign layer0_outputs[6415] = 1'b1;
    assign layer0_outputs[6416] = inputs[879];
    assign layer0_outputs[6417] = inputs[979];
    assign layer0_outputs[6418] = ~(inputs[683]) | (inputs[803]);
    assign layer0_outputs[6419] = ~((inputs[306]) | (inputs[341]));
    assign layer0_outputs[6420] = inputs[831];
    assign layer0_outputs[6421] = inputs[178];
    assign layer0_outputs[6422] = (inputs[903]) & ~(inputs[18]);
    assign layer0_outputs[6423] = ~(inputs[487]);
    assign layer0_outputs[6424] = inputs[293];
    assign layer0_outputs[6425] = (inputs[376]) | (inputs[486]);
    assign layer0_outputs[6426] = ~(inputs[464]);
    assign layer0_outputs[6427] = ~((inputs[164]) | (inputs[288]));
    assign layer0_outputs[6428] = ~((inputs[124]) ^ (inputs[759]));
    assign layer0_outputs[6429] = 1'b1;
    assign layer0_outputs[6430] = (inputs[199]) & ~(inputs[358]);
    assign layer0_outputs[6431] = ~(inputs[756]);
    assign layer0_outputs[6432] = ~((inputs[515]) | (inputs[263]));
    assign layer0_outputs[6433] = (inputs[236]) & (inputs[446]);
    assign layer0_outputs[6434] = (inputs[974]) & ~(inputs[135]);
    assign layer0_outputs[6435] = inputs[848];
    assign layer0_outputs[6436] = ~(inputs[163]) | (inputs[328]);
    assign layer0_outputs[6437] = (inputs[485]) | (inputs[289]);
    assign layer0_outputs[6438] = ~(inputs[674]) | (inputs[964]);
    assign layer0_outputs[6439] = ~(inputs[904]) | (inputs[638]);
    assign layer0_outputs[6440] = ~((inputs[766]) | (inputs[620]));
    assign layer0_outputs[6441] = ~(inputs[185]) | (inputs[894]);
    assign layer0_outputs[6442] = inputs[315];
    assign layer0_outputs[6443] = inputs[154];
    assign layer0_outputs[6444] = inputs[360];
    assign layer0_outputs[6445] = ~(inputs[836]);
    assign layer0_outputs[6446] = (inputs[885]) & (inputs[885]);
    assign layer0_outputs[6447] = ~(inputs[59]);
    assign layer0_outputs[6448] = 1'b0;
    assign layer0_outputs[6449] = (inputs[984]) & ~(inputs[895]);
    assign layer0_outputs[6450] = ~((inputs[967]) | (inputs[720]));
    assign layer0_outputs[6451] = (inputs[503]) | (inputs[802]);
    assign layer0_outputs[6452] = inputs[42];
    assign layer0_outputs[6453] = (inputs[635]) & (inputs[929]);
    assign layer0_outputs[6454] = ~((inputs[135]) & (inputs[476]));
    assign layer0_outputs[6455] = (inputs[403]) | (inputs[614]);
    assign layer0_outputs[6456] = ~(inputs[756]);
    assign layer0_outputs[6457] = ~(inputs[571]);
    assign layer0_outputs[6458] = ~(inputs[436]);
    assign layer0_outputs[6459] = inputs[473];
    assign layer0_outputs[6460] = 1'b1;
    assign layer0_outputs[6461] = inputs[818];
    assign layer0_outputs[6462] = ~(inputs[693]) | (inputs[895]);
    assign layer0_outputs[6463] = inputs[587];
    assign layer0_outputs[6464] = ~(inputs[680]) | (inputs[921]);
    assign layer0_outputs[6465] = (inputs[616]) & ~(inputs[379]);
    assign layer0_outputs[6466] = ~(inputs[748]);
    assign layer0_outputs[6467] = ~(inputs[521]);
    assign layer0_outputs[6468] = ~((inputs[396]) ^ (inputs[728]));
    assign layer0_outputs[6469] = inputs[850];
    assign layer0_outputs[6470] = ~(inputs[142]);
    assign layer0_outputs[6471] = 1'b1;
    assign layer0_outputs[6472] = 1'b0;
    assign layer0_outputs[6473] = ~((inputs[474]) ^ (inputs[119]));
    assign layer0_outputs[6474] = (inputs[732]) & ~(inputs[179]);
    assign layer0_outputs[6475] = ~(inputs[485]);
    assign layer0_outputs[6476] = (inputs[465]) ^ (inputs[153]);
    assign layer0_outputs[6477] = ~((inputs[1005]) | (inputs[683]));
    assign layer0_outputs[6478] = (inputs[369]) ^ (inputs[319]);
    assign layer0_outputs[6479] = (inputs[333]) ^ (inputs[52]);
    assign layer0_outputs[6480] = ~((inputs[799]) | (inputs[825]));
    assign layer0_outputs[6481] = inputs[463];
    assign layer0_outputs[6482] = (inputs[485]) | (inputs[887]);
    assign layer0_outputs[6483] = inputs[715];
    assign layer0_outputs[6484] = (inputs[680]) ^ (inputs[332]);
    assign layer0_outputs[6485] = (inputs[434]) & ~(inputs[441]);
    assign layer0_outputs[6486] = (inputs[29]) | (inputs[723]);
    assign layer0_outputs[6487] = ~((inputs[30]) ^ (inputs[837]));
    assign layer0_outputs[6488] = inputs[849];
    assign layer0_outputs[6489] = 1'b1;
    assign layer0_outputs[6490] = (inputs[533]) ^ (inputs[179]);
    assign layer0_outputs[6491] = inputs[113];
    assign layer0_outputs[6492] = ~((inputs[633]) | (inputs[320]));
    assign layer0_outputs[6493] = ~(inputs[687]) | (inputs[356]);
    assign layer0_outputs[6494] = ~((inputs[938]) | (inputs[914]));
    assign layer0_outputs[6495] = ~(inputs[0]) | (inputs[783]);
    assign layer0_outputs[6496] = ~((inputs[879]) | (inputs[267]));
    assign layer0_outputs[6497] = ~((inputs[851]) | (inputs[554]));
    assign layer0_outputs[6498] = (inputs[714]) & ~(inputs[1008]);
    assign layer0_outputs[6499] = (inputs[791]) | (inputs[824]);
    assign layer0_outputs[6500] = ~((inputs[199]) | (inputs[200]));
    assign layer0_outputs[6501] = (inputs[637]) | (inputs[20]);
    assign layer0_outputs[6502] = ~((inputs[400]) ^ (inputs[66]));
    assign layer0_outputs[6503] = ~((inputs[579]) ^ (inputs[690]));
    assign layer0_outputs[6504] = ~(inputs[885]) | (inputs[895]);
    assign layer0_outputs[6505] = ~((inputs[57]) | (inputs[531]));
    assign layer0_outputs[6506] = ~(inputs[533]);
    assign layer0_outputs[6507] = ~(inputs[804]) | (inputs[873]);
    assign layer0_outputs[6508] = ~(inputs[593]) | (inputs[891]);
    assign layer0_outputs[6509] = (inputs[406]) | (inputs[505]);
    assign layer0_outputs[6510] = ~(inputs[78]);
    assign layer0_outputs[6511] = (inputs[161]) ^ (inputs[144]);
    assign layer0_outputs[6512] = ~((inputs[680]) ^ (inputs[694]));
    assign layer0_outputs[6513] = ~(inputs[3]);
    assign layer0_outputs[6514] = ~(inputs[445]) | (inputs[674]);
    assign layer0_outputs[6515] = ~((inputs[972]) | (inputs[216]));
    assign layer0_outputs[6516] = ~(inputs[861]) | (inputs[270]);
    assign layer0_outputs[6517] = ~(inputs[634]) | (inputs[484]);
    assign layer0_outputs[6518] = ~((inputs[846]) ^ (inputs[227]));
    assign layer0_outputs[6519] = ~(inputs[481]) | (inputs[559]);
    assign layer0_outputs[6520] = 1'b1;
    assign layer0_outputs[6521] = (inputs[522]) | (inputs[223]);
    assign layer0_outputs[6522] = (inputs[553]) & ~(inputs[803]);
    assign layer0_outputs[6523] = ~(inputs[245]) | (inputs[921]);
    assign layer0_outputs[6524] = (inputs[395]) & ~(inputs[515]);
    assign layer0_outputs[6525] = ~(inputs[957]);
    assign layer0_outputs[6526] = (inputs[440]) | (inputs[349]);
    assign layer0_outputs[6527] = ~((inputs[99]) | (inputs[164]));
    assign layer0_outputs[6528] = inputs[881];
    assign layer0_outputs[6529] = (inputs[764]) ^ (inputs[688]);
    assign layer0_outputs[6530] = inputs[334];
    assign layer0_outputs[6531] = (inputs[677]) ^ (inputs[499]);
    assign layer0_outputs[6532] = (inputs[64]) ^ (inputs[843]);
    assign layer0_outputs[6533] = inputs[654];
    assign layer0_outputs[6534] = inputs[850];
    assign layer0_outputs[6535] = (inputs[351]) & (inputs[962]);
    assign layer0_outputs[6536] = (inputs[1002]) ^ (inputs[647]);
    assign layer0_outputs[6537] = ~((inputs[1015]) ^ (inputs[691]));
    assign layer0_outputs[6538] = ~(inputs[658]) | (inputs[378]);
    assign layer0_outputs[6539] = (inputs[258]) & ~(inputs[24]);
    assign layer0_outputs[6540] = ~(inputs[719]) | (inputs[315]);
    assign layer0_outputs[6541] = inputs[864];
    assign layer0_outputs[6542] = (inputs[854]) & ~(inputs[701]);
    assign layer0_outputs[6543] = ~((inputs[830]) ^ (inputs[881]));
    assign layer0_outputs[6544] = inputs[70];
    assign layer0_outputs[6545] = (inputs[371]) | (inputs[888]);
    assign layer0_outputs[6546] = (inputs[676]) & (inputs[14]);
    assign layer0_outputs[6547] = (inputs[590]) | (inputs[204]);
    assign layer0_outputs[6548] = (inputs[873]) | (inputs[570]);
    assign layer0_outputs[6549] = ~((inputs[747]) ^ (inputs[198]));
    assign layer0_outputs[6550] = ~((inputs[138]) | (inputs[875]));
    assign layer0_outputs[6551] = ~((inputs[887]) | (inputs[189]));
    assign layer0_outputs[6552] = (inputs[409]) | (inputs[174]);
    assign layer0_outputs[6553] = (inputs[820]) | (inputs[827]);
    assign layer0_outputs[6554] = ~(inputs[495]);
    assign layer0_outputs[6555] = (inputs[841]) & ~(inputs[193]);
    assign layer0_outputs[6556] = ~((inputs[502]) & (inputs[658]));
    assign layer0_outputs[6557] = (inputs[328]) ^ (inputs[552]);
    assign layer0_outputs[6558] = 1'b1;
    assign layer0_outputs[6559] = ~(inputs[902]) | (inputs[199]);
    assign layer0_outputs[6560] = (inputs[70]) & (inputs[639]);
    assign layer0_outputs[6561] = (inputs[275]) & ~(inputs[60]);
    assign layer0_outputs[6562] = ~(inputs[622]);
    assign layer0_outputs[6563] = ~(inputs[831]);
    assign layer0_outputs[6564] = ~(inputs[325]);
    assign layer0_outputs[6565] = (inputs[884]) & ~(inputs[874]);
    assign layer0_outputs[6566] = (inputs[818]) & ~(inputs[944]);
    assign layer0_outputs[6567] = ~(inputs[813]) | (inputs[127]);
    assign layer0_outputs[6568] = (inputs[810]) & ~(inputs[26]);
    assign layer0_outputs[6569] = (inputs[118]) & (inputs[35]);
    assign layer0_outputs[6570] = ~(inputs[1014]);
    assign layer0_outputs[6571] = ~((inputs[99]) ^ (inputs[993]));
    assign layer0_outputs[6572] = inputs[563];
    assign layer0_outputs[6573] = ~((inputs[905]) | (inputs[954]));
    assign layer0_outputs[6574] = ~(inputs[263]) | (inputs[46]);
    assign layer0_outputs[6575] = ~(inputs[127]) | (inputs[357]);
    assign layer0_outputs[6576] = (inputs[914]) ^ (inputs[1020]);
    assign layer0_outputs[6577] = ~(inputs[928]) | (inputs[734]);
    assign layer0_outputs[6578] = ~((inputs[171]) ^ (inputs[606]));
    assign layer0_outputs[6579] = (inputs[396]) | (inputs[564]);
    assign layer0_outputs[6580] = ~((inputs[1005]) | (inputs[361]));
    assign layer0_outputs[6581] = ~((inputs[827]) | (inputs[942]));
    assign layer0_outputs[6582] = ~(inputs[203]) | (inputs[323]);
    assign layer0_outputs[6583] = ~(inputs[424]);
    assign layer0_outputs[6584] = ~((inputs[890]) & (inputs[4]));
    assign layer0_outputs[6585] = (inputs[790]) & ~(inputs[719]);
    assign layer0_outputs[6586] = (inputs[760]) | (inputs[6]);
    assign layer0_outputs[6587] = ~((inputs[630]) | (inputs[9]));
    assign layer0_outputs[6588] = ~(inputs[388]) | (inputs[325]);
    assign layer0_outputs[6589] = inputs[927];
    assign layer0_outputs[6590] = ~(inputs[781]);
    assign layer0_outputs[6591] = (inputs[420]) & ~(inputs[862]);
    assign layer0_outputs[6592] = ~((inputs[696]) | (inputs[292]));
    assign layer0_outputs[6593] = 1'b0;
    assign layer0_outputs[6594] = 1'b1;
    assign layer0_outputs[6595] = ~((inputs[237]) ^ (inputs[807]));
    assign layer0_outputs[6596] = ~((inputs[723]) | (inputs[699]));
    assign layer0_outputs[6597] = ~((inputs[599]) & (inputs[617]));
    assign layer0_outputs[6598] = (inputs[676]) & ~(inputs[210]);
    assign layer0_outputs[6599] = ~((inputs[697]) | (inputs[305]));
    assign layer0_outputs[6600] = 1'b1;
    assign layer0_outputs[6601] = ~((inputs[960]) & (inputs[951]));
    assign layer0_outputs[6602] = (inputs[835]) ^ (inputs[586]);
    assign layer0_outputs[6603] = inputs[206];
    assign layer0_outputs[6604] = ~(inputs[583]);
    assign layer0_outputs[6605] = (inputs[63]) | (inputs[145]);
    assign layer0_outputs[6606] = (inputs[421]) | (inputs[880]);
    assign layer0_outputs[6607] = inputs[650];
    assign layer0_outputs[6608] = (inputs[771]) & (inputs[615]);
    assign layer0_outputs[6609] = ~((inputs[288]) | (inputs[52]));
    assign layer0_outputs[6610] = ~((inputs[583]) | (inputs[8]));
    assign layer0_outputs[6611] = ~((inputs[289]) & (inputs[400]));
    assign layer0_outputs[6612] = (inputs[571]) & ~(inputs[961]);
    assign layer0_outputs[6613] = (inputs[769]) ^ (inputs[766]);
    assign layer0_outputs[6614] = inputs[1012];
    assign layer0_outputs[6615] = (inputs[634]) & ~(inputs[967]);
    assign layer0_outputs[6616] = inputs[223];
    assign layer0_outputs[6617] = inputs[739];
    assign layer0_outputs[6618] = ~(inputs[457]);
    assign layer0_outputs[6619] = (inputs[559]) & ~(inputs[219]);
    assign layer0_outputs[6620] = (inputs[129]) & ~(inputs[867]);
    assign layer0_outputs[6621] = ~((inputs[215]) ^ (inputs[481]));
    assign layer0_outputs[6622] = ~(inputs[551]) | (inputs[741]);
    assign layer0_outputs[6623] = (inputs[498]) & ~(inputs[744]);
    assign layer0_outputs[6624] = (inputs[736]) | (inputs[850]);
    assign layer0_outputs[6625] = (inputs[564]) | (inputs[463]);
    assign layer0_outputs[6626] = inputs[905];
    assign layer0_outputs[6627] = ~((inputs[276]) ^ (inputs[881]));
    assign layer0_outputs[6628] = inputs[330];
    assign layer0_outputs[6629] = ~(inputs[339]) | (inputs[181]);
    assign layer0_outputs[6630] = (inputs[681]) & ~(inputs[952]);
    assign layer0_outputs[6631] = ~((inputs[366]) ^ (inputs[459]));
    assign layer0_outputs[6632] = ~((inputs[6]) | (inputs[241]));
    assign layer0_outputs[6633] = ~(inputs[744]) | (inputs[944]);
    assign layer0_outputs[6634] = (inputs[755]) & ~(inputs[701]);
    assign layer0_outputs[6635] = ~(inputs[212]);
    assign layer0_outputs[6636] = (inputs[713]) & ~(inputs[951]);
    assign layer0_outputs[6637] = (inputs[67]) & (inputs[865]);
    assign layer0_outputs[6638] = 1'b1;
    assign layer0_outputs[6639] = ~(inputs[562]) | (inputs[234]);
    assign layer0_outputs[6640] = (inputs[337]) ^ (inputs[710]);
    assign layer0_outputs[6641] = ~(inputs[6]);
    assign layer0_outputs[6642] = (inputs[996]) ^ (inputs[314]);
    assign layer0_outputs[6643] = ~((inputs[646]) | (inputs[310]));
    assign layer0_outputs[6644] = ~(inputs[614]);
    assign layer0_outputs[6645] = ~(inputs[870]);
    assign layer0_outputs[6646] = ~((inputs[295]) ^ (inputs[603]));
    assign layer0_outputs[6647] = ~(inputs[496]);
    assign layer0_outputs[6648] = (inputs[496]) | (inputs[350]);
    assign layer0_outputs[6649] = (inputs[180]) & ~(inputs[508]);
    assign layer0_outputs[6650] = ~((inputs[908]) | (inputs[246]));
    assign layer0_outputs[6651] = (inputs[877]) ^ (inputs[869]);
    assign layer0_outputs[6652] = inputs[506];
    assign layer0_outputs[6653] = (inputs[738]) | (inputs[39]);
    assign layer0_outputs[6654] = inputs[942];
    assign layer0_outputs[6655] = ~(inputs[955]) | (inputs[736]);
    assign layer0_outputs[6656] = ~(inputs[392]) | (inputs[105]);
    assign layer0_outputs[6657] = ~((inputs[309]) | (inputs[535]));
    assign layer0_outputs[6658] = ~((inputs[489]) | (inputs[518]));
    assign layer0_outputs[6659] = ~((inputs[352]) ^ (inputs[765]));
    assign layer0_outputs[6660] = ~(inputs[396]);
    assign layer0_outputs[6661] = 1'b1;
    assign layer0_outputs[6662] = inputs[619];
    assign layer0_outputs[6663] = ~((inputs[312]) | (inputs[937]));
    assign layer0_outputs[6664] = inputs[395];
    assign layer0_outputs[6665] = ~(inputs[515]) | (inputs[485]);
    assign layer0_outputs[6666] = ~(inputs[496]) | (inputs[930]);
    assign layer0_outputs[6667] = ~(inputs[782]) | (inputs[836]);
    assign layer0_outputs[6668] = inputs[748];
    assign layer0_outputs[6669] = ~((inputs[739]) ^ (inputs[42]));
    assign layer0_outputs[6670] = ~(inputs[744]);
    assign layer0_outputs[6671] = ~(inputs[176]) | (inputs[65]);
    assign layer0_outputs[6672] = ~((inputs[677]) | (inputs[59]));
    assign layer0_outputs[6673] = (inputs[235]) | (inputs[323]);
    assign layer0_outputs[6674] = ~((inputs[131]) ^ (inputs[571]));
    assign layer0_outputs[6675] = (inputs[600]) & ~(inputs[329]);
    assign layer0_outputs[6676] = ~(inputs[844]) | (inputs[976]);
    assign layer0_outputs[6677] = ~(inputs[556]);
    assign layer0_outputs[6678] = ~(inputs[715]);
    assign layer0_outputs[6679] = ~((inputs[868]) | (inputs[610]));
    assign layer0_outputs[6680] = ~(inputs[64]);
    assign layer0_outputs[6681] = inputs[331];
    assign layer0_outputs[6682] = ~(inputs[727]);
    assign layer0_outputs[6683] = ~(inputs[18]) | (inputs[584]);
    assign layer0_outputs[6684] = inputs[892];
    assign layer0_outputs[6685] = ~(inputs[586]) | (inputs[858]);
    assign layer0_outputs[6686] = (inputs[682]) & ~(inputs[511]);
    assign layer0_outputs[6687] = ~((inputs[329]) | (inputs[1009]));
    assign layer0_outputs[6688] = ~((inputs[734]) ^ (inputs[528]));
    assign layer0_outputs[6689] = (inputs[773]) & ~(inputs[937]);
    assign layer0_outputs[6690] = ~((inputs[355]) ^ (inputs[401]));
    assign layer0_outputs[6691] = (inputs[839]) & (inputs[34]);
    assign layer0_outputs[6692] = ~(inputs[455]) | (inputs[932]);
    assign layer0_outputs[6693] = (inputs[826]) | (inputs[460]);
    assign layer0_outputs[6694] = inputs[811];
    assign layer0_outputs[6695] = ~(inputs[437]);
    assign layer0_outputs[6696] = inputs[238];
    assign layer0_outputs[6697] = ~(inputs[731]);
    assign layer0_outputs[6698] = ~((inputs[442]) | (inputs[843]));
    assign layer0_outputs[6699] = inputs[744];
    assign layer0_outputs[6700] = inputs[188];
    assign layer0_outputs[6701] = (inputs[281]) | (inputs[912]);
    assign layer0_outputs[6702] = 1'b1;
    assign layer0_outputs[6703] = ~((inputs[841]) | (inputs[227]));
    assign layer0_outputs[6704] = ~(inputs[651]);
    assign layer0_outputs[6705] = inputs[932];
    assign layer0_outputs[6706] = (inputs[162]) & (inputs[625]);
    assign layer0_outputs[6707] = ~((inputs[73]) ^ (inputs[399]));
    assign layer0_outputs[6708] = (inputs[733]) & ~(inputs[916]);
    assign layer0_outputs[6709] = ~((inputs[703]) | (inputs[749]));
    assign layer0_outputs[6710] = (inputs[763]) | (inputs[321]);
    assign layer0_outputs[6711] = (inputs[859]) & ~(inputs[149]);
    assign layer0_outputs[6712] = ~((inputs[717]) | (inputs[966]));
    assign layer0_outputs[6713] = 1'b1;
    assign layer0_outputs[6714] = (inputs[745]) & ~(inputs[589]);
    assign layer0_outputs[6715] = ~((inputs[435]) & (inputs[788]));
    assign layer0_outputs[6716] = ~((inputs[970]) | (inputs[294]));
    assign layer0_outputs[6717] = inputs[133];
    assign layer0_outputs[6718] = ~(inputs[93]) | (inputs[123]);
    assign layer0_outputs[6719] = ~(inputs[202]);
    assign layer0_outputs[6720] = ~((inputs[105]) | (inputs[135]));
    assign layer0_outputs[6721] = (inputs[452]) | (inputs[150]);
    assign layer0_outputs[6722] = 1'b0;
    assign layer0_outputs[6723] = ~(inputs[756]) | (inputs[342]);
    assign layer0_outputs[6724] = (inputs[123]) | (inputs[189]);
    assign layer0_outputs[6725] = (inputs[899]) & ~(inputs[738]);
    assign layer0_outputs[6726] = inputs[622];
    assign layer0_outputs[6727] = (inputs[697]) | (inputs[893]);
    assign layer0_outputs[6728] = ~((inputs[509]) | (inputs[888]));
    assign layer0_outputs[6729] = ~(inputs[932]) | (inputs[263]);
    assign layer0_outputs[6730] = ~((inputs[474]) | (inputs[307]));
    assign layer0_outputs[6731] = (inputs[244]) & ~(inputs[930]);
    assign layer0_outputs[6732] = ~((inputs[762]) | (inputs[884]));
    assign layer0_outputs[6733] = (inputs[276]) & ~(inputs[99]);
    assign layer0_outputs[6734] = (inputs[293]) ^ (inputs[679]);
    assign layer0_outputs[6735] = (inputs[330]) & ~(inputs[145]);
    assign layer0_outputs[6736] = ~(inputs[462]) | (inputs[1009]);
    assign layer0_outputs[6737] = (inputs[49]) & ~(inputs[139]);
    assign layer0_outputs[6738] = 1'b0;
    assign layer0_outputs[6739] = inputs[521];
    assign layer0_outputs[6740] = ~((inputs[382]) ^ (inputs[55]));
    assign layer0_outputs[6741] = (inputs[290]) | (inputs[647]);
    assign layer0_outputs[6742] = ~((inputs[116]) | (inputs[341]));
    assign layer0_outputs[6743] = ~(inputs[323]);
    assign layer0_outputs[6744] = inputs[890];
    assign layer0_outputs[6745] = ~(inputs[495]);
    assign layer0_outputs[6746] = ~((inputs[39]) ^ (inputs[503]));
    assign layer0_outputs[6747] = (inputs[543]) ^ (inputs[346]);
    assign layer0_outputs[6748] = inputs[576];
    assign layer0_outputs[6749] = ~(inputs[854]);
    assign layer0_outputs[6750] = (inputs[113]) & ~(inputs[83]);
    assign layer0_outputs[6751] = (inputs[408]) | (inputs[886]);
    assign layer0_outputs[6752] = 1'b1;
    assign layer0_outputs[6753] = (inputs[270]) | (inputs[455]);
    assign layer0_outputs[6754] = ~((inputs[690]) | (inputs[867]));
    assign layer0_outputs[6755] = ~(inputs[29]) | (inputs[122]);
    assign layer0_outputs[6756] = inputs[281];
    assign layer0_outputs[6757] = (inputs[432]) ^ (inputs[640]);
    assign layer0_outputs[6758] = ~((inputs[517]) ^ (inputs[465]));
    assign layer0_outputs[6759] = ~(inputs[524]);
    assign layer0_outputs[6760] = (inputs[248]) ^ (inputs[482]);
    assign layer0_outputs[6761] = ~((inputs[488]) ^ (inputs[666]));
    assign layer0_outputs[6762] = (inputs[558]) & (inputs[1016]);
    assign layer0_outputs[6763] = ~((inputs[636]) ^ (inputs[964]));
    assign layer0_outputs[6764] = ~((inputs[197]) ^ (inputs[684]));
    assign layer0_outputs[6765] = (inputs[530]) & (inputs[242]);
    assign layer0_outputs[6766] = (inputs[178]) | (inputs[625]);
    assign layer0_outputs[6767] = (inputs[14]) | (inputs[377]);
    assign layer0_outputs[6768] = (inputs[896]) ^ (inputs[258]);
    assign layer0_outputs[6769] = ~(inputs[688]) | (inputs[423]);
    assign layer0_outputs[6770] = ~(inputs[374]) | (inputs[995]);
    assign layer0_outputs[6771] = (inputs[498]) & ~(inputs[219]);
    assign layer0_outputs[6772] = ~((inputs[110]) | (inputs[681]));
    assign layer0_outputs[6773] = ~((inputs[254]) & (inputs[387]));
    assign layer0_outputs[6774] = ~(inputs[166]) | (inputs[785]);
    assign layer0_outputs[6775] = ~(inputs[817]) | (inputs[892]);
    assign layer0_outputs[6776] = (inputs[757]) | (inputs[152]);
    assign layer0_outputs[6777] = (inputs[592]) & ~(inputs[1005]);
    assign layer0_outputs[6778] = ~((inputs[677]) | (inputs[808]));
    assign layer0_outputs[6779] = inputs[407];
    assign layer0_outputs[6780] = inputs[411];
    assign layer0_outputs[6781] = ~((inputs[1007]) | (inputs[621]));
    assign layer0_outputs[6782] = ~((inputs[642]) | (inputs[742]));
    assign layer0_outputs[6783] = ~((inputs[648]) | (inputs[597]));
    assign layer0_outputs[6784] = ~((inputs[606]) ^ (inputs[585]));
    assign layer0_outputs[6785] = ~((inputs[714]) | (inputs[118]));
    assign layer0_outputs[6786] = (inputs[128]) ^ (inputs[747]);
    assign layer0_outputs[6787] = ~((inputs[461]) | (inputs[148]));
    assign layer0_outputs[6788] = (inputs[125]) ^ (inputs[464]);
    assign layer0_outputs[6789] = ~((inputs[231]) ^ (inputs[944]));
    assign layer0_outputs[6790] = inputs[844];
    assign layer0_outputs[6791] = ~((inputs[365]) | (inputs[304]));
    assign layer0_outputs[6792] = ~((inputs[32]) ^ (inputs[748]));
    assign layer0_outputs[6793] = (inputs[305]) & ~(inputs[609]);
    assign layer0_outputs[6794] = inputs[374];
    assign layer0_outputs[6795] = inputs[137];
    assign layer0_outputs[6796] = inputs[291];
    assign layer0_outputs[6797] = ~((inputs[137]) & (inputs[541]));
    assign layer0_outputs[6798] = ~(inputs[810]);
    assign layer0_outputs[6799] = ~(inputs[655]) | (inputs[8]);
    assign layer0_outputs[6800] = ~(inputs[510]);
    assign layer0_outputs[6801] = (inputs[306]) | (inputs[277]);
    assign layer0_outputs[6802] = (inputs[933]) | (inputs[302]);
    assign layer0_outputs[6803] = inputs[252];
    assign layer0_outputs[6804] = (inputs[928]) | (inputs[852]);
    assign layer0_outputs[6805] = ~((inputs[954]) ^ (inputs[196]));
    assign layer0_outputs[6806] = ~((inputs[926]) | (inputs[381]));
    assign layer0_outputs[6807] = ~(inputs[522]);
    assign layer0_outputs[6808] = (inputs[647]) | (inputs[355]);
    assign layer0_outputs[6809] = ~(inputs[98]);
    assign layer0_outputs[6810] = ~(inputs[225]) | (inputs[226]);
    assign layer0_outputs[6811] = (inputs[790]) & ~(inputs[485]);
    assign layer0_outputs[6812] = ~((inputs[635]) ^ (inputs[307]));
    assign layer0_outputs[6813] = (inputs[534]) & ~(inputs[423]);
    assign layer0_outputs[6814] = ~(inputs[877]);
    assign layer0_outputs[6815] = ~(inputs[201]);
    assign layer0_outputs[6816] = 1'b0;
    assign layer0_outputs[6817] = ~(inputs[893]) | (inputs[119]);
    assign layer0_outputs[6818] = ~(inputs[213]) | (inputs[61]);
    assign layer0_outputs[6819] = inputs[258];
    assign layer0_outputs[6820] = 1'b1;
    assign layer0_outputs[6821] = ~(inputs[587]) | (inputs[931]);
    assign layer0_outputs[6822] = ~((inputs[146]) | (inputs[99]));
    assign layer0_outputs[6823] = (inputs[648]) | (inputs[264]);
    assign layer0_outputs[6824] = ~(inputs[595]);
    assign layer0_outputs[6825] = (inputs[671]) & ~(inputs[343]);
    assign layer0_outputs[6826] = ~(inputs[548]) | (inputs[562]);
    assign layer0_outputs[6827] = (inputs[329]) | (inputs[332]);
    assign layer0_outputs[6828] = (inputs[654]) & ~(inputs[2]);
    assign layer0_outputs[6829] = 1'b0;
    assign layer0_outputs[6830] = (inputs[519]) & ~(inputs[575]);
    assign layer0_outputs[6831] = ~(inputs[821]);
    assign layer0_outputs[6832] = ~(inputs[987]);
    assign layer0_outputs[6833] = ~(inputs[375]) | (inputs[959]);
    assign layer0_outputs[6834] = inputs[736];
    assign layer0_outputs[6835] = ~(inputs[270]) | (inputs[421]);
    assign layer0_outputs[6836] = (inputs[962]) | (inputs[750]);
    assign layer0_outputs[6837] = ~((inputs[787]) ^ (inputs[142]));
    assign layer0_outputs[6838] = inputs[156];
    assign layer0_outputs[6839] = (inputs[846]) & ~(inputs[261]);
    assign layer0_outputs[6840] = ~((inputs[417]) ^ (inputs[48]));
    assign layer0_outputs[6841] = (inputs[703]) | (inputs[497]);
    assign layer0_outputs[6842] = ~(inputs[492]) | (inputs[204]);
    assign layer0_outputs[6843] = ~((inputs[967]) ^ (inputs[359]));
    assign layer0_outputs[6844] = ~((inputs[69]) | (inputs[45]));
    assign layer0_outputs[6845] = ~(inputs[239]);
    assign layer0_outputs[6846] = ~((inputs[682]) | (inputs[176]));
    assign layer0_outputs[6847] = inputs[462];
    assign layer0_outputs[6848] = (inputs[102]) & ~(inputs[762]);
    assign layer0_outputs[6849] = ~((inputs[480]) & (inputs[86]));
    assign layer0_outputs[6850] = ~((inputs[260]) | (inputs[678]));
    assign layer0_outputs[6851] = ~(inputs[280]) | (inputs[580]);
    assign layer0_outputs[6852] = (inputs[123]) ^ (inputs[244]);
    assign layer0_outputs[6853] = (inputs[753]) & ~(inputs[120]);
    assign layer0_outputs[6854] = ~((inputs[462]) ^ (inputs[200]));
    assign layer0_outputs[6855] = inputs[987];
    assign layer0_outputs[6856] = (inputs[785]) & ~(inputs[996]);
    assign layer0_outputs[6857] = ~(inputs[665]) | (inputs[155]);
    assign layer0_outputs[6858] = ~((inputs[795]) & (inputs[673]));
    assign layer0_outputs[6859] = inputs[333];
    assign layer0_outputs[6860] = ~(inputs[65]);
    assign layer0_outputs[6861] = inputs[588];
    assign layer0_outputs[6862] = (inputs[95]) | (inputs[520]);
    assign layer0_outputs[6863] = ~((inputs[1018]) & (inputs[553]));
    assign layer0_outputs[6864] = ~(inputs[988]) | (inputs[989]);
    assign layer0_outputs[6865] = (inputs[410]) | (inputs[261]);
    assign layer0_outputs[6866] = (inputs[419]) ^ (inputs[720]);
    assign layer0_outputs[6867] = (inputs[982]) & ~(inputs[957]);
    assign layer0_outputs[6868] = 1'b0;
    assign layer0_outputs[6869] = ~(inputs[591]) | (inputs[388]);
    assign layer0_outputs[6870] = (inputs[1021]) | (inputs[435]);
    assign layer0_outputs[6871] = (inputs[769]) ^ (inputs[576]);
    assign layer0_outputs[6872] = (inputs[264]) & ~(inputs[74]);
    assign layer0_outputs[6873] = ~((inputs[839]) | (inputs[679]));
    assign layer0_outputs[6874] = inputs[272];
    assign layer0_outputs[6875] = (inputs[71]) ^ (inputs[370]);
    assign layer0_outputs[6876] = 1'b0;
    assign layer0_outputs[6877] = (inputs[695]) & ~(inputs[401]);
    assign layer0_outputs[6878] = (inputs[628]) ^ (inputs[28]);
    assign layer0_outputs[6879] = ~(inputs[283]) | (inputs[475]);
    assign layer0_outputs[6880] = (inputs[568]) | (inputs[993]);
    assign layer0_outputs[6881] = (inputs[925]) | (inputs[551]);
    assign layer0_outputs[6882] = ~((inputs[472]) | (inputs[889]));
    assign layer0_outputs[6883] = (inputs[874]) & ~(inputs[207]);
    assign layer0_outputs[6884] = 1'b1;
    assign layer0_outputs[6885] = ~((inputs[417]) | (inputs[946]));
    assign layer0_outputs[6886] = ~(inputs[401]);
    assign layer0_outputs[6887] = (inputs[687]) | (inputs[652]);
    assign layer0_outputs[6888] = (inputs[690]) ^ (inputs[625]);
    assign layer0_outputs[6889] = (inputs[1004]) ^ (inputs[533]);
    assign layer0_outputs[6890] = (inputs[670]) & (inputs[65]);
    assign layer0_outputs[6891] = ~(inputs[315]);
    assign layer0_outputs[6892] = inputs[652];
    assign layer0_outputs[6893] = ~(inputs[489]);
    assign layer0_outputs[6894] = ~(inputs[861]) | (inputs[46]);
    assign layer0_outputs[6895] = ~(inputs[651]) | (inputs[65]);
    assign layer0_outputs[6896] = inputs[688];
    assign layer0_outputs[6897] = (inputs[556]) & ~(inputs[961]);
    assign layer0_outputs[6898] = ~((inputs[706]) ^ (inputs[34]));
    assign layer0_outputs[6899] = ~(inputs[534]);
    assign layer0_outputs[6900] = ~((inputs[38]) ^ (inputs[524]));
    assign layer0_outputs[6901] = (inputs[245]) & ~(inputs[150]);
    assign layer0_outputs[6902] = (inputs[803]) | (inputs[323]);
    assign layer0_outputs[6903] = (inputs[722]) ^ (inputs[660]);
    assign layer0_outputs[6904] = inputs[142];
    assign layer0_outputs[6905] = (inputs[136]) & ~(inputs[542]);
    assign layer0_outputs[6906] = ~((inputs[236]) | (inputs[564]));
    assign layer0_outputs[6907] = ~((inputs[451]) | (inputs[366]));
    assign layer0_outputs[6908] = ~(inputs[532]);
    assign layer0_outputs[6909] = (inputs[244]) & (inputs[978]);
    assign layer0_outputs[6910] = ~(inputs[917]);
    assign layer0_outputs[6911] = (inputs[751]) & ~(inputs[612]);
    assign layer0_outputs[6912] = ~((inputs[39]) ^ (inputs[746]));
    assign layer0_outputs[6913] = (inputs[409]) & ~(inputs[46]);
    assign layer0_outputs[6914] = inputs[162];
    assign layer0_outputs[6915] = (inputs[553]) | (inputs[985]);
    assign layer0_outputs[6916] = ~((inputs[762]) | (inputs[841]));
    assign layer0_outputs[6917] = inputs[646];
    assign layer0_outputs[6918] = ~(inputs[426]) | (inputs[112]);
    assign layer0_outputs[6919] = ~(inputs[340]) | (inputs[520]);
    assign layer0_outputs[6920] = (inputs[401]) & (inputs[341]);
    assign layer0_outputs[6921] = (inputs[911]) | (inputs[421]);
    assign layer0_outputs[6922] = ~((inputs[220]) & (inputs[328]));
    assign layer0_outputs[6923] = ~((inputs[572]) | (inputs[848]));
    assign layer0_outputs[6924] = ~((inputs[661]) | (inputs[566]));
    assign layer0_outputs[6925] = ~((inputs[280]) | (inputs[246]));
    assign layer0_outputs[6926] = ~((inputs[235]) | (inputs[835]));
    assign layer0_outputs[6927] = (inputs[554]) & ~(inputs[463]);
    assign layer0_outputs[6928] = (inputs[217]) & ~(inputs[442]);
    assign layer0_outputs[6929] = ~((inputs[894]) ^ (inputs[203]));
    assign layer0_outputs[6930] = 1'b0;
    assign layer0_outputs[6931] = ~(inputs[278]);
    assign layer0_outputs[6932] = ~((inputs[504]) | (inputs[635]));
    assign layer0_outputs[6933] = ~((inputs[314]) | (inputs[171]));
    assign layer0_outputs[6934] = ~(inputs[207]) | (inputs[474]);
    assign layer0_outputs[6935] = (inputs[301]) | (inputs[809]);
    assign layer0_outputs[6936] = ~(inputs[742]) | (inputs[765]);
    assign layer0_outputs[6937] = (inputs[13]) & ~(inputs[152]);
    assign layer0_outputs[6938] = ~(inputs[438]) | (inputs[966]);
    assign layer0_outputs[6939] = (inputs[406]) & (inputs[587]);
    assign layer0_outputs[6940] = 1'b1;
    assign layer0_outputs[6941] = (inputs[332]) ^ (inputs[702]);
    assign layer0_outputs[6942] = ~(inputs[500]) | (inputs[697]);
    assign layer0_outputs[6943] = ~((inputs[608]) & (inputs[135]));
    assign layer0_outputs[6944] = (inputs[830]) & ~(inputs[970]);
    assign layer0_outputs[6945] = ~(inputs[316]) | (inputs[442]);
    assign layer0_outputs[6946] = ~(inputs[664]) | (inputs[384]);
    assign layer0_outputs[6947] = (inputs[320]) ^ (inputs[558]);
    assign layer0_outputs[6948] = ~((inputs[503]) | (inputs[968]));
    assign layer0_outputs[6949] = inputs[467];
    assign layer0_outputs[6950] = 1'b0;
    assign layer0_outputs[6951] = ~(inputs[427]);
    assign layer0_outputs[6952] = ~(inputs[725]);
    assign layer0_outputs[6953] = 1'b0;
    assign layer0_outputs[6954] = inputs[657];
    assign layer0_outputs[6955] = (inputs[847]) & ~(inputs[1008]);
    assign layer0_outputs[6956] = (inputs[317]) | (inputs[949]);
    assign layer0_outputs[6957] = (inputs[645]) ^ (inputs[581]);
    assign layer0_outputs[6958] = 1'b1;
    assign layer0_outputs[6959] = (inputs[907]) | (inputs[432]);
    assign layer0_outputs[6960] = (inputs[39]) ^ (inputs[709]);
    assign layer0_outputs[6961] = (inputs[765]) ^ (inputs[407]);
    assign layer0_outputs[6962] = (inputs[308]) ^ (inputs[185]);
    assign layer0_outputs[6963] = ~(inputs[375]) | (inputs[25]);
    assign layer0_outputs[6964] = inputs[470];
    assign layer0_outputs[6965] = (inputs[463]) & ~(inputs[991]);
    assign layer0_outputs[6966] = (inputs[898]) & ~(inputs[470]);
    assign layer0_outputs[6967] = ~(inputs[317]);
    assign layer0_outputs[6968] = (inputs[60]) | (inputs[695]);
    assign layer0_outputs[6969] = ~(inputs[434]);
    assign layer0_outputs[6970] = ~(inputs[621]) | (inputs[968]);
    assign layer0_outputs[6971] = inputs[725];
    assign layer0_outputs[6972] = (inputs[952]) & (inputs[982]);
    assign layer0_outputs[6973] = (inputs[782]) ^ (inputs[111]);
    assign layer0_outputs[6974] = ~((inputs[778]) | (inputs[742]));
    assign layer0_outputs[6975] = inputs[134];
    assign layer0_outputs[6976] = ~((inputs[821]) & (inputs[577]));
    assign layer0_outputs[6977] = ~(inputs[752]) | (inputs[382]);
    assign layer0_outputs[6978] = ~(inputs[15]) | (inputs[42]);
    assign layer0_outputs[6979] = 1'b1;
    assign layer0_outputs[6980] = ~(inputs[108]);
    assign layer0_outputs[6981] = ~(inputs[629]) | (inputs[878]);
    assign layer0_outputs[6982] = (inputs[350]) & (inputs[669]);
    assign layer0_outputs[6983] = ~((inputs[20]) ^ (inputs[561]));
    assign layer0_outputs[6984] = inputs[686];
    assign layer0_outputs[6985] = 1'b1;
    assign layer0_outputs[6986] = (inputs[248]) & ~(inputs[611]);
    assign layer0_outputs[6987] = (inputs[378]) | (inputs[943]);
    assign layer0_outputs[6988] = ~(inputs[25]);
    assign layer0_outputs[6989] = (inputs[438]) ^ (inputs[604]);
    assign layer0_outputs[6990] = (inputs[385]) | (inputs[316]);
    assign layer0_outputs[6991] = ~(inputs[628]) | (inputs[19]);
    assign layer0_outputs[6992] = inputs[371];
    assign layer0_outputs[6993] = (inputs[97]) | (inputs[771]);
    assign layer0_outputs[6994] = ~((inputs[369]) | (inputs[642]));
    assign layer0_outputs[6995] = ~(inputs[938]);
    assign layer0_outputs[6996] = (inputs[626]) & ~(inputs[799]);
    assign layer0_outputs[6997] = ~(inputs[918]);
    assign layer0_outputs[6998] = (inputs[932]) ^ (inputs[672]);
    assign layer0_outputs[6999] = ~(inputs[389]) | (inputs[258]);
    assign layer0_outputs[7000] = ~(inputs[521]) | (inputs[859]);
    assign layer0_outputs[7001] = inputs[465];
    assign layer0_outputs[7002] = ~((inputs[319]) | (inputs[190]));
    assign layer0_outputs[7003] = ~((inputs[774]) | (inputs[208]));
    assign layer0_outputs[7004] = ~(inputs[479]);
    assign layer0_outputs[7005] = (inputs[249]) & ~(inputs[873]);
    assign layer0_outputs[7006] = (inputs[519]) | (inputs[333]);
    assign layer0_outputs[7007] = ~((inputs[928]) | (inputs[618]));
    assign layer0_outputs[7008] = ~((inputs[201]) | (inputs[149]));
    assign layer0_outputs[7009] = 1'b0;
    assign layer0_outputs[7010] = ~((inputs[412]) | (inputs[782]));
    assign layer0_outputs[7011] = ~((inputs[191]) | (inputs[883]));
    assign layer0_outputs[7012] = (inputs[502]) | (inputs[359]);
    assign layer0_outputs[7013] = 1'b0;
    assign layer0_outputs[7014] = (inputs[644]) | (inputs[157]);
    assign layer0_outputs[7015] = ~(inputs[329]) | (inputs[826]);
    assign layer0_outputs[7016] = ~((inputs[753]) ^ (inputs[788]));
    assign layer0_outputs[7017] = (inputs[149]) & (inputs[955]);
    assign layer0_outputs[7018] = ~(inputs[456]) | (inputs[216]);
    assign layer0_outputs[7019] = ~(inputs[308]);
    assign layer0_outputs[7020] = 1'b0;
    assign layer0_outputs[7021] = inputs[690];
    assign layer0_outputs[7022] = inputs[241];
    assign layer0_outputs[7023] = ~((inputs[495]) ^ (inputs[859]));
    assign layer0_outputs[7024] = ~((inputs[817]) ^ (inputs[842]));
    assign layer0_outputs[7025] = (inputs[113]) & ~(inputs[446]);
    assign layer0_outputs[7026] = (inputs[630]) ^ (inputs[479]);
    assign layer0_outputs[7027] = inputs[236];
    assign layer0_outputs[7028] = (inputs[268]) & ~(inputs[659]);
    assign layer0_outputs[7029] = ~((inputs[518]) & (inputs[669]));
    assign layer0_outputs[7030] = (inputs[751]) & ~(inputs[768]);
    assign layer0_outputs[7031] = (inputs[498]) & ~(inputs[299]);
    assign layer0_outputs[7032] = ~(inputs[562]) | (inputs[970]);
    assign layer0_outputs[7033] = inputs[462];
    assign layer0_outputs[7034] = (inputs[705]) | (inputs[139]);
    assign layer0_outputs[7035] = (inputs[24]) & (inputs[320]);
    assign layer0_outputs[7036] = 1'b1;
    assign layer0_outputs[7037] = ~(inputs[26]);
    assign layer0_outputs[7038] = 1'b0;
    assign layer0_outputs[7039] = ~(inputs[845]) | (inputs[126]);
    assign layer0_outputs[7040] = ~(inputs[984]) | (inputs[888]);
    assign layer0_outputs[7041] = ~((inputs[515]) ^ (inputs[270]));
    assign layer0_outputs[7042] = ~(inputs[729]) | (inputs[224]);
    assign layer0_outputs[7043] = inputs[339];
    assign layer0_outputs[7044] = (inputs[82]) & ~(inputs[753]);
    assign layer0_outputs[7045] = ~(inputs[684]);
    assign layer0_outputs[7046] = 1'b0;
    assign layer0_outputs[7047] = inputs[448];
    assign layer0_outputs[7048] = (inputs[244]) | (inputs[378]);
    assign layer0_outputs[7049] = ~((inputs[74]) & (inputs[420]));
    assign layer0_outputs[7050] = ~(inputs[339]);
    assign layer0_outputs[7051] = ~((inputs[565]) | (inputs[706]));
    assign layer0_outputs[7052] = ~(inputs[893]);
    assign layer0_outputs[7053] = (inputs[743]) & (inputs[168]);
    assign layer0_outputs[7054] = inputs[239];
    assign layer0_outputs[7055] = ~(inputs[364]);
    assign layer0_outputs[7056] = inputs[837];
    assign layer0_outputs[7057] = (inputs[785]) | (inputs[474]);
    assign layer0_outputs[7058] = inputs[275];
    assign layer0_outputs[7059] = (inputs[516]) & (inputs[34]);
    assign layer0_outputs[7060] = (inputs[336]) ^ (inputs[773]);
    assign layer0_outputs[7061] = (inputs[957]) ^ (inputs[176]);
    assign layer0_outputs[7062] = ~(inputs[657]) | (inputs[74]);
    assign layer0_outputs[7063] = (inputs[47]) & ~(inputs[627]);
    assign layer0_outputs[7064] = ~(inputs[755]);
    assign layer0_outputs[7065] = inputs[174];
    assign layer0_outputs[7066] = (inputs[632]) & ~(inputs[197]);
    assign layer0_outputs[7067] = (inputs[1001]) & (inputs[482]);
    assign layer0_outputs[7068] = ~(inputs[911]) | (inputs[872]);
    assign layer0_outputs[7069] = inputs[340];
    assign layer0_outputs[7070] = ~(inputs[361]);
    assign layer0_outputs[7071] = (inputs[33]) & (inputs[504]);
    assign layer0_outputs[7072] = (inputs[27]) ^ (inputs[959]);
    assign layer0_outputs[7073] = ~((inputs[551]) ^ (inputs[415]));
    assign layer0_outputs[7074] = ~(inputs[680]);
    assign layer0_outputs[7075] = ~(inputs[880]) | (inputs[102]);
    assign layer0_outputs[7076] = (inputs[358]) | (inputs[228]);
    assign layer0_outputs[7077] = ~(inputs[589]) | (inputs[864]);
    assign layer0_outputs[7078] = ~((inputs[600]) | (inputs[901]));
    assign layer0_outputs[7079] = (inputs[124]) & (inputs[545]);
    assign layer0_outputs[7080] = 1'b1;
    assign layer0_outputs[7081] = (inputs[631]) & ~(inputs[237]);
    assign layer0_outputs[7082] = ~(inputs[468]);
    assign layer0_outputs[7083] = ~(inputs[313]);
    assign layer0_outputs[7084] = ~(inputs[278]) | (inputs[189]);
    assign layer0_outputs[7085] = inputs[146];
    assign layer0_outputs[7086] = ~(inputs[469]);
    assign layer0_outputs[7087] = (inputs[274]) | (inputs[939]);
    assign layer0_outputs[7088] = ~(inputs[438]);
    assign layer0_outputs[7089] = ~((inputs[370]) ^ (inputs[133]));
    assign layer0_outputs[7090] = (inputs[308]) ^ (inputs[889]);
    assign layer0_outputs[7091] = ~((inputs[80]) | (inputs[26]));
    assign layer0_outputs[7092] = 1'b1;
    assign layer0_outputs[7093] = (inputs[670]) & ~(inputs[733]);
    assign layer0_outputs[7094] = 1'b1;
    assign layer0_outputs[7095] = (inputs[205]) & ~(inputs[974]);
    assign layer0_outputs[7096] = (inputs[873]) & ~(inputs[886]);
    assign layer0_outputs[7097] = inputs[423];
    assign layer0_outputs[7098] = ~(inputs[87]) | (inputs[765]);
    assign layer0_outputs[7099] = (inputs[423]) | (inputs[139]);
    assign layer0_outputs[7100] = ~(inputs[101]) | (inputs[165]);
    assign layer0_outputs[7101] = ~((inputs[313]) | (inputs[233]));
    assign layer0_outputs[7102] = ~(inputs[619]) | (inputs[343]);
    assign layer0_outputs[7103] = ~(inputs[776]) | (inputs[229]);
    assign layer0_outputs[7104] = ~(inputs[721]);
    assign layer0_outputs[7105] = ~(inputs[330]) | (inputs[442]);
    assign layer0_outputs[7106] = (inputs[345]) ^ (inputs[319]);
    assign layer0_outputs[7107] = inputs[876];
    assign layer0_outputs[7108] = (inputs[272]) & (inputs[302]);
    assign layer0_outputs[7109] = ~(inputs[811]);
    assign layer0_outputs[7110] = ~((inputs[360]) | (inputs[982]));
    assign layer0_outputs[7111] = (inputs[8]) ^ (inputs[579]);
    assign layer0_outputs[7112] = (inputs[774]) | (inputs[855]);
    assign layer0_outputs[7113] = 1'b0;
    assign layer0_outputs[7114] = inputs[147];
    assign layer0_outputs[7115] = ~((inputs[867]) ^ (inputs[563]));
    assign layer0_outputs[7116] = ~((inputs[70]) | (inputs[214]));
    assign layer0_outputs[7117] = (inputs[442]) ^ (inputs[212]);
    assign layer0_outputs[7118] = ~(inputs[187]);
    assign layer0_outputs[7119] = (inputs[300]) ^ (inputs[256]);
    assign layer0_outputs[7120] = inputs[238];
    assign layer0_outputs[7121] = ~(inputs[478]) | (inputs[638]);
    assign layer0_outputs[7122] = (inputs[359]) & ~(inputs[611]);
    assign layer0_outputs[7123] = (inputs[879]) | (inputs[924]);
    assign layer0_outputs[7124] = (inputs[1016]) ^ (inputs[819]);
    assign layer0_outputs[7125] = (inputs[990]) ^ (inputs[427]);
    assign layer0_outputs[7126] = ~(inputs[876]);
    assign layer0_outputs[7127] = ~((inputs[672]) ^ (inputs[47]));
    assign layer0_outputs[7128] = (inputs[297]) ^ (inputs[928]);
    assign layer0_outputs[7129] = inputs[955];
    assign layer0_outputs[7130] = ~(inputs[199]);
    assign layer0_outputs[7131] = ~(inputs[927]) | (inputs[374]);
    assign layer0_outputs[7132] = (inputs[635]) | (inputs[651]);
    assign layer0_outputs[7133] = (inputs[67]) | (inputs[623]);
    assign layer0_outputs[7134] = ~(inputs[554]) | (inputs[958]);
    assign layer0_outputs[7135] = (inputs[465]) & ~(inputs[587]);
    assign layer0_outputs[7136] = (inputs[791]) & ~(inputs[555]);
    assign layer0_outputs[7137] = inputs[719];
    assign layer0_outputs[7138] = ~((inputs[719]) | (inputs[686]));
    assign layer0_outputs[7139] = ~(inputs[64]) | (inputs[637]);
    assign layer0_outputs[7140] = inputs[912];
    assign layer0_outputs[7141] = ~((inputs[119]) ^ (inputs[444]));
    assign layer0_outputs[7142] = (inputs[250]) & ~(inputs[552]);
    assign layer0_outputs[7143] = (inputs[960]) ^ (inputs[448]);
    assign layer0_outputs[7144] = 1'b1;
    assign layer0_outputs[7145] = ~(inputs[627]);
    assign layer0_outputs[7146] = 1'b0;
    assign layer0_outputs[7147] = ~(inputs[364]) | (inputs[143]);
    assign layer0_outputs[7148] = ~(inputs[93]);
    assign layer0_outputs[7149] = ~((inputs[575]) | (inputs[776]));
    assign layer0_outputs[7150] = inputs[212];
    assign layer0_outputs[7151] = inputs[882];
    assign layer0_outputs[7152] = (inputs[322]) & (inputs[865]);
    assign layer0_outputs[7153] = ~(inputs[776]) | (inputs[324]);
    assign layer0_outputs[7154] = ~(inputs[108]);
    assign layer0_outputs[7155] = ~((inputs[265]) | (inputs[236]));
    assign layer0_outputs[7156] = ~(inputs[887]) | (inputs[804]);
    assign layer0_outputs[7157] = ~(inputs[282]) | (inputs[35]);
    assign layer0_outputs[7158] = ~(inputs[936]) | (inputs[894]);
    assign layer0_outputs[7159] = ~(inputs[568]) | (inputs[890]);
    assign layer0_outputs[7160] = ~(inputs[819]);
    assign layer0_outputs[7161] = (inputs[825]) | (inputs[220]);
    assign layer0_outputs[7162] = ~((inputs[351]) ^ (inputs[898]));
    assign layer0_outputs[7163] = ~((inputs[979]) ^ (inputs[190]));
    assign layer0_outputs[7164] = inputs[566];
    assign layer0_outputs[7165] = inputs[532];
    assign layer0_outputs[7166] = ~((inputs[121]) | (inputs[210]));
    assign layer0_outputs[7167] = ~((inputs[282]) ^ (inputs[194]));
    assign layer0_outputs[7168] = ~(inputs[666]) | (inputs[230]);
    assign layer0_outputs[7169] = (inputs[912]) & ~(inputs[311]);
    assign layer0_outputs[7170] = (inputs[410]) | (inputs[1004]);
    assign layer0_outputs[7171] = (inputs[222]) & ~(inputs[581]);
    assign layer0_outputs[7172] = (inputs[561]) ^ (inputs[667]);
    assign layer0_outputs[7173] = inputs[559];
    assign layer0_outputs[7174] = ~((inputs[264]) | (inputs[318]));
    assign layer0_outputs[7175] = ~(inputs[321]) | (inputs[642]);
    assign layer0_outputs[7176] = inputs[569];
    assign layer0_outputs[7177] = inputs[712];
    assign layer0_outputs[7178] = (inputs[687]) & ~(inputs[328]);
    assign layer0_outputs[7179] = (inputs[415]) | (inputs[938]);
    assign layer0_outputs[7180] = (inputs[762]) & ~(inputs[925]);
    assign layer0_outputs[7181] = inputs[753];
    assign layer0_outputs[7182] = ~((inputs[899]) ^ (inputs[250]));
    assign layer0_outputs[7183] = (inputs[789]) & ~(inputs[917]);
    assign layer0_outputs[7184] = ~(inputs[829]) | (inputs[351]);
    assign layer0_outputs[7185] = ~(inputs[641]);
    assign layer0_outputs[7186] = (inputs[705]) | (inputs[93]);
    assign layer0_outputs[7187] = ~(inputs[723]) | (inputs[805]);
    assign layer0_outputs[7188] = ~(inputs[160]);
    assign layer0_outputs[7189] = (inputs[157]) & ~(inputs[932]);
    assign layer0_outputs[7190] = ~(inputs[116]) | (inputs[576]);
    assign layer0_outputs[7191] = (inputs[265]) ^ (inputs[409]);
    assign layer0_outputs[7192] = ~(inputs[402]);
    assign layer0_outputs[7193] = (inputs[505]) & ~(inputs[802]);
    assign layer0_outputs[7194] = (inputs[712]) ^ (inputs[995]);
    assign layer0_outputs[7195] = ~(inputs[528]) | (inputs[7]);
    assign layer0_outputs[7196] = (inputs[297]) & ~(inputs[577]);
    assign layer0_outputs[7197] = inputs[911];
    assign layer0_outputs[7198] = ~(inputs[50]);
    assign layer0_outputs[7199] = inputs[933];
    assign layer0_outputs[7200] = ~(inputs[580]);
    assign layer0_outputs[7201] = (inputs[565]) | (inputs[981]);
    assign layer0_outputs[7202] = (inputs[220]) ^ (inputs[828]);
    assign layer0_outputs[7203] = (inputs[17]) & ~(inputs[482]);
    assign layer0_outputs[7204] = 1'b1;
    assign layer0_outputs[7205] = ~((inputs[509]) | (inputs[115]));
    assign layer0_outputs[7206] = inputs[664];
    assign layer0_outputs[7207] = inputs[961];
    assign layer0_outputs[7208] = ~((inputs[59]) | (inputs[430]));
    assign layer0_outputs[7209] = ~((inputs[675]) ^ (inputs[776]));
    assign layer0_outputs[7210] = (inputs[762]) & (inputs[263]);
    assign layer0_outputs[7211] = (inputs[677]) | (inputs[582]);
    assign layer0_outputs[7212] = ~((inputs[557]) | (inputs[60]));
    assign layer0_outputs[7213] = ~((inputs[240]) | (inputs[620]));
    assign layer0_outputs[7214] = (inputs[440]) & ~(inputs[316]);
    assign layer0_outputs[7215] = (inputs[707]) ^ (inputs[748]);
    assign layer0_outputs[7216] = inputs[886];
    assign layer0_outputs[7217] = ~((inputs[348]) ^ (inputs[394]));
    assign layer0_outputs[7218] = ~((inputs[568]) | (inputs[292]));
    assign layer0_outputs[7219] = (inputs[674]) | (inputs[206]);
    assign layer0_outputs[7220] = inputs[315];
    assign layer0_outputs[7221] = ~((inputs[573]) | (inputs[125]));
    assign layer0_outputs[7222] = ~((inputs[670]) ^ (inputs[414]));
    assign layer0_outputs[7223] = 1'b1;
    assign layer0_outputs[7224] = ~(inputs[682]);
    assign layer0_outputs[7225] = ~(inputs[126]) | (inputs[31]);
    assign layer0_outputs[7226] = inputs[398];
    assign layer0_outputs[7227] = 1'b1;
    assign layer0_outputs[7228] = (inputs[740]) | (inputs[976]);
    assign layer0_outputs[7229] = ~((inputs[151]) | (inputs[274]));
    assign layer0_outputs[7230] = ~(inputs[153]);
    assign layer0_outputs[7231] = ~(inputs[623]) | (inputs[768]);
    assign layer0_outputs[7232] = inputs[808];
    assign layer0_outputs[7233] = (inputs[259]) & ~(inputs[829]);
    assign layer0_outputs[7234] = (inputs[896]) & ~(inputs[71]);
    assign layer0_outputs[7235] = (inputs[311]) ^ (inputs[578]);
    assign layer0_outputs[7236] = (inputs[922]) & ~(inputs[608]);
    assign layer0_outputs[7237] = ~(inputs[345]);
    assign layer0_outputs[7238] = ~(inputs[150]) | (inputs[225]);
    assign layer0_outputs[7239] = ~(inputs[503]);
    assign layer0_outputs[7240] = (inputs[698]) & ~(inputs[221]);
    assign layer0_outputs[7241] = ~(inputs[617]);
    assign layer0_outputs[7242] = (inputs[497]) ^ (inputs[57]);
    assign layer0_outputs[7243] = ~((inputs[578]) ^ (inputs[425]));
    assign layer0_outputs[7244] = ~(inputs[289]) | (inputs[71]);
    assign layer0_outputs[7245] = ~(inputs[294]);
    assign layer0_outputs[7246] = inputs[596];
    assign layer0_outputs[7247] = ~(inputs[434]) | (inputs[92]);
    assign layer0_outputs[7248] = (inputs[73]) | (inputs[232]);
    assign layer0_outputs[7249] = ~(inputs[658]) | (inputs[545]);
    assign layer0_outputs[7250] = (inputs[658]) & ~(inputs[105]);
    assign layer0_outputs[7251] = ~((inputs[992]) ^ (inputs[480]));
    assign layer0_outputs[7252] = ~((inputs[8]) & (inputs[503]));
    assign layer0_outputs[7253] = ~((inputs[361]) | (inputs[693]));
    assign layer0_outputs[7254] = (inputs[500]) & ~(inputs[966]);
    assign layer0_outputs[7255] = ~(inputs[157]);
    assign layer0_outputs[7256] = (inputs[978]) & ~(inputs[97]);
    assign layer0_outputs[7257] = ~(inputs[688]);
    assign layer0_outputs[7258] = (inputs[759]) | (inputs[695]);
    assign layer0_outputs[7259] = ~((inputs[1013]) | (inputs[855]));
    assign layer0_outputs[7260] = (inputs[326]) | (inputs[192]);
    assign layer0_outputs[7261] = (inputs[940]) ^ (inputs[601]);
    assign layer0_outputs[7262] = ~((inputs[149]) | (inputs[756]));
    assign layer0_outputs[7263] = (inputs[672]) & (inputs[29]);
    assign layer0_outputs[7264] = ~((inputs[507]) | (inputs[858]));
    assign layer0_outputs[7265] = (inputs[320]) & ~(inputs[885]);
    assign layer0_outputs[7266] = (inputs[564]) ^ (inputs[964]);
    assign layer0_outputs[7267] = ~((inputs[496]) ^ (inputs[566]));
    assign layer0_outputs[7268] = inputs[293];
    assign layer0_outputs[7269] = 1'b0;
    assign layer0_outputs[7270] = (inputs[787]) & ~(inputs[81]);
    assign layer0_outputs[7271] = (inputs[24]) | (inputs[922]);
    assign layer0_outputs[7272] = ~(inputs[439]) | (inputs[732]);
    assign layer0_outputs[7273] = ~((inputs[26]) & (inputs[476]));
    assign layer0_outputs[7274] = ~((inputs[544]) | (inputs[753]));
    assign layer0_outputs[7275] = inputs[463];
    assign layer0_outputs[7276] = (inputs[373]) ^ (inputs[369]);
    assign layer0_outputs[7277] = (inputs[620]) | (inputs[97]);
    assign layer0_outputs[7278] = 1'b0;
    assign layer0_outputs[7279] = ~((inputs[586]) ^ (inputs[808]));
    assign layer0_outputs[7280] = (inputs[919]) & ~(inputs[441]);
    assign layer0_outputs[7281] = (inputs[303]) ^ (inputs[484]);
    assign layer0_outputs[7282] = (inputs[530]) & ~(inputs[248]);
    assign layer0_outputs[7283] = ~((inputs[285]) ^ (inputs[434]));
    assign layer0_outputs[7284] = ~((inputs[366]) ^ (inputs[1002]));
    assign layer0_outputs[7285] = ~((inputs[982]) | (inputs[475]));
    assign layer0_outputs[7286] = ~((inputs[802]) | (inputs[749]));
    assign layer0_outputs[7287] = ~((inputs[101]) | (inputs[843]));
    assign layer0_outputs[7288] = (inputs[493]) ^ (inputs[797]);
    assign layer0_outputs[7289] = inputs[702];
    assign layer0_outputs[7290] = (inputs[397]) | (inputs[967]);
    assign layer0_outputs[7291] = ~((inputs[181]) | (inputs[117]));
    assign layer0_outputs[7292] = 1'b0;
    assign layer0_outputs[7293] = (inputs[816]) & ~(inputs[543]);
    assign layer0_outputs[7294] = (inputs[397]) | (inputs[104]);
    assign layer0_outputs[7295] = (inputs[64]) & ~(inputs[641]);
    assign layer0_outputs[7296] = ~(inputs[618]) | (inputs[165]);
    assign layer0_outputs[7297] = (inputs[740]) & ~(inputs[59]);
    assign layer0_outputs[7298] = ~(inputs[728]);
    assign layer0_outputs[7299] = (inputs[758]) ^ (inputs[673]);
    assign layer0_outputs[7300] = ~(inputs[207]) | (inputs[220]);
    assign layer0_outputs[7301] = ~(inputs[534]);
    assign layer0_outputs[7302] = ~(inputs[936]);
    assign layer0_outputs[7303] = (inputs[413]) | (inputs[722]);
    assign layer0_outputs[7304] = inputs[792];
    assign layer0_outputs[7305] = (inputs[732]) | (inputs[330]);
    assign layer0_outputs[7306] = ~(inputs[828]) | (inputs[140]);
    assign layer0_outputs[7307] = ~((inputs[819]) ^ (inputs[820]));
    assign layer0_outputs[7308] = ~(inputs[500]);
    assign layer0_outputs[7309] = ~((inputs[633]) | (inputs[875]));
    assign layer0_outputs[7310] = (inputs[970]) | (inputs[145]);
    assign layer0_outputs[7311] = ~((inputs[455]) ^ (inputs[170]));
    assign layer0_outputs[7312] = 1'b1;
    assign layer0_outputs[7313] = (inputs[11]) & ~(inputs[542]);
    assign layer0_outputs[7314] = inputs[525];
    assign layer0_outputs[7315] = (inputs[741]) | (inputs[709]);
    assign layer0_outputs[7316] = (inputs[620]) ^ (inputs[280]);
    assign layer0_outputs[7317] = ~(inputs[918]) | (inputs[655]);
    assign layer0_outputs[7318] = ~((inputs[944]) ^ (inputs[150]));
    assign layer0_outputs[7319] = ~(inputs[207]);
    assign layer0_outputs[7320] = (inputs[723]) | (inputs[455]);
    assign layer0_outputs[7321] = (inputs[174]) | (inputs[464]);
    assign layer0_outputs[7322] = ~((inputs[38]) & (inputs[286]));
    assign layer0_outputs[7323] = ~(inputs[633]) | (inputs[544]);
    assign layer0_outputs[7324] = ~(inputs[273]);
    assign layer0_outputs[7325] = (inputs[265]) | (inputs[735]);
    assign layer0_outputs[7326] = ~((inputs[195]) | (inputs[1001]));
    assign layer0_outputs[7327] = ~(inputs[212]) | (inputs[158]);
    assign layer0_outputs[7328] = ~((inputs[734]) ^ (inputs[854]));
    assign layer0_outputs[7329] = inputs[785];
    assign layer0_outputs[7330] = (inputs[777]) & ~(inputs[85]);
    assign layer0_outputs[7331] = ~((inputs[441]) ^ (inputs[466]));
    assign layer0_outputs[7332] = ~((inputs[738]) ^ (inputs[467]));
    assign layer0_outputs[7333] = (inputs[973]) | (inputs[303]);
    assign layer0_outputs[7334] = ~((inputs[193]) ^ (inputs[450]));
    assign layer0_outputs[7335] = ~(inputs[380]) | (inputs[735]);
    assign layer0_outputs[7336] = ~((inputs[97]) | (inputs[895]));
    assign layer0_outputs[7337] = (inputs[894]) ^ (inputs[337]);
    assign layer0_outputs[7338] = ~(inputs[482]);
    assign layer0_outputs[7339] = ~(inputs[148]) | (inputs[881]);
    assign layer0_outputs[7340] = (inputs[538]) | (inputs[804]);
    assign layer0_outputs[7341] = ~(inputs[617]);
    assign layer0_outputs[7342] = ~(inputs[554]);
    assign layer0_outputs[7343] = ~((inputs[705]) | (inputs[437]));
    assign layer0_outputs[7344] = ~(inputs[912]) | (inputs[189]);
    assign layer0_outputs[7345] = (inputs[54]) ^ (inputs[925]);
    assign layer0_outputs[7346] = (inputs[723]) | (inputs[107]);
    assign layer0_outputs[7347] = (inputs[584]) & ~(inputs[176]);
    assign layer0_outputs[7348] = inputs[654];
    assign layer0_outputs[7349] = (inputs[531]) & ~(inputs[512]);
    assign layer0_outputs[7350] = 1'b0;
    assign layer0_outputs[7351] = (inputs[606]) & (inputs[967]);
    assign layer0_outputs[7352] = inputs[977];
    assign layer0_outputs[7353] = inputs[70];
    assign layer0_outputs[7354] = (inputs[395]) & ~(inputs[658]);
    assign layer0_outputs[7355] = ~(inputs[832]) | (inputs[12]);
    assign layer0_outputs[7356] = ~((inputs[676]) | (inputs[172]));
    assign layer0_outputs[7357] = inputs[945];
    assign layer0_outputs[7358] = inputs[795];
    assign layer0_outputs[7359] = (inputs[335]) & ~(inputs[283]);
    assign layer0_outputs[7360] = ~((inputs[367]) ^ (inputs[747]));
    assign layer0_outputs[7361] = ~(inputs[590]);
    assign layer0_outputs[7362] = ~(inputs[661]);
    assign layer0_outputs[7363] = ~(inputs[992]);
    assign layer0_outputs[7364] = inputs[607];
    assign layer0_outputs[7365] = 1'b1;
    assign layer0_outputs[7366] = ~((inputs[968]) | (inputs[244]));
    assign layer0_outputs[7367] = ~(inputs[902]);
    assign layer0_outputs[7368] = (inputs[617]) ^ (inputs[652]);
    assign layer0_outputs[7369] = (inputs[745]) & ~(inputs[366]);
    assign layer0_outputs[7370] = ~((inputs[652]) | (inputs[78]));
    assign layer0_outputs[7371] = (inputs[484]) | (inputs[372]);
    assign layer0_outputs[7372] = (inputs[166]) ^ (inputs[574]);
    assign layer0_outputs[7373] = ~(inputs[598]);
    assign layer0_outputs[7374] = (inputs[243]) & ~(inputs[952]);
    assign layer0_outputs[7375] = ~(inputs[921]) | (inputs[605]);
    assign layer0_outputs[7376] = ~(inputs[506]);
    assign layer0_outputs[7377] = ~(inputs[338]);
    assign layer0_outputs[7378] = ~(inputs[562]);
    assign layer0_outputs[7379] = (inputs[201]) ^ (inputs[967]);
    assign layer0_outputs[7380] = ~((inputs[944]) | (inputs[514]));
    assign layer0_outputs[7381] = (inputs[460]) & ~(inputs[260]);
    assign layer0_outputs[7382] = ~(inputs[718]) | (inputs[990]);
    assign layer0_outputs[7383] = ~(inputs[679]);
    assign layer0_outputs[7384] = (inputs[24]) & ~(inputs[962]);
    assign layer0_outputs[7385] = ~((inputs[662]) ^ (inputs[725]));
    assign layer0_outputs[7386] = (inputs[751]) | (inputs[141]);
    assign layer0_outputs[7387] = (inputs[567]) | (inputs[823]);
    assign layer0_outputs[7388] = ~(inputs[101]);
    assign layer0_outputs[7389] = (inputs[755]) ^ (inputs[651]);
    assign layer0_outputs[7390] = ~(inputs[492]);
    assign layer0_outputs[7391] = ~(inputs[648]);
    assign layer0_outputs[7392] = inputs[420];
    assign layer0_outputs[7393] = (inputs[466]) & ~(inputs[106]);
    assign layer0_outputs[7394] = (inputs[132]) | (inputs[531]);
    assign layer0_outputs[7395] = ~(inputs[310]);
    assign layer0_outputs[7396] = (inputs[359]) & ~(inputs[159]);
    assign layer0_outputs[7397] = inputs[300];
    assign layer0_outputs[7398] = ~(inputs[80]);
    assign layer0_outputs[7399] = inputs[826];
    assign layer0_outputs[7400] = ~((inputs[416]) | (inputs[192]));
    assign layer0_outputs[7401] = (inputs[852]) | (inputs[851]);
    assign layer0_outputs[7402] = inputs[207];
    assign layer0_outputs[7403] = ~((inputs[71]) | (inputs[245]));
    assign layer0_outputs[7404] = ~((inputs[45]) ^ (inputs[644]));
    assign layer0_outputs[7405] = ~(inputs[1004]) | (inputs[947]);
    assign layer0_outputs[7406] = ~(inputs[303]) | (inputs[130]);
    assign layer0_outputs[7407] = (inputs[111]) & ~(inputs[413]);
    assign layer0_outputs[7408] = (inputs[562]) & ~(inputs[987]);
    assign layer0_outputs[7409] = ~((inputs[429]) | (inputs[195]));
    assign layer0_outputs[7410] = ~((inputs[63]) ^ (inputs[305]));
    assign layer0_outputs[7411] = inputs[386];
    assign layer0_outputs[7412] = ~(inputs[535]);
    assign layer0_outputs[7413] = ~(inputs[793]);
    assign layer0_outputs[7414] = ~(inputs[62]);
    assign layer0_outputs[7415] = ~(inputs[178]);
    assign layer0_outputs[7416] = (inputs[581]) ^ (inputs[446]);
    assign layer0_outputs[7417] = inputs[497];
    assign layer0_outputs[7418] = ~((inputs[521]) | (inputs[510]));
    assign layer0_outputs[7419] = ~(inputs[629]) | (inputs[938]);
    assign layer0_outputs[7420] = (inputs[551]) | (inputs[986]);
    assign layer0_outputs[7421] = (inputs[357]) ^ (inputs[541]);
    assign layer0_outputs[7422] = ~((inputs[701]) | (inputs[698]));
    assign layer0_outputs[7423] = (inputs[979]) | (inputs[987]);
    assign layer0_outputs[7424] = 1'b1;
    assign layer0_outputs[7425] = (inputs[299]) & ~(inputs[154]);
    assign layer0_outputs[7426] = ~(inputs[822]) | (inputs[208]);
    assign layer0_outputs[7427] = ~((inputs[449]) | (inputs[596]));
    assign layer0_outputs[7428] = (inputs[710]) | (inputs[812]);
    assign layer0_outputs[7429] = ~((inputs[977]) | (inputs[340]));
    assign layer0_outputs[7430] = ~((inputs[614]) | (inputs[277]));
    assign layer0_outputs[7431] = inputs[395];
    assign layer0_outputs[7432] = ~(inputs[689]) | (inputs[182]);
    assign layer0_outputs[7433] = inputs[856];
    assign layer0_outputs[7434] = (inputs[339]) | (inputs[582]);
    assign layer0_outputs[7435] = 1'b0;
    assign layer0_outputs[7436] = (inputs[984]) | (inputs[233]);
    assign layer0_outputs[7437] = (inputs[624]) | (inputs[162]);
    assign layer0_outputs[7438] = 1'b1;
    assign layer0_outputs[7439] = (inputs[461]) & ~(inputs[197]);
    assign layer0_outputs[7440] = ~((inputs[408]) ^ (inputs[225]));
    assign layer0_outputs[7441] = ~((inputs[548]) ^ (inputs[458]));
    assign layer0_outputs[7442] = (inputs[999]) & (inputs[163]);
    assign layer0_outputs[7443] = inputs[340];
    assign layer0_outputs[7444] = inputs[584];
    assign layer0_outputs[7445] = ~((inputs[826]) | (inputs[848]));
    assign layer0_outputs[7446] = (inputs[152]) & ~(inputs[644]);
    assign layer0_outputs[7447] = inputs[609];
    assign layer0_outputs[7448] = (inputs[343]) & ~(inputs[334]);
    assign layer0_outputs[7449] = ~((inputs[237]) ^ (inputs[36]));
    assign layer0_outputs[7450] = ~(inputs[120]);
    assign layer0_outputs[7451] = ~((inputs[89]) ^ (inputs[506]));
    assign layer0_outputs[7452] = inputs[387];
    assign layer0_outputs[7453] = inputs[979];
    assign layer0_outputs[7454] = inputs[213];
    assign layer0_outputs[7455] = ~((inputs[225]) ^ (inputs[308]));
    assign layer0_outputs[7456] = ~(inputs[547]);
    assign layer0_outputs[7457] = (inputs[516]) ^ (inputs[544]);
    assign layer0_outputs[7458] = ~(inputs[682]);
    assign layer0_outputs[7459] = (inputs[465]) | (inputs[1017]);
    assign layer0_outputs[7460] = ~(inputs[400]);
    assign layer0_outputs[7461] = ~((inputs[685]) ^ (inputs[568]));
    assign layer0_outputs[7462] = ~((inputs[223]) | (inputs[849]));
    assign layer0_outputs[7463] = ~((inputs[97]) ^ (inputs[18]));
    assign layer0_outputs[7464] = inputs[527];
    assign layer0_outputs[7465] = inputs[711];
    assign layer0_outputs[7466] = (inputs[218]) | (inputs[489]);
    assign layer0_outputs[7467] = (inputs[175]) & ~(inputs[35]);
    assign layer0_outputs[7468] = inputs[939];
    assign layer0_outputs[7469] = ~(inputs[273]) | (inputs[636]);
    assign layer0_outputs[7470] = ~(inputs[558]);
    assign layer0_outputs[7471] = ~(inputs[17]);
    assign layer0_outputs[7472] = inputs[366];
    assign layer0_outputs[7473] = ~((inputs[559]) | (inputs[109]));
    assign layer0_outputs[7474] = inputs[747];
    assign layer0_outputs[7475] = ~(inputs[298]) | (inputs[47]);
    assign layer0_outputs[7476] = (inputs[754]) & ~(inputs[637]);
    assign layer0_outputs[7477] = ~(inputs[781]);
    assign layer0_outputs[7478] = ~(inputs[529]);
    assign layer0_outputs[7479] = (inputs[687]) & ~(inputs[150]);
    assign layer0_outputs[7480] = ~(inputs[927]) | (inputs[170]);
    assign layer0_outputs[7481] = (inputs[651]) | (inputs[472]);
    assign layer0_outputs[7482] = (inputs[358]) ^ (inputs[447]);
    assign layer0_outputs[7483] = (inputs[789]) | (inputs[914]);
    assign layer0_outputs[7484] = ~((inputs[338]) & (inputs[54]));
    assign layer0_outputs[7485] = (inputs[38]) & (inputs[893]);
    assign layer0_outputs[7486] = (inputs[850]) | (inputs[710]);
    assign layer0_outputs[7487] = ~((inputs[575]) ^ (inputs[219]));
    assign layer0_outputs[7488] = inputs[277];
    assign layer0_outputs[7489] = ~((inputs[203]) | (inputs[783]));
    assign layer0_outputs[7490] = (inputs[200]) ^ (inputs[711]);
    assign layer0_outputs[7491] = ~((inputs[814]) | (inputs[128]));
    assign layer0_outputs[7492] = (inputs[423]) | (inputs[32]);
    assign layer0_outputs[7493] = inputs[282];
    assign layer0_outputs[7494] = ~((inputs[712]) | (inputs[604]));
    assign layer0_outputs[7495] = ~((inputs[150]) ^ (inputs[204]));
    assign layer0_outputs[7496] = (inputs[373]) & ~(inputs[121]);
    assign layer0_outputs[7497] = ~((inputs[801]) ^ (inputs[385]));
    assign layer0_outputs[7498] = inputs[635];
    assign layer0_outputs[7499] = ~(inputs[910]);
    assign layer0_outputs[7500] = (inputs[1015]) ^ (inputs[278]);
    assign layer0_outputs[7501] = ~(inputs[961]) | (inputs[62]);
    assign layer0_outputs[7502] = inputs[504];
    assign layer0_outputs[7503] = ~(inputs[205]);
    assign layer0_outputs[7504] = ~((inputs[869]) | (inputs[761]));
    assign layer0_outputs[7505] = ~(inputs[499]);
    assign layer0_outputs[7506] = (inputs[45]) | (inputs[224]);
    assign layer0_outputs[7507] = ~(inputs[745]);
    assign layer0_outputs[7508] = ~(inputs[1019]);
    assign layer0_outputs[7509] = inputs[415];
    assign layer0_outputs[7510] = (inputs[17]) & ~(inputs[422]);
    assign layer0_outputs[7511] = ~(inputs[207]);
    assign layer0_outputs[7512] = ~((inputs[730]) | (inputs[381]));
    assign layer0_outputs[7513] = (inputs[768]) & ~(inputs[787]);
    assign layer0_outputs[7514] = ~((inputs[226]) ^ (inputs[248]));
    assign layer0_outputs[7515] = (inputs[834]) ^ (inputs[307]);
    assign layer0_outputs[7516] = (inputs[877]) & ~(inputs[295]);
    assign layer0_outputs[7517] = ~((inputs[327]) ^ (inputs[711]));
    assign layer0_outputs[7518] = ~((inputs[39]) & (inputs[858]));
    assign layer0_outputs[7519] = (inputs[848]) | (inputs[909]);
    assign layer0_outputs[7520] = ~(inputs[502]);
    assign layer0_outputs[7521] = (inputs[815]) ^ (inputs[609]);
    assign layer0_outputs[7522] = ~(inputs[994]) | (inputs[857]);
    assign layer0_outputs[7523] = (inputs[625]) & ~(inputs[969]);
    assign layer0_outputs[7524] = (inputs[678]) & ~(inputs[192]);
    assign layer0_outputs[7525] = ~((inputs[850]) | (inputs[30]));
    assign layer0_outputs[7526] = ~((inputs[742]) ^ (inputs[792]));
    assign layer0_outputs[7527] = ~((inputs[709]) ^ (inputs[896]));
    assign layer0_outputs[7528] = (inputs[915]) & ~(inputs[139]);
    assign layer0_outputs[7529] = ~(inputs[374]) | (inputs[46]);
    assign layer0_outputs[7530] = (inputs[984]) & (inputs[356]);
    assign layer0_outputs[7531] = ~(inputs[588]);
    assign layer0_outputs[7532] = ~(inputs[467]) | (inputs[346]);
    assign layer0_outputs[7533] = 1'b1;
    assign layer0_outputs[7534] = ~(inputs[823]);
    assign layer0_outputs[7535] = ~(inputs[587]) | (inputs[1010]);
    assign layer0_outputs[7536] = ~((inputs[733]) & (inputs[25]));
    assign layer0_outputs[7537] = (inputs[1018]) & ~(inputs[231]);
    assign layer0_outputs[7538] = (inputs[146]) | (inputs[794]);
    assign layer0_outputs[7539] = ~((inputs[530]) | (inputs[983]));
    assign layer0_outputs[7540] = (inputs[1014]) & (inputs[833]);
    assign layer0_outputs[7541] = (inputs[655]) & ~(inputs[169]);
    assign layer0_outputs[7542] = (inputs[234]) ^ (inputs[226]);
    assign layer0_outputs[7543] = ~((inputs[477]) | (inputs[274]));
    assign layer0_outputs[7544] = ~((inputs[496]) ^ (inputs[773]));
    assign layer0_outputs[7545] = (inputs[375]) & (inputs[275]);
    assign layer0_outputs[7546] = (inputs[590]) & ~(inputs[1001]);
    assign layer0_outputs[7547] = inputs[171];
    assign layer0_outputs[7548] = ~((inputs[626]) ^ (inputs[385]));
    assign layer0_outputs[7549] = ~((inputs[158]) | (inputs[838]));
    assign layer0_outputs[7550] = ~((inputs[228]) | (inputs[0]));
    assign layer0_outputs[7551] = ~((inputs[824]) ^ (inputs[833]));
    assign layer0_outputs[7552] = ~((inputs[1006]) | (inputs[547]));
    assign layer0_outputs[7553] = ~(inputs[336]);
    assign layer0_outputs[7554] = inputs[366];
    assign layer0_outputs[7555] = 1'b0;
    assign layer0_outputs[7556] = 1'b0;
    assign layer0_outputs[7557] = ~((inputs[103]) | (inputs[845]));
    assign layer0_outputs[7558] = ~((inputs[683]) ^ (inputs[149]));
    assign layer0_outputs[7559] = ~(inputs[38]);
    assign layer0_outputs[7560] = 1'b0;
    assign layer0_outputs[7561] = ~(inputs[215]) | (inputs[162]);
    assign layer0_outputs[7562] = inputs[728];
    assign layer0_outputs[7563] = ~((inputs[252]) ^ (inputs[377]));
    assign layer0_outputs[7564] = inputs[327];
    assign layer0_outputs[7565] = (inputs[758]) & ~(inputs[962]);
    assign layer0_outputs[7566] = (inputs[128]) ^ (inputs[790]);
    assign layer0_outputs[7567] = ~(inputs[570]) | (inputs[224]);
    assign layer0_outputs[7568] = inputs[134];
    assign layer0_outputs[7569] = ~((inputs[140]) | (inputs[447]));
    assign layer0_outputs[7570] = (inputs[556]) & ~(inputs[443]);
    assign layer0_outputs[7571] = (inputs[251]) | (inputs[710]);
    assign layer0_outputs[7572] = (inputs[209]) | (inputs[610]);
    assign layer0_outputs[7573] = ~((inputs[776]) ^ (inputs[57]));
    assign layer0_outputs[7574] = ~((inputs[405]) | (inputs[178]));
    assign layer0_outputs[7575] = inputs[668];
    assign layer0_outputs[7576] = (inputs[33]) & ~(inputs[747]);
    assign layer0_outputs[7577] = ~(inputs[404]);
    assign layer0_outputs[7578] = (inputs[810]) & ~(inputs[647]);
    assign layer0_outputs[7579] = ~(inputs[688]) | (inputs[516]);
    assign layer0_outputs[7580] = ~((inputs[403]) ^ (inputs[767]));
    assign layer0_outputs[7581] = inputs[864];
    assign layer0_outputs[7582] = ~(inputs[625]);
    assign layer0_outputs[7583] = ~(inputs[624]) | (inputs[934]);
    assign layer0_outputs[7584] = (inputs[519]) ^ (inputs[427]);
    assign layer0_outputs[7585] = (inputs[902]) ^ (inputs[12]);
    assign layer0_outputs[7586] = (inputs[49]) | (inputs[462]);
    assign layer0_outputs[7587] = ~((inputs[209]) | (inputs[144]));
    assign layer0_outputs[7588] = ~(inputs[267]);
    assign layer0_outputs[7589] = ~((inputs[933]) | (inputs[445]));
    assign layer0_outputs[7590] = ~(inputs[861]);
    assign layer0_outputs[7591] = (inputs[664]) & (inputs[638]);
    assign layer0_outputs[7592] = inputs[191];
    assign layer0_outputs[7593] = inputs[715];
    assign layer0_outputs[7594] = (inputs[605]) | (inputs[560]);
    assign layer0_outputs[7595] = ~((inputs[200]) & (inputs[414]));
    assign layer0_outputs[7596] = ~(inputs[349]) | (inputs[572]);
    assign layer0_outputs[7597] = inputs[432];
    assign layer0_outputs[7598] = inputs[597];
    assign layer0_outputs[7599] = ~((inputs[345]) | (inputs[798]));
    assign layer0_outputs[7600] = ~((inputs[656]) | (inputs[32]));
    assign layer0_outputs[7601] = inputs[558];
    assign layer0_outputs[7602] = ~(inputs[98]);
    assign layer0_outputs[7603] = inputs[389];
    assign layer0_outputs[7604] = ~((inputs[583]) | (inputs[338]));
    assign layer0_outputs[7605] = (inputs[125]) | (inputs[918]);
    assign layer0_outputs[7606] = (inputs[351]) & ~(inputs[259]);
    assign layer0_outputs[7607] = (inputs[779]) & (inputs[376]);
    assign layer0_outputs[7608] = (inputs[527]) & ~(inputs[37]);
    assign layer0_outputs[7609] = ~(inputs[159]);
    assign layer0_outputs[7610] = (inputs[796]) ^ (inputs[747]);
    assign layer0_outputs[7611] = (inputs[926]) | (inputs[524]);
    assign layer0_outputs[7612] = ~((inputs[550]) ^ (inputs[553]));
    assign layer0_outputs[7613] = ~((inputs[911]) | (inputs[4]));
    assign layer0_outputs[7614] = ~(inputs[763]);
    assign layer0_outputs[7615] = ~((inputs[382]) ^ (inputs[184]));
    assign layer0_outputs[7616] = (inputs[794]) | (inputs[240]);
    assign layer0_outputs[7617] = (inputs[127]) ^ (inputs[326]);
    assign layer0_outputs[7618] = (inputs[998]) ^ (inputs[704]);
    assign layer0_outputs[7619] = (inputs[779]) | (inputs[580]);
    assign layer0_outputs[7620] = (inputs[595]) & ~(inputs[462]);
    assign layer0_outputs[7621] = ~(inputs[375]) | (inputs[147]);
    assign layer0_outputs[7622] = ~(inputs[88]) | (inputs[993]);
    assign layer0_outputs[7623] = ~(inputs[780]) | (inputs[990]);
    assign layer0_outputs[7624] = (inputs[359]) ^ (inputs[649]);
    assign layer0_outputs[7625] = inputs[401];
    assign layer0_outputs[7626] = (inputs[645]) ^ (inputs[769]);
    assign layer0_outputs[7627] = (inputs[480]) & ~(inputs[502]);
    assign layer0_outputs[7628] = ~(inputs[403]) | (inputs[698]);
    assign layer0_outputs[7629] = ~((inputs[911]) | (inputs[844]));
    assign layer0_outputs[7630] = inputs[527];
    assign layer0_outputs[7631] = ~(inputs[230]) | (inputs[1021]);
    assign layer0_outputs[7632] = ~((inputs[523]) ^ (inputs[549]));
    assign layer0_outputs[7633] = ~((inputs[856]) | (inputs[876]));
    assign layer0_outputs[7634] = ~(inputs[316]) | (inputs[1011]);
    assign layer0_outputs[7635] = 1'b0;
    assign layer0_outputs[7636] = (inputs[393]) | (inputs[713]);
    assign layer0_outputs[7637] = inputs[714];
    assign layer0_outputs[7638] = (inputs[235]) ^ (inputs[344]);
    assign layer0_outputs[7639] = (inputs[974]) & ~(inputs[865]);
    assign layer0_outputs[7640] = ~(inputs[384]) | (inputs[104]);
    assign layer0_outputs[7641] = inputs[430];
    assign layer0_outputs[7642] = ~(inputs[743]);
    assign layer0_outputs[7643] = (inputs[555]) | (inputs[767]);
    assign layer0_outputs[7644] = ~(inputs[868]) | (inputs[890]);
    assign layer0_outputs[7645] = ~(inputs[689]) | (inputs[818]);
    assign layer0_outputs[7646] = (inputs[10]) ^ (inputs[295]);
    assign layer0_outputs[7647] = ~(inputs[171]) | (inputs[330]);
    assign layer0_outputs[7648] = (inputs[864]) ^ (inputs[744]);
    assign layer0_outputs[7649] = inputs[588];
    assign layer0_outputs[7650] = ~((inputs[507]) | (inputs[828]));
    assign layer0_outputs[7651] = ~((inputs[548]) | (inputs[739]));
    assign layer0_outputs[7652] = ~((inputs[402]) ^ (inputs[800]));
    assign layer0_outputs[7653] = inputs[316];
    assign layer0_outputs[7654] = (inputs[1005]) & (inputs[773]);
    assign layer0_outputs[7655] = 1'b1;
    assign layer0_outputs[7656] = (inputs[613]) | (inputs[241]);
    assign layer0_outputs[7657] = (inputs[478]) ^ (inputs[338]);
    assign layer0_outputs[7658] = inputs[326];
    assign layer0_outputs[7659] = ~((inputs[176]) | (inputs[920]));
    assign layer0_outputs[7660] = inputs[425];
    assign layer0_outputs[7661] = ~(inputs[361]) | (inputs[886]);
    assign layer0_outputs[7662] = (inputs[476]) | (inputs[357]);
    assign layer0_outputs[7663] = ~((inputs[897]) | (inputs[247]));
    assign layer0_outputs[7664] = (inputs[643]) & ~(inputs[12]);
    assign layer0_outputs[7665] = ~((inputs[786]) ^ (inputs[370]));
    assign layer0_outputs[7666] = ~((inputs[461]) ^ (inputs[385]));
    assign layer0_outputs[7667] = (inputs[170]) | (inputs[973]);
    assign layer0_outputs[7668] = inputs[879];
    assign layer0_outputs[7669] = (inputs[295]) | (inputs[268]);
    assign layer0_outputs[7670] = ~(inputs[415]) | (inputs[930]);
    assign layer0_outputs[7671] = (inputs[164]) ^ (inputs[590]);
    assign layer0_outputs[7672] = 1'b1;
    assign layer0_outputs[7673] = (inputs[712]) ^ (inputs[37]);
    assign layer0_outputs[7674] = (inputs[352]) & ~(inputs[1013]);
    assign layer0_outputs[7675] = ~((inputs[293]) | (inputs[71]));
    assign layer0_outputs[7676] = 1'b1;
    assign layer0_outputs[7677] = ~(inputs[426]);
    assign layer0_outputs[7678] = (inputs[771]) | (inputs[82]);
    assign layer0_outputs[7679] = inputs[889];
    assign layer0_outputs[7680] = ~((inputs[665]) | (inputs[206]));
    assign layer0_outputs[7681] = (inputs[236]) ^ (inputs[239]);
    assign layer0_outputs[7682] = ~(inputs[522]) | (inputs[140]);
    assign layer0_outputs[7683] = (inputs[560]) & ~(inputs[992]);
    assign layer0_outputs[7684] = (inputs[577]) & ~(inputs[182]);
    assign layer0_outputs[7685] = (inputs[836]) & (inputs[946]);
    assign layer0_outputs[7686] = (inputs[832]) ^ (inputs[625]);
    assign layer0_outputs[7687] = ~((inputs[36]) | (inputs[930]));
    assign layer0_outputs[7688] = inputs[752];
    assign layer0_outputs[7689] = ~(inputs[482]);
    assign layer0_outputs[7690] = inputs[999];
    assign layer0_outputs[7691] = ~((inputs[32]) ^ (inputs[918]));
    assign layer0_outputs[7692] = ~((inputs[394]) | (inputs[36]));
    assign layer0_outputs[7693] = ~(inputs[273]) | (inputs[71]);
    assign layer0_outputs[7694] = ~(inputs[927]) | (inputs[612]);
    assign layer0_outputs[7695] = (inputs[917]) & ~(inputs[79]);
    assign layer0_outputs[7696] = ~((inputs[854]) | (inputs[206]));
    assign layer0_outputs[7697] = inputs[567];
    assign layer0_outputs[7698] = ~(inputs[657]);
    assign layer0_outputs[7699] = ~(inputs[938]) | (inputs[153]);
    assign layer0_outputs[7700] = inputs[305];
    assign layer0_outputs[7701] = ~(inputs[754]) | (inputs[262]);
    assign layer0_outputs[7702] = 1'b0;
    assign layer0_outputs[7703] = (inputs[661]) ^ (inputs[164]);
    assign layer0_outputs[7704] = (inputs[880]) | (inputs[981]);
    assign layer0_outputs[7705] = (inputs[863]) & (inputs[734]);
    assign layer0_outputs[7706] = ~((inputs[362]) | (inputs[15]));
    assign layer0_outputs[7707] = ~(inputs[547]) | (inputs[106]);
    assign layer0_outputs[7708] = (inputs[630]) & ~(inputs[828]);
    assign layer0_outputs[7709] = (inputs[10]) | (inputs[214]);
    assign layer0_outputs[7710] = ~(inputs[175]);
    assign layer0_outputs[7711] = ~(inputs[570]);
    assign layer0_outputs[7712] = ~((inputs[42]) | (inputs[132]));
    assign layer0_outputs[7713] = ~(inputs[688]);
    assign layer0_outputs[7714] = ~(inputs[781]);
    assign layer0_outputs[7715] = (inputs[194]) & (inputs[954]);
    assign layer0_outputs[7716] = (inputs[397]) & ~(inputs[573]);
    assign layer0_outputs[7717] = (inputs[522]) ^ (inputs[141]);
    assign layer0_outputs[7718] = inputs[369];
    assign layer0_outputs[7719] = inputs[573];
    assign layer0_outputs[7720] = ~(inputs[729]);
    assign layer0_outputs[7721] = inputs[636];
    assign layer0_outputs[7722] = ~((inputs[422]) ^ (inputs[639]));
    assign layer0_outputs[7723] = inputs[118];
    assign layer0_outputs[7724] = (inputs[776]) & ~(inputs[46]);
    assign layer0_outputs[7725] = ~(inputs[996]);
    assign layer0_outputs[7726] = ~(inputs[685]);
    assign layer0_outputs[7727] = ~((inputs[890]) ^ (inputs[583]));
    assign layer0_outputs[7728] = ~((inputs[299]) & (inputs[447]));
    assign layer0_outputs[7729] = inputs[570];
    assign layer0_outputs[7730] = ~((inputs[879]) | (inputs[451]));
    assign layer0_outputs[7731] = (inputs[327]) & ~(inputs[613]);
    assign layer0_outputs[7732] = inputs[850];
    assign layer0_outputs[7733] = inputs[619];
    assign layer0_outputs[7734] = ~(inputs[281]);
    assign layer0_outputs[7735] = (inputs[846]) & ~(inputs[132]);
    assign layer0_outputs[7736] = ~((inputs[685]) ^ (inputs[697]));
    assign layer0_outputs[7737] = ~(inputs[712]);
    assign layer0_outputs[7738] = ~(inputs[170]) | (inputs[511]);
    assign layer0_outputs[7739] = ~((inputs[75]) & (inputs[703]));
    assign layer0_outputs[7740] = ~(inputs[291]) | (inputs[407]);
    assign layer0_outputs[7741] = ~(inputs[236]) | (inputs[319]);
    assign layer0_outputs[7742] = (inputs[327]) ^ (inputs[426]);
    assign layer0_outputs[7743] = inputs[814];
    assign layer0_outputs[7744] = (inputs[607]) & ~(inputs[721]);
    assign layer0_outputs[7745] = ~(inputs[365]);
    assign layer0_outputs[7746] = (inputs[165]) & (inputs[1000]);
    assign layer0_outputs[7747] = ~((inputs[583]) ^ (inputs[257]));
    assign layer0_outputs[7748] = ~(inputs[898]) | (inputs[958]);
    assign layer0_outputs[7749] = ~((inputs[738]) ^ (inputs[51]));
    assign layer0_outputs[7750] = (inputs[773]) & ~(inputs[84]);
    assign layer0_outputs[7751] = inputs[912];
    assign layer0_outputs[7752] = ~(inputs[302]);
    assign layer0_outputs[7753] = ~(inputs[479]) | (inputs[81]);
    assign layer0_outputs[7754] = (inputs[782]) & ~(inputs[859]);
    assign layer0_outputs[7755] = ~((inputs[441]) ^ (inputs[313]));
    assign layer0_outputs[7756] = ~(inputs[1]);
    assign layer0_outputs[7757] = (inputs[136]) & ~(inputs[103]);
    assign layer0_outputs[7758] = ~((inputs[229]) | (inputs[827]));
    assign layer0_outputs[7759] = ~(inputs[378]);
    assign layer0_outputs[7760] = ~((inputs[343]) ^ (inputs[1019]));
    assign layer0_outputs[7761] = inputs[997];
    assign layer0_outputs[7762] = ~(inputs[491]) | (inputs[361]);
    assign layer0_outputs[7763] = ~(inputs[566]) | (inputs[1009]);
    assign layer0_outputs[7764] = (inputs[208]) | (inputs[1009]);
    assign layer0_outputs[7765] = inputs[393];
    assign layer0_outputs[7766] = ~((inputs[787]) | (inputs[801]));
    assign layer0_outputs[7767] = ~(inputs[76]);
    assign layer0_outputs[7768] = inputs[440];
    assign layer0_outputs[7769] = ~((inputs[617]) | (inputs[612]));
    assign layer0_outputs[7770] = inputs[844];
    assign layer0_outputs[7771] = ~(inputs[149]) | (inputs[965]);
    assign layer0_outputs[7772] = (inputs[0]) | (inputs[791]);
    assign layer0_outputs[7773] = inputs[22];
    assign layer0_outputs[7774] = (inputs[58]) ^ (inputs[765]);
    assign layer0_outputs[7775] = (inputs[137]) | (inputs[155]);
    assign layer0_outputs[7776] = ~(inputs[903]) | (inputs[821]);
    assign layer0_outputs[7777] = (inputs[54]) & ~(inputs[899]);
    assign layer0_outputs[7778] = ~((inputs[664]) ^ (inputs[741]));
    assign layer0_outputs[7779] = ~((inputs[160]) & (inputs[719]));
    assign layer0_outputs[7780] = ~(inputs[813]);
    assign layer0_outputs[7781] = (inputs[261]) ^ (inputs[165]);
    assign layer0_outputs[7782] = (inputs[59]) & ~(inputs[993]);
    assign layer0_outputs[7783] = ~((inputs[1021]) | (inputs[671]));
    assign layer0_outputs[7784] = ~(inputs[755]) | (inputs[1017]);
    assign layer0_outputs[7785] = ~(inputs[881]) | (inputs[315]);
    assign layer0_outputs[7786] = (inputs[939]) | (inputs[163]);
    assign layer0_outputs[7787] = (inputs[101]) ^ (inputs[28]);
    assign layer0_outputs[7788] = (inputs[529]) & ~(inputs[76]);
    assign layer0_outputs[7789] = (inputs[298]) | (inputs[188]);
    assign layer0_outputs[7790] = inputs[759];
    assign layer0_outputs[7791] = (inputs[499]) & ~(inputs[794]);
    assign layer0_outputs[7792] = ~((inputs[172]) ^ (inputs[560]));
    assign layer0_outputs[7793] = ~(inputs[902]);
    assign layer0_outputs[7794] = inputs[208];
    assign layer0_outputs[7795] = inputs[900];
    assign layer0_outputs[7796] = ~(inputs[862]);
    assign layer0_outputs[7797] = (inputs[799]) & ~(inputs[834]);
    assign layer0_outputs[7798] = 1'b0;
    assign layer0_outputs[7799] = ~(inputs[437]) | (inputs[665]);
    assign layer0_outputs[7800] = ~((inputs[695]) & (inputs[567]));
    assign layer0_outputs[7801] = (inputs[662]) & ~(inputs[547]);
    assign layer0_outputs[7802] = inputs[776];
    assign layer0_outputs[7803] = ~((inputs[581]) | (inputs[631]));
    assign layer0_outputs[7804] = (inputs[798]) ^ (inputs[171]);
    assign layer0_outputs[7805] = inputs[929];
    assign layer0_outputs[7806] = ~(inputs[10]) | (inputs[168]);
    assign layer0_outputs[7807] = ~(inputs[787]);
    assign layer0_outputs[7808] = ~((inputs[387]) ^ (inputs[496]));
    assign layer0_outputs[7809] = ~(inputs[564]);
    assign layer0_outputs[7810] = (inputs[890]) & ~(inputs[784]);
    assign layer0_outputs[7811] = ~((inputs[736]) & (inputs[94]));
    assign layer0_outputs[7812] = inputs[172];
    assign layer0_outputs[7813] = ~((inputs[190]) ^ (inputs[637]));
    assign layer0_outputs[7814] = (inputs[2]) | (inputs[949]);
    assign layer0_outputs[7815] = ~((inputs[402]) ^ (inputs[31]));
    assign layer0_outputs[7816] = ~(inputs[9]);
    assign layer0_outputs[7817] = (inputs[847]) & ~(inputs[111]);
    assign layer0_outputs[7818] = ~(inputs[447]);
    assign layer0_outputs[7819] = ~(inputs[698]);
    assign layer0_outputs[7820] = ~(inputs[650]) | (inputs[744]);
    assign layer0_outputs[7821] = (inputs[1022]) ^ (inputs[826]);
    assign layer0_outputs[7822] = ~((inputs[323]) ^ (inputs[784]));
    assign layer0_outputs[7823] = ~((inputs[134]) ^ (inputs[837]));
    assign layer0_outputs[7824] = ~(inputs[998]);
    assign layer0_outputs[7825] = (inputs[709]) ^ (inputs[477]);
    assign layer0_outputs[7826] = (inputs[567]) | (inputs[531]);
    assign layer0_outputs[7827] = ~(inputs[884]);
    assign layer0_outputs[7828] = inputs[144];
    assign layer0_outputs[7829] = ~(inputs[835]) | (inputs[854]);
    assign layer0_outputs[7830] = inputs[696];
    assign layer0_outputs[7831] = (inputs[296]) ^ (inputs[373]);
    assign layer0_outputs[7832] = ~(inputs[731]);
    assign layer0_outputs[7833] = ~(inputs[430]);
    assign layer0_outputs[7834] = 1'b1;
    assign layer0_outputs[7835] = ~((inputs[556]) | (inputs[233]));
    assign layer0_outputs[7836] = ~((inputs[468]) | (inputs[971]));
    assign layer0_outputs[7837] = (inputs[121]) & (inputs[994]);
    assign layer0_outputs[7838] = ~(inputs[149]);
    assign layer0_outputs[7839] = ~(inputs[597]) | (inputs[31]);
    assign layer0_outputs[7840] = 1'b0;
    assign layer0_outputs[7841] = (inputs[335]) & ~(inputs[699]);
    assign layer0_outputs[7842] = inputs[916];
    assign layer0_outputs[7843] = inputs[201];
    assign layer0_outputs[7844] = ~(inputs[618]) | (inputs[793]);
    assign layer0_outputs[7845] = (inputs[909]) | (inputs[306]);
    assign layer0_outputs[7846] = ~(inputs[550]);
    assign layer0_outputs[7847] = ~((inputs[976]) | (inputs[661]));
    assign layer0_outputs[7848] = (inputs[365]) & ~(inputs[41]);
    assign layer0_outputs[7849] = ~(inputs[24]);
    assign layer0_outputs[7850] = ~(inputs[437]) | (inputs[635]);
    assign layer0_outputs[7851] = ~(inputs[260]) | (inputs[254]);
    assign layer0_outputs[7852] = ~(inputs[761]);
    assign layer0_outputs[7853] = (inputs[388]) & ~(inputs[380]);
    assign layer0_outputs[7854] = ~((inputs[694]) | (inputs[479]));
    assign layer0_outputs[7855] = (inputs[853]) & (inputs[908]);
    assign layer0_outputs[7856] = (inputs[638]) ^ (inputs[98]);
    assign layer0_outputs[7857] = ~(inputs[630]);
    assign layer0_outputs[7858] = ~(inputs[598]) | (inputs[837]);
    assign layer0_outputs[7859] = (inputs[753]) & ~(inputs[336]);
    assign layer0_outputs[7860] = ~(inputs[314]) | (inputs[449]);
    assign layer0_outputs[7861] = (inputs[771]) & ~(inputs[875]);
    assign layer0_outputs[7862] = ~((inputs[979]) | (inputs[635]));
    assign layer0_outputs[7863] = inputs[923];
    assign layer0_outputs[7864] = ~(inputs[158]) | (inputs[516]);
    assign layer0_outputs[7865] = ~(inputs[584]);
    assign layer0_outputs[7866] = ~((inputs[163]) ^ (inputs[482]));
    assign layer0_outputs[7867] = ~(inputs[264]);
    assign layer0_outputs[7868] = (inputs[303]) & ~(inputs[829]);
    assign layer0_outputs[7869] = inputs[813];
    assign layer0_outputs[7870] = inputs[413];
    assign layer0_outputs[7871] = (inputs[994]) ^ (inputs[619]);
    assign layer0_outputs[7872] = ~(inputs[441]) | (inputs[896]);
    assign layer0_outputs[7873] = ~((inputs[441]) ^ (inputs[799]));
    assign layer0_outputs[7874] = ~(inputs[440]);
    assign layer0_outputs[7875] = ~((inputs[358]) | (inputs[548]));
    assign layer0_outputs[7876] = inputs[369];
    assign layer0_outputs[7877] = ~((inputs[553]) | (inputs[583]));
    assign layer0_outputs[7878] = (inputs[488]) | (inputs[346]);
    assign layer0_outputs[7879] = (inputs[530]) ^ (inputs[740]);
    assign layer0_outputs[7880] = inputs[422];
    assign layer0_outputs[7881] = ~((inputs[656]) | (inputs[150]));
    assign layer0_outputs[7882] = ~((inputs[860]) | (inputs[486]));
    assign layer0_outputs[7883] = inputs[755];
    assign layer0_outputs[7884] = ~((inputs[290]) & (inputs[735]));
    assign layer0_outputs[7885] = ~(inputs[983]) | (inputs[418]);
    assign layer0_outputs[7886] = ~(inputs[26]) | (inputs[381]);
    assign layer0_outputs[7887] = ~(inputs[420]);
    assign layer0_outputs[7888] = inputs[913];
    assign layer0_outputs[7889] = 1'b0;
    assign layer0_outputs[7890] = ~((inputs[758]) | (inputs[772]));
    assign layer0_outputs[7891] = inputs[530];
    assign layer0_outputs[7892] = inputs[847];
    assign layer0_outputs[7893] = ~((inputs[396]) ^ (inputs[948]));
    assign layer0_outputs[7894] = ~(inputs[241]) | (inputs[833]);
    assign layer0_outputs[7895] = ~((inputs[371]) | (inputs[105]));
    assign layer0_outputs[7896] = ~(inputs[654]);
    assign layer0_outputs[7897] = 1'b0;
    assign layer0_outputs[7898] = 1'b1;
    assign layer0_outputs[7899] = inputs[623];
    assign layer0_outputs[7900] = ~(inputs[653]) | (inputs[697]);
    assign layer0_outputs[7901] = (inputs[59]) | (inputs[549]);
    assign layer0_outputs[7902] = (inputs[886]) | (inputs[335]);
    assign layer0_outputs[7903] = inputs[852];
    assign layer0_outputs[7904] = 1'b1;
    assign layer0_outputs[7905] = ~(inputs[393]);
    assign layer0_outputs[7906] = (inputs[913]) & ~(inputs[192]);
    assign layer0_outputs[7907] = ~(inputs[399]) | (inputs[90]);
    assign layer0_outputs[7908] = (inputs[37]) & ~(inputs[802]);
    assign layer0_outputs[7909] = ~((inputs[300]) | (inputs[563]));
    assign layer0_outputs[7910] = ~(inputs[677]);
    assign layer0_outputs[7911] = ~(inputs[748]);
    assign layer0_outputs[7912] = inputs[472];
    assign layer0_outputs[7913] = ~(inputs[437]);
    assign layer0_outputs[7914] = ~(inputs[427]);
    assign layer0_outputs[7915] = inputs[23];
    assign layer0_outputs[7916] = ~(inputs[214]) | (inputs[601]);
    assign layer0_outputs[7917] = (inputs[813]) & ~(inputs[390]);
    assign layer0_outputs[7918] = (inputs[555]) & ~(inputs[971]);
    assign layer0_outputs[7919] = inputs[653];
    assign layer0_outputs[7920] = ~((inputs[563]) | (inputs[310]));
    assign layer0_outputs[7921] = ~(inputs[200]) | (inputs[354]);
    assign layer0_outputs[7922] = ~(inputs[202]);
    assign layer0_outputs[7923] = ~((inputs[417]) ^ (inputs[754]));
    assign layer0_outputs[7924] = 1'b0;
    assign layer0_outputs[7925] = ~(inputs[966]) | (inputs[270]);
    assign layer0_outputs[7926] = inputs[699];
    assign layer0_outputs[7927] = (inputs[685]) ^ (inputs[431]);
    assign layer0_outputs[7928] = ~((inputs[904]) | (inputs[394]));
    assign layer0_outputs[7929] = ~(inputs[650]);
    assign layer0_outputs[7930] = inputs[884];
    assign layer0_outputs[7931] = ~(inputs[784]) | (inputs[252]);
    assign layer0_outputs[7932] = ~((inputs[138]) ^ (inputs[581]));
    assign layer0_outputs[7933] = ~(inputs[583]);
    assign layer0_outputs[7934] = ~(inputs[889]);
    assign layer0_outputs[7935] = (inputs[503]) & ~(inputs[157]);
    assign layer0_outputs[7936] = 1'b1;
    assign layer0_outputs[7937] = ~((inputs[715]) | (inputs[802]));
    assign layer0_outputs[7938] = (inputs[468]) ^ (inputs[386]);
    assign layer0_outputs[7939] = (inputs[748]) & ~(inputs[861]);
    assign layer0_outputs[7940] = ~((inputs[141]) | (inputs[172]));
    assign layer0_outputs[7941] = ~((inputs[880]) | (inputs[405]));
    assign layer0_outputs[7942] = ~(inputs[242]) | (inputs[506]);
    assign layer0_outputs[7943] = ~((inputs[626]) | (inputs[137]));
    assign layer0_outputs[7944] = (inputs[788]) ^ (inputs[321]);
    assign layer0_outputs[7945] = (inputs[453]) | (inputs[571]);
    assign layer0_outputs[7946] = ~(inputs[738]) | (inputs[642]);
    assign layer0_outputs[7947] = ~(inputs[618]);
    assign layer0_outputs[7948] = (inputs[804]) | (inputs[785]);
    assign layer0_outputs[7949] = ~(inputs[439]);
    assign layer0_outputs[7950] = inputs[569];
    assign layer0_outputs[7951] = (inputs[509]) | (inputs[243]);
    assign layer0_outputs[7952] = (inputs[397]) & ~(inputs[206]);
    assign layer0_outputs[7953] = inputs[420];
    assign layer0_outputs[7954] = ~(inputs[822]) | (inputs[570]);
    assign layer0_outputs[7955] = ~((inputs[920]) ^ (inputs[251]));
    assign layer0_outputs[7956] = (inputs[172]) ^ (inputs[933]);
    assign layer0_outputs[7957] = ~(inputs[38]);
    assign layer0_outputs[7958] = inputs[572];
    assign layer0_outputs[7959] = inputs[398];
    assign layer0_outputs[7960] = ~((inputs[986]) ^ (inputs[486]));
    assign layer0_outputs[7961] = ~((inputs[852]) | (inputs[825]));
    assign layer0_outputs[7962] = ~(inputs[885]) | (inputs[226]);
    assign layer0_outputs[7963] = (inputs[542]) & ~(inputs[9]);
    assign layer0_outputs[7964] = 1'b0;
    assign layer0_outputs[7965] = (inputs[931]) & ~(inputs[67]);
    assign layer0_outputs[7966] = (inputs[12]) | (inputs[425]);
    assign layer0_outputs[7967] = (inputs[284]) | (inputs[694]);
    assign layer0_outputs[7968] = inputs[465];
    assign layer0_outputs[7969] = (inputs[405]) & ~(inputs[206]);
    assign layer0_outputs[7970] = (inputs[822]) & ~(inputs[57]);
    assign layer0_outputs[7971] = (inputs[523]) & ~(inputs[841]);
    assign layer0_outputs[7972] = ~(inputs[560]) | (inputs[1011]);
    assign layer0_outputs[7973] = ~(inputs[236]);
    assign layer0_outputs[7974] = (inputs[724]) & ~(inputs[221]);
    assign layer0_outputs[7975] = ~((inputs[995]) & (inputs[190]));
    assign layer0_outputs[7976] = ~(inputs[469]) | (inputs[777]);
    assign layer0_outputs[7977] = inputs[36];
    assign layer0_outputs[7978] = (inputs[171]) | (inputs[856]);
    assign layer0_outputs[7979] = ~(inputs[746]) | (inputs[129]);
    assign layer0_outputs[7980] = inputs[371];
    assign layer0_outputs[7981] = ~(inputs[461]);
    assign layer0_outputs[7982] = ~(inputs[208]) | (inputs[946]);
    assign layer0_outputs[7983] = inputs[212];
    assign layer0_outputs[7984] = inputs[242];
    assign layer0_outputs[7985] = (inputs[1]) & ~(inputs[351]);
    assign layer0_outputs[7986] = ~(inputs[574]);
    assign layer0_outputs[7987] = ~(inputs[618]) | (inputs[780]);
    assign layer0_outputs[7988] = ~(inputs[645]) | (inputs[1004]);
    assign layer0_outputs[7989] = ~(inputs[331]);
    assign layer0_outputs[7990] = inputs[873];
    assign layer0_outputs[7991] = ~((inputs[932]) ^ (inputs[691]));
    assign layer0_outputs[7992] = (inputs[665]) & ~(inputs[32]);
    assign layer0_outputs[7993] = ~((inputs[525]) | (inputs[253]));
    assign layer0_outputs[7994] = 1'b0;
    assign layer0_outputs[7995] = ~(inputs[401]) | (inputs[572]);
    assign layer0_outputs[7996] = inputs[389];
    assign layer0_outputs[7997] = (inputs[118]) & ~(inputs[19]);
    assign layer0_outputs[7998] = ~((inputs[297]) | (inputs[312]));
    assign layer0_outputs[7999] = 1'b1;
    assign layer0_outputs[8000] = inputs[462];
    assign layer0_outputs[8001] = (inputs[101]) ^ (inputs[216]);
    assign layer0_outputs[8002] = (inputs[659]) & ~(inputs[433]);
    assign layer0_outputs[8003] = inputs[785];
    assign layer0_outputs[8004] = inputs[506];
    assign layer0_outputs[8005] = 1'b1;
    assign layer0_outputs[8006] = ~((inputs[923]) | (inputs[621]));
    assign layer0_outputs[8007] = ~(inputs[577]);
    assign layer0_outputs[8008] = (inputs[649]) | (inputs[999]);
    assign layer0_outputs[8009] = (inputs[470]) ^ (inputs[299]);
    assign layer0_outputs[8010] = (inputs[590]) & ~(inputs[844]);
    assign layer0_outputs[8011] = inputs[951];
    assign layer0_outputs[8012] = (inputs[170]) | (inputs[662]);
    assign layer0_outputs[8013] = ~((inputs[39]) ^ (inputs[310]));
    assign layer0_outputs[8014] = ~(inputs[390]) | (inputs[919]);
    assign layer0_outputs[8015] = (inputs[815]) & ~(inputs[89]);
    assign layer0_outputs[8016] = inputs[719];
    assign layer0_outputs[8017] = inputs[502];
    assign layer0_outputs[8018] = ~((inputs[294]) ^ (inputs[648]));
    assign layer0_outputs[8019] = (inputs[727]) | (inputs[710]);
    assign layer0_outputs[8020] = (inputs[597]) & ~(inputs[75]);
    assign layer0_outputs[8021] = (inputs[129]) | (inputs[901]);
    assign layer0_outputs[8022] = ~(inputs[658]) | (inputs[805]);
    assign layer0_outputs[8023] = 1'b1;
    assign layer0_outputs[8024] = (inputs[523]) & ~(inputs[118]);
    assign layer0_outputs[8025] = inputs[679];
    assign layer0_outputs[8026] = ~((inputs[72]) | (inputs[913]));
    assign layer0_outputs[8027] = (inputs[586]) | (inputs[470]);
    assign layer0_outputs[8028] = (inputs[944]) ^ (inputs[905]);
    assign layer0_outputs[8029] = (inputs[289]) | (inputs[50]);
    assign layer0_outputs[8030] = ~(inputs[342]) | (inputs[892]);
    assign layer0_outputs[8031] = ~(inputs[5]);
    assign layer0_outputs[8032] = (inputs[559]) | (inputs[259]);
    assign layer0_outputs[8033] = inputs[275];
    assign layer0_outputs[8034] = ~((inputs[680]) | (inputs[939]));
    assign layer0_outputs[8035] = inputs[735];
    assign layer0_outputs[8036] = ~((inputs[635]) ^ (inputs[1021]));
    assign layer0_outputs[8037] = ~(inputs[753]);
    assign layer0_outputs[8038] = ~(inputs[722]);
    assign layer0_outputs[8039] = 1'b1;
    assign layer0_outputs[8040] = ~(inputs[191]) | (inputs[95]);
    assign layer0_outputs[8041] = ~((inputs[117]) ^ (inputs[335]));
    assign layer0_outputs[8042] = (inputs[421]) | (inputs[433]);
    assign layer0_outputs[8043] = inputs[456];
    assign layer0_outputs[8044] = (inputs[600]) & ~(inputs[382]);
    assign layer0_outputs[8045] = ~(inputs[570]);
    assign layer0_outputs[8046] = ~(inputs[241]);
    assign layer0_outputs[8047] = (inputs[869]) & (inputs[385]);
    assign layer0_outputs[8048] = ~(inputs[201]);
    assign layer0_outputs[8049] = (inputs[356]) | (inputs[110]);
    assign layer0_outputs[8050] = ~(inputs[302]);
    assign layer0_outputs[8051] = inputs[679];
    assign layer0_outputs[8052] = (inputs[742]) & ~(inputs[857]);
    assign layer0_outputs[8053] = ~(inputs[808]) | (inputs[127]);
    assign layer0_outputs[8054] = ~((inputs[988]) & (inputs[254]));
    assign layer0_outputs[8055] = ~(inputs[809]);
    assign layer0_outputs[8056] = 1'b1;
    assign layer0_outputs[8057] = inputs[456];
    assign layer0_outputs[8058] = ~(inputs[685]);
    assign layer0_outputs[8059] = ~((inputs[328]) ^ (inputs[147]));
    assign layer0_outputs[8060] = ~(inputs[913]) | (inputs[859]);
    assign layer0_outputs[8061] = ~((inputs[589]) ^ (inputs[634]));
    assign layer0_outputs[8062] = inputs[885];
    assign layer0_outputs[8063] = ~((inputs[943]) & (inputs[596]));
    assign layer0_outputs[8064] = inputs[212];
    assign layer0_outputs[8065] = ~((inputs[787]) & (inputs[356]));
    assign layer0_outputs[8066] = (inputs[840]) ^ (inputs[684]);
    assign layer0_outputs[8067] = (inputs[33]) & ~(inputs[829]);
    assign layer0_outputs[8068] = (inputs[181]) ^ (inputs[211]);
    assign layer0_outputs[8069] = inputs[267];
    assign layer0_outputs[8070] = (inputs[703]) | (inputs[514]);
    assign layer0_outputs[8071] = ~((inputs[623]) & (inputs[479]));
    assign layer0_outputs[8072] = ~(inputs[182]) | (inputs[293]);
    assign layer0_outputs[8073] = ~(inputs[88]);
    assign layer0_outputs[8074] = ~(inputs[512]) | (inputs[197]);
    assign layer0_outputs[8075] = ~((inputs[891]) ^ (inputs[566]));
    assign layer0_outputs[8076] = (inputs[752]) & ~(inputs[472]);
    assign layer0_outputs[8077] = inputs[638];
    assign layer0_outputs[8078] = ~((inputs[218]) & (inputs[70]));
    assign layer0_outputs[8079] = ~(inputs[52]) | (inputs[834]);
    assign layer0_outputs[8080] = (inputs[461]) & ~(inputs[1007]);
    assign layer0_outputs[8081] = ~(inputs[646]) | (inputs[580]);
    assign layer0_outputs[8082] = ~(inputs[391]);
    assign layer0_outputs[8083] = (inputs[550]) ^ (inputs[979]);
    assign layer0_outputs[8084] = (inputs[974]) | (inputs[508]);
    assign layer0_outputs[8085] = ~((inputs[69]) | (inputs[455]));
    assign layer0_outputs[8086] = ~(inputs[590]) | (inputs[158]);
    assign layer0_outputs[8087] = ~(inputs[745]) | (inputs[910]);
    assign layer0_outputs[8088] = 1'b0;
    assign layer0_outputs[8089] = ~((inputs[600]) ^ (inputs[992]));
    assign layer0_outputs[8090] = ~((inputs[483]) | (inputs[886]));
    assign layer0_outputs[8091] = ~((inputs[240]) | (inputs[85]));
    assign layer0_outputs[8092] = inputs[677];
    assign layer0_outputs[8093] = 1'b1;
    assign layer0_outputs[8094] = ~(inputs[880]);
    assign layer0_outputs[8095] = ~((inputs[291]) | (inputs[288]));
    assign layer0_outputs[8096] = ~((inputs[545]) | (inputs[428]));
    assign layer0_outputs[8097] = ~(inputs[274]);
    assign layer0_outputs[8098] = (inputs[72]) ^ (inputs[697]);
    assign layer0_outputs[8099] = (inputs[725]) & ~(inputs[424]);
    assign layer0_outputs[8100] = (inputs[30]) & (inputs[917]);
    assign layer0_outputs[8101] = (inputs[76]) ^ (inputs[239]);
    assign layer0_outputs[8102] = ~(inputs[696]) | (inputs[190]);
    assign layer0_outputs[8103] = (inputs[236]) | (inputs[616]);
    assign layer0_outputs[8104] = inputs[788];
    assign layer0_outputs[8105] = inputs[655];
    assign layer0_outputs[8106] = ~((inputs[710]) | (inputs[339]));
    assign layer0_outputs[8107] = ~((inputs[384]) | (inputs[678]));
    assign layer0_outputs[8108] = ~((inputs[175]) ^ (inputs[712]));
    assign layer0_outputs[8109] = 1'b1;
    assign layer0_outputs[8110] = (inputs[457]) | (inputs[124]);
    assign layer0_outputs[8111] = (inputs[1012]) | (inputs[522]);
    assign layer0_outputs[8112] = (inputs[537]) | (inputs[997]);
    assign layer0_outputs[8113] = inputs[407];
    assign layer0_outputs[8114] = ~(inputs[973]);
    assign layer0_outputs[8115] = ~(inputs[401]);
    assign layer0_outputs[8116] = ~(inputs[419]);
    assign layer0_outputs[8117] = ~((inputs[851]) | (inputs[45]));
    assign layer0_outputs[8118] = (inputs[899]) | (inputs[614]);
    assign layer0_outputs[8119] = ~((inputs[845]) ^ (inputs[637]));
    assign layer0_outputs[8120] = ~(inputs[806]);
    assign layer0_outputs[8121] = 1'b1;
    assign layer0_outputs[8122] = ~(inputs[966]) | (inputs[77]);
    assign layer0_outputs[8123] = inputs[564];
    assign layer0_outputs[8124] = ~(inputs[994]);
    assign layer0_outputs[8125] = ~(inputs[515]);
    assign layer0_outputs[8126] = ~(inputs[463]);
    assign layer0_outputs[8127] = inputs[767];
    assign layer0_outputs[8128] = ~(inputs[911]);
    assign layer0_outputs[8129] = ~((inputs[297]) | (inputs[718]));
    assign layer0_outputs[8130] = (inputs[486]) & ~(inputs[991]);
    assign layer0_outputs[8131] = ~(inputs[193]) | (inputs[477]);
    assign layer0_outputs[8132] = (inputs[774]) | (inputs[909]);
    assign layer0_outputs[8133] = inputs[873];
    assign layer0_outputs[8134] = ~(inputs[19]);
    assign layer0_outputs[8135] = inputs[701];
    assign layer0_outputs[8136] = ~(inputs[965]) | (inputs[151]);
    assign layer0_outputs[8137] = ~(inputs[508]);
    assign layer0_outputs[8138] = inputs[112];
    assign layer0_outputs[8139] = ~((inputs[202]) | (inputs[612]));
    assign layer0_outputs[8140] = inputs[243];
    assign layer0_outputs[8141] = (inputs[18]) & ~(inputs[1003]);
    assign layer0_outputs[8142] = (inputs[632]) ^ (inputs[534]);
    assign layer0_outputs[8143] = ~(inputs[662]);
    assign layer0_outputs[8144] = ~((inputs[546]) & (inputs[973]));
    assign layer0_outputs[8145] = ~((inputs[739]) | (inputs[669]));
    assign layer0_outputs[8146] = ~((inputs[942]) ^ (inputs[238]));
    assign layer0_outputs[8147] = (inputs[467]) & ~(inputs[114]);
    assign layer0_outputs[8148] = ~((inputs[668]) ^ (inputs[855]));
    assign layer0_outputs[8149] = ~(inputs[204]) | (inputs[617]);
    assign layer0_outputs[8150] = (inputs[1013]) ^ (inputs[720]);
    assign layer0_outputs[8151] = ~(inputs[198]);
    assign layer0_outputs[8152] = 1'b0;
    assign layer0_outputs[8153] = ~((inputs[909]) | (inputs[119]));
    assign layer0_outputs[8154] = 1'b1;
    assign layer0_outputs[8155] = ~((inputs[822]) ^ (inputs[789]));
    assign layer0_outputs[8156] = (inputs[358]) | (inputs[229]);
    assign layer0_outputs[8157] = ~(inputs[620]);
    assign layer0_outputs[8158] = ~((inputs[218]) & (inputs[288]));
    assign layer0_outputs[8159] = (inputs[21]) ^ (inputs[144]);
    assign layer0_outputs[8160] = (inputs[834]) ^ (inputs[856]);
    assign layer0_outputs[8161] = ~((inputs[616]) ^ (inputs[9]));
    assign layer0_outputs[8162] = (inputs[678]) & ~(inputs[86]);
    assign layer0_outputs[8163] = ~(inputs[282]);
    assign layer0_outputs[8164] = (inputs[242]) & ~(inputs[578]);
    assign layer0_outputs[8165] = (inputs[405]) & ~(inputs[826]);
    assign layer0_outputs[8166] = inputs[784];
    assign layer0_outputs[8167] = ~((inputs[808]) ^ (inputs[419]));
    assign layer0_outputs[8168] = ~(inputs[398]);
    assign layer0_outputs[8169] = ~(inputs[485]) | (inputs[848]);
    assign layer0_outputs[8170] = inputs[115];
    assign layer0_outputs[8171] = (inputs[203]) | (inputs[649]);
    assign layer0_outputs[8172] = ~(inputs[342]);
    assign layer0_outputs[8173] = inputs[306];
    assign layer0_outputs[8174] = (inputs[883]) | (inputs[744]);
    assign layer0_outputs[8175] = (inputs[584]) ^ (inputs[287]);
    assign layer0_outputs[8176] = (inputs[866]) | (inputs[362]);
    assign layer0_outputs[8177] = ~(inputs[662]);
    assign layer0_outputs[8178] = inputs[1003];
    assign layer0_outputs[8179] = ~(inputs[644]) | (inputs[857]);
    assign layer0_outputs[8180] = ~((inputs[443]) ^ (inputs[465]));
    assign layer0_outputs[8181] = inputs[87];
    assign layer0_outputs[8182] = ~(inputs[347]) | (inputs[969]);
    assign layer0_outputs[8183] = ~(inputs[982]);
    assign layer0_outputs[8184] = (inputs[409]) & ~(inputs[449]);
    assign layer0_outputs[8185] = ~((inputs[79]) ^ (inputs[292]));
    assign layer0_outputs[8186] = ~((inputs[1010]) | (inputs[933]));
    assign layer0_outputs[8187] = (inputs[925]) ^ (inputs[947]);
    assign layer0_outputs[8188] = ~(inputs[848]) | (inputs[307]);
    assign layer0_outputs[8189] = ~((inputs[881]) | (inputs[390]));
    assign layer0_outputs[8190] = (inputs[561]) & ~(inputs[264]);
    assign layer0_outputs[8191] = ~((inputs[671]) ^ (inputs[516]));
    assign layer0_outputs[8192] = ~(inputs[46]);
    assign layer0_outputs[8193] = (inputs[134]) ^ (inputs[846]);
    assign layer0_outputs[8194] = ~((inputs[347]) | (inputs[1007]));
    assign layer0_outputs[8195] = (inputs[558]) & ~(inputs[195]);
    assign layer0_outputs[8196] = inputs[306];
    assign layer0_outputs[8197] = inputs[477];
    assign layer0_outputs[8198] = (inputs[615]) & ~(inputs[285]);
    assign layer0_outputs[8199] = ~((inputs[699]) ^ (inputs[653]));
    assign layer0_outputs[8200] = (inputs[424]) | (inputs[77]);
    assign layer0_outputs[8201] = (inputs[96]) & ~(inputs[326]);
    assign layer0_outputs[8202] = ~(inputs[211]);
    assign layer0_outputs[8203] = ~(inputs[778]);
    assign layer0_outputs[8204] = ~((inputs[266]) ^ (inputs[92]));
    assign layer0_outputs[8205] = inputs[292];
    assign layer0_outputs[8206] = ~(inputs[314]) | (inputs[966]);
    assign layer0_outputs[8207] = ~(inputs[346]) | (inputs[983]);
    assign layer0_outputs[8208] = (inputs[933]) & ~(inputs[759]);
    assign layer0_outputs[8209] = (inputs[234]) & ~(inputs[81]);
    assign layer0_outputs[8210] = (inputs[883]) & ~(inputs[256]);
    assign layer0_outputs[8211] = (inputs[374]) | (inputs[887]);
    assign layer0_outputs[8212] = (inputs[946]) & ~(inputs[377]);
    assign layer0_outputs[8213] = ~((inputs[678]) | (inputs[111]));
    assign layer0_outputs[8214] = 1'b0;
    assign layer0_outputs[8215] = (inputs[196]) | (inputs[237]);
    assign layer0_outputs[8216] = ~(inputs[15]) | (inputs[191]);
    assign layer0_outputs[8217] = (inputs[685]) & ~(inputs[1015]);
    assign layer0_outputs[8218] = ~(inputs[343]);
    assign layer0_outputs[8219] = ~((inputs[492]) | (inputs[1000]));
    assign layer0_outputs[8220] = inputs[750];
    assign layer0_outputs[8221] = ~(inputs[598]) | (inputs[381]);
    assign layer0_outputs[8222] = ~(inputs[302]) | (inputs[48]);
    assign layer0_outputs[8223] = ~((inputs[447]) & (inputs[170]));
    assign layer0_outputs[8224] = ~(inputs[117]) | (inputs[856]);
    assign layer0_outputs[8225] = inputs[333];
    assign layer0_outputs[8226] = 1'b1;
    assign layer0_outputs[8227] = ~(inputs[437]);
    assign layer0_outputs[8228] = ~(inputs[255]) | (inputs[450]);
    assign layer0_outputs[8229] = (inputs[875]) & ~(inputs[249]);
    assign layer0_outputs[8230] = ~((inputs[30]) & (inputs[122]));
    assign layer0_outputs[8231] = ~((inputs[602]) | (inputs[266]));
    assign layer0_outputs[8232] = ~((inputs[35]) ^ (inputs[109]));
    assign layer0_outputs[8233] = 1'b1;
    assign layer0_outputs[8234] = ~(inputs[630]);
    assign layer0_outputs[8235] = (inputs[908]) & ~(inputs[344]);
    assign layer0_outputs[8236] = ~((inputs[852]) | (inputs[352]));
    assign layer0_outputs[8237] = ~(inputs[234]) | (inputs[412]);
    assign layer0_outputs[8238] = ~(inputs[952]);
    assign layer0_outputs[8239] = ~(inputs[408]);
    assign layer0_outputs[8240] = 1'b0;
    assign layer0_outputs[8241] = inputs[20];
    assign layer0_outputs[8242] = ~((inputs[696]) | (inputs[772]));
    assign layer0_outputs[8243] = (inputs[426]) & ~(inputs[638]);
    assign layer0_outputs[8244] = (inputs[805]) | (inputs[239]);
    assign layer0_outputs[8245] = ~(inputs[527]);
    assign layer0_outputs[8246] = (inputs[232]) | (inputs[758]);
    assign layer0_outputs[8247] = 1'b1;
    assign layer0_outputs[8248] = (inputs[879]) | (inputs[936]);
    assign layer0_outputs[8249] = 1'b0;
    assign layer0_outputs[8250] = (inputs[131]) | (inputs[257]);
    assign layer0_outputs[8251] = ~((inputs[142]) | (inputs[722]));
    assign layer0_outputs[8252] = ~((inputs[289]) | (inputs[512]));
    assign layer0_outputs[8253] = inputs[280];
    assign layer0_outputs[8254] = (inputs[335]) ^ (inputs[63]);
    assign layer0_outputs[8255] = inputs[143];
    assign layer0_outputs[8256] = (inputs[90]) & (inputs[963]);
    assign layer0_outputs[8257] = ~((inputs[69]) | (inputs[917]));
    assign layer0_outputs[8258] = inputs[777];
    assign layer0_outputs[8259] = ~(inputs[562]);
    assign layer0_outputs[8260] = (inputs[352]) ^ (inputs[873]);
    assign layer0_outputs[8261] = ~(inputs[548]);
    assign layer0_outputs[8262] = inputs[783];
    assign layer0_outputs[8263] = (inputs[618]) & ~(inputs[979]);
    assign layer0_outputs[8264] = ~((inputs[685]) ^ (inputs[75]));
    assign layer0_outputs[8265] = ~(inputs[240]) | (inputs[350]);
    assign layer0_outputs[8266] = (inputs[951]) | (inputs[765]);
    assign layer0_outputs[8267] = ~(inputs[813]);
    assign layer0_outputs[8268] = ~(inputs[593]) | (inputs[650]);
    assign layer0_outputs[8269] = (inputs[734]) | (inputs[861]);
    assign layer0_outputs[8270] = ~(inputs[724]);
    assign layer0_outputs[8271] = ~((inputs[217]) | (inputs[568]));
    assign layer0_outputs[8272] = ~((inputs[199]) ^ (inputs[138]));
    assign layer0_outputs[8273] = ~(inputs[952]);
    assign layer0_outputs[8274] = inputs[349];
    assign layer0_outputs[8275] = ~(inputs[587]) | (inputs[856]);
    assign layer0_outputs[8276] = ~((inputs[755]) | (inputs[514]));
    assign layer0_outputs[8277] = inputs[775];
    assign layer0_outputs[8278] = (inputs[957]) | (inputs[592]);
    assign layer0_outputs[8279] = inputs[943];
    assign layer0_outputs[8280] = (inputs[849]) | (inputs[378]);
    assign layer0_outputs[8281] = ~(inputs[514]) | (inputs[16]);
    assign layer0_outputs[8282] = inputs[370];
    assign layer0_outputs[8283] = (inputs[284]) ^ (inputs[955]);
    assign layer0_outputs[8284] = (inputs[368]) ^ (inputs[95]);
    assign layer0_outputs[8285] = inputs[661];
    assign layer0_outputs[8286] = (inputs[526]) | (inputs[446]);
    assign layer0_outputs[8287] = 1'b1;
    assign layer0_outputs[8288] = ~(inputs[300]);
    assign layer0_outputs[8289] = ~(inputs[237]) | (inputs[642]);
    assign layer0_outputs[8290] = ~(inputs[461]) | (inputs[820]);
    assign layer0_outputs[8291] = (inputs[369]) ^ (inputs[130]);
    assign layer0_outputs[8292] = ~(inputs[621]);
    assign layer0_outputs[8293] = (inputs[142]) & ~(inputs[574]);
    assign layer0_outputs[8294] = ~(inputs[843]);
    assign layer0_outputs[8295] = ~(inputs[169]);
    assign layer0_outputs[8296] = ~(inputs[942]) | (inputs[867]);
    assign layer0_outputs[8297] = 1'b1;
    assign layer0_outputs[8298] = ~(inputs[458]);
    assign layer0_outputs[8299] = (inputs[577]) & ~(inputs[222]);
    assign layer0_outputs[8300] = (inputs[395]) & (inputs[424]);
    assign layer0_outputs[8301] = ~(inputs[19]) | (inputs[982]);
    assign layer0_outputs[8302] = (inputs[787]) & ~(inputs[383]);
    assign layer0_outputs[8303] = ~(inputs[36]);
    assign layer0_outputs[8304] = (inputs[460]) & ~(inputs[1010]);
    assign layer0_outputs[8305] = (inputs[69]) & ~(inputs[611]);
    assign layer0_outputs[8306] = ~((inputs[518]) | (inputs[446]));
    assign layer0_outputs[8307] = inputs[311];
    assign layer0_outputs[8308] = ~((inputs[595]) | (inputs[16]));
    assign layer0_outputs[8309] = (inputs[512]) | (inputs[185]);
    assign layer0_outputs[8310] = (inputs[107]) ^ (inputs[140]);
    assign layer0_outputs[8311] = ~(inputs[632]);
    assign layer0_outputs[8312] = (inputs[384]) & (inputs[935]);
    assign layer0_outputs[8313] = 1'b1;
    assign layer0_outputs[8314] = (inputs[817]) ^ (inputs[445]);
    assign layer0_outputs[8315] = ~(inputs[592]);
    assign layer0_outputs[8316] = (inputs[250]) & ~(inputs[48]);
    assign layer0_outputs[8317] = ~(inputs[337]);
    assign layer0_outputs[8318] = ~(inputs[463]);
    assign layer0_outputs[8319] = 1'b1;
    assign layer0_outputs[8320] = ~(inputs[481]);
    assign layer0_outputs[8321] = (inputs[607]) | (inputs[270]);
    assign layer0_outputs[8322] = ~((inputs[824]) ^ (inputs[848]));
    assign layer0_outputs[8323] = ~((inputs[758]) ^ (inputs[595]));
    assign layer0_outputs[8324] = (inputs[534]) & ~(inputs[700]);
    assign layer0_outputs[8325] = (inputs[547]) | (inputs[462]);
    assign layer0_outputs[8326] = 1'b0;
    assign layer0_outputs[8327] = ~((inputs[282]) ^ (inputs[672]));
    assign layer0_outputs[8328] = (inputs[360]) & ~(inputs[419]);
    assign layer0_outputs[8329] = (inputs[731]) | (inputs[334]);
    assign layer0_outputs[8330] = (inputs[195]) ^ (inputs[465]);
    assign layer0_outputs[8331] = (inputs[891]) & ~(inputs[837]);
    assign layer0_outputs[8332] = inputs[561];
    assign layer0_outputs[8333] = 1'b0;
    assign layer0_outputs[8334] = ~(inputs[597]) | (inputs[1006]);
    assign layer0_outputs[8335] = ~(inputs[470]);
    assign layer0_outputs[8336] = ~(inputs[441]) | (inputs[997]);
    assign layer0_outputs[8337] = ~(inputs[532]);
    assign layer0_outputs[8338] = ~((inputs[812]) | (inputs[45]));
    assign layer0_outputs[8339] = ~((inputs[563]) & (inputs[931]));
    assign layer0_outputs[8340] = (inputs[397]) ^ (inputs[602]);
    assign layer0_outputs[8341] = ~(inputs[111]);
    assign layer0_outputs[8342] = (inputs[694]) | (inputs[853]);
    assign layer0_outputs[8343] = inputs[532];
    assign layer0_outputs[8344] = (inputs[692]) | (inputs[975]);
    assign layer0_outputs[8345] = (inputs[232]) | (inputs[499]);
    assign layer0_outputs[8346] = inputs[599];
    assign layer0_outputs[8347] = ~((inputs[372]) | (inputs[772]));
    assign layer0_outputs[8348] = ~(inputs[495]) | (inputs[87]);
    assign layer0_outputs[8349] = (inputs[667]) ^ (inputs[684]);
    assign layer0_outputs[8350] = (inputs[385]) | (inputs[437]);
    assign layer0_outputs[8351] = (inputs[429]) & ~(inputs[829]);
    assign layer0_outputs[8352] = (inputs[657]) | (inputs[909]);
    assign layer0_outputs[8353] = ~((inputs[320]) | (inputs[819]));
    assign layer0_outputs[8354] = 1'b0;
    assign layer0_outputs[8355] = inputs[780];
    assign layer0_outputs[8356] = ~(inputs[468]);
    assign layer0_outputs[8357] = ~((inputs[778]) & (inputs[610]));
    assign layer0_outputs[8358] = ~((inputs[447]) & (inputs[72]));
    assign layer0_outputs[8359] = ~(inputs[426]);
    assign layer0_outputs[8360] = inputs[615];
    assign layer0_outputs[8361] = (inputs[823]) ^ (inputs[794]);
    assign layer0_outputs[8362] = (inputs[955]) | (inputs[166]);
    assign layer0_outputs[8363] = (inputs[321]) & ~(inputs[604]);
    assign layer0_outputs[8364] = (inputs[526]) | (inputs[168]);
    assign layer0_outputs[8365] = ~(inputs[780]);
    assign layer0_outputs[8366] = ~(inputs[876]) | (inputs[958]);
    assign layer0_outputs[8367] = ~(inputs[429]);
    assign layer0_outputs[8368] = ~(inputs[845]) | (inputs[81]);
    assign layer0_outputs[8369] = ~(inputs[402]) | (inputs[255]);
    assign layer0_outputs[8370] = ~((inputs[256]) & (inputs[561]));
    assign layer0_outputs[8371] = ~(inputs[593]);
    assign layer0_outputs[8372] = ~((inputs[997]) & (inputs[1006]));
    assign layer0_outputs[8373] = ~(inputs[869]) | (inputs[677]);
    assign layer0_outputs[8374] = ~(inputs[721]);
    assign layer0_outputs[8375] = ~((inputs[359]) | (inputs[166]));
    assign layer0_outputs[8376] = (inputs[610]) & (inputs[738]);
    assign layer0_outputs[8377] = 1'b0;
    assign layer0_outputs[8378] = (inputs[35]) ^ (inputs[947]);
    assign layer0_outputs[8379] = (inputs[459]) | (inputs[930]);
    assign layer0_outputs[8380] = ~(inputs[102]);
    assign layer0_outputs[8381] = ~(inputs[899]) | (inputs[222]);
    assign layer0_outputs[8382] = 1'b0;
    assign layer0_outputs[8383] = ~((inputs[696]) | (inputs[210]));
    assign layer0_outputs[8384] = ~(inputs[897]) | (inputs[49]);
    assign layer0_outputs[8385] = inputs[456];
    assign layer0_outputs[8386] = ~(inputs[500]);
    assign layer0_outputs[8387] = ~(inputs[778]) | (inputs[389]);
    assign layer0_outputs[8388] = ~((inputs[929]) | (inputs[90]));
    assign layer0_outputs[8389] = ~(inputs[340]) | (inputs[852]);
    assign layer0_outputs[8390] = (inputs[586]) & ~(inputs[4]);
    assign layer0_outputs[8391] = ~((inputs[923]) | (inputs[7]));
    assign layer0_outputs[8392] = (inputs[343]) & ~(inputs[514]);
    assign layer0_outputs[8393] = inputs[711];
    assign layer0_outputs[8394] = (inputs[950]) | (inputs[854]);
    assign layer0_outputs[8395] = (inputs[814]) ^ (inputs[90]);
    assign layer0_outputs[8396] = (inputs[292]) | (inputs[946]);
    assign layer0_outputs[8397] = ~(inputs[929]) | (inputs[76]);
    assign layer0_outputs[8398] = ~(inputs[487]);
    assign layer0_outputs[8399] = ~(inputs[309]);
    assign layer0_outputs[8400] = ~((inputs[396]) | (inputs[195]));
    assign layer0_outputs[8401] = ~((inputs[934]) | (inputs[650]));
    assign layer0_outputs[8402] = inputs[665];
    assign layer0_outputs[8403] = inputs[215];
    assign layer0_outputs[8404] = ~((inputs[69]) & (inputs[706]));
    assign layer0_outputs[8405] = (inputs[858]) & ~(inputs[649]);
    assign layer0_outputs[8406] = inputs[690];
    assign layer0_outputs[8407] = 1'b1;
    assign layer0_outputs[8408] = (inputs[266]) | (inputs[792]);
    assign layer0_outputs[8409] = 1'b0;
    assign layer0_outputs[8410] = inputs[399];
    assign layer0_outputs[8411] = ~(inputs[994]);
    assign layer0_outputs[8412] = inputs[57];
    assign layer0_outputs[8413] = (inputs[705]) | (inputs[835]);
    assign layer0_outputs[8414] = ~(inputs[370]) | (inputs[776]);
    assign layer0_outputs[8415] = ~(inputs[551]) | (inputs[118]);
    assign layer0_outputs[8416] = ~(inputs[460]) | (inputs[293]);
    assign layer0_outputs[8417] = inputs[335];
    assign layer0_outputs[8418] = inputs[657];
    assign layer0_outputs[8419] = (inputs[622]) & ~(inputs[191]);
    assign layer0_outputs[8420] = (inputs[366]) & ~(inputs[912]);
    assign layer0_outputs[8421] = ~((inputs[699]) ^ (inputs[192]));
    assign layer0_outputs[8422] = (inputs[995]) | (inputs[428]);
    assign layer0_outputs[8423] = (inputs[210]) | (inputs[243]);
    assign layer0_outputs[8424] = inputs[292];
    assign layer0_outputs[8425] = inputs[868];
    assign layer0_outputs[8426] = (inputs[291]) & ~(inputs[617]);
    assign layer0_outputs[8427] = (inputs[882]) & ~(inputs[136]);
    assign layer0_outputs[8428] = inputs[344];
    assign layer0_outputs[8429] = 1'b1;
    assign layer0_outputs[8430] = ~(inputs[981]) | (inputs[157]);
    assign layer0_outputs[8431] = ~((inputs[705]) | (inputs[625]));
    assign layer0_outputs[8432] = ~(inputs[529]);
    assign layer0_outputs[8433] = (inputs[656]) | (inputs[586]);
    assign layer0_outputs[8434] = ~(inputs[912]) | (inputs[107]);
    assign layer0_outputs[8435] = ~(inputs[817]) | (inputs[575]);
    assign layer0_outputs[8436] = 1'b1;
    assign layer0_outputs[8437] = ~((inputs[944]) | (inputs[876]));
    assign layer0_outputs[8438] = inputs[330];
    assign layer0_outputs[8439] = ~((inputs[641]) ^ (inputs[172]));
    assign layer0_outputs[8440] = (inputs[43]) & ~(inputs[226]);
    assign layer0_outputs[8441] = (inputs[420]) ^ (inputs[612]);
    assign layer0_outputs[8442] = inputs[494];
    assign layer0_outputs[8443] = ~((inputs[457]) | (inputs[321]));
    assign layer0_outputs[8444] = (inputs[153]) | (inputs[437]);
    assign layer0_outputs[8445] = ~(inputs[746]);
    assign layer0_outputs[8446] = ~(inputs[820]) | (inputs[980]);
    assign layer0_outputs[8447] = (inputs[948]) & (inputs[184]);
    assign layer0_outputs[8448] = ~((inputs[480]) | (inputs[125]));
    assign layer0_outputs[8449] = ~((inputs[170]) | (inputs[180]));
    assign layer0_outputs[8450] = ~((inputs[398]) | (inputs[882]));
    assign layer0_outputs[8451] = (inputs[562]) & ~(inputs[732]);
    assign layer0_outputs[8452] = ~((inputs[540]) ^ (inputs[750]));
    assign layer0_outputs[8453] = (inputs[780]) & ~(inputs[56]);
    assign layer0_outputs[8454] = (inputs[291]) & ~(inputs[123]);
    assign layer0_outputs[8455] = inputs[323];
    assign layer0_outputs[8456] = (inputs[530]) & ~(inputs[709]);
    assign layer0_outputs[8457] = inputs[553];
    assign layer0_outputs[8458] = ~(inputs[726]);
    assign layer0_outputs[8459] = inputs[935];
    assign layer0_outputs[8460] = ~(inputs[533]);
    assign layer0_outputs[8461] = ~((inputs[365]) | (inputs[961]));
    assign layer0_outputs[8462] = ~((inputs[117]) | (inputs[398]));
    assign layer0_outputs[8463] = inputs[685];
    assign layer0_outputs[8464] = ~(inputs[296]) | (inputs[40]);
    assign layer0_outputs[8465] = ~((inputs[650]) ^ (inputs[948]));
    assign layer0_outputs[8466] = (inputs[404]) | (inputs[545]);
    assign layer0_outputs[8467] = ~(inputs[8]) | (inputs[1019]);
    assign layer0_outputs[8468] = (inputs[324]) & (inputs[88]);
    assign layer0_outputs[8469] = inputs[734];
    assign layer0_outputs[8470] = (inputs[314]) | (inputs[978]);
    assign layer0_outputs[8471] = (inputs[240]) | (inputs[709]);
    assign layer0_outputs[8472] = inputs[233];
    assign layer0_outputs[8473] = (inputs[147]) | (inputs[715]);
    assign layer0_outputs[8474] = ~((inputs[191]) ^ (inputs[488]));
    assign layer0_outputs[8475] = ~((inputs[132]) ^ (inputs[206]));
    assign layer0_outputs[8476] = 1'b0;
    assign layer0_outputs[8477] = (inputs[878]) & ~(inputs[795]);
    assign layer0_outputs[8478] = ~(inputs[470]);
    assign layer0_outputs[8479] = ~(inputs[494]);
    assign layer0_outputs[8480] = ~((inputs[818]) ^ (inputs[660]));
    assign layer0_outputs[8481] = (inputs[118]) ^ (inputs[441]);
    assign layer0_outputs[8482] = (inputs[404]) & ~(inputs[385]);
    assign layer0_outputs[8483] = ~(inputs[52]);
    assign layer0_outputs[8484] = ~((inputs[24]) | (inputs[1015]));
    assign layer0_outputs[8485] = (inputs[178]) | (inputs[656]);
    assign layer0_outputs[8486] = (inputs[382]) ^ (inputs[686]);
    assign layer0_outputs[8487] = ~(inputs[532]);
    assign layer0_outputs[8488] = inputs[311];
    assign layer0_outputs[8489] = ~(inputs[613]);
    assign layer0_outputs[8490] = 1'b1;
    assign layer0_outputs[8491] = ~(inputs[282]);
    assign layer0_outputs[8492] = (inputs[64]) & (inputs[41]);
    assign layer0_outputs[8493] = ~(inputs[502]) | (inputs[354]);
    assign layer0_outputs[8494] = (inputs[398]) ^ (inputs[539]);
    assign layer0_outputs[8495] = (inputs[267]) ^ (inputs[831]);
    assign layer0_outputs[8496] = inputs[982];
    assign layer0_outputs[8497] = ~((inputs[413]) | (inputs[1010]));
    assign layer0_outputs[8498] = inputs[583];
    assign layer0_outputs[8499] = (inputs[368]) & (inputs[523]);
    assign layer0_outputs[8500] = 1'b1;
    assign layer0_outputs[8501] = inputs[372];
    assign layer0_outputs[8502] = (inputs[602]) ^ (inputs[839]);
    assign layer0_outputs[8503] = inputs[315];
    assign layer0_outputs[8504] = 1'b0;
    assign layer0_outputs[8505] = (inputs[171]) & ~(inputs[475]);
    assign layer0_outputs[8506] = 1'b1;
    assign layer0_outputs[8507] = inputs[394];
    assign layer0_outputs[8508] = ~(inputs[265]);
    assign layer0_outputs[8509] = inputs[187];
    assign layer0_outputs[8510] = 1'b0;
    assign layer0_outputs[8511] = 1'b1;
    assign layer0_outputs[8512] = (inputs[244]) | (inputs[112]);
    assign layer0_outputs[8513] = 1'b1;
    assign layer0_outputs[8514] = ~((inputs[277]) ^ (inputs[471]));
    assign layer0_outputs[8515] = ~((inputs[633]) ^ (inputs[415]));
    assign layer0_outputs[8516] = ~(inputs[728]);
    assign layer0_outputs[8517] = ~(inputs[463]) | (inputs[410]);
    assign layer0_outputs[8518] = ~((inputs[14]) ^ (inputs[121]));
    assign layer0_outputs[8519] = inputs[399];
    assign layer0_outputs[8520] = (inputs[890]) ^ (inputs[560]);
    assign layer0_outputs[8521] = ~((inputs[457]) ^ (inputs[452]));
    assign layer0_outputs[8522] = ~(inputs[344]);
    assign layer0_outputs[8523] = (inputs[969]) | (inputs[581]);
    assign layer0_outputs[8524] = (inputs[278]) ^ (inputs[865]);
    assign layer0_outputs[8525] = ~(inputs[434]);
    assign layer0_outputs[8526] = ~(inputs[36]);
    assign layer0_outputs[8527] = ~((inputs[187]) | (inputs[718]));
    assign layer0_outputs[8528] = 1'b0;
    assign layer0_outputs[8529] = inputs[570];
    assign layer0_outputs[8530] = (inputs[17]) ^ (inputs[191]);
    assign layer0_outputs[8531] = ~(inputs[967]);
    assign layer0_outputs[8532] = inputs[881];
    assign layer0_outputs[8533] = ~((inputs[529]) ^ (inputs[895]));
    assign layer0_outputs[8534] = ~(inputs[718]);
    assign layer0_outputs[8535] = inputs[315];
    assign layer0_outputs[8536] = ~(inputs[446]) | (inputs[998]);
    assign layer0_outputs[8537] = (inputs[559]) & ~(inputs[449]);
    assign layer0_outputs[8538] = (inputs[497]) & ~(inputs[763]);
    assign layer0_outputs[8539] = ~(inputs[267]) | (inputs[137]);
    assign layer0_outputs[8540] = ~((inputs[425]) | (inputs[41]));
    assign layer0_outputs[8541] = ~((inputs[764]) | (inputs[450]));
    assign layer0_outputs[8542] = ~((inputs[662]) & (inputs[390]));
    assign layer0_outputs[8543] = (inputs[395]) & ~(inputs[638]);
    assign layer0_outputs[8544] = inputs[718];
    assign layer0_outputs[8545] = (inputs[306]) & ~(inputs[34]);
    assign layer0_outputs[8546] = (inputs[792]) & ~(inputs[2]);
    assign layer0_outputs[8547] = ~((inputs[336]) | (inputs[1001]));
    assign layer0_outputs[8548] = ~((inputs[675]) | (inputs[921]));
    assign layer0_outputs[8549] = (inputs[1005]) | (inputs[772]);
    assign layer0_outputs[8550] = ~((inputs[754]) ^ (inputs[932]));
    assign layer0_outputs[8551] = (inputs[339]) & ~(inputs[112]);
    assign layer0_outputs[8552] = ~((inputs[686]) & (inputs[574]));
    assign layer0_outputs[8553] = ~((inputs[473]) | (inputs[495]));
    assign layer0_outputs[8554] = (inputs[408]) | (inputs[21]);
    assign layer0_outputs[8555] = (inputs[650]) & ~(inputs[34]);
    assign layer0_outputs[8556] = (inputs[259]) ^ (inputs[278]);
    assign layer0_outputs[8557] = 1'b1;
    assign layer0_outputs[8558] = (inputs[36]) & ~(inputs[284]);
    assign layer0_outputs[8559] = (inputs[598]) & ~(inputs[605]);
    assign layer0_outputs[8560] = ~(inputs[814]);
    assign layer0_outputs[8561] = (inputs[1020]) ^ (inputs[15]);
    assign layer0_outputs[8562] = (inputs[65]) | (inputs[705]);
    assign layer0_outputs[8563] = (inputs[842]) | (inputs[95]);
    assign layer0_outputs[8564] = (inputs[181]) ^ (inputs[329]);
    assign layer0_outputs[8565] = ~(inputs[555]) | (inputs[181]);
    assign layer0_outputs[8566] = (inputs[727]) & ~(inputs[360]);
    assign layer0_outputs[8567] = ~(inputs[473]);
    assign layer0_outputs[8568] = inputs[556];
    assign layer0_outputs[8569] = ~((inputs[71]) ^ (inputs[402]));
    assign layer0_outputs[8570] = (inputs[830]) & ~(inputs[545]);
    assign layer0_outputs[8571] = (inputs[504]) | (inputs[503]);
    assign layer0_outputs[8572] = (inputs[997]) & ~(inputs[508]);
    assign layer0_outputs[8573] = inputs[99];
    assign layer0_outputs[8574] = ~(inputs[707]) | (inputs[705]);
    assign layer0_outputs[8575] = ~(inputs[422]);
    assign layer0_outputs[8576] = ~(inputs[190]) | (inputs[800]);
    assign layer0_outputs[8577] = (inputs[760]) | (inputs[600]);
    assign layer0_outputs[8578] = ~((inputs[135]) | (inputs[238]));
    assign layer0_outputs[8579] = ~((inputs[680]) | (inputs[348]));
    assign layer0_outputs[8580] = inputs[755];
    assign layer0_outputs[8581] = ~(inputs[552]) | (inputs[921]);
    assign layer0_outputs[8582] = (inputs[378]) & ~(inputs[869]);
    assign layer0_outputs[8583] = ~((inputs[677]) ^ (inputs[31]));
    assign layer0_outputs[8584] = ~(inputs[508]);
    assign layer0_outputs[8585] = ~(inputs[112]);
    assign layer0_outputs[8586] = ~(inputs[500]) | (inputs[126]);
    assign layer0_outputs[8587] = (inputs[857]) ^ (inputs[117]);
    assign layer0_outputs[8588] = (inputs[67]) ^ (inputs[560]);
    assign layer0_outputs[8589] = inputs[530];
    assign layer0_outputs[8590] = (inputs[659]) | (inputs[885]);
    assign layer0_outputs[8591] = inputs[518];
    assign layer0_outputs[8592] = 1'b0;
    assign layer0_outputs[8593] = ~(inputs[627]) | (inputs[452]);
    assign layer0_outputs[8594] = ~(inputs[717]);
    assign layer0_outputs[8595] = 1'b0;
    assign layer0_outputs[8596] = ~(inputs[915]);
    assign layer0_outputs[8597] = inputs[560];
    assign layer0_outputs[8598] = (inputs[286]) | (inputs[449]);
    assign layer0_outputs[8599] = ~(inputs[641]);
    assign layer0_outputs[8600] = ~(inputs[758]);
    assign layer0_outputs[8601] = inputs[438];
    assign layer0_outputs[8602] = (inputs[170]) & ~(inputs[311]);
    assign layer0_outputs[8603] = inputs[784];
    assign layer0_outputs[8604] = (inputs[315]) ^ (inputs[342]);
    assign layer0_outputs[8605] = ~((inputs[809]) | (inputs[643]));
    assign layer0_outputs[8606] = (inputs[673]) & ~(inputs[294]);
    assign layer0_outputs[8607] = (inputs[298]) & ~(inputs[772]);
    assign layer0_outputs[8608] = (inputs[898]) | (inputs[400]);
    assign layer0_outputs[8609] = ~(inputs[871]) | (inputs[545]);
    assign layer0_outputs[8610] = ~((inputs[534]) | (inputs[550]));
    assign layer0_outputs[8611] = ~(inputs[786]) | (inputs[982]);
    assign layer0_outputs[8612] = (inputs[134]) ^ (inputs[185]);
    assign layer0_outputs[8613] = (inputs[409]) & ~(inputs[995]);
    assign layer0_outputs[8614] = ~(inputs[620]);
    assign layer0_outputs[8615] = inputs[885];
    assign layer0_outputs[8616] = inputs[603];
    assign layer0_outputs[8617] = ~(inputs[441]);
    assign layer0_outputs[8618] = (inputs[363]) & ~(inputs[833]);
    assign layer0_outputs[8619] = (inputs[469]) ^ (inputs[140]);
    assign layer0_outputs[8620] = ~((inputs[514]) | (inputs[864]));
    assign layer0_outputs[8621] = (inputs[83]) & ~(inputs[958]);
    assign layer0_outputs[8622] = inputs[836];
    assign layer0_outputs[8623] = (inputs[579]) & (inputs[83]);
    assign layer0_outputs[8624] = (inputs[970]) & ~(inputs[573]);
    assign layer0_outputs[8625] = ~(inputs[359]);
    assign layer0_outputs[8626] = ~((inputs[855]) | (inputs[425]));
    assign layer0_outputs[8627] = ~(inputs[504]);
    assign layer0_outputs[8628] = ~(inputs[1012]);
    assign layer0_outputs[8629] = (inputs[543]) & (inputs[900]);
    assign layer0_outputs[8630] = ~(inputs[1000]);
    assign layer0_outputs[8631] = inputs[784];
    assign layer0_outputs[8632] = ~(inputs[316]);
    assign layer0_outputs[8633] = ~((inputs[449]) | (inputs[94]));
    assign layer0_outputs[8634] = ~((inputs[122]) & (inputs[230]));
    assign layer0_outputs[8635] = ~(inputs[342]);
    assign layer0_outputs[8636] = ~((inputs[647]) ^ (inputs[554]));
    assign layer0_outputs[8637] = 1'b0;
    assign layer0_outputs[8638] = 1'b1;
    assign layer0_outputs[8639] = (inputs[227]) & ~(inputs[423]);
    assign layer0_outputs[8640] = 1'b0;
    assign layer0_outputs[8641] = (inputs[395]) ^ (inputs[269]);
    assign layer0_outputs[8642] = ~((inputs[202]) | (inputs[1002]));
    assign layer0_outputs[8643] = ~(inputs[749]) | (inputs[68]);
    assign layer0_outputs[8644] = (inputs[251]) | (inputs[72]);
    assign layer0_outputs[8645] = ~(inputs[347]);
    assign layer0_outputs[8646] = 1'b0;
    assign layer0_outputs[8647] = ~(inputs[975]);
    assign layer0_outputs[8648] = ~((inputs[872]) ^ (inputs[746]));
    assign layer0_outputs[8649] = ~(inputs[950]) | (inputs[936]);
    assign layer0_outputs[8650] = ~(inputs[340]);
    assign layer0_outputs[8651] = 1'b1;
    assign layer0_outputs[8652] = (inputs[426]) ^ (inputs[879]);
    assign layer0_outputs[8653] = (inputs[497]) & ~(inputs[454]);
    assign layer0_outputs[8654] = (inputs[264]) | (inputs[234]);
    assign layer0_outputs[8655] = (inputs[381]) ^ (inputs[381]);
    assign layer0_outputs[8656] = ~((inputs[590]) | (inputs[761]));
    assign layer0_outputs[8657] = (inputs[373]) & ~(inputs[849]);
    assign layer0_outputs[8658] = inputs[341];
    assign layer0_outputs[8659] = ~(inputs[322]);
    assign layer0_outputs[8660] = ~((inputs[924]) | (inputs[968]));
    assign layer0_outputs[8661] = ~(inputs[565]);
    assign layer0_outputs[8662] = ~(inputs[590]);
    assign layer0_outputs[8663] = ~((inputs[787]) & (inputs[134]));
    assign layer0_outputs[8664] = (inputs[679]) ^ (inputs[63]);
    assign layer0_outputs[8665] = ~(inputs[122]) | (inputs[889]);
    assign layer0_outputs[8666] = ~((inputs[295]) | (inputs[872]));
    assign layer0_outputs[8667] = (inputs[625]) ^ (inputs[864]);
    assign layer0_outputs[8668] = (inputs[96]) | (inputs[468]);
    assign layer0_outputs[8669] = ~(inputs[244]);
    assign layer0_outputs[8670] = (inputs[635]) & ~(inputs[963]);
    assign layer0_outputs[8671] = ~((inputs[242]) ^ (inputs[569]));
    assign layer0_outputs[8672] = (inputs[120]) | (inputs[458]);
    assign layer0_outputs[8673] = (inputs[325]) & ~(inputs[317]);
    assign layer0_outputs[8674] = 1'b1;
    assign layer0_outputs[8675] = ~((inputs[122]) ^ (inputs[641]));
    assign layer0_outputs[8676] = ~(inputs[98]) | (inputs[645]);
    assign layer0_outputs[8677] = (inputs[697]) ^ (inputs[875]);
    assign layer0_outputs[8678] = inputs[998];
    assign layer0_outputs[8679] = ~((inputs[939]) ^ (inputs[525]));
    assign layer0_outputs[8680] = ~(inputs[820]);
    assign layer0_outputs[8681] = ~((inputs[437]) ^ (inputs[14]));
    assign layer0_outputs[8682] = ~(inputs[365]);
    assign layer0_outputs[8683] = ~(inputs[431]) | (inputs[913]);
    assign layer0_outputs[8684] = (inputs[896]) ^ (inputs[279]);
    assign layer0_outputs[8685] = (inputs[884]) ^ (inputs[258]);
    assign layer0_outputs[8686] = ~(inputs[336]);
    assign layer0_outputs[8687] = (inputs[713]) | (inputs[542]);
    assign layer0_outputs[8688] = (inputs[526]) | (inputs[85]);
    assign layer0_outputs[8689] = ~(inputs[754]);
    assign layer0_outputs[8690] = (inputs[187]) ^ (inputs[1002]);
    assign layer0_outputs[8691] = ~(inputs[905]) | (inputs[576]);
    assign layer0_outputs[8692] = (inputs[946]) | (inputs[759]);
    assign layer0_outputs[8693] = (inputs[128]) | (inputs[94]);
    assign layer0_outputs[8694] = (inputs[785]) & ~(inputs[498]);
    assign layer0_outputs[8695] = (inputs[214]) & ~(inputs[977]);
    assign layer0_outputs[8696] = ~(inputs[550]) | (inputs[754]);
    assign layer0_outputs[8697] = ~(inputs[257]) | (inputs[353]);
    assign layer0_outputs[8698] = (inputs[308]) & ~(inputs[326]);
    assign layer0_outputs[8699] = ~(inputs[589]) | (inputs[335]);
    assign layer0_outputs[8700] = ~(inputs[625]) | (inputs[845]);
    assign layer0_outputs[8701] = ~(inputs[561]);
    assign layer0_outputs[8702] = (inputs[901]) & ~(inputs[1016]);
    assign layer0_outputs[8703] = ~(inputs[139]);
    assign layer0_outputs[8704] = (inputs[41]) ^ (inputs[588]);
    assign layer0_outputs[8705] = (inputs[560]) & ~(inputs[450]);
    assign layer0_outputs[8706] = ~(inputs[624]);
    assign layer0_outputs[8707] = ~(inputs[134]) | (inputs[1]);
    assign layer0_outputs[8708] = (inputs[761]) & ~(inputs[362]);
    assign layer0_outputs[8709] = 1'b1;
    assign layer0_outputs[8710] = ~(inputs[335]);
    assign layer0_outputs[8711] = ~((inputs[110]) & (inputs[56]));
    assign layer0_outputs[8712] = ~(inputs[524]);
    assign layer0_outputs[8713] = inputs[566];
    assign layer0_outputs[8714] = inputs[778];
    assign layer0_outputs[8715] = ~(inputs[707]) | (inputs[551]);
    assign layer0_outputs[8716] = ~(inputs[398]);
    assign layer0_outputs[8717] = inputs[241];
    assign layer0_outputs[8718] = inputs[259];
    assign layer0_outputs[8719] = (inputs[266]) | (inputs[728]);
    assign layer0_outputs[8720] = (inputs[316]) ^ (inputs[746]);
    assign layer0_outputs[8721] = ~(inputs[77]);
    assign layer0_outputs[8722] = 1'b0;
    assign layer0_outputs[8723] = (inputs[223]) & ~(inputs[979]);
    assign layer0_outputs[8724] = ~(inputs[247]) | (inputs[868]);
    assign layer0_outputs[8725] = (inputs[75]) & ~(inputs[669]);
    assign layer0_outputs[8726] = ~((inputs[411]) | (inputs[589]));
    assign layer0_outputs[8727] = ~(inputs[202]) | (inputs[53]);
    assign layer0_outputs[8728] = (inputs[177]) | (inputs[731]);
    assign layer0_outputs[8729] = (inputs[516]) ^ (inputs[281]);
    assign layer0_outputs[8730] = inputs[495];
    assign layer0_outputs[8731] = inputs[653];
    assign layer0_outputs[8732] = ~(inputs[204]) | (inputs[323]);
    assign layer0_outputs[8733] = (inputs[775]) & ~(inputs[951]);
    assign layer0_outputs[8734] = inputs[692];
    assign layer0_outputs[8735] = ~(inputs[589]);
    assign layer0_outputs[8736] = ~((inputs[84]) ^ (inputs[79]));
    assign layer0_outputs[8737] = (inputs[220]) | (inputs[330]);
    assign layer0_outputs[8738] = ~((inputs[221]) ^ (inputs[855]));
    assign layer0_outputs[8739] = ~(inputs[454]);
    assign layer0_outputs[8740] = (inputs[235]) & ~(inputs[577]);
    assign layer0_outputs[8741] = 1'b0;
    assign layer0_outputs[8742] = (inputs[895]) ^ (inputs[262]);
    assign layer0_outputs[8743] = ~(inputs[173]) | (inputs[368]);
    assign layer0_outputs[8744] = (inputs[396]) & ~(inputs[838]);
    assign layer0_outputs[8745] = ~((inputs[367]) ^ (inputs[328]));
    assign layer0_outputs[8746] = (inputs[444]) | (inputs[746]);
    assign layer0_outputs[8747] = (inputs[1022]) ^ (inputs[899]);
    assign layer0_outputs[8748] = ~((inputs[551]) & (inputs[537]));
    assign layer0_outputs[8749] = ~(inputs[103]) | (inputs[303]);
    assign layer0_outputs[8750] = ~((inputs[708]) ^ (inputs[130]));
    assign layer0_outputs[8751] = ~(inputs[465]);
    assign layer0_outputs[8752] = (inputs[168]) ^ (inputs[144]);
    assign layer0_outputs[8753] = ~(inputs[751]) | (inputs[260]);
    assign layer0_outputs[8754] = ~(inputs[922]);
    assign layer0_outputs[8755] = ~(inputs[303]);
    assign layer0_outputs[8756] = ~((inputs[464]) | (inputs[757]));
    assign layer0_outputs[8757] = (inputs[338]) & ~(inputs[407]);
    assign layer0_outputs[8758] = inputs[181];
    assign layer0_outputs[8759] = 1'b1;
    assign layer0_outputs[8760] = (inputs[402]) ^ (inputs[9]);
    assign layer0_outputs[8761] = (inputs[659]) | (inputs[294]);
    assign layer0_outputs[8762] = (inputs[235]) & ~(inputs[91]);
    assign layer0_outputs[8763] = (inputs[454]) ^ (inputs[893]);
    assign layer0_outputs[8764] = (inputs[363]) & ~(inputs[458]);
    assign layer0_outputs[8765] = ~((inputs[329]) & (inputs[480]));
    assign layer0_outputs[8766] = ~((inputs[777]) | (inputs[749]));
    assign layer0_outputs[8767] = ~(inputs[692]);
    assign layer0_outputs[8768] = ~(inputs[551]);
    assign layer0_outputs[8769] = (inputs[493]) | (inputs[495]);
    assign layer0_outputs[8770] = (inputs[985]) & ~(inputs[601]);
    assign layer0_outputs[8771] = ~(inputs[616]);
    assign layer0_outputs[8772] = inputs[249];
    assign layer0_outputs[8773] = (inputs[687]) & ~(inputs[887]);
    assign layer0_outputs[8774] = ~(inputs[678]) | (inputs[454]);
    assign layer0_outputs[8775] = ~(inputs[175]) | (inputs[575]);
    assign layer0_outputs[8776] = ~((inputs[571]) | (inputs[407]));
    assign layer0_outputs[8777] = ~((inputs[803]) ^ (inputs[782]));
    assign layer0_outputs[8778] = inputs[494];
    assign layer0_outputs[8779] = ~(inputs[565]) | (inputs[510]);
    assign layer0_outputs[8780] = inputs[912];
    assign layer0_outputs[8781] = ~((inputs[236]) & (inputs[244]));
    assign layer0_outputs[8782] = (inputs[399]) ^ (inputs[421]);
    assign layer0_outputs[8783] = (inputs[668]) | (inputs[978]);
    assign layer0_outputs[8784] = ~(inputs[814]) | (inputs[226]);
    assign layer0_outputs[8785] = ~(inputs[842]);
    assign layer0_outputs[8786] = ~((inputs[735]) & (inputs[25]));
    assign layer0_outputs[8787] = inputs[812];
    assign layer0_outputs[8788] = inputs[439];
    assign layer0_outputs[8789] = ~(inputs[970]);
    assign layer0_outputs[8790] = 1'b1;
    assign layer0_outputs[8791] = inputs[457];
    assign layer0_outputs[8792] = inputs[361];
    assign layer0_outputs[8793] = (inputs[976]) | (inputs[103]);
    assign layer0_outputs[8794] = inputs[557];
    assign layer0_outputs[8795] = ~((inputs[696]) | (inputs[467]));
    assign layer0_outputs[8796] = (inputs[673]) ^ (inputs[34]);
    assign layer0_outputs[8797] = 1'b1;
    assign layer0_outputs[8798] = (inputs[120]) | (inputs[467]);
    assign layer0_outputs[8799] = ~(inputs[218]) | (inputs[73]);
    assign layer0_outputs[8800] = ~(inputs[320]) | (inputs[607]);
    assign layer0_outputs[8801] = ~(inputs[727]) | (inputs[538]);
    assign layer0_outputs[8802] = ~(inputs[275]);
    assign layer0_outputs[8803] = (inputs[90]) ^ (inputs[717]);
    assign layer0_outputs[8804] = ~(inputs[139]);
    assign layer0_outputs[8805] = inputs[649];
    assign layer0_outputs[8806] = ~(inputs[858]) | (inputs[865]);
    assign layer0_outputs[8807] = ~(inputs[331]) | (inputs[934]);
    assign layer0_outputs[8808] = (inputs[7]) ^ (inputs[547]);
    assign layer0_outputs[8809] = ~((inputs[934]) & (inputs[960]));
    assign layer0_outputs[8810] = ~(inputs[209]);
    assign layer0_outputs[8811] = (inputs[795]) & ~(inputs[708]);
    assign layer0_outputs[8812] = ~((inputs[118]) | (inputs[596]));
    assign layer0_outputs[8813] = (inputs[205]) & ~(inputs[491]);
    assign layer0_outputs[8814] = 1'b1;
    assign layer0_outputs[8815] = (inputs[239]) & ~(inputs[506]);
    assign layer0_outputs[8816] = (inputs[849]) | (inputs[484]);
    assign layer0_outputs[8817] = (inputs[272]) ^ (inputs[309]);
    assign layer0_outputs[8818] = (inputs[983]) & (inputs[602]);
    assign layer0_outputs[8819] = (inputs[242]) & (inputs[684]);
    assign layer0_outputs[8820] = (inputs[686]) | (inputs[999]);
    assign layer0_outputs[8821] = (inputs[252]) & (inputs[844]);
    assign layer0_outputs[8822] = (inputs[464]) | (inputs[496]);
    assign layer0_outputs[8823] = ~(inputs[600]) | (inputs[58]);
    assign layer0_outputs[8824] = inputs[405];
    assign layer0_outputs[8825] = ~((inputs[0]) & (inputs[604]));
    assign layer0_outputs[8826] = (inputs[104]) | (inputs[114]);
    assign layer0_outputs[8827] = (inputs[901]) ^ (inputs[119]);
    assign layer0_outputs[8828] = inputs[593];
    assign layer0_outputs[8829] = ~((inputs[553]) | (inputs[290]));
    assign layer0_outputs[8830] = ~((inputs[642]) ^ (inputs[103]));
    assign layer0_outputs[8831] = ~(inputs[617]);
    assign layer0_outputs[8832] = (inputs[660]) ^ (inputs[940]);
    assign layer0_outputs[8833] = ~((inputs[338]) | (inputs[325]));
    assign layer0_outputs[8834] = (inputs[938]) & ~(inputs[577]);
    assign layer0_outputs[8835] = ~((inputs[739]) | (inputs[439]));
    assign layer0_outputs[8836] = (inputs[26]) | (inputs[33]);
    assign layer0_outputs[8837] = (inputs[417]) | (inputs[822]);
    assign layer0_outputs[8838] = (inputs[105]) | (inputs[459]);
    assign layer0_outputs[8839] = (inputs[563]) & ~(inputs[507]);
    assign layer0_outputs[8840] = inputs[519];
    assign layer0_outputs[8841] = (inputs[2]) & ~(inputs[484]);
    assign layer0_outputs[8842] = ~(inputs[798]) | (inputs[935]);
    assign layer0_outputs[8843] = ~(inputs[180]);
    assign layer0_outputs[8844] = ~((inputs[272]) ^ (inputs[126]));
    assign layer0_outputs[8845] = (inputs[549]) & ~(inputs[255]);
    assign layer0_outputs[8846] = ~(inputs[368]) | (inputs[794]);
    assign layer0_outputs[8847] = (inputs[341]) | (inputs[580]);
    assign layer0_outputs[8848] = inputs[490];
    assign layer0_outputs[8849] = (inputs[352]) ^ (inputs[505]);
    assign layer0_outputs[8850] = ~(inputs[999]) | (inputs[804]);
    assign layer0_outputs[8851] = (inputs[546]) | (inputs[400]);
    assign layer0_outputs[8852] = (inputs[891]) & (inputs[557]);
    assign layer0_outputs[8853] = (inputs[780]) & ~(inputs[23]);
    assign layer0_outputs[8854] = ~((inputs[341]) ^ (inputs[419]));
    assign layer0_outputs[8855] = inputs[745];
    assign layer0_outputs[8856] = ~(inputs[626]) | (inputs[48]);
    assign layer0_outputs[8857] = (inputs[662]) & ~(inputs[444]);
    assign layer0_outputs[8858] = ~((inputs[121]) ^ (inputs[63]));
    assign layer0_outputs[8859] = ~(inputs[839]) | (inputs[821]);
    assign layer0_outputs[8860] = (inputs[368]) ^ (inputs[53]);
    assign layer0_outputs[8861] = (inputs[284]) ^ (inputs[441]);
    assign layer0_outputs[8862] = ~((inputs[906]) ^ (inputs[254]));
    assign layer0_outputs[8863] = ~((inputs[332]) | (inputs[292]));
    assign layer0_outputs[8864] = ~(inputs[845]);
    assign layer0_outputs[8865] = inputs[423];
    assign layer0_outputs[8866] = ~((inputs[720]) ^ (inputs[209]));
    assign layer0_outputs[8867] = ~(inputs[685]);
    assign layer0_outputs[8868] = (inputs[589]) ^ (inputs[802]);
    assign layer0_outputs[8869] = ~((inputs[782]) ^ (inputs[133]));
    assign layer0_outputs[8870] = (inputs[48]) | (inputs[732]);
    assign layer0_outputs[8871] = (inputs[765]) & ~(inputs[650]);
    assign layer0_outputs[8872] = inputs[756];
    assign layer0_outputs[8873] = inputs[404];
    assign layer0_outputs[8874] = inputs[396];
    assign layer0_outputs[8875] = ~((inputs[345]) ^ (inputs[900]));
    assign layer0_outputs[8876] = (inputs[542]) & (inputs[927]);
    assign layer0_outputs[8877] = ~(inputs[495]);
    assign layer0_outputs[8878] = ~(inputs[206]) | (inputs[120]);
    assign layer0_outputs[8879] = ~(inputs[131]) | (inputs[163]);
    assign layer0_outputs[8880] = ~((inputs[892]) ^ (inputs[834]));
    assign layer0_outputs[8881] = ~(inputs[456]);
    assign layer0_outputs[8882] = inputs[775];
    assign layer0_outputs[8883] = ~((inputs[789]) ^ (inputs[179]));
    assign layer0_outputs[8884] = ~(inputs[209]) | (inputs[760]);
    assign layer0_outputs[8885] = (inputs[654]) & ~(inputs[224]);
    assign layer0_outputs[8886] = (inputs[795]) ^ (inputs[687]);
    assign layer0_outputs[8887] = (inputs[563]) | (inputs[507]);
    assign layer0_outputs[8888] = ~(inputs[617]) | (inputs[26]);
    assign layer0_outputs[8889] = (inputs[210]) | (inputs[452]);
    assign layer0_outputs[8890] = ~(inputs[136]) | (inputs[187]);
    assign layer0_outputs[8891] = (inputs[203]) | (inputs[3]);
    assign layer0_outputs[8892] = inputs[727];
    assign layer0_outputs[8893] = ~((inputs[810]) | (inputs[102]));
    assign layer0_outputs[8894] = ~(inputs[591]) | (inputs[424]);
    assign layer0_outputs[8895] = inputs[561];
    assign layer0_outputs[8896] = inputs[333];
    assign layer0_outputs[8897] = ~((inputs[472]) ^ (inputs[598]));
    assign layer0_outputs[8898] = (inputs[853]) | (inputs[42]);
    assign layer0_outputs[8899] = inputs[176];
    assign layer0_outputs[8900] = inputs[436];
    assign layer0_outputs[8901] = ~((inputs[102]) & (inputs[802]));
    assign layer0_outputs[8902] = ~(inputs[356]);
    assign layer0_outputs[8903] = ~((inputs[232]) & (inputs[669]));
    assign layer0_outputs[8904] = inputs[603];
    assign layer0_outputs[8905] = ~(inputs[528]);
    assign layer0_outputs[8906] = ~(inputs[835]) | (inputs[674]);
    assign layer0_outputs[8907] = (inputs[213]) | (inputs[619]);
    assign layer0_outputs[8908] = ~(inputs[27]);
    assign layer0_outputs[8909] = ~(inputs[724]) | (inputs[609]);
    assign layer0_outputs[8910] = (inputs[896]) & ~(inputs[18]);
    assign layer0_outputs[8911] = (inputs[942]) ^ (inputs[673]);
    assign layer0_outputs[8912] = (inputs[898]) | (inputs[915]);
    assign layer0_outputs[8913] = ~((inputs[511]) & (inputs[410]));
    assign layer0_outputs[8914] = ~(inputs[368]) | (inputs[973]);
    assign layer0_outputs[8915] = ~(inputs[432]);
    assign layer0_outputs[8916] = ~(inputs[664]) | (inputs[359]);
    assign layer0_outputs[8917] = ~((inputs[557]) ^ (inputs[876]));
    assign layer0_outputs[8918] = (inputs[175]) & (inputs[112]);
    assign layer0_outputs[8919] = ~((inputs[364]) ^ (inputs[377]));
    assign layer0_outputs[8920] = ~(inputs[295]);
    assign layer0_outputs[8921] = 1'b0;
    assign layer0_outputs[8922] = ~(inputs[181]);
    assign layer0_outputs[8923] = ~((inputs[542]) | (inputs[211]));
    assign layer0_outputs[8924] = ~((inputs[86]) | (inputs[652]));
    assign layer0_outputs[8925] = (inputs[514]) & ~(inputs[687]);
    assign layer0_outputs[8926] = ~(inputs[407]);
    assign layer0_outputs[8927] = inputs[680];
    assign layer0_outputs[8928] = ~(inputs[35]) | (inputs[322]);
    assign layer0_outputs[8929] = ~(inputs[78]);
    assign layer0_outputs[8930] = ~((inputs[851]) ^ (inputs[980]));
    assign layer0_outputs[8931] = ~((inputs[742]) ^ (inputs[838]));
    assign layer0_outputs[8932] = ~((inputs[756]) ^ (inputs[641]));
    assign layer0_outputs[8933] = ~(inputs[230]);
    assign layer0_outputs[8934] = ~(inputs[912]);
    assign layer0_outputs[8935] = inputs[100];
    assign layer0_outputs[8936] = inputs[680];
    assign layer0_outputs[8937] = inputs[73];
    assign layer0_outputs[8938] = ~((inputs[735]) ^ (inputs[134]));
    assign layer0_outputs[8939] = ~((inputs[67]) ^ (inputs[592]));
    assign layer0_outputs[8940] = (inputs[154]) & ~(inputs[858]);
    assign layer0_outputs[8941] = ~((inputs[699]) ^ (inputs[379]));
    assign layer0_outputs[8942] = ~((inputs[254]) | (inputs[344]));
    assign layer0_outputs[8943] = (inputs[406]) & ~(inputs[133]);
    assign layer0_outputs[8944] = ~(inputs[719]) | (inputs[345]);
    assign layer0_outputs[8945] = ~((inputs[541]) ^ (inputs[263]));
    assign layer0_outputs[8946] = ~((inputs[121]) ^ (inputs[594]));
    assign layer0_outputs[8947] = ~(inputs[247]);
    assign layer0_outputs[8948] = ~((inputs[252]) | (inputs[415]));
    assign layer0_outputs[8949] = ~((inputs[54]) | (inputs[300]));
    assign layer0_outputs[8950] = ~(inputs[591]);
    assign layer0_outputs[8951] = ~((inputs[926]) | (inputs[559]));
    assign layer0_outputs[8952] = inputs[917];
    assign layer0_outputs[8953] = ~(inputs[595]);
    assign layer0_outputs[8954] = ~(inputs[492]) | (inputs[667]);
    assign layer0_outputs[8955] = (inputs[288]) ^ (inputs[654]);
    assign layer0_outputs[8956] = inputs[47];
    assign layer0_outputs[8957] = ~((inputs[59]) | (inputs[114]));
    assign layer0_outputs[8958] = ~((inputs[198]) | (inputs[980]));
    assign layer0_outputs[8959] = ~(inputs[529]);
    assign layer0_outputs[8960] = (inputs[485]) & ~(inputs[63]);
    assign layer0_outputs[8961] = (inputs[916]) | (inputs[498]);
    assign layer0_outputs[8962] = ~((inputs[773]) ^ (inputs[28]));
    assign layer0_outputs[8963] = ~(inputs[276]);
    assign layer0_outputs[8964] = ~(inputs[111]);
    assign layer0_outputs[8965] = ~(inputs[481]) | (inputs[109]);
    assign layer0_outputs[8966] = ~(inputs[812]);
    assign layer0_outputs[8967] = ~((inputs[701]) ^ (inputs[500]));
    assign layer0_outputs[8968] = ~(inputs[112]) | (inputs[94]);
    assign layer0_outputs[8969] = inputs[889];
    assign layer0_outputs[8970] = (inputs[1016]) & (inputs[516]);
    assign layer0_outputs[8971] = (inputs[917]) & ~(inputs[442]);
    assign layer0_outputs[8972] = ~((inputs[207]) ^ (inputs[296]));
    assign layer0_outputs[8973] = 1'b0;
    assign layer0_outputs[8974] = (inputs[245]) | (inputs[93]);
    assign layer0_outputs[8975] = ~((inputs[179]) | (inputs[443]));
    assign layer0_outputs[8976] = ~((inputs[87]) ^ (inputs[850]));
    assign layer0_outputs[8977] = (inputs[626]) | (inputs[933]);
    assign layer0_outputs[8978] = 1'b1;
    assign layer0_outputs[8979] = ~(inputs[694]) | (inputs[84]);
    assign layer0_outputs[8980] = (inputs[208]) | (inputs[985]);
    assign layer0_outputs[8981] = (inputs[983]) & ~(inputs[864]);
    assign layer0_outputs[8982] = inputs[969];
    assign layer0_outputs[8983] = ~((inputs[927]) ^ (inputs[855]));
    assign layer0_outputs[8984] = ~(inputs[399]) | (inputs[110]);
    assign layer0_outputs[8985] = inputs[715];
    assign layer0_outputs[8986] = inputs[614];
    assign layer0_outputs[8987] = (inputs[818]) ^ (inputs[29]);
    assign layer0_outputs[8988] = (inputs[894]) | (inputs[90]);
    assign layer0_outputs[8989] = ~((inputs[628]) ^ (inputs[985]));
    assign layer0_outputs[8990] = ~(inputs[670]) | (inputs[842]);
    assign layer0_outputs[8991] = ~(inputs[680]);
    assign layer0_outputs[8992] = ~((inputs[107]) | (inputs[242]));
    assign layer0_outputs[8993] = (inputs[556]) & (inputs[491]);
    assign layer0_outputs[8994] = ~(inputs[906]);
    assign layer0_outputs[8995] = ~((inputs[454]) | (inputs[878]));
    assign layer0_outputs[8996] = ~(inputs[177]);
    assign layer0_outputs[8997] = ~(inputs[348]);
    assign layer0_outputs[8998] = ~(inputs[373]) | (inputs[25]);
    assign layer0_outputs[8999] = inputs[782];
    assign layer0_outputs[9000] = (inputs[582]) & ~(inputs[244]);
    assign layer0_outputs[9001] = ~(inputs[5]);
    assign layer0_outputs[9002] = 1'b0;
    assign layer0_outputs[9003] = ~(inputs[947]);
    assign layer0_outputs[9004] = (inputs[257]) & (inputs[68]);
    assign layer0_outputs[9005] = inputs[770];
    assign layer0_outputs[9006] = (inputs[841]) ^ (inputs[98]);
    assign layer0_outputs[9007] = ~(inputs[735]) | (inputs[632]);
    assign layer0_outputs[9008] = inputs[753];
    assign layer0_outputs[9009] = (inputs[807]) & ~(inputs[251]);
    assign layer0_outputs[9010] = ~(inputs[967]);
    assign layer0_outputs[9011] = ~(inputs[249]);
    assign layer0_outputs[9012] = (inputs[853]) & (inputs[580]);
    assign layer0_outputs[9013] = (inputs[830]) ^ (inputs[382]);
    assign layer0_outputs[9014] = ~((inputs[54]) | (inputs[483]));
    assign layer0_outputs[9015] = 1'b1;
    assign layer0_outputs[9016] = (inputs[726]) & ~(inputs[230]);
    assign layer0_outputs[9017] = ~((inputs[7]) | (inputs[461]));
    assign layer0_outputs[9018] = ~((inputs[31]) ^ (inputs[634]));
    assign layer0_outputs[9019] = ~(inputs[52]) | (inputs[825]);
    assign layer0_outputs[9020] = ~((inputs[740]) | (inputs[739]));
    assign layer0_outputs[9021] = (inputs[718]) | (inputs[199]);
    assign layer0_outputs[9022] = inputs[234];
    assign layer0_outputs[9023] = ~((inputs[114]) | (inputs[199]));
    assign layer0_outputs[9024] = ~((inputs[866]) | (inputs[839]));
    assign layer0_outputs[9025] = (inputs[139]) & ~(inputs[517]);
    assign layer0_outputs[9026] = (inputs[52]) & (inputs[196]);
    assign layer0_outputs[9027] = (inputs[49]) ^ (inputs[646]);
    assign layer0_outputs[9028] = ~((inputs[372]) & (inputs[435]));
    assign layer0_outputs[9029] = inputs[209];
    assign layer0_outputs[9030] = (inputs[408]) | (inputs[705]);
    assign layer0_outputs[9031] = ~((inputs[423]) & (inputs[503]));
    assign layer0_outputs[9032] = 1'b0;
    assign layer0_outputs[9033] = ~(inputs[793]);
    assign layer0_outputs[9034] = 1'b1;
    assign layer0_outputs[9035] = ~((inputs[611]) | (inputs[493]));
    assign layer0_outputs[9036] = 1'b1;
    assign layer0_outputs[9037] = ~(inputs[182]);
    assign layer0_outputs[9038] = ~(inputs[273]) | (inputs[335]);
    assign layer0_outputs[9039] = ~(inputs[839]) | (inputs[513]);
    assign layer0_outputs[9040] = ~((inputs[563]) | (inputs[407]));
    assign layer0_outputs[9041] = ~((inputs[219]) | (inputs[65]));
    assign layer0_outputs[9042] = (inputs[56]) | (inputs[650]);
    assign layer0_outputs[9043] = (inputs[879]) & ~(inputs[854]);
    assign layer0_outputs[9044] = (inputs[961]) & ~(inputs[183]);
    assign layer0_outputs[9045] = ~(inputs[710]) | (inputs[28]);
    assign layer0_outputs[9046] = (inputs[992]) ^ (inputs[234]);
    assign layer0_outputs[9047] = (inputs[891]) & ~(inputs[153]);
    assign layer0_outputs[9048] = ~((inputs[198]) | (inputs[569]));
    assign layer0_outputs[9049] = ~((inputs[700]) ^ (inputs[990]));
    assign layer0_outputs[9050] = ~((inputs[978]) | (inputs[304]));
    assign layer0_outputs[9051] = ~(inputs[764]);
    assign layer0_outputs[9052] = inputs[661];
    assign layer0_outputs[9053] = ~(inputs[368]);
    assign layer0_outputs[9054] = (inputs[731]) ^ (inputs[138]);
    assign layer0_outputs[9055] = ~(inputs[537]) | (inputs[798]);
    assign layer0_outputs[9056] = (inputs[620]) & (inputs[896]);
    assign layer0_outputs[9057] = inputs[12];
    assign layer0_outputs[9058] = inputs[79];
    assign layer0_outputs[9059] = (inputs[506]) | (inputs[754]);
    assign layer0_outputs[9060] = inputs[911];
    assign layer0_outputs[9061] = ~(inputs[358]) | (inputs[589]);
    assign layer0_outputs[9062] = inputs[715];
    assign layer0_outputs[9063] = ~(inputs[217]);
    assign layer0_outputs[9064] = ~((inputs[531]) | (inputs[870]));
    assign layer0_outputs[9065] = 1'b1;
    assign layer0_outputs[9066] = inputs[871];
    assign layer0_outputs[9067] = ~((inputs[500]) | (inputs[494]));
    assign layer0_outputs[9068] = inputs[584];
    assign layer0_outputs[9069] = ~((inputs[991]) | (inputs[532]));
    assign layer0_outputs[9070] = (inputs[534]) | (inputs[569]);
    assign layer0_outputs[9071] = ~((inputs[81]) | (inputs[223]));
    assign layer0_outputs[9072] = ~(inputs[317]) | (inputs[733]);
    assign layer0_outputs[9073] = (inputs[890]) | (inputs[392]);
    assign layer0_outputs[9074] = inputs[745];
    assign layer0_outputs[9075] = 1'b0;
    assign layer0_outputs[9076] = (inputs[248]) ^ (inputs[188]);
    assign layer0_outputs[9077] = ~(inputs[565]) | (inputs[1023]);
    assign layer0_outputs[9078] = ~((inputs[351]) ^ (inputs[369]));
    assign layer0_outputs[9079] = (inputs[484]) ^ (inputs[644]);
    assign layer0_outputs[9080] = ~((inputs[863]) | (inputs[515]));
    assign layer0_outputs[9081] = (inputs[330]) & ~(inputs[67]);
    assign layer0_outputs[9082] = 1'b1;
    assign layer0_outputs[9083] = (inputs[111]) | (inputs[787]);
    assign layer0_outputs[9084] = ~((inputs[606]) & (inputs[669]));
    assign layer0_outputs[9085] = ~(inputs[209]);
    assign layer0_outputs[9086] = inputs[242];
    assign layer0_outputs[9087] = ~(inputs[855]);
    assign layer0_outputs[9088] = (inputs[427]) & ~(inputs[201]);
    assign layer0_outputs[9089] = ~(inputs[486]);
    assign layer0_outputs[9090] = ~(inputs[930]);
    assign layer0_outputs[9091] = ~((inputs[232]) | (inputs[436]));
    assign layer0_outputs[9092] = ~(inputs[283]) | (inputs[676]);
    assign layer0_outputs[9093] = ~((inputs[230]) | (inputs[494]));
    assign layer0_outputs[9094] = 1'b0;
    assign layer0_outputs[9095] = (inputs[944]) ^ (inputs[1007]);
    assign layer0_outputs[9096] = (inputs[702]) & ~(inputs[202]);
    assign layer0_outputs[9097] = (inputs[686]) | (inputs[996]);
    assign layer0_outputs[9098] = ~((inputs[403]) ^ (inputs[30]));
    assign layer0_outputs[9099] = inputs[866];
    assign layer0_outputs[9100] = inputs[600];
    assign layer0_outputs[9101] = 1'b0;
    assign layer0_outputs[9102] = inputs[818];
    assign layer0_outputs[9103] = ~(inputs[323]) | (inputs[944]);
    assign layer0_outputs[9104] = ~(inputs[364]);
    assign layer0_outputs[9105] = inputs[205];
    assign layer0_outputs[9106] = ~(inputs[87]) | (inputs[350]);
    assign layer0_outputs[9107] = ~((inputs[14]) | (inputs[976]));
    assign layer0_outputs[9108] = (inputs[303]) | (inputs[1007]);
    assign layer0_outputs[9109] = 1'b0;
    assign layer0_outputs[9110] = 1'b1;
    assign layer0_outputs[9111] = (inputs[624]) | (inputs[11]);
    assign layer0_outputs[9112] = (inputs[535]) | (inputs[568]);
    assign layer0_outputs[9113] = (inputs[839]) & ~(inputs[795]);
    assign layer0_outputs[9114] = ~((inputs[249]) ^ (inputs[333]));
    assign layer0_outputs[9115] = inputs[50];
    assign layer0_outputs[9116] = ~(inputs[376]);
    assign layer0_outputs[9117] = (inputs[293]) & ~(inputs[575]);
    assign layer0_outputs[9118] = (inputs[766]) ^ (inputs[634]);
    assign layer0_outputs[9119] = (inputs[653]) | (inputs[991]);
    assign layer0_outputs[9120] = inputs[730];
    assign layer0_outputs[9121] = ~(inputs[174]);
    assign layer0_outputs[9122] = ~(inputs[344]) | (inputs[269]);
    assign layer0_outputs[9123] = (inputs[175]) & ~(inputs[432]);
    assign layer0_outputs[9124] = ~((inputs[188]) | (inputs[169]));
    assign layer0_outputs[9125] = ~(inputs[351]) | (inputs[543]);
    assign layer0_outputs[9126] = ~(inputs[471]) | (inputs[995]);
    assign layer0_outputs[9127] = (inputs[137]) | (inputs[928]);
    assign layer0_outputs[9128] = ~((inputs[477]) ^ (inputs[587]));
    assign layer0_outputs[9129] = ~(inputs[998]) | (inputs[903]);
    assign layer0_outputs[9130] = ~(inputs[717]) | (inputs[302]);
    assign layer0_outputs[9131] = 1'b0;
    assign layer0_outputs[9132] = (inputs[550]) ^ (inputs[3]);
    assign layer0_outputs[9133] = ~((inputs[992]) | (inputs[185]));
    assign layer0_outputs[9134] = (inputs[21]) | (inputs[7]);
    assign layer0_outputs[9135] = inputs[657];
    assign layer0_outputs[9136] = (inputs[36]) & (inputs[26]);
    assign layer0_outputs[9137] = ~(inputs[800]) | (inputs[856]);
    assign layer0_outputs[9138] = inputs[525];
    assign layer0_outputs[9139] = (inputs[911]) | (inputs[866]);
    assign layer0_outputs[9140] = inputs[439];
    assign layer0_outputs[9141] = ~(inputs[600]) | (inputs[410]);
    assign layer0_outputs[9142] = (inputs[746]) & (inputs[924]);
    assign layer0_outputs[9143] = ~(inputs[910]);
    assign layer0_outputs[9144] = inputs[403];
    assign layer0_outputs[9145] = inputs[846];
    assign layer0_outputs[9146] = inputs[567];
    assign layer0_outputs[9147] = (inputs[169]) | (inputs[474]);
    assign layer0_outputs[9148] = 1'b0;
    assign layer0_outputs[9149] = inputs[240];
    assign layer0_outputs[9150] = 1'b1;
    assign layer0_outputs[9151] = inputs[376];
    assign layer0_outputs[9152] = (inputs[956]) & ~(inputs[143]);
    assign layer0_outputs[9153] = ~(inputs[175]) | (inputs[256]);
    assign layer0_outputs[9154] = ~((inputs[98]) | (inputs[250]));
    assign layer0_outputs[9155] = ~(inputs[650]) | (inputs[763]);
    assign layer0_outputs[9156] = ~((inputs[339]) ^ (inputs[39]));
    assign layer0_outputs[9157] = inputs[918];
    assign layer0_outputs[9158] = 1'b0;
    assign layer0_outputs[9159] = (inputs[274]) | (inputs[337]);
    assign layer0_outputs[9160] = ~((inputs[122]) | (inputs[792]));
    assign layer0_outputs[9161] = inputs[490];
    assign layer0_outputs[9162] = ~(inputs[372]);
    assign layer0_outputs[9163] = inputs[493];
    assign layer0_outputs[9164] = ~(inputs[907]);
    assign layer0_outputs[9165] = (inputs[523]) & ~(inputs[792]);
    assign layer0_outputs[9166] = (inputs[152]) ^ (inputs[236]);
    assign layer0_outputs[9167] = ~((inputs[180]) ^ (inputs[160]));
    assign layer0_outputs[9168] = ~(inputs[684]);
    assign layer0_outputs[9169] = ~(inputs[1009]);
    assign layer0_outputs[9170] = ~((inputs[362]) | (inputs[729]));
    assign layer0_outputs[9171] = (inputs[319]) & ~(inputs[823]);
    assign layer0_outputs[9172] = (inputs[912]) ^ (inputs[882]);
    assign layer0_outputs[9173] = (inputs[135]) | (inputs[747]);
    assign layer0_outputs[9174] = ~(inputs[333]) | (inputs[480]);
    assign layer0_outputs[9175] = (inputs[428]) & ~(inputs[150]);
    assign layer0_outputs[9176] = ~(inputs[608]);
    assign layer0_outputs[9177] = 1'b0;
    assign layer0_outputs[9178] = (inputs[211]) & ~(inputs[420]);
    assign layer0_outputs[9179] = ~(inputs[786]);
    assign layer0_outputs[9180] = (inputs[929]) ^ (inputs[742]);
    assign layer0_outputs[9181] = inputs[922];
    assign layer0_outputs[9182] = (inputs[871]) | (inputs[436]);
    assign layer0_outputs[9183] = ~((inputs[241]) | (inputs[734]));
    assign layer0_outputs[9184] = ~((inputs[870]) ^ (inputs[1015]));
    assign layer0_outputs[9185] = (inputs[578]) ^ (inputs[487]);
    assign layer0_outputs[9186] = ~(inputs[682]);
    assign layer0_outputs[9187] = ~(inputs[458]) | (inputs[546]);
    assign layer0_outputs[9188] = inputs[245];
    assign layer0_outputs[9189] = ~((inputs[173]) | (inputs[761]));
    assign layer0_outputs[9190] = ~((inputs[722]) ^ (inputs[543]));
    assign layer0_outputs[9191] = (inputs[148]) ^ (inputs[237]);
    assign layer0_outputs[9192] = ~(inputs[276]) | (inputs[78]);
    assign layer0_outputs[9193] = (inputs[245]) | (inputs[238]);
    assign layer0_outputs[9194] = ~((inputs[5]) | (inputs[523]));
    assign layer0_outputs[9195] = (inputs[437]) & ~(inputs[605]);
    assign layer0_outputs[9196] = ~(inputs[360]) | (inputs[992]);
    assign layer0_outputs[9197] = ~(inputs[523]);
    assign layer0_outputs[9198] = 1'b1;
    assign layer0_outputs[9199] = (inputs[824]) & ~(inputs[695]);
    assign layer0_outputs[9200] = ~(inputs[41]);
    assign layer0_outputs[9201] = ~((inputs[6]) | (inputs[999]));
    assign layer0_outputs[9202] = (inputs[1016]) & ~(inputs[1013]);
    assign layer0_outputs[9203] = ~(inputs[384]) | (inputs[540]);
    assign layer0_outputs[9204] = (inputs[265]) ^ (inputs[889]);
    assign layer0_outputs[9205] = inputs[254];
    assign layer0_outputs[9206] = ~((inputs[535]) | (inputs[283]));
    assign layer0_outputs[9207] = ~(inputs[854]) | (inputs[184]);
    assign layer0_outputs[9208] = ~((inputs[253]) | (inputs[810]));
    assign layer0_outputs[9209] = ~(inputs[778]) | (inputs[948]);
    assign layer0_outputs[9210] = (inputs[424]) & ~(inputs[143]);
    assign layer0_outputs[9211] = (inputs[185]) & ~(inputs[955]);
    assign layer0_outputs[9212] = (inputs[487]) | (inputs[200]);
    assign layer0_outputs[9213] = inputs[489];
    assign layer0_outputs[9214] = (inputs[10]) & ~(inputs[479]);
    assign layer0_outputs[9215] = (inputs[328]) | (inputs[796]);
    assign layer0_outputs[9216] = inputs[559];
    assign layer0_outputs[9217] = (inputs[782]) | (inputs[206]);
    assign layer0_outputs[9218] = inputs[558];
    assign layer0_outputs[9219] = (inputs[178]) & ~(inputs[7]);
    assign layer0_outputs[9220] = ~((inputs[527]) | (inputs[228]));
    assign layer0_outputs[9221] = ~((inputs[1016]) | (inputs[344]));
    assign layer0_outputs[9222] = (inputs[664]) | (inputs[201]);
    assign layer0_outputs[9223] = (inputs[324]) & ~(inputs[506]);
    assign layer0_outputs[9224] = ~((inputs[685]) ^ (inputs[353]));
    assign layer0_outputs[9225] = (inputs[164]) & (inputs[322]);
    assign layer0_outputs[9226] = ~((inputs[78]) | (inputs[1002]));
    assign layer0_outputs[9227] = (inputs[246]) ^ (inputs[130]);
    assign layer0_outputs[9228] = (inputs[446]) & (inputs[180]);
    assign layer0_outputs[9229] = inputs[814];
    assign layer0_outputs[9230] = ~(inputs[424]);
    assign layer0_outputs[9231] = ~((inputs[206]) | (inputs[496]));
    assign layer0_outputs[9232] = ~((inputs[647]) | (inputs[982]));
    assign layer0_outputs[9233] = ~(inputs[751]);
    assign layer0_outputs[9234] = inputs[501];
    assign layer0_outputs[9235] = inputs[850];
    assign layer0_outputs[9236] = ~(inputs[648]) | (inputs[708]);
    assign layer0_outputs[9237] = inputs[67];
    assign layer0_outputs[9238] = inputs[622];
    assign layer0_outputs[9239] = inputs[80];
    assign layer0_outputs[9240] = (inputs[373]) | (inputs[76]);
    assign layer0_outputs[9241] = ~((inputs[274]) | (inputs[815]));
    assign layer0_outputs[9242] = ~((inputs[943]) | (inputs[761]));
    assign layer0_outputs[9243] = 1'b1;
    assign layer0_outputs[9244] = ~(inputs[852]) | (inputs[362]);
    assign layer0_outputs[9245] = ~(inputs[240]) | (inputs[283]);
    assign layer0_outputs[9246] = (inputs[573]) ^ (inputs[922]);
    assign layer0_outputs[9247] = inputs[79];
    assign layer0_outputs[9248] = inputs[241];
    assign layer0_outputs[9249] = (inputs[192]) & ~(inputs[991]);
    assign layer0_outputs[9250] = ~((inputs[612]) | (inputs[781]));
    assign layer0_outputs[9251] = (inputs[270]) ^ (inputs[268]);
    assign layer0_outputs[9252] = ~((inputs[197]) ^ (inputs[757]));
    assign layer0_outputs[9253] = (inputs[957]) | (inputs[111]);
    assign layer0_outputs[9254] = ~(inputs[426]);
    assign layer0_outputs[9255] = ~(inputs[459]);
    assign layer0_outputs[9256] = inputs[758];
    assign layer0_outputs[9257] = ~((inputs[631]) ^ (inputs[54]));
    assign layer0_outputs[9258] = ~((inputs[22]) ^ (inputs[155]));
    assign layer0_outputs[9259] = ~(inputs[130]);
    assign layer0_outputs[9260] = (inputs[714]) & ~(inputs[571]);
    assign layer0_outputs[9261] = (inputs[614]) | (inputs[490]);
    assign layer0_outputs[9262] = ~((inputs[106]) & (inputs[106]));
    assign layer0_outputs[9263] = inputs[711];
    assign layer0_outputs[9264] = ~(inputs[889]) | (inputs[864]);
    assign layer0_outputs[9265] = ~((inputs[131]) | (inputs[690]));
    assign layer0_outputs[9266] = (inputs[988]) & ~(inputs[110]);
    assign layer0_outputs[9267] = (inputs[336]) | (inputs[241]);
    assign layer0_outputs[9268] = inputs[451];
    assign layer0_outputs[9269] = inputs[532];
    assign layer0_outputs[9270] = ~(inputs[273]);
    assign layer0_outputs[9271] = inputs[325];
    assign layer0_outputs[9272] = (inputs[247]) & ~(inputs[25]);
    assign layer0_outputs[9273] = 1'b0;
    assign layer0_outputs[9274] = ~(inputs[915]);
    assign layer0_outputs[9275] = ~(inputs[0]) | (inputs[178]);
    assign layer0_outputs[9276] = ~((inputs[267]) | (inputs[903]));
    assign layer0_outputs[9277] = (inputs[563]) & ~(inputs[83]);
    assign layer0_outputs[9278] = (inputs[1007]) & ~(inputs[941]);
    assign layer0_outputs[9279] = ~((inputs[422]) | (inputs[848]));
    assign layer0_outputs[9280] = ~((inputs[960]) ^ (inputs[411]));
    assign layer0_outputs[9281] = (inputs[620]) & ~(inputs[948]);
    assign layer0_outputs[9282] = (inputs[294]) & ~(inputs[318]);
    assign layer0_outputs[9283] = ~((inputs[298]) ^ (inputs[505]));
    assign layer0_outputs[9284] = (inputs[12]) ^ (inputs[882]);
    assign layer0_outputs[9285] = inputs[943];
    assign layer0_outputs[9286] = (inputs[903]) ^ (inputs[405]);
    assign layer0_outputs[9287] = ~((inputs[532]) | (inputs[499]));
    assign layer0_outputs[9288] = (inputs[1011]) | (inputs[559]);
    assign layer0_outputs[9289] = (inputs[771]) & ~(inputs[58]);
    assign layer0_outputs[9290] = ~(inputs[624]);
    assign layer0_outputs[9291] = inputs[455];
    assign layer0_outputs[9292] = ~(inputs[199]);
    assign layer0_outputs[9293] = (inputs[451]) | (inputs[975]);
    assign layer0_outputs[9294] = (inputs[507]) | (inputs[536]);
    assign layer0_outputs[9295] = ~(inputs[812]);
    assign layer0_outputs[9296] = (inputs[794]) & (inputs[928]);
    assign layer0_outputs[9297] = ~(inputs[246]) | (inputs[223]);
    assign layer0_outputs[9298] = ~(inputs[612]) | (inputs[13]);
    assign layer0_outputs[9299] = (inputs[34]) | (inputs[459]);
    assign layer0_outputs[9300] = ~(inputs[598]) | (inputs[187]);
    assign layer0_outputs[9301] = inputs[827];
    assign layer0_outputs[9302] = inputs[633];
    assign layer0_outputs[9303] = inputs[85];
    assign layer0_outputs[9304] = (inputs[757]) | (inputs[262]);
    assign layer0_outputs[9305] = inputs[96];
    assign layer0_outputs[9306] = ~(inputs[554]) | (inputs[321]);
    assign layer0_outputs[9307] = ~((inputs[162]) & (inputs[833]));
    assign layer0_outputs[9308] = ~(inputs[368]);
    assign layer0_outputs[9309] = inputs[686];
    assign layer0_outputs[9310] = (inputs[497]) & ~(inputs[656]);
    assign layer0_outputs[9311] = (inputs[664]) & ~(inputs[28]);
    assign layer0_outputs[9312] = ~((inputs[863]) ^ (inputs[147]));
    assign layer0_outputs[9313] = inputs[470];
    assign layer0_outputs[9314] = ~((inputs[438]) | (inputs[394]));
    assign layer0_outputs[9315] = (inputs[847]) & ~(inputs[122]);
    assign layer0_outputs[9316] = inputs[371];
    assign layer0_outputs[9317] = inputs[527];
    assign layer0_outputs[9318] = ~((inputs[359]) | (inputs[432]));
    assign layer0_outputs[9319] = (inputs[398]) & ~(inputs[807]);
    assign layer0_outputs[9320] = ~(inputs[432]) | (inputs[989]);
    assign layer0_outputs[9321] = (inputs[234]) | (inputs[99]);
    assign layer0_outputs[9322] = (inputs[357]) ^ (inputs[271]);
    assign layer0_outputs[9323] = (inputs[759]) | (inputs[583]);
    assign layer0_outputs[9324] = ~((inputs[779]) ^ (inputs[646]));
    assign layer0_outputs[9325] = (inputs[716]) ^ (inputs[615]);
    assign layer0_outputs[9326] = inputs[654];
    assign layer0_outputs[9327] = ~((inputs[136]) ^ (inputs[297]));
    assign layer0_outputs[9328] = ~(inputs[154]) | (inputs[421]);
    assign layer0_outputs[9329] = ~((inputs[790]) | (inputs[521]));
    assign layer0_outputs[9330] = (inputs[630]) | (inputs[601]);
    assign layer0_outputs[9331] = ~((inputs[388]) ^ (inputs[603]));
    assign layer0_outputs[9332] = ~(inputs[801]) | (inputs[14]);
    assign layer0_outputs[9333] = inputs[520];
    assign layer0_outputs[9334] = ~(inputs[679]);
    assign layer0_outputs[9335] = (inputs[138]) & ~(inputs[46]);
    assign layer0_outputs[9336] = ~((inputs[805]) & (inputs[758]));
    assign layer0_outputs[9337] = ~((inputs[42]) & (inputs[677]));
    assign layer0_outputs[9338] = (inputs[698]) & ~(inputs[606]);
    assign layer0_outputs[9339] = 1'b0;
    assign layer0_outputs[9340] = ~(inputs[434]);
    assign layer0_outputs[9341] = ~(inputs[916]);
    assign layer0_outputs[9342] = (inputs[708]) | (inputs[509]);
    assign layer0_outputs[9343] = ~((inputs[565]) | (inputs[906]));
    assign layer0_outputs[9344] = ~((inputs[43]) ^ (inputs[413]));
    assign layer0_outputs[9345] = ~(inputs[157]);
    assign layer0_outputs[9346] = inputs[553];
    assign layer0_outputs[9347] = ~((inputs[551]) ^ (inputs[620]));
    assign layer0_outputs[9348] = ~(inputs[493]) | (inputs[935]);
    assign layer0_outputs[9349] = ~(inputs[219]);
    assign layer0_outputs[9350] = inputs[308];
    assign layer0_outputs[9351] = (inputs[882]) ^ (inputs[43]);
    assign layer0_outputs[9352] = inputs[426];
    assign layer0_outputs[9353] = (inputs[361]) & ~(inputs[934]);
    assign layer0_outputs[9354] = (inputs[618]) & (inputs[721]);
    assign layer0_outputs[9355] = (inputs[392]) & ~(inputs[348]);
    assign layer0_outputs[9356] = ~(inputs[280]) | (inputs[286]);
    assign layer0_outputs[9357] = ~((inputs[595]) ^ (inputs[645]));
    assign layer0_outputs[9358] = 1'b0;
    assign layer0_outputs[9359] = ~(inputs[953]);
    assign layer0_outputs[9360] = (inputs[75]) ^ (inputs[502]);
    assign layer0_outputs[9361] = (inputs[730]) ^ (inputs[908]);
    assign layer0_outputs[9362] = ~(inputs[704]) | (inputs[418]);
    assign layer0_outputs[9363] = ~(inputs[627]) | (inputs[292]);
    assign layer0_outputs[9364] = (inputs[790]) | (inputs[200]);
    assign layer0_outputs[9365] = 1'b1;
    assign layer0_outputs[9366] = ~(inputs[587]) | (inputs[741]);
    assign layer0_outputs[9367] = ~((inputs[708]) ^ (inputs[142]));
    assign layer0_outputs[9368] = ~(inputs[808]);
    assign layer0_outputs[9369] = (inputs[37]) & (inputs[977]);
    assign layer0_outputs[9370] = ~((inputs[966]) | (inputs[192]));
    assign layer0_outputs[9371] = ~(inputs[594]) | (inputs[296]);
    assign layer0_outputs[9372] = ~((inputs[930]) & (inputs[783]));
    assign layer0_outputs[9373] = ~((inputs[869]) & (inputs[629]));
    assign layer0_outputs[9374] = ~(inputs[690]);
    assign layer0_outputs[9375] = ~((inputs[271]) | (inputs[919]));
    assign layer0_outputs[9376] = (inputs[589]) & ~(inputs[613]);
    assign layer0_outputs[9377] = ~((inputs[926]) ^ (inputs[213]));
    assign layer0_outputs[9378] = inputs[174];
    assign layer0_outputs[9379] = (inputs[110]) & ~(inputs[869]);
    assign layer0_outputs[9380] = ~(inputs[801]) | (inputs[705]);
    assign layer0_outputs[9381] = (inputs[680]) | (inputs[80]);
    assign layer0_outputs[9382] = ~((inputs[976]) & (inputs[390]));
    assign layer0_outputs[9383] = 1'b1;
    assign layer0_outputs[9384] = (inputs[705]) | (inputs[10]);
    assign layer0_outputs[9385] = (inputs[831]) | (inputs[642]);
    assign layer0_outputs[9386] = ~(inputs[469]) | (inputs[135]);
    assign layer0_outputs[9387] = (inputs[492]) & ~(inputs[984]);
    assign layer0_outputs[9388] = ~((inputs[199]) ^ (inputs[340]));
    assign layer0_outputs[9389] = ~(inputs[166]) | (inputs[582]);
    assign layer0_outputs[9390] = ~((inputs[321]) | (inputs[51]));
    assign layer0_outputs[9391] = ~((inputs[814]) & (inputs[1008]));
    assign layer0_outputs[9392] = (inputs[923]) | (inputs[410]);
    assign layer0_outputs[9393] = inputs[757];
    assign layer0_outputs[9394] = ~((inputs[161]) ^ (inputs[711]));
    assign layer0_outputs[9395] = (inputs[443]) & ~(inputs[88]);
    assign layer0_outputs[9396] = ~((inputs[591]) | (inputs[318]));
    assign layer0_outputs[9397] = ~(inputs[1005]) | (inputs[870]);
    assign layer0_outputs[9398] = ~((inputs[449]) & (inputs[769]));
    assign layer0_outputs[9399] = ~((inputs[484]) & (inputs[75]));
    assign layer0_outputs[9400] = (inputs[715]) ^ (inputs[841]);
    assign layer0_outputs[9401] = (inputs[593]) ^ (inputs[8]);
    assign layer0_outputs[9402] = inputs[690];
    assign layer0_outputs[9403] = ~(inputs[552]);
    assign layer0_outputs[9404] = (inputs[148]) & ~(inputs[1016]);
    assign layer0_outputs[9405] = inputs[238];
    assign layer0_outputs[9406] = ~(inputs[590]);
    assign layer0_outputs[9407] = (inputs[517]) & ~(inputs[31]);
    assign layer0_outputs[9408] = ~(inputs[340]) | (inputs[551]);
    assign layer0_outputs[9409] = ~((inputs[933]) ^ (inputs[574]));
    assign layer0_outputs[9410] = (inputs[187]) ^ (inputs[263]);
    assign layer0_outputs[9411] = ~(inputs[454]) | (inputs[740]);
    assign layer0_outputs[9412] = inputs[69];
    assign layer0_outputs[9413] = ~((inputs[122]) | (inputs[456]));
    assign layer0_outputs[9414] = (inputs[713]) & ~(inputs[862]);
    assign layer0_outputs[9415] = ~(inputs[346]);
    assign layer0_outputs[9416] = inputs[77];
    assign layer0_outputs[9417] = ~((inputs[32]) ^ (inputs[302]));
    assign layer0_outputs[9418] = ~(inputs[803]);
    assign layer0_outputs[9419] = ~((inputs[486]) | (inputs[23]));
    assign layer0_outputs[9420] = (inputs[783]) & ~(inputs[390]);
    assign layer0_outputs[9421] = (inputs[714]) ^ (inputs[338]);
    assign layer0_outputs[9422] = ~(inputs[218]) | (inputs[448]);
    assign layer0_outputs[9423] = (inputs[84]) & ~(inputs[1009]);
    assign layer0_outputs[9424] = ~(inputs[184]);
    assign layer0_outputs[9425] = inputs[741];
    assign layer0_outputs[9426] = 1'b1;
    assign layer0_outputs[9427] = (inputs[461]) & ~(inputs[606]);
    assign layer0_outputs[9428] = ~(inputs[441]);
    assign layer0_outputs[9429] = inputs[94];
    assign layer0_outputs[9430] = (inputs[16]) | (inputs[101]);
    assign layer0_outputs[9431] = ~((inputs[962]) | (inputs[558]));
    assign layer0_outputs[9432] = inputs[948];
    assign layer0_outputs[9433] = (inputs[527]) ^ (inputs[419]);
    assign layer0_outputs[9434] = (inputs[623]) | (inputs[925]);
    assign layer0_outputs[9435] = 1'b0;
    assign layer0_outputs[9436] = (inputs[681]) | (inputs[640]);
    assign layer0_outputs[9437] = 1'b0;
    assign layer0_outputs[9438] = (inputs[227]) | (inputs[511]);
    assign layer0_outputs[9439] = ~((inputs[494]) ^ (inputs[24]));
    assign layer0_outputs[9440] = (inputs[578]) & ~(inputs[391]);
    assign layer0_outputs[9441] = (inputs[816]) ^ (inputs[28]);
    assign layer0_outputs[9442] = ~(inputs[312]);
    assign layer0_outputs[9443] = (inputs[77]) & ~(inputs[930]);
    assign layer0_outputs[9444] = ~(inputs[250]);
    assign layer0_outputs[9445] = ~((inputs[909]) | (inputs[1]));
    assign layer0_outputs[9446] = inputs[591];
    assign layer0_outputs[9447] = (inputs[872]) & (inputs[595]);
    assign layer0_outputs[9448] = ~((inputs[268]) | (inputs[334]));
    assign layer0_outputs[9449] = (inputs[326]) & ~(inputs[940]);
    assign layer0_outputs[9450] = inputs[643];
    assign layer0_outputs[9451] = inputs[339];
    assign layer0_outputs[9452] = ~((inputs[839]) | (inputs[419]));
    assign layer0_outputs[9453] = ~((inputs[189]) | (inputs[967]));
    assign layer0_outputs[9454] = 1'b0;
    assign layer0_outputs[9455] = inputs[588];
    assign layer0_outputs[9456] = ~((inputs[108]) ^ (inputs[316]));
    assign layer0_outputs[9457] = inputs[436];
    assign layer0_outputs[9458] = ~(inputs[750]) | (inputs[164]);
    assign layer0_outputs[9459] = inputs[298];
    assign layer0_outputs[9460] = (inputs[370]) | (inputs[577]);
    assign layer0_outputs[9461] = (inputs[903]) | (inputs[403]);
    assign layer0_outputs[9462] = ~((inputs[440]) ^ (inputs[227]));
    assign layer0_outputs[9463] = (inputs[418]) | (inputs[171]);
    assign layer0_outputs[9464] = (inputs[907]) & ~(inputs[386]);
    assign layer0_outputs[9465] = ~(inputs[419]) | (inputs[772]);
    assign layer0_outputs[9466] = (inputs[807]) ^ (inputs[604]);
    assign layer0_outputs[9467] = (inputs[357]) & ~(inputs[102]);
    assign layer0_outputs[9468] = ~(inputs[717]);
    assign layer0_outputs[9469] = (inputs[1012]) ^ (inputs[40]);
    assign layer0_outputs[9470] = ~((inputs[1006]) | (inputs[125]));
    assign layer0_outputs[9471] = ~(inputs[712]) | (inputs[187]);
    assign layer0_outputs[9472] = ~((inputs[876]) | (inputs[920]));
    assign layer0_outputs[9473] = inputs[628];
    assign layer0_outputs[9474] = (inputs[791]) & ~(inputs[126]);
    assign layer0_outputs[9475] = ~((inputs[773]) ^ (inputs[217]));
    assign layer0_outputs[9476] = ~(inputs[711]);
    assign layer0_outputs[9477] = (inputs[382]) & (inputs[980]);
    assign layer0_outputs[9478] = ~(inputs[188]);
    assign layer0_outputs[9479] = inputs[592];
    assign layer0_outputs[9480] = inputs[766];
    assign layer0_outputs[9481] = ~(inputs[922]);
    assign layer0_outputs[9482] = (inputs[859]) ^ (inputs[916]);
    assign layer0_outputs[9483] = (inputs[533]) & ~(inputs[203]);
    assign layer0_outputs[9484] = inputs[633];
    assign layer0_outputs[9485] = (inputs[796]) ^ (inputs[346]);
    assign layer0_outputs[9486] = ~((inputs[478]) & (inputs[73]));
    assign layer0_outputs[9487] = ~(inputs[370]);
    assign layer0_outputs[9488] = ~(inputs[655]) | (inputs[762]);
    assign layer0_outputs[9489] = ~((inputs[243]) | (inputs[959]));
    assign layer0_outputs[9490] = ~(inputs[145]) | (inputs[326]);
    assign layer0_outputs[9491] = ~((inputs[524]) | (inputs[576]));
    assign layer0_outputs[9492] = inputs[256];
    assign layer0_outputs[9493] = ~((inputs[325]) | (inputs[431]));
    assign layer0_outputs[9494] = ~((inputs[901]) | (inputs[1014]));
    assign layer0_outputs[9495] = 1'b1;
    assign layer0_outputs[9496] = ~((inputs[701]) & (inputs[901]));
    assign layer0_outputs[9497] = (inputs[208]) & ~(inputs[706]);
    assign layer0_outputs[9498] = ~((inputs[30]) & (inputs[444]));
    assign layer0_outputs[9499] = ~(inputs[816]) | (inputs[481]);
    assign layer0_outputs[9500] = ~((inputs[1015]) | (inputs[62]));
    assign layer0_outputs[9501] = ~((inputs[595]) ^ (inputs[450]));
    assign layer0_outputs[9502] = (inputs[687]) & ~(inputs[547]);
    assign layer0_outputs[9503] = (inputs[122]) ^ (inputs[201]);
    assign layer0_outputs[9504] = ~((inputs[379]) | (inputs[588]));
    assign layer0_outputs[9505] = ~((inputs[554]) | (inputs[488]));
    assign layer0_outputs[9506] = ~((inputs[81]) | (inputs[905]));
    assign layer0_outputs[9507] = inputs[359];
    assign layer0_outputs[9508] = (inputs[156]) | (inputs[904]);
    assign layer0_outputs[9509] = ~(inputs[364]) | (inputs[693]);
    assign layer0_outputs[9510] = ~(inputs[250]) | (inputs[412]);
    assign layer0_outputs[9511] = ~(inputs[462]) | (inputs[921]);
    assign layer0_outputs[9512] = ~((inputs[536]) ^ (inputs[4]));
    assign layer0_outputs[9513] = (inputs[198]) | (inputs[696]);
    assign layer0_outputs[9514] = ~((inputs[737]) ^ (inputs[606]));
    assign layer0_outputs[9515] = (inputs[647]) & ~(inputs[988]);
    assign layer0_outputs[9516] = (inputs[33]) ^ (inputs[106]);
    assign layer0_outputs[9517] = (inputs[499]) & ~(inputs[842]);
    assign layer0_outputs[9518] = inputs[539];
    assign layer0_outputs[9519] = (inputs[664]) & ~(inputs[472]);
    assign layer0_outputs[9520] = ~(inputs[622]) | (inputs[584]);
    assign layer0_outputs[9521] = (inputs[288]) | (inputs[164]);
    assign layer0_outputs[9522] = ~((inputs[666]) | (inputs[84]));
    assign layer0_outputs[9523] = inputs[681];
    assign layer0_outputs[9524] = ~((inputs[122]) | (inputs[80]));
    assign layer0_outputs[9525] = ~((inputs[222]) ^ (inputs[426]));
    assign layer0_outputs[9526] = ~(inputs[842]) | (inputs[700]);
    assign layer0_outputs[9527] = (inputs[767]) | (inputs[28]);
    assign layer0_outputs[9528] = ~(inputs[867]);
    assign layer0_outputs[9529] = 1'b0;
    assign layer0_outputs[9530] = ~((inputs[625]) ^ (inputs[465]));
    assign layer0_outputs[9531] = inputs[664];
    assign layer0_outputs[9532] = 1'b1;
    assign layer0_outputs[9533] = ~(inputs[703]);
    assign layer0_outputs[9534] = ~(inputs[566]);
    assign layer0_outputs[9535] = (inputs[275]) | (inputs[843]);
    assign layer0_outputs[9536] = ~(inputs[908]) | (inputs[266]);
    assign layer0_outputs[9537] = ~(inputs[562]);
    assign layer0_outputs[9538] = (inputs[737]) & ~(inputs[542]);
    assign layer0_outputs[9539] = ~(inputs[457]) | (inputs[975]);
    assign layer0_outputs[9540] = ~((inputs[279]) | (inputs[1006]));
    assign layer0_outputs[9541] = ~(inputs[53]) | (inputs[162]);
    assign layer0_outputs[9542] = (inputs[1001]) & ~(inputs[222]);
    assign layer0_outputs[9543] = (inputs[497]) | (inputs[219]);
    assign layer0_outputs[9544] = ~((inputs[938]) | (inputs[241]));
    assign layer0_outputs[9545] = ~((inputs[780]) ^ (inputs[985]));
    assign layer0_outputs[9546] = inputs[499];
    assign layer0_outputs[9547] = ~((inputs[784]) | (inputs[266]));
    assign layer0_outputs[9548] = ~((inputs[287]) | (inputs[96]));
    assign layer0_outputs[9549] = ~(inputs[968]) | (inputs[197]);
    assign layer0_outputs[9550] = ~(inputs[434]);
    assign layer0_outputs[9551] = (inputs[235]) ^ (inputs[440]);
    assign layer0_outputs[9552] = ~((inputs[37]) ^ (inputs[266]));
    assign layer0_outputs[9553] = ~((inputs[142]) | (inputs[594]));
    assign layer0_outputs[9554] = ~((inputs[142]) ^ (inputs[1009]));
    assign layer0_outputs[9555] = (inputs[598]) | (inputs[420]);
    assign layer0_outputs[9556] = (inputs[510]) | (inputs[766]);
    assign layer0_outputs[9557] = ~(inputs[429]) | (inputs[714]);
    assign layer0_outputs[9558] = inputs[277];
    assign layer0_outputs[9559] = ~((inputs[473]) ^ (inputs[535]));
    assign layer0_outputs[9560] = (inputs[121]) & ~(inputs[797]);
    assign layer0_outputs[9561] = (inputs[118]) | (inputs[675]);
    assign layer0_outputs[9562] = ~(inputs[947]);
    assign layer0_outputs[9563] = ~(inputs[368]);
    assign layer0_outputs[9564] = (inputs[784]) & (inputs[668]);
    assign layer0_outputs[9565] = inputs[507];
    assign layer0_outputs[9566] = ~(inputs[399]);
    assign layer0_outputs[9567] = (inputs[171]) | (inputs[238]);
    assign layer0_outputs[9568] = (inputs[746]) | (inputs[970]);
    assign layer0_outputs[9569] = ~((inputs[46]) & (inputs[308]));
    assign layer0_outputs[9570] = ~(inputs[579]);
    assign layer0_outputs[9571] = (inputs[646]) | (inputs[593]);
    assign layer0_outputs[9572] = (inputs[772]) & ~(inputs[696]);
    assign layer0_outputs[9573] = (inputs[92]) & (inputs[485]);
    assign layer0_outputs[9574] = (inputs[75]) & (inputs[389]);
    assign layer0_outputs[9575] = ~(inputs[613]);
    assign layer0_outputs[9576] = ~((inputs[315]) | (inputs[491]));
    assign layer0_outputs[9577] = (inputs[971]) & ~(inputs[741]);
    assign layer0_outputs[9578] = ~(inputs[615]);
    assign layer0_outputs[9579] = ~(inputs[0]);
    assign layer0_outputs[9580] = (inputs[746]) & ~(inputs[854]);
    assign layer0_outputs[9581] = (inputs[843]) & ~(inputs[763]);
    assign layer0_outputs[9582] = ~((inputs[317]) ^ (inputs[252]));
    assign layer0_outputs[9583] = (inputs[2]) ^ (inputs[963]);
    assign layer0_outputs[9584] = ~(inputs[906]) | (inputs[153]);
    assign layer0_outputs[9585] = ~(inputs[848]) | (inputs[800]);
    assign layer0_outputs[9586] = ~((inputs[745]) ^ (inputs[410]));
    assign layer0_outputs[9587] = (inputs[726]) ^ (inputs[60]);
    assign layer0_outputs[9588] = inputs[87];
    assign layer0_outputs[9589] = (inputs[512]) | (inputs[863]);
    assign layer0_outputs[9590] = inputs[214];
    assign layer0_outputs[9591] = (inputs[260]) | (inputs[785]);
    assign layer0_outputs[9592] = inputs[743];
    assign layer0_outputs[9593] = ~(inputs[701]);
    assign layer0_outputs[9594] = ~(inputs[948]) | (inputs[446]);
    assign layer0_outputs[9595] = ~((inputs[874]) | (inputs[929]));
    assign layer0_outputs[9596] = ~(inputs[811]);
    assign layer0_outputs[9597] = 1'b0;
    assign layer0_outputs[9598] = (inputs[255]) | (inputs[832]);
    assign layer0_outputs[9599] = ~(inputs[433]);
    assign layer0_outputs[9600] = inputs[524];
    assign layer0_outputs[9601] = ~(inputs[585]);
    assign layer0_outputs[9602] = (inputs[313]) ^ (inputs[467]);
    assign layer0_outputs[9603] = (inputs[975]) & ~(inputs[644]);
    assign layer0_outputs[9604] = ~((inputs[675]) | (inputs[817]));
    assign layer0_outputs[9605] = (inputs[646]) | (inputs[95]);
    assign layer0_outputs[9606] = (inputs[873]) | (inputs[262]);
    assign layer0_outputs[9607] = ~((inputs[22]) | (inputs[169]));
    assign layer0_outputs[9608] = (inputs[217]) ^ (inputs[932]);
    assign layer0_outputs[9609] = ~(inputs[524]);
    assign layer0_outputs[9610] = inputs[274];
    assign layer0_outputs[9611] = (inputs[925]) | (inputs[813]);
    assign layer0_outputs[9612] = (inputs[290]) & ~(inputs[17]);
    assign layer0_outputs[9613] = ~((inputs[248]) | (inputs[127]));
    assign layer0_outputs[9614] = ~((inputs[1013]) | (inputs[463]));
    assign layer0_outputs[9615] = inputs[716];
    assign layer0_outputs[9616] = (inputs[975]) & ~(inputs[914]);
    assign layer0_outputs[9617] = ~(inputs[584]);
    assign layer0_outputs[9618] = ~((inputs[671]) & (inputs[85]));
    assign layer0_outputs[9619] = inputs[493];
    assign layer0_outputs[9620] = ~((inputs[209]) & (inputs[237]));
    assign layer0_outputs[9621] = inputs[940];
    assign layer0_outputs[9622] = inputs[166];
    assign layer0_outputs[9623] = ~(inputs[451]) | (inputs[1021]);
    assign layer0_outputs[9624] = ~(inputs[527]);
    assign layer0_outputs[9625] = (inputs[99]) ^ (inputs[211]);
    assign layer0_outputs[9626] = inputs[277];
    assign layer0_outputs[9627] = ~(inputs[795]) | (inputs[476]);
    assign layer0_outputs[9628] = ~((inputs[214]) & (inputs[213]));
    assign layer0_outputs[9629] = ~(inputs[822]);
    assign layer0_outputs[9630] = (inputs[539]) | (inputs[505]);
    assign layer0_outputs[9631] = ~((inputs[956]) | (inputs[980]));
    assign layer0_outputs[9632] = (inputs[350]) & ~(inputs[19]);
    assign layer0_outputs[9633] = ~(inputs[762]) | (inputs[390]);
    assign layer0_outputs[9634] = (inputs[282]) & ~(inputs[925]);
    assign layer0_outputs[9635] = ~((inputs[285]) | (inputs[404]));
    assign layer0_outputs[9636] = ~((inputs[768]) ^ (inputs[626]));
    assign layer0_outputs[9637] = (inputs[602]) & ~(inputs[131]);
    assign layer0_outputs[9638] = ~((inputs[400]) | (inputs[400]));
    assign layer0_outputs[9639] = (inputs[193]) & (inputs[50]);
    assign layer0_outputs[9640] = (inputs[722]) & ~(inputs[898]);
    assign layer0_outputs[9641] = (inputs[349]) ^ (inputs[901]);
    assign layer0_outputs[9642] = (inputs[655]) | (inputs[356]);
    assign layer0_outputs[9643] = (inputs[640]) ^ (inputs[804]);
    assign layer0_outputs[9644] = (inputs[733]) | (inputs[974]);
    assign layer0_outputs[9645] = inputs[540];
    assign layer0_outputs[9646] = (inputs[35]) | (inputs[79]);
    assign layer0_outputs[9647] = ~(inputs[263]) | (inputs[704]);
    assign layer0_outputs[9648] = ~(inputs[524]);
    assign layer0_outputs[9649] = ~(inputs[528]) | (inputs[973]);
    assign layer0_outputs[9650] = ~((inputs[202]) | (inputs[454]));
    assign layer0_outputs[9651] = (inputs[447]) ^ (inputs[622]);
    assign layer0_outputs[9652] = 1'b0;
    assign layer0_outputs[9653] = (inputs[705]) ^ (inputs[265]);
    assign layer0_outputs[9654] = ~((inputs[214]) | (inputs[412]));
    assign layer0_outputs[9655] = ~((inputs[737]) & (inputs[566]));
    assign layer0_outputs[9656] = inputs[500];
    assign layer0_outputs[9657] = inputs[531];
    assign layer0_outputs[9658] = ~(inputs[272]) | (inputs[813]);
    assign layer0_outputs[9659] = 1'b0;
    assign layer0_outputs[9660] = ~((inputs[377]) | (inputs[391]));
    assign layer0_outputs[9661] = 1'b0;
    assign layer0_outputs[9662] = ~(inputs[622]) | (inputs[317]);
    assign layer0_outputs[9663] = inputs[102];
    assign layer0_outputs[9664] = ~(inputs[567]);
    assign layer0_outputs[9665] = 1'b0;
    assign layer0_outputs[9666] = ~(inputs[510]) | (inputs[777]);
    assign layer0_outputs[9667] = 1'b0;
    assign layer0_outputs[9668] = ~(inputs[626]);
    assign layer0_outputs[9669] = (inputs[28]) & ~(inputs[8]);
    assign layer0_outputs[9670] = (inputs[456]) & ~(inputs[539]);
    assign layer0_outputs[9671] = (inputs[903]) ^ (inputs[575]);
    assign layer0_outputs[9672] = (inputs[1021]) & ~(inputs[623]);
    assign layer0_outputs[9673] = ~(inputs[269]) | (inputs[517]);
    assign layer0_outputs[9674] = (inputs[870]) ^ (inputs[576]);
    assign layer0_outputs[9675] = ~((inputs[96]) & (inputs[291]));
    assign layer0_outputs[9676] = ~(inputs[94]) | (inputs[636]);
    assign layer0_outputs[9677] = (inputs[880]) & ~(inputs[242]);
    assign layer0_outputs[9678] = inputs[895];
    assign layer0_outputs[9679] = (inputs[14]) ^ (inputs[527]);
    assign layer0_outputs[9680] = ~((inputs[523]) & (inputs[274]));
    assign layer0_outputs[9681] = (inputs[927]) ^ (inputs[682]);
    assign layer0_outputs[9682] = inputs[427];
    assign layer0_outputs[9683] = inputs[792];
    assign layer0_outputs[9684] = (inputs[910]) | (inputs[915]);
    assign layer0_outputs[9685] = 1'b1;
    assign layer0_outputs[9686] = ~(inputs[272]);
    assign layer0_outputs[9687] = (inputs[61]) & (inputs[528]);
    assign layer0_outputs[9688] = (inputs[733]) ^ (inputs[64]);
    assign layer0_outputs[9689] = inputs[387];
    assign layer0_outputs[9690] = inputs[763];
    assign layer0_outputs[9691] = (inputs[395]) & ~(inputs[827]);
    assign layer0_outputs[9692] = (inputs[910]) ^ (inputs[263]);
    assign layer0_outputs[9693] = inputs[532];
    assign layer0_outputs[9694] = ~((inputs[608]) & (inputs[384]));
    assign layer0_outputs[9695] = inputs[404];
    assign layer0_outputs[9696] = ~(inputs[919]);
    assign layer0_outputs[9697] = ~(inputs[317]) | (inputs[604]);
    assign layer0_outputs[9698] = inputs[781];
    assign layer0_outputs[9699] = ~((inputs[862]) | (inputs[470]));
    assign layer0_outputs[9700] = ~((inputs[707]) | (inputs[698]));
    assign layer0_outputs[9701] = ~(inputs[816]);
    assign layer0_outputs[9702] = ~(inputs[697]) | (inputs[37]);
    assign layer0_outputs[9703] = ~((inputs[869]) ^ (inputs[876]));
    assign layer0_outputs[9704] = ~((inputs[841]) | (inputs[623]));
    assign layer0_outputs[9705] = ~(inputs[538]);
    assign layer0_outputs[9706] = ~((inputs[695]) | (inputs[833]));
    assign layer0_outputs[9707] = ~((inputs[824]) | (inputs[924]));
    assign layer0_outputs[9708] = (inputs[426]) & ~(inputs[223]);
    assign layer0_outputs[9709] = inputs[162];
    assign layer0_outputs[9710] = ~((inputs[617]) & (inputs[586]));
    assign layer0_outputs[9711] = ~((inputs[486]) ^ (inputs[302]));
    assign layer0_outputs[9712] = ~(inputs[830]) | (inputs[828]);
    assign layer0_outputs[9713] = (inputs[6]) & ~(inputs[103]);
    assign layer0_outputs[9714] = ~(inputs[1008]);
    assign layer0_outputs[9715] = ~((inputs[296]) | (inputs[375]));
    assign layer0_outputs[9716] = ~((inputs[265]) | (inputs[410]));
    assign layer0_outputs[9717] = (inputs[910]) & ~(inputs[152]);
    assign layer0_outputs[9718] = (inputs[658]) & ~(inputs[179]);
    assign layer0_outputs[9719] = (inputs[356]) & ~(inputs[121]);
    assign layer0_outputs[9720] = inputs[319];
    assign layer0_outputs[9721] = (inputs[180]) ^ (inputs[319]);
    assign layer0_outputs[9722] = 1'b1;
    assign layer0_outputs[9723] = inputs[540];
    assign layer0_outputs[9724] = ~((inputs[775]) | (inputs[395]));
    assign layer0_outputs[9725] = (inputs[693]) & ~(inputs[143]);
    assign layer0_outputs[9726] = (inputs[613]) & (inputs[195]);
    assign layer0_outputs[9727] = 1'b1;
    assign layer0_outputs[9728] = inputs[281];
    assign layer0_outputs[9729] = ~(inputs[334]);
    assign layer0_outputs[9730] = (inputs[164]) ^ (inputs[502]);
    assign layer0_outputs[9731] = inputs[29];
    assign layer0_outputs[9732] = ~(inputs[455]);
    assign layer0_outputs[9733] = inputs[988];
    assign layer0_outputs[9734] = ~((inputs[1017]) ^ (inputs[340]));
    assign layer0_outputs[9735] = (inputs[580]) & ~(inputs[410]);
    assign layer0_outputs[9736] = ~((inputs[423]) ^ (inputs[395]));
    assign layer0_outputs[9737] = (inputs[806]) | (inputs[634]);
    assign layer0_outputs[9738] = inputs[897];
    assign layer0_outputs[9739] = (inputs[83]) | (inputs[512]);
    assign layer0_outputs[9740] = ~((inputs[73]) | (inputs[949]));
    assign layer0_outputs[9741] = ~((inputs[200]) | (inputs[946]));
    assign layer0_outputs[9742] = ~((inputs[76]) & (inputs[872]));
    assign layer0_outputs[9743] = ~((inputs[431]) | (inputs[966]));
    assign layer0_outputs[9744] = inputs[560];
    assign layer0_outputs[9745] = ~(inputs[316]);
    assign layer0_outputs[9746] = ~((inputs[152]) | (inputs[123]));
    assign layer0_outputs[9747] = ~(inputs[492]);
    assign layer0_outputs[9748] = ~((inputs[217]) ^ (inputs[0]));
    assign layer0_outputs[9749] = (inputs[453]) | (inputs[499]);
    assign layer0_outputs[9750] = (inputs[896]) & ~(inputs[132]);
    assign layer0_outputs[9751] = ~((inputs[117]) | (inputs[190]));
    assign layer0_outputs[9752] = ~((inputs[136]) | (inputs[745]));
    assign layer0_outputs[9753] = (inputs[86]) | (inputs[453]);
    assign layer0_outputs[9754] = (inputs[103]) & (inputs[830]);
    assign layer0_outputs[9755] = 1'b0;
    assign layer0_outputs[9756] = ~(inputs[416]) | (inputs[921]);
    assign layer0_outputs[9757] = (inputs[891]) & ~(inputs[865]);
    assign layer0_outputs[9758] = ~(inputs[245]) | (inputs[192]);
    assign layer0_outputs[9759] = ~(inputs[26]) | (inputs[444]);
    assign layer0_outputs[9760] = (inputs[666]) ^ (inputs[1]);
    assign layer0_outputs[9761] = (inputs[964]) | (inputs[40]);
    assign layer0_outputs[9762] = ~(inputs[709]);
    assign layer0_outputs[9763] = (inputs[791]) ^ (inputs[897]);
    assign layer0_outputs[9764] = ~(inputs[386]);
    assign layer0_outputs[9765] = ~((inputs[308]) | (inputs[422]));
    assign layer0_outputs[9766] = (inputs[856]) | (inputs[363]);
    assign layer0_outputs[9767] = (inputs[21]) | (inputs[315]);
    assign layer0_outputs[9768] = ~(inputs[943]);
    assign layer0_outputs[9769] = ~((inputs[488]) & (inputs[505]));
    assign layer0_outputs[9770] = inputs[907];
    assign layer0_outputs[9771] = ~(inputs[112]);
    assign layer0_outputs[9772] = (inputs[120]) | (inputs[343]);
    assign layer0_outputs[9773] = ~(inputs[776]) | (inputs[1004]);
    assign layer0_outputs[9774] = ~((inputs[499]) ^ (inputs[507]));
    assign layer0_outputs[9775] = ~(inputs[174]);
    assign layer0_outputs[9776] = inputs[725];
    assign layer0_outputs[9777] = 1'b1;
    assign layer0_outputs[9778] = (inputs[314]) & ~(inputs[446]);
    assign layer0_outputs[9779] = inputs[950];
    assign layer0_outputs[9780] = ~((inputs[805]) | (inputs[433]));
    assign layer0_outputs[9781] = inputs[813];
    assign layer0_outputs[9782] = ~((inputs[1014]) ^ (inputs[77]));
    assign layer0_outputs[9783] = ~((inputs[394]) | (inputs[694]));
    assign layer0_outputs[9784] = (inputs[853]) & ~(inputs[674]);
    assign layer0_outputs[9785] = ~(inputs[113]) | (inputs[960]);
    assign layer0_outputs[9786] = inputs[599];
    assign layer0_outputs[9787] = (inputs[179]) | (inputs[180]);
    assign layer0_outputs[9788] = (inputs[416]) & ~(inputs[913]);
    assign layer0_outputs[9789] = (inputs[143]) | (inputs[976]);
    assign layer0_outputs[9790] = ~((inputs[412]) | (inputs[490]));
    assign layer0_outputs[9791] = ~(inputs[962]);
    assign layer0_outputs[9792] = (inputs[4]) | (inputs[803]);
    assign layer0_outputs[9793] = ~(inputs[761]) | (inputs[991]);
    assign layer0_outputs[9794] = ~(inputs[74]);
    assign layer0_outputs[9795] = (inputs[141]) | (inputs[239]);
    assign layer0_outputs[9796] = ~((inputs[37]) & (inputs[636]));
    assign layer0_outputs[9797] = ~((inputs[687]) | (inputs[145]));
    assign layer0_outputs[9798] = ~(inputs[392]);
    assign layer0_outputs[9799] = (inputs[204]) & ~(inputs[627]);
    assign layer0_outputs[9800] = (inputs[136]) ^ (inputs[892]);
    assign layer0_outputs[9801] = ~((inputs[105]) | (inputs[681]));
    assign layer0_outputs[9802] = (inputs[915]) ^ (inputs[909]);
    assign layer0_outputs[9803] = inputs[591];
    assign layer0_outputs[9804] = ~((inputs[193]) ^ (inputs[889]));
    assign layer0_outputs[9805] = (inputs[3]) & ~(inputs[892]);
    assign layer0_outputs[9806] = ~((inputs[769]) | (inputs[0]));
    assign layer0_outputs[9807] = (inputs[691]) | (inputs[605]);
    assign layer0_outputs[9808] = ~(inputs[922]) | (inputs[994]);
    assign layer0_outputs[9809] = (inputs[765]) | (inputs[576]);
    assign layer0_outputs[9810] = ~((inputs[431]) | (inputs[748]));
    assign layer0_outputs[9811] = ~(inputs[684]);
    assign layer0_outputs[9812] = (inputs[340]) | (inputs[378]);
    assign layer0_outputs[9813] = ~((inputs[426]) ^ (inputs[728]));
    assign layer0_outputs[9814] = ~((inputs[601]) | (inputs[802]));
    assign layer0_outputs[9815] = ~((inputs[924]) ^ (inputs[345]));
    assign layer0_outputs[9816] = ~((inputs[671]) ^ (inputs[238]));
    assign layer0_outputs[9817] = inputs[475];
    assign layer0_outputs[9818] = (inputs[754]) | (inputs[677]);
    assign layer0_outputs[9819] = ~(inputs[915]) | (inputs[762]);
    assign layer0_outputs[9820] = ~((inputs[342]) | (inputs[761]));
    assign layer0_outputs[9821] = inputs[22];
    assign layer0_outputs[9822] = (inputs[660]) | (inputs[936]);
    assign layer0_outputs[9823] = (inputs[211]) & ~(inputs[661]);
    assign layer0_outputs[9824] = inputs[238];
    assign layer0_outputs[9825] = (inputs[922]) | (inputs[755]);
    assign layer0_outputs[9826] = ~(inputs[657]);
    assign layer0_outputs[9827] = ~(inputs[468]);
    assign layer0_outputs[9828] = ~(inputs[201]);
    assign layer0_outputs[9829] = 1'b1;
    assign layer0_outputs[9830] = (inputs[434]) | (inputs[14]);
    assign layer0_outputs[9831] = ~(inputs[394]) | (inputs[658]);
    assign layer0_outputs[9832] = inputs[1018];
    assign layer0_outputs[9833] = (inputs[832]) & ~(inputs[9]);
    assign layer0_outputs[9834] = ~(inputs[666]);
    assign layer0_outputs[9835] = (inputs[649]) & ~(inputs[40]);
    assign layer0_outputs[9836] = ~(inputs[250]);
    assign layer0_outputs[9837] = ~(inputs[442]) | (inputs[960]);
    assign layer0_outputs[9838] = ~(inputs[646]);
    assign layer0_outputs[9839] = ~((inputs[526]) ^ (inputs[693]));
    assign layer0_outputs[9840] = (inputs[297]) ^ (inputs[379]);
    assign layer0_outputs[9841] = ~(inputs[30]);
    assign layer0_outputs[9842] = ~(inputs[740]) | (inputs[1015]);
    assign layer0_outputs[9843] = (inputs[125]) | (inputs[499]);
    assign layer0_outputs[9844] = ~((inputs[269]) ^ (inputs[536]));
    assign layer0_outputs[9845] = ~((inputs[48]) | (inputs[520]));
    assign layer0_outputs[9846] = inputs[296];
    assign layer0_outputs[9847] = (inputs[461]) & ~(inputs[39]);
    assign layer0_outputs[9848] = ~((inputs[831]) | (inputs[227]));
    assign layer0_outputs[9849] = ~(inputs[440]);
    assign layer0_outputs[9850] = ~((inputs[928]) & (inputs[930]));
    assign layer0_outputs[9851] = (inputs[857]) & (inputs[883]);
    assign layer0_outputs[9852] = ~((inputs[9]) & (inputs[620]));
    assign layer0_outputs[9853] = ~((inputs[917]) | (inputs[914]));
    assign layer0_outputs[9854] = ~((inputs[76]) ^ (inputs[540]));
    assign layer0_outputs[9855] = ~((inputs[847]) | (inputs[253]));
    assign layer0_outputs[9856] = (inputs[529]) & ~(inputs[202]);
    assign layer0_outputs[9857] = (inputs[14]) & (inputs[286]);
    assign layer0_outputs[9858] = (inputs[455]) & ~(inputs[157]);
    assign layer0_outputs[9859] = (inputs[37]) & ~(inputs[276]);
    assign layer0_outputs[9860] = (inputs[916]) & ~(inputs[1016]);
    assign layer0_outputs[9861] = ~(inputs[425]) | (inputs[516]);
    assign layer0_outputs[9862] = inputs[786];
    assign layer0_outputs[9863] = (inputs[743]) ^ (inputs[43]);
    assign layer0_outputs[9864] = (inputs[610]) & ~(inputs[168]);
    assign layer0_outputs[9865] = ~((inputs[601]) ^ (inputs[129]));
    assign layer0_outputs[9866] = ~(inputs[683]) | (inputs[863]);
    assign layer0_outputs[9867] = ~((inputs[417]) | (inputs[11]));
    assign layer0_outputs[9868] = 1'b1;
    assign layer0_outputs[9869] = (inputs[141]) | (inputs[437]);
    assign layer0_outputs[9870] = (inputs[986]) | (inputs[653]);
    assign layer0_outputs[9871] = (inputs[369]) & ~(inputs[153]);
    assign layer0_outputs[9872] = inputs[431];
    assign layer0_outputs[9873] = (inputs[990]) ^ (inputs[466]);
    assign layer0_outputs[9874] = ~((inputs[943]) | (inputs[693]));
    assign layer0_outputs[9875] = (inputs[828]) | (inputs[850]);
    assign layer0_outputs[9876] = ~((inputs[969]) ^ (inputs[983]));
    assign layer0_outputs[9877] = ~(inputs[376]);
    assign layer0_outputs[9878] = (inputs[216]) ^ (inputs[737]);
    assign layer0_outputs[9879] = ~((inputs[64]) ^ (inputs[691]));
    assign layer0_outputs[9880] = ~((inputs[313]) ^ (inputs[214]));
    assign layer0_outputs[9881] = (inputs[747]) | (inputs[842]);
    assign layer0_outputs[9882] = (inputs[145]) & ~(inputs[13]);
    assign layer0_outputs[9883] = (inputs[175]) ^ (inputs[864]);
    assign layer0_outputs[9884] = 1'b1;
    assign layer0_outputs[9885] = (inputs[229]) & ~(inputs[97]);
    assign layer0_outputs[9886] = 1'b1;
    assign layer0_outputs[9887] = inputs[662];
    assign layer0_outputs[9888] = ~((inputs[574]) ^ (inputs[487]));
    assign layer0_outputs[9889] = 1'b0;
    assign layer0_outputs[9890] = inputs[538];
    assign layer0_outputs[9891] = ~(inputs[16]);
    assign layer0_outputs[9892] = 1'b0;
    assign layer0_outputs[9893] = (inputs[746]) & ~(inputs[320]);
    assign layer0_outputs[9894] = ~(inputs[405]);
    assign layer0_outputs[9895] = ~((inputs[369]) | (inputs[1020]));
    assign layer0_outputs[9896] = (inputs[216]) & ~(inputs[833]);
    assign layer0_outputs[9897] = (inputs[1002]) ^ (inputs[319]);
    assign layer0_outputs[9898] = ~(inputs[364]) | (inputs[811]);
    assign layer0_outputs[9899] = (inputs[820]) | (inputs[443]);
    assign layer0_outputs[9900] = 1'b0;
    assign layer0_outputs[9901] = ~(inputs[596]) | (inputs[904]);
    assign layer0_outputs[9902] = ~(inputs[121]) | (inputs[743]);
    assign layer0_outputs[9903] = (inputs[984]) & ~(inputs[166]);
    assign layer0_outputs[9904] = (inputs[814]) | (inputs[421]);
    assign layer0_outputs[9905] = (inputs[924]) | (inputs[289]);
    assign layer0_outputs[9906] = (inputs[141]) | (inputs[676]);
    assign layer0_outputs[9907] = (inputs[920]) & ~(inputs[1013]);
    assign layer0_outputs[9908] = (inputs[168]) ^ (inputs[503]);
    assign layer0_outputs[9909] = 1'b0;
    assign layer0_outputs[9910] = ~((inputs[66]) & (inputs[977]));
    assign layer0_outputs[9911] = ~(inputs[338]);
    assign layer0_outputs[9912] = inputs[555];
    assign layer0_outputs[9913] = (inputs[257]) & ~(inputs[732]);
    assign layer0_outputs[9914] = (inputs[678]) & (inputs[964]);
    assign layer0_outputs[9915] = (inputs[240]) & ~(inputs[462]);
    assign layer0_outputs[9916] = ~((inputs[70]) & (inputs[137]));
    assign layer0_outputs[9917] = ~((inputs[574]) ^ (inputs[602]));
    assign layer0_outputs[9918] = ~((inputs[259]) ^ (inputs[485]));
    assign layer0_outputs[9919] = ~((inputs[448]) ^ (inputs[692]));
    assign layer0_outputs[9920] = 1'b0;
    assign layer0_outputs[9921] = (inputs[86]) ^ (inputs[396]);
    assign layer0_outputs[9922] = ~((inputs[165]) ^ (inputs[875]));
    assign layer0_outputs[9923] = ~((inputs[877]) | (inputs[423]));
    assign layer0_outputs[9924] = (inputs[945]) & ~(inputs[16]);
    assign layer0_outputs[9925] = 1'b1;
    assign layer0_outputs[9926] = ~(inputs[424]);
    assign layer0_outputs[9927] = ~(inputs[976]);
    assign layer0_outputs[9928] = ~(inputs[767]);
    assign layer0_outputs[9929] = ~((inputs[417]) ^ (inputs[774]));
    assign layer0_outputs[9930] = 1'b1;
    assign layer0_outputs[9931] = (inputs[473]) | (inputs[389]);
    assign layer0_outputs[9932] = ~(inputs[498]);
    assign layer0_outputs[9933] = ~((inputs[159]) | (inputs[895]));
    assign layer0_outputs[9934] = ~((inputs[627]) | (inputs[223]));
    assign layer0_outputs[9935] = ~((inputs[744]) | (inputs[374]));
    assign layer0_outputs[9936] = ~(inputs[1008]);
    assign layer0_outputs[9937] = ~(inputs[693]) | (inputs[1003]);
    assign layer0_outputs[9938] = ~((inputs[638]) | (inputs[127]));
    assign layer0_outputs[9939] = ~((inputs[581]) ^ (inputs[733]));
    assign layer0_outputs[9940] = (inputs[195]) | (inputs[325]);
    assign layer0_outputs[9941] = (inputs[659]) & ~(inputs[185]);
    assign layer0_outputs[9942] = ~(inputs[840]) | (inputs[981]);
    assign layer0_outputs[9943] = ~(inputs[777]);
    assign layer0_outputs[9944] = (inputs[251]) ^ (inputs[914]);
    assign layer0_outputs[9945] = (inputs[981]) | (inputs[623]);
    assign layer0_outputs[9946] = (inputs[409]) & ~(inputs[19]);
    assign layer0_outputs[9947] = ~((inputs[363]) ^ (inputs[876]));
    assign layer0_outputs[9948] = (inputs[781]) | (inputs[676]);
    assign layer0_outputs[9949] = ~(inputs[966]);
    assign layer0_outputs[9950] = inputs[464];
    assign layer0_outputs[9951] = inputs[409];
    assign layer0_outputs[9952] = ~(inputs[1019]);
    assign layer0_outputs[9953] = (inputs[494]) | (inputs[668]);
    assign layer0_outputs[9954] = (inputs[266]) | (inputs[808]);
    assign layer0_outputs[9955] = ~(inputs[282]);
    assign layer0_outputs[9956] = ~((inputs[661]) | (inputs[89]));
    assign layer0_outputs[9957] = ~(inputs[743]);
    assign layer0_outputs[9958] = ~((inputs[348]) | (inputs[91]));
    assign layer0_outputs[9959] = ~((inputs[427]) | (inputs[712]));
    assign layer0_outputs[9960] = 1'b0;
    assign layer0_outputs[9961] = ~(inputs[756]) | (inputs[970]);
    assign layer0_outputs[9962] = (inputs[429]) & ~(inputs[173]);
    assign layer0_outputs[9963] = (inputs[25]) & ~(inputs[72]);
    assign layer0_outputs[9964] = ~((inputs[327]) ^ (inputs[726]));
    assign layer0_outputs[9965] = 1'b1;
    assign layer0_outputs[9966] = ~(inputs[393]) | (inputs[582]);
    assign layer0_outputs[9967] = (inputs[937]) | (inputs[95]);
    assign layer0_outputs[9968] = ~((inputs[80]) & (inputs[81]));
    assign layer0_outputs[9969] = ~(inputs[870]);
    assign layer0_outputs[9970] = (inputs[947]) | (inputs[188]);
    assign layer0_outputs[9971] = ~(inputs[367]);
    assign layer0_outputs[9972] = (inputs[355]) & ~(inputs[706]);
    assign layer0_outputs[9973] = (inputs[582]) | (inputs[146]);
    assign layer0_outputs[9974] = (inputs[563]) ^ (inputs[200]);
    assign layer0_outputs[9975] = inputs[980];
    assign layer0_outputs[9976] = ~(inputs[415]);
    assign layer0_outputs[9977] = ~((inputs[507]) | (inputs[652]));
    assign layer0_outputs[9978] = ~(inputs[347]) | (inputs[60]);
    assign layer0_outputs[9979] = ~(inputs[868]) | (inputs[80]);
    assign layer0_outputs[9980] = inputs[338];
    assign layer0_outputs[9981] = ~((inputs[320]) | (inputs[814]));
    assign layer0_outputs[9982] = (inputs[822]) & ~(inputs[570]);
    assign layer0_outputs[9983] = ~((inputs[850]) | (inputs[1019]));
    assign layer0_outputs[9984] = ~((inputs[21]) ^ (inputs[442]));
    assign layer0_outputs[9985] = ~(inputs[791]);
    assign layer0_outputs[9986] = ~((inputs[852]) | (inputs[947]));
    assign layer0_outputs[9987] = (inputs[323]) ^ (inputs[434]);
    assign layer0_outputs[9988] = ~((inputs[353]) ^ (inputs[878]));
    assign layer0_outputs[9989] = ~(inputs[229]);
    assign layer0_outputs[9990] = (inputs[377]) & (inputs[164]);
    assign layer0_outputs[9991] = ~(inputs[1000]);
    assign layer0_outputs[9992] = ~((inputs[785]) & (inputs[846]));
    assign layer0_outputs[9993] = ~(inputs[490]);
    assign layer0_outputs[9994] = inputs[165];
    assign layer0_outputs[9995] = ~(inputs[370]);
    assign layer0_outputs[9996] = ~((inputs[643]) ^ (inputs[240]));
    assign layer0_outputs[9997] = (inputs[269]) & ~(inputs[1002]);
    assign layer0_outputs[9998] = (inputs[839]) | (inputs[479]);
    assign layer0_outputs[9999] = ~(inputs[560]);
    assign layer0_outputs[10000] = ~((inputs[397]) ^ (inputs[823]));
    assign layer0_outputs[10001] = inputs[785];
    assign layer0_outputs[10002] = ~(inputs[164]);
    assign layer0_outputs[10003] = ~(inputs[339]);
    assign layer0_outputs[10004] = ~(inputs[399]) | (inputs[207]);
    assign layer0_outputs[10005] = inputs[743];
    assign layer0_outputs[10006] = ~((inputs[392]) | (inputs[887]));
    assign layer0_outputs[10007] = ~(inputs[713]) | (inputs[543]);
    assign layer0_outputs[10008] = (inputs[695]) | (inputs[680]);
    assign layer0_outputs[10009] = inputs[214];
    assign layer0_outputs[10010] = (inputs[888]) ^ (inputs[623]);
    assign layer0_outputs[10011] = (inputs[868]) | (inputs[444]);
    assign layer0_outputs[10012] = (inputs[477]) & (inputs[381]);
    assign layer0_outputs[10013] = (inputs[126]) ^ (inputs[949]);
    assign layer0_outputs[10014] = ~((inputs[366]) ^ (inputs[272]));
    assign layer0_outputs[10015] = ~((inputs[344]) | (inputs[695]));
    assign layer0_outputs[10016] = ~(inputs[449]);
    assign layer0_outputs[10017] = (inputs[947]) & ~(inputs[771]);
    assign layer0_outputs[10018] = (inputs[126]) ^ (inputs[250]);
    assign layer0_outputs[10019] = ~((inputs[720]) ^ (inputs[420]));
    assign layer0_outputs[10020] = ~((inputs[913]) | (inputs[271]));
    assign layer0_outputs[10021] = ~((inputs[771]) ^ (inputs[287]));
    assign layer0_outputs[10022] = ~((inputs[896]) ^ (inputs[237]));
    assign layer0_outputs[10023] = 1'b1;
    assign layer0_outputs[10024] = inputs[475];
    assign layer0_outputs[10025] = ~(inputs[392]);
    assign layer0_outputs[10026] = inputs[198];
    assign layer0_outputs[10027] = (inputs[597]) ^ (inputs[72]);
    assign layer0_outputs[10028] = ~(inputs[106]) | (inputs[861]);
    assign layer0_outputs[10029] = (inputs[871]) | (inputs[938]);
    assign layer0_outputs[10030] = (inputs[301]) & ~(inputs[186]);
    assign layer0_outputs[10031] = (inputs[676]) | (inputs[925]);
    assign layer0_outputs[10032] = (inputs[180]) | (inputs[533]);
    assign layer0_outputs[10033] = (inputs[159]) & (inputs[52]);
    assign layer0_outputs[10034] = ~((inputs[718]) | (inputs[97]));
    assign layer0_outputs[10035] = ~((inputs[198]) | (inputs[481]));
    assign layer0_outputs[10036] = ~((inputs[816]) ^ (inputs[971]));
    assign layer0_outputs[10037] = ~((inputs[122]) ^ (inputs[116]));
    assign layer0_outputs[10038] = ~(inputs[207]);
    assign layer0_outputs[10039] = ~(inputs[752]) | (inputs[990]);
    assign layer0_outputs[10040] = (inputs[942]) | (inputs[21]);
    assign layer0_outputs[10041] = (inputs[434]) & ~(inputs[778]);
    assign layer0_outputs[10042] = ~(inputs[220]) | (inputs[110]);
    assign layer0_outputs[10043] = ~(inputs[530]) | (inputs[183]);
    assign layer0_outputs[10044] = ~((inputs[466]) | (inputs[954]));
    assign layer0_outputs[10045] = (inputs[776]) | (inputs[50]);
    assign layer0_outputs[10046] = ~((inputs[594]) ^ (inputs[551]));
    assign layer0_outputs[10047] = ~(inputs[277]);
    assign layer0_outputs[10048] = (inputs[718]) | (inputs[872]);
    assign layer0_outputs[10049] = inputs[583];
    assign layer0_outputs[10050] = ~(inputs[425]);
    assign layer0_outputs[10051] = ~(inputs[43]);
    assign layer0_outputs[10052] = (inputs[647]) & ~(inputs[485]);
    assign layer0_outputs[10053] = (inputs[108]) & (inputs[638]);
    assign layer0_outputs[10054] = (inputs[633]) & (inputs[440]);
    assign layer0_outputs[10055] = ~((inputs[229]) | (inputs[286]));
    assign layer0_outputs[10056] = ~((inputs[500]) ^ (inputs[560]));
    assign layer0_outputs[10057] = ~(inputs[591]);
    assign layer0_outputs[10058] = (inputs[168]) | (inputs[650]);
    assign layer0_outputs[10059] = (inputs[823]) ^ (inputs[539]);
    assign layer0_outputs[10060] = (inputs[720]) & ~(inputs[151]);
    assign layer0_outputs[10061] = (inputs[525]) & ~(inputs[667]);
    assign layer0_outputs[10062] = ~((inputs[121]) | (inputs[611]));
    assign layer0_outputs[10063] = ~((inputs[668]) & (inputs[173]));
    assign layer0_outputs[10064] = inputs[194];
    assign layer0_outputs[10065] = (inputs[758]) ^ (inputs[195]);
    assign layer0_outputs[10066] = (inputs[1019]) ^ (inputs[226]);
    assign layer0_outputs[10067] = ~((inputs[656]) ^ (inputs[606]));
    assign layer0_outputs[10068] = ~(inputs[427]) | (inputs[774]);
    assign layer0_outputs[10069] = ~((inputs[963]) & (inputs[99]));
    assign layer0_outputs[10070] = ~(inputs[431]) | (inputs[966]);
    assign layer0_outputs[10071] = ~(inputs[724]);
    assign layer0_outputs[10072] = ~(inputs[723]);
    assign layer0_outputs[10073] = ~(inputs[514]);
    assign layer0_outputs[10074] = ~(inputs[399]);
    assign layer0_outputs[10075] = ~((inputs[1021]) | (inputs[742]));
    assign layer0_outputs[10076] = inputs[976];
    assign layer0_outputs[10077] = ~((inputs[583]) | (inputs[729]));
    assign layer0_outputs[10078] = ~(inputs[278]) | (inputs[601]);
    assign layer0_outputs[10079] = ~(inputs[877]);
    assign layer0_outputs[10080] = ~((inputs[412]) & (inputs[968]));
    assign layer0_outputs[10081] = inputs[118];
    assign layer0_outputs[10082] = ~((inputs[210]) | (inputs[250]));
    assign layer0_outputs[10083] = (inputs[84]) | (inputs[268]);
    assign layer0_outputs[10084] = ~(inputs[378]) | (inputs[314]);
    assign layer0_outputs[10085] = inputs[996];
    assign layer0_outputs[10086] = inputs[728];
    assign layer0_outputs[10087] = ~((inputs[536]) | (inputs[120]));
    assign layer0_outputs[10088] = (inputs[92]) & ~(inputs[83]);
    assign layer0_outputs[10089] = ~(inputs[302]) | (inputs[1016]);
    assign layer0_outputs[10090] = ~((inputs[545]) | (inputs[231]));
    assign layer0_outputs[10091] = ~(inputs[811]) | (inputs[829]);
    assign layer0_outputs[10092] = (inputs[400]) | (inputs[784]);
    assign layer0_outputs[10093] = ~((inputs[109]) | (inputs[649]));
    assign layer0_outputs[10094] = (inputs[204]) | (inputs[440]);
    assign layer0_outputs[10095] = (inputs[394]) & ~(inputs[479]);
    assign layer0_outputs[10096] = 1'b1;
    assign layer0_outputs[10097] = ~(inputs[376]) | (inputs[634]);
    assign layer0_outputs[10098] = (inputs[357]) ^ (inputs[267]);
    assign layer0_outputs[10099] = (inputs[937]) | (inputs[659]);
    assign layer0_outputs[10100] = ~(inputs[746]) | (inputs[441]);
    assign layer0_outputs[10101] = (inputs[163]) & ~(inputs[739]);
    assign layer0_outputs[10102] = 1'b0;
    assign layer0_outputs[10103] = (inputs[882]) | (inputs[189]);
    assign layer0_outputs[10104] = (inputs[734]) ^ (inputs[235]);
    assign layer0_outputs[10105] = (inputs[346]) & ~(inputs[707]);
    assign layer0_outputs[10106] = ~(inputs[485]);
    assign layer0_outputs[10107] = (inputs[548]) & (inputs[225]);
    assign layer0_outputs[10108] = ~((inputs[268]) | (inputs[637]));
    assign layer0_outputs[10109] = ~((inputs[781]) | (inputs[11]));
    assign layer0_outputs[10110] = (inputs[427]) & ~(inputs[872]);
    assign layer0_outputs[10111] = ~(inputs[588]) | (inputs[572]);
    assign layer0_outputs[10112] = ~((inputs[892]) ^ (inputs[492]));
    assign layer0_outputs[10113] = 1'b0;
    assign layer0_outputs[10114] = (inputs[374]) & ~(inputs[934]);
    assign layer0_outputs[10115] = inputs[549];
    assign layer0_outputs[10116] = ~(inputs[402]) | (inputs[797]);
    assign layer0_outputs[10117] = (inputs[682]) | (inputs[855]);
    assign layer0_outputs[10118] = inputs[747];
    assign layer0_outputs[10119] = (inputs[593]) & (inputs[688]);
    assign layer0_outputs[10120] = ~((inputs[14]) ^ (inputs[575]));
    assign layer0_outputs[10121] = ~(inputs[535]) | (inputs[296]);
    assign layer0_outputs[10122] = ~((inputs[1016]) ^ (inputs[1022]));
    assign layer0_outputs[10123] = (inputs[545]) ^ (inputs[183]);
    assign layer0_outputs[10124] = ~(inputs[333]);
    assign layer0_outputs[10125] = (inputs[894]) ^ (inputs[208]);
    assign layer0_outputs[10126] = ~((inputs[405]) ^ (inputs[646]));
    assign layer0_outputs[10127] = ~(inputs[563]) | (inputs[743]);
    assign layer0_outputs[10128] = (inputs[240]) | (inputs[870]);
    assign layer0_outputs[10129] = (inputs[364]) | (inputs[33]);
    assign layer0_outputs[10130] = ~(inputs[215]);
    assign layer0_outputs[10131] = ~(inputs[752]);
    assign layer0_outputs[10132] = (inputs[79]) & ~(inputs[161]);
    assign layer0_outputs[10133] = 1'b1;
    assign layer0_outputs[10134] = (inputs[261]) | (inputs[204]);
    assign layer0_outputs[10135] = (inputs[555]) ^ (inputs[379]);
    assign layer0_outputs[10136] = (inputs[740]) & ~(inputs[231]);
    assign layer0_outputs[10137] = ~((inputs[715]) | (inputs[112]));
    assign layer0_outputs[10138] = (inputs[331]) & ~(inputs[579]);
    assign layer0_outputs[10139] = (inputs[530]) & ~(inputs[683]);
    assign layer0_outputs[10140] = inputs[253];
    assign layer0_outputs[10141] = (inputs[143]) | (inputs[732]);
    assign layer0_outputs[10142] = ~((inputs[128]) ^ (inputs[388]));
    assign layer0_outputs[10143] = (inputs[961]) ^ (inputs[684]);
    assign layer0_outputs[10144] = ~((inputs[809]) & (inputs[267]));
    assign layer0_outputs[10145] = (inputs[565]) & ~(inputs[705]);
    assign layer0_outputs[10146] = inputs[838];
    assign layer0_outputs[10147] = ~((inputs[620]) ^ (inputs[6]));
    assign layer0_outputs[10148] = ~((inputs[693]) | (inputs[1000]));
    assign layer0_outputs[10149] = inputs[521];
    assign layer0_outputs[10150] = 1'b0;
    assign layer0_outputs[10151] = (inputs[166]) & ~(inputs[173]);
    assign layer0_outputs[10152] = ~(inputs[673]);
    assign layer0_outputs[10153] = 1'b0;
    assign layer0_outputs[10154] = (inputs[868]) & (inputs[569]);
    assign layer0_outputs[10155] = ~(inputs[646]) | (inputs[186]);
    assign layer0_outputs[10156] = ~((inputs[172]) ^ (inputs[267]));
    assign layer0_outputs[10157] = (inputs[377]) | (inputs[814]);
    assign layer0_outputs[10158] = 1'b0;
    assign layer0_outputs[10159] = ~(inputs[527]) | (inputs[575]);
    assign layer0_outputs[10160] = inputs[677];
    assign layer0_outputs[10161] = (inputs[96]) | (inputs[301]);
    assign layer0_outputs[10162] = ~(inputs[160]) | (inputs[95]);
    assign layer0_outputs[10163] = ~(inputs[755]) | (inputs[699]);
    assign layer0_outputs[10164] = ~(inputs[954]);
    assign layer0_outputs[10165] = ~(inputs[497]) | (inputs[538]);
    assign layer0_outputs[10166] = (inputs[501]) ^ (inputs[509]);
    assign layer0_outputs[10167] = 1'b1;
    assign layer0_outputs[10168] = ~(inputs[812]);
    assign layer0_outputs[10169] = inputs[535];
    assign layer0_outputs[10170] = inputs[198];
    assign layer0_outputs[10171] = ~(inputs[212]) | (inputs[883]);
    assign layer0_outputs[10172] = (inputs[308]) | (inputs[904]);
    assign layer0_outputs[10173] = (inputs[343]) & (inputs[797]);
    assign layer0_outputs[10174] = (inputs[444]) ^ (inputs[196]);
    assign layer0_outputs[10175] = (inputs[74]) & ~(inputs[354]);
    assign layer0_outputs[10176] = ~(inputs[475]);
    assign layer0_outputs[10177] = 1'b1;
    assign layer0_outputs[10178] = ~((inputs[546]) & (inputs[474]));
    assign layer0_outputs[10179] = (inputs[180]) | (inputs[513]);
    assign layer0_outputs[10180] = ~((inputs[139]) | (inputs[428]));
    assign layer0_outputs[10181] = ~((inputs[308]) ^ (inputs[31]));
    assign layer0_outputs[10182] = ~(inputs[683]) | (inputs[318]);
    assign layer0_outputs[10183] = (inputs[285]) | (inputs[961]);
    assign layer0_outputs[10184] = (inputs[763]) | (inputs[342]);
    assign layer0_outputs[10185] = (inputs[734]) ^ (inputs[235]);
    assign layer0_outputs[10186] = ~(inputs[502]);
    assign layer0_outputs[10187] = (inputs[279]) | (inputs[240]);
    assign layer0_outputs[10188] = (inputs[174]) | (inputs[314]);
    assign layer0_outputs[10189] = ~((inputs[332]) | (inputs[16]));
    assign layer0_outputs[10190] = ~(inputs[177]) | (inputs[904]);
    assign layer0_outputs[10191] = ~((inputs[616]) | (inputs[2]));
    assign layer0_outputs[10192] = (inputs[862]) ^ (inputs[83]);
    assign layer0_outputs[10193] = (inputs[191]) | (inputs[967]);
    assign layer0_outputs[10194] = (inputs[547]) & ~(inputs[491]);
    assign layer0_outputs[10195] = ~(inputs[962]);
    assign layer0_outputs[10196] = (inputs[599]) & ~(inputs[813]);
    assign layer0_outputs[10197] = (inputs[970]) ^ (inputs[497]);
    assign layer0_outputs[10198] = ~((inputs[193]) | (inputs[851]));
    assign layer0_outputs[10199] = ~((inputs[702]) ^ (inputs[375]));
    assign layer0_outputs[10200] = ~(inputs[468]) | (inputs[365]);
    assign layer0_outputs[10201] = inputs[567];
    assign layer0_outputs[10202] = inputs[122];
    assign layer0_outputs[10203] = inputs[181];
    assign layer0_outputs[10204] = (inputs[913]) & ~(inputs[751]);
    assign layer0_outputs[10205] = (inputs[137]) ^ (inputs[820]);
    assign layer0_outputs[10206] = inputs[55];
    assign layer0_outputs[10207] = (inputs[313]) & ~(inputs[30]);
    assign layer0_outputs[10208] = (inputs[758]) ^ (inputs[967]);
    assign layer0_outputs[10209] = ~(inputs[754]);
    assign layer0_outputs[10210] = inputs[682];
    assign layer0_outputs[10211] = (inputs[821]) & ~(inputs[648]);
    assign layer0_outputs[10212] = ~((inputs[677]) ^ (inputs[306]));
    assign layer0_outputs[10213] = inputs[451];
    assign layer0_outputs[10214] = ~(inputs[751]) | (inputs[536]);
    assign layer0_outputs[10215] = ~((inputs[425]) | (inputs[904]));
    assign layer0_outputs[10216] = ~((inputs[586]) ^ (inputs[872]));
    assign layer0_outputs[10217] = 1'b1;
    assign layer0_outputs[10218] = (inputs[183]) ^ (inputs[497]);
    assign layer0_outputs[10219] = ~(inputs[251]) | (inputs[154]);
    assign layer0_outputs[10220] = (inputs[33]) | (inputs[771]);
    assign layer0_outputs[10221] = 1'b1;
    assign layer0_outputs[10222] = ~(inputs[559]);
    assign layer0_outputs[10223] = inputs[687];
    assign layer0_outputs[10224] = ~(inputs[200]);
    assign layer0_outputs[10225] = ~(inputs[586]);
    assign layer0_outputs[10226] = ~(inputs[693]) | (inputs[764]);
    assign layer0_outputs[10227] = (inputs[890]) ^ (inputs[495]);
    assign layer0_outputs[10228] = ~((inputs[431]) ^ (inputs[193]));
    assign layer0_outputs[10229] = (inputs[176]) & ~(inputs[935]);
    assign layer0_outputs[10230] = ~((inputs[670]) ^ (inputs[391]));
    assign layer0_outputs[10231] = ~((inputs[920]) | (inputs[410]));
    assign layer0_outputs[10232] = ~(inputs[279]) | (inputs[406]);
    assign layer0_outputs[10233] = ~(inputs[350]);
    assign layer0_outputs[10234] = ~((inputs[188]) ^ (inputs[349]));
    assign layer0_outputs[10235] = ~((inputs[98]) & (inputs[823]));
    assign layer0_outputs[10236] = 1'b1;
    assign layer0_outputs[10237] = (inputs[814]) | (inputs[346]);
    assign layer0_outputs[10238] = inputs[117];
    assign layer0_outputs[10239] = ~((inputs[410]) ^ (inputs[380]));
    assign outputs[0] = layer0_outputs[9891];
    assign outputs[1] = layer0_outputs[5752];
    assign outputs[2] = ~(layer0_outputs[385]);
    assign outputs[3] = ~((layer0_outputs[8082]) ^ (layer0_outputs[8527]));
    assign outputs[4] = ~(layer0_outputs[1537]);
    assign outputs[5] = ~(layer0_outputs[9186]) | (layer0_outputs[6724]);
    assign outputs[6] = (layer0_outputs[8555]) & ~(layer0_outputs[1701]);
    assign outputs[7] = ~((layer0_outputs[6148]) ^ (layer0_outputs[3738]));
    assign outputs[8] = ~(layer0_outputs[1886]) | (layer0_outputs[2157]);
    assign outputs[9] = 1'b1;
    assign outputs[10] = ~(layer0_outputs[7286]);
    assign outputs[11] = ~((layer0_outputs[7922]) ^ (layer0_outputs[9798]));
    assign outputs[12] = ~(layer0_outputs[1246]);
    assign outputs[13] = layer0_outputs[2246];
    assign outputs[14] = ~((layer0_outputs[9933]) ^ (layer0_outputs[8680]));
    assign outputs[15] = ~((layer0_outputs[8145]) ^ (layer0_outputs[6272]));
    assign outputs[16] = (layer0_outputs[6415]) ^ (layer0_outputs[1225]);
    assign outputs[17] = layer0_outputs[69];
    assign outputs[18] = (layer0_outputs[670]) & (layer0_outputs[2446]);
    assign outputs[19] = ~(layer0_outputs[6785]);
    assign outputs[20] = layer0_outputs[9599];
    assign outputs[21] = ~(layer0_outputs[9194]);
    assign outputs[22] = layer0_outputs[9721];
    assign outputs[23] = layer0_outputs[8371];
    assign outputs[24] = layer0_outputs[6939];
    assign outputs[25] = ~(layer0_outputs[2645]);
    assign outputs[26] = ~((layer0_outputs[5435]) & (layer0_outputs[9664]));
    assign outputs[27] = ~(layer0_outputs[10139]);
    assign outputs[28] = (layer0_outputs[3253]) ^ (layer0_outputs[6691]);
    assign outputs[29] = (layer0_outputs[2556]) ^ (layer0_outputs[310]);
    assign outputs[30] = ~(layer0_outputs[7778]) | (layer0_outputs[6675]);
    assign outputs[31] = (layer0_outputs[2855]) & (layer0_outputs[286]);
    assign outputs[32] = ~((layer0_outputs[1435]) ^ (layer0_outputs[6032]));
    assign outputs[33] = ~(layer0_outputs[8740]);
    assign outputs[34] = (layer0_outputs[8967]) & ~(layer0_outputs[4190]);
    assign outputs[35] = (layer0_outputs[3632]) & ~(layer0_outputs[1936]);
    assign outputs[36] = ~(layer0_outputs[6490]);
    assign outputs[37] = ~(layer0_outputs[7154]) | (layer0_outputs[3033]);
    assign outputs[38] = layer0_outputs[10162];
    assign outputs[39] = layer0_outputs[6331];
    assign outputs[40] = ~((layer0_outputs[10113]) ^ (layer0_outputs[1721]));
    assign outputs[41] = layer0_outputs[5577];
    assign outputs[42] = ~(layer0_outputs[1815]);
    assign outputs[43] = ~((layer0_outputs[801]) | (layer0_outputs[9135]));
    assign outputs[44] = ~(layer0_outputs[4103]);
    assign outputs[45] = layer0_outputs[8502];
    assign outputs[46] = layer0_outputs[6262];
    assign outputs[47] = ~(layer0_outputs[10145]);
    assign outputs[48] = layer0_outputs[164];
    assign outputs[49] = ~(layer0_outputs[6643]);
    assign outputs[50] = layer0_outputs[2807];
    assign outputs[51] = (layer0_outputs[7027]) ^ (layer0_outputs[3034]);
    assign outputs[52] = ~(layer0_outputs[2633]) | (layer0_outputs[2357]);
    assign outputs[53] = ~((layer0_outputs[7199]) ^ (layer0_outputs[4660]));
    assign outputs[54] = ~((layer0_outputs[9784]) ^ (layer0_outputs[10238]));
    assign outputs[55] = ~(layer0_outputs[184]);
    assign outputs[56] = ~(layer0_outputs[4419]);
    assign outputs[57] = (layer0_outputs[3638]) & ~(layer0_outputs[1015]);
    assign outputs[58] = ~((layer0_outputs[9791]) ^ (layer0_outputs[7302]));
    assign outputs[59] = (layer0_outputs[1089]) & ~(layer0_outputs[3690]);
    assign outputs[60] = ~(layer0_outputs[2166]);
    assign outputs[61] = ~(layer0_outputs[172]);
    assign outputs[62] = ~((layer0_outputs[3012]) | (layer0_outputs[7653]));
    assign outputs[63] = ~(layer0_outputs[8895]);
    assign outputs[64] = ~(layer0_outputs[4423]);
    assign outputs[65] = (layer0_outputs[4553]) ^ (layer0_outputs[5763]);
    assign outputs[66] = layer0_outputs[879];
    assign outputs[67] = ~((layer0_outputs[3427]) & (layer0_outputs[130]));
    assign outputs[68] = ~((layer0_outputs[5354]) ^ (layer0_outputs[2122]));
    assign outputs[69] = ~(layer0_outputs[3942]);
    assign outputs[70] = (layer0_outputs[553]) ^ (layer0_outputs[3973]);
    assign outputs[71] = ~((layer0_outputs[9523]) ^ (layer0_outputs[6181]));
    assign outputs[72] = ~(layer0_outputs[8137]);
    assign outputs[73] = layer0_outputs[6662];
    assign outputs[74] = layer0_outputs[4898];
    assign outputs[75] = ~(layer0_outputs[8383]) | (layer0_outputs[7022]);
    assign outputs[76] = ~(layer0_outputs[413]);
    assign outputs[77] = layer0_outputs[7735];
    assign outputs[78] = layer0_outputs[3533];
    assign outputs[79] = layer0_outputs[7743];
    assign outputs[80] = ~(layer0_outputs[3565]);
    assign outputs[81] = layer0_outputs[9624];
    assign outputs[82] = ~((layer0_outputs[6454]) & (layer0_outputs[9232]));
    assign outputs[83] = ~(layer0_outputs[9534]);
    assign outputs[84] = layer0_outputs[1798];
    assign outputs[85] = layer0_outputs[1657];
    assign outputs[86] = (layer0_outputs[4653]) & ~(layer0_outputs[5476]);
    assign outputs[87] = (layer0_outputs[3968]) & (layer0_outputs[3076]);
    assign outputs[88] = ~(layer0_outputs[9114]);
    assign outputs[89] = (layer0_outputs[1662]) & ~(layer0_outputs[10151]);
    assign outputs[90] = (layer0_outputs[1283]) & (layer0_outputs[8872]);
    assign outputs[91] = ~(layer0_outputs[4191]);
    assign outputs[92] = ~((layer0_outputs[4890]) ^ (layer0_outputs[1940]));
    assign outputs[93] = ~(layer0_outputs[2491]);
    assign outputs[94] = layer0_outputs[7428];
    assign outputs[95] = ~(layer0_outputs[9216]) | (layer0_outputs[926]);
    assign outputs[96] = (layer0_outputs[5101]) ^ (layer0_outputs[7097]);
    assign outputs[97] = ~((layer0_outputs[2399]) & (layer0_outputs[5790]));
    assign outputs[98] = ~(layer0_outputs[4164]);
    assign outputs[99] = (layer0_outputs[3722]) & (layer0_outputs[7544]);
    assign outputs[100] = layer0_outputs[1417];
    assign outputs[101] = ~(layer0_outputs[1580]) | (layer0_outputs[1504]);
    assign outputs[102] = (layer0_outputs[7653]) ^ (layer0_outputs[4537]);
    assign outputs[103] = ~(layer0_outputs[9394]);
    assign outputs[104] = ~(layer0_outputs[5492]);
    assign outputs[105] = ~((layer0_outputs[4263]) | (layer0_outputs[8378]));
    assign outputs[106] = 1'b1;
    assign outputs[107] = ~((layer0_outputs[3252]) | (layer0_outputs[2052]));
    assign outputs[108] = (layer0_outputs[6498]) ^ (layer0_outputs[8892]);
    assign outputs[109] = ~(layer0_outputs[4947]);
    assign outputs[110] = (layer0_outputs[170]) ^ (layer0_outputs[7201]);
    assign outputs[111] = ~(layer0_outputs[1286]);
    assign outputs[112] = ~((layer0_outputs[4443]) & (layer0_outputs[6312]));
    assign outputs[113] = ~(layer0_outputs[6260]) | (layer0_outputs[1457]);
    assign outputs[114] = ~((layer0_outputs[9539]) ^ (layer0_outputs[4567]));
    assign outputs[115] = (layer0_outputs[1136]) ^ (layer0_outputs[6781]);
    assign outputs[116] = (layer0_outputs[3418]) ^ (layer0_outputs[5390]);
    assign outputs[117] = layer0_outputs[179];
    assign outputs[118] = ~(layer0_outputs[3358]);
    assign outputs[119] = ~(layer0_outputs[6678]);
    assign outputs[120] = (layer0_outputs[2609]) & ~(layer0_outputs[6912]);
    assign outputs[121] = ~((layer0_outputs[6373]) ^ (layer0_outputs[5276]));
    assign outputs[122] = ~(layer0_outputs[4842]);
    assign outputs[123] = 1'b1;
    assign outputs[124] = (layer0_outputs[4417]) ^ (layer0_outputs[4274]);
    assign outputs[125] = ~(layer0_outputs[5293]);
    assign outputs[126] = (layer0_outputs[6292]) & ~(layer0_outputs[8921]);
    assign outputs[127] = (layer0_outputs[373]) ^ (layer0_outputs[6357]);
    assign outputs[128] = ~((layer0_outputs[8823]) | (layer0_outputs[8969]));
    assign outputs[129] = ~(layer0_outputs[4485]);
    assign outputs[130] = ~(layer0_outputs[4923]);
    assign outputs[131] = ~((layer0_outputs[6672]) ^ (layer0_outputs[8471]));
    assign outputs[132] = layer0_outputs[3163];
    assign outputs[133] = (layer0_outputs[5318]) ^ (layer0_outputs[2403]);
    assign outputs[134] = ~((layer0_outputs[2852]) ^ (layer0_outputs[8435]));
    assign outputs[135] = (layer0_outputs[8699]) & ~(layer0_outputs[1790]);
    assign outputs[136] = layer0_outputs[607];
    assign outputs[137] = layer0_outputs[5232];
    assign outputs[138] = ~(layer0_outputs[8926]);
    assign outputs[139] = ~(layer0_outputs[6049]) | (layer0_outputs[9100]);
    assign outputs[140] = ~(layer0_outputs[2169]);
    assign outputs[141] = layer0_outputs[8679];
    assign outputs[142] = ~((layer0_outputs[5850]) ^ (layer0_outputs[8080]));
    assign outputs[143] = (layer0_outputs[1213]) ^ (layer0_outputs[2724]);
    assign outputs[144] = ~(layer0_outputs[7019]);
    assign outputs[145] = layer0_outputs[253];
    assign outputs[146] = ~(layer0_outputs[6625]);
    assign outputs[147] = ~(layer0_outputs[1906]);
    assign outputs[148] = ~(layer0_outputs[7947]);
    assign outputs[149] = (layer0_outputs[3469]) | (layer0_outputs[5584]);
    assign outputs[150] = layer0_outputs[1852];
    assign outputs[151] = ~(layer0_outputs[8705]);
    assign outputs[152] = layer0_outputs[5224];
    assign outputs[153] = layer0_outputs[2850];
    assign outputs[154] = ~(layer0_outputs[4170]);
    assign outputs[155] = layer0_outputs[5240];
    assign outputs[156] = layer0_outputs[1027];
    assign outputs[157] = ~(layer0_outputs[7491]);
    assign outputs[158] = (layer0_outputs[7261]) ^ (layer0_outputs[10145]);
    assign outputs[159] = 1'b1;
    assign outputs[160] = ~(layer0_outputs[4807]);
    assign outputs[161] = ~(layer0_outputs[275]);
    assign outputs[162] = layer0_outputs[2167];
    assign outputs[163] = layer0_outputs[1958];
    assign outputs[164] = ~(layer0_outputs[9563]);
    assign outputs[165] = ~(layer0_outputs[2354]);
    assign outputs[166] = layer0_outputs[1317];
    assign outputs[167] = ~(layer0_outputs[5767]);
    assign outputs[168] = 1'b1;
    assign outputs[169] = (layer0_outputs[1851]) & ~(layer0_outputs[3122]);
    assign outputs[170] = ~((layer0_outputs[5392]) | (layer0_outputs[6140]));
    assign outputs[171] = (layer0_outputs[4920]) & ~(layer0_outputs[848]);
    assign outputs[172] = ~((layer0_outputs[1753]) & (layer0_outputs[1196]));
    assign outputs[173] = ~(layer0_outputs[807]);
    assign outputs[174] = ~((layer0_outputs[4213]) ^ (layer0_outputs[8048]));
    assign outputs[175] = (layer0_outputs[7946]) ^ (layer0_outputs[6676]);
    assign outputs[176] = ~(layer0_outputs[1199]);
    assign outputs[177] = (layer0_outputs[6537]) ^ (layer0_outputs[9108]);
    assign outputs[178] = ~((layer0_outputs[4032]) ^ (layer0_outputs[6377]));
    assign outputs[179] = (layer0_outputs[212]) & (layer0_outputs[2101]);
    assign outputs[180] = ~(layer0_outputs[7001]);
    assign outputs[181] = layer0_outputs[10044];
    assign outputs[182] = layer0_outputs[8488];
    assign outputs[183] = ~(layer0_outputs[9402]);
    assign outputs[184] = ~(layer0_outputs[6301]) | (layer0_outputs[10102]);
    assign outputs[185] = (layer0_outputs[1352]) | (layer0_outputs[9542]);
    assign outputs[186] = ~(layer0_outputs[5138]);
    assign outputs[187] = ~(layer0_outputs[7601]);
    assign outputs[188] = ~((layer0_outputs[6542]) ^ (layer0_outputs[5256]));
    assign outputs[189] = ~(layer0_outputs[8108]);
    assign outputs[190] = ~(layer0_outputs[8109]) | (layer0_outputs[2133]);
    assign outputs[191] = (layer0_outputs[205]) ^ (layer0_outputs[1244]);
    assign outputs[192] = (layer0_outputs[7581]) ^ (layer0_outputs[4074]);
    assign outputs[193] = (layer0_outputs[6127]) & ~(layer0_outputs[1530]);
    assign outputs[194] = ~((layer0_outputs[7639]) ^ (layer0_outputs[1596]));
    assign outputs[195] = layer0_outputs[7200];
    assign outputs[196] = (layer0_outputs[1838]) ^ (layer0_outputs[8744]);
    assign outputs[197] = layer0_outputs[743];
    assign outputs[198] = (layer0_outputs[8318]) ^ (layer0_outputs[6113]);
    assign outputs[199] = layer0_outputs[544];
    assign outputs[200] = layer0_outputs[8958];
    assign outputs[201] = ~((layer0_outputs[7848]) ^ (layer0_outputs[6971]));
    assign outputs[202] = ~(layer0_outputs[5157]);
    assign outputs[203] = (layer0_outputs[7119]) & ~(layer0_outputs[9892]);
    assign outputs[204] = layer0_outputs[6];
    assign outputs[205] = layer0_outputs[8529];
    assign outputs[206] = ~((layer0_outputs[87]) ^ (layer0_outputs[9714]));
    assign outputs[207] = (layer0_outputs[4656]) ^ (layer0_outputs[5145]);
    assign outputs[208] = (layer0_outputs[4814]) | (layer0_outputs[5111]);
    assign outputs[209] = ~(layer0_outputs[4895]);
    assign outputs[210] = (layer0_outputs[5907]) ^ (layer0_outputs[8387]);
    assign outputs[211] = ~((layer0_outputs[751]) ^ (layer0_outputs[2391]));
    assign outputs[212] = ~(layer0_outputs[2704]);
    assign outputs[213] = layer0_outputs[3645];
    assign outputs[214] = layer0_outputs[353];
    assign outputs[215] = (layer0_outputs[870]) & ~(layer0_outputs[2754]);
    assign outputs[216] = (layer0_outputs[9267]) ^ (layer0_outputs[4176]);
    assign outputs[217] = ~((layer0_outputs[5990]) & (layer0_outputs[4529]));
    assign outputs[218] = (layer0_outputs[4542]) ^ (layer0_outputs[6903]);
    assign outputs[219] = layer0_outputs[6397];
    assign outputs[220] = ~(layer0_outputs[579]);
    assign outputs[221] = (layer0_outputs[1309]) ^ (layer0_outputs[5699]);
    assign outputs[222] = (layer0_outputs[487]) ^ (layer0_outputs[2702]);
    assign outputs[223] = (layer0_outputs[6979]) & ~(layer0_outputs[7810]);
    assign outputs[224] = layer0_outputs[721];
    assign outputs[225] = layer0_outputs[6745];
    assign outputs[226] = (layer0_outputs[2739]) & ~(layer0_outputs[5469]);
    assign outputs[227] = layer0_outputs[4141];
    assign outputs[228] = ~((layer0_outputs[3038]) ^ (layer0_outputs[2396]));
    assign outputs[229] = (layer0_outputs[3035]) & ~(layer0_outputs[2758]);
    assign outputs[230] = layer0_outputs[2501];
    assign outputs[231] = (layer0_outputs[1664]) | (layer0_outputs[5730]);
    assign outputs[232] = ~((layer0_outputs[4119]) & (layer0_outputs[8920]));
    assign outputs[233] = ~(layer0_outputs[9744]);
    assign outputs[234] = ~(layer0_outputs[1493]);
    assign outputs[235] = ~(layer0_outputs[2612]);
    assign outputs[236] = layer0_outputs[3790];
    assign outputs[237] = (layer0_outputs[1170]) & ~(layer0_outputs[7299]);
    assign outputs[238] = (layer0_outputs[2907]) ^ (layer0_outputs[7510]);
    assign outputs[239] = ~((layer0_outputs[6517]) & (layer0_outputs[9481]));
    assign outputs[240] = ~(layer0_outputs[5587]);
    assign outputs[241] = ~(layer0_outputs[6601]) | (layer0_outputs[189]);
    assign outputs[242] = ~((layer0_outputs[5575]) | (layer0_outputs[8345]));
    assign outputs[243] = ~(layer0_outputs[5490]) | (layer0_outputs[7657]);
    assign outputs[244] = (layer0_outputs[4919]) ^ (layer0_outputs[7493]);
    assign outputs[245] = ~((layer0_outputs[8733]) ^ (layer0_outputs[2575]));
    assign outputs[246] = ~((layer0_outputs[1257]) ^ (layer0_outputs[1351]));
    assign outputs[247] = ~((layer0_outputs[9056]) & (layer0_outputs[2883]));
    assign outputs[248] = ~(layer0_outputs[1368]);
    assign outputs[249] = layer0_outputs[4532];
    assign outputs[250] = ~(layer0_outputs[8416]);
    assign outputs[251] = ~(layer0_outputs[3083]) | (layer0_outputs[6805]);
    assign outputs[252] = (layer0_outputs[1506]) ^ (layer0_outputs[1859]);
    assign outputs[253] = layer0_outputs[9315];
    assign outputs[254] = ~(layer0_outputs[9410]);
    assign outputs[255] = ~((layer0_outputs[2548]) ^ (layer0_outputs[5997]));
    assign outputs[256] = (layer0_outputs[5473]) & ~(layer0_outputs[7715]);
    assign outputs[257] = layer0_outputs[2024];
    assign outputs[258] = ~(layer0_outputs[8579]);
    assign outputs[259] = ~((layer0_outputs[152]) & (layer0_outputs[7759]));
    assign outputs[260] = layer0_outputs[4748];
    assign outputs[261] = (layer0_outputs[4813]) & ~(layer0_outputs[52]);
    assign outputs[262] = ~(layer0_outputs[1833]);
    assign outputs[263] = ~((layer0_outputs[6225]) & (layer0_outputs[10126]));
    assign outputs[264] = layer0_outputs[7717];
    assign outputs[265] = ~((layer0_outputs[864]) ^ (layer0_outputs[924]));
    assign outputs[266] = (layer0_outputs[2600]) | (layer0_outputs[5036]);
    assign outputs[267] = (layer0_outputs[2786]) ^ (layer0_outputs[2614]);
    assign outputs[268] = layer0_outputs[1702];
    assign outputs[269] = ~(layer0_outputs[4340]);
    assign outputs[270] = ~((layer0_outputs[1338]) ^ (layer0_outputs[8937]));
    assign outputs[271] = ~((layer0_outputs[8858]) & (layer0_outputs[4980]));
    assign outputs[272] = layer0_outputs[9746];
    assign outputs[273] = (layer0_outputs[1507]) ^ (layer0_outputs[4464]);
    assign outputs[274] = ~((layer0_outputs[6990]) ^ (layer0_outputs[7797]));
    assign outputs[275] = layer0_outputs[891];
    assign outputs[276] = ~(layer0_outputs[7423]);
    assign outputs[277] = layer0_outputs[5377];
    assign outputs[278] = ~((layer0_outputs[7877]) | (layer0_outputs[3914]));
    assign outputs[279] = layer0_outputs[6879];
    assign outputs[280] = ~(layer0_outputs[2063]);
    assign outputs[281] = ~((layer0_outputs[7661]) ^ (layer0_outputs[2893]));
    assign outputs[282] = (layer0_outputs[6853]) ^ (layer0_outputs[6034]);
    assign outputs[283] = layer0_outputs[9901];
    assign outputs[284] = ~(layer0_outputs[7879]);
    assign outputs[285] = ~(layer0_outputs[4449]);
    assign outputs[286] = (layer0_outputs[5652]) ^ (layer0_outputs[777]);
    assign outputs[287] = ~(layer0_outputs[7774]) | (layer0_outputs[2500]);
    assign outputs[288] = ~((layer0_outputs[9434]) | (layer0_outputs[8581]));
    assign outputs[289] = ~(layer0_outputs[4991]);
    assign outputs[290] = layer0_outputs[10092];
    assign outputs[291] = ~(layer0_outputs[2512]);
    assign outputs[292] = (layer0_outputs[3089]) | (layer0_outputs[6158]);
    assign outputs[293] = ~(layer0_outputs[2229]);
    assign outputs[294] = ~(layer0_outputs[5065]);
    assign outputs[295] = ~(layer0_outputs[6730]);
    assign outputs[296] = ~(layer0_outputs[7982]);
    assign outputs[297] = layer0_outputs[1241];
    assign outputs[298] = layer0_outputs[6836];
    assign outputs[299] = ~(layer0_outputs[8018]);
    assign outputs[300] = ~(layer0_outputs[4338]);
    assign outputs[301] = layer0_outputs[6498];
    assign outputs[302] = ~(layer0_outputs[2771]);
    assign outputs[303] = (layer0_outputs[360]) & ~(layer0_outputs[1628]);
    assign outputs[304] = layer0_outputs[2110];
    assign outputs[305] = ~(layer0_outputs[2063]);
    assign outputs[306] = ~(layer0_outputs[2472]);
    assign outputs[307] = layer0_outputs[3534];
    assign outputs[308] = (layer0_outputs[1255]) & ~(layer0_outputs[7538]);
    assign outputs[309] = ~(layer0_outputs[2437]);
    assign outputs[310] = (layer0_outputs[6283]) ^ (layer0_outputs[1587]);
    assign outputs[311] = 1'b1;
    assign outputs[312] = (layer0_outputs[1787]) ^ (layer0_outputs[336]);
    assign outputs[313] = layer0_outputs[1869];
    assign outputs[314] = (layer0_outputs[9404]) ^ (layer0_outputs[5345]);
    assign outputs[315] = layer0_outputs[8856];
    assign outputs[316] = layer0_outputs[910];
    assign outputs[317] = ~(layer0_outputs[3116]);
    assign outputs[318] = layer0_outputs[3530];
    assign outputs[319] = ~(layer0_outputs[1684]);
    assign outputs[320] = ~(layer0_outputs[5547]);
    assign outputs[321] = layer0_outputs[7473];
    assign outputs[322] = ~((layer0_outputs[9301]) & (layer0_outputs[226]));
    assign outputs[323] = ~(layer0_outputs[9843]);
    assign outputs[324] = (layer0_outputs[9023]) & ~(layer0_outputs[3873]);
    assign outputs[325] = (layer0_outputs[1633]) | (layer0_outputs[7013]);
    assign outputs[326] = layer0_outputs[1345];
    assign outputs[327] = (layer0_outputs[7305]) ^ (layer0_outputs[4812]);
    assign outputs[328] = (layer0_outputs[6593]) ^ (layer0_outputs[8323]);
    assign outputs[329] = layer0_outputs[9638];
    assign outputs[330] = (layer0_outputs[3890]) ^ (layer0_outputs[3579]);
    assign outputs[331] = (layer0_outputs[1244]) & ~(layer0_outputs[5621]);
    assign outputs[332] = ~((layer0_outputs[6416]) ^ (layer0_outputs[1186]));
    assign outputs[333] = ~(layer0_outputs[8884]);
    assign outputs[334] = ~(layer0_outputs[9769]) | (layer0_outputs[6630]);
    assign outputs[335] = ~(layer0_outputs[5913]);
    assign outputs[336] = ~(layer0_outputs[4124]);
    assign outputs[337] = layer0_outputs[2055];
    assign outputs[338] = ~(layer0_outputs[2953]);
    assign outputs[339] = ~((layer0_outputs[6287]) ^ (layer0_outputs[8157]));
    assign outputs[340] = layer0_outputs[5431];
    assign outputs[341] = (layer0_outputs[9902]) ^ (layer0_outputs[1966]);
    assign outputs[342] = layer0_outputs[8315];
    assign outputs[343] = ~(layer0_outputs[6355]);
    assign outputs[344] = ~((layer0_outputs[2337]) ^ (layer0_outputs[289]));
    assign outputs[345] = (layer0_outputs[4510]) ^ (layer0_outputs[7074]);
    assign outputs[346] = ~(layer0_outputs[3779]) | (layer0_outputs[4026]);
    assign outputs[347] = layer0_outputs[5309];
    assign outputs[348] = layer0_outputs[9795];
    assign outputs[349] = (layer0_outputs[6450]) & ~(layer0_outputs[9767]);
    assign outputs[350] = ~(layer0_outputs[639]);
    assign outputs[351] = ~(layer0_outputs[5081]);
    assign outputs[352] = ~((layer0_outputs[1173]) & (layer0_outputs[7706]));
    assign outputs[353] = ~(layer0_outputs[3634]);
    assign outputs[354] = (layer0_outputs[5837]) & (layer0_outputs[471]);
    assign outputs[355] = ~(layer0_outputs[85]);
    assign outputs[356] = ~(layer0_outputs[8260]);
    assign outputs[357] = layer0_outputs[3207];
    assign outputs[358] = ~(layer0_outputs[6996]);
    assign outputs[359] = ~((layer0_outputs[7969]) ^ (layer0_outputs[4015]));
    assign outputs[360] = layer0_outputs[5784];
    assign outputs[361] = layer0_outputs[5942];
    assign outputs[362] = (layer0_outputs[8727]) | (layer0_outputs[6394]);
    assign outputs[363] = (layer0_outputs[1534]) & ~(layer0_outputs[7857]);
    assign outputs[364] = (layer0_outputs[179]) ^ (layer0_outputs[645]);
    assign outputs[365] = ~(layer0_outputs[2989]) | (layer0_outputs[4931]);
    assign outputs[366] = ~(layer0_outputs[3928]);
    assign outputs[367] = (layer0_outputs[7876]) | (layer0_outputs[2156]);
    assign outputs[368] = ~(layer0_outputs[6156]);
    assign outputs[369] = ~(layer0_outputs[8614]);
    assign outputs[370] = (layer0_outputs[6731]) & ~(layer0_outputs[8239]);
    assign outputs[371] = ~(layer0_outputs[7927]);
    assign outputs[372] = layer0_outputs[3206];
    assign outputs[373] = ~(layer0_outputs[5178]);
    assign outputs[374] = (layer0_outputs[2131]) ^ (layer0_outputs[2544]);
    assign outputs[375] = (layer0_outputs[2140]) & ~(layer0_outputs[5669]);
    assign outputs[376] = ~(layer0_outputs[5818]);
    assign outputs[377] = ~(layer0_outputs[1167]);
    assign outputs[378] = (layer0_outputs[9048]) ^ (layer0_outputs[6217]);
    assign outputs[379] = ~(layer0_outputs[4547]);
    assign outputs[380] = ~((layer0_outputs[1628]) ^ (layer0_outputs[9574]));
    assign outputs[381] = layer0_outputs[1311];
    assign outputs[382] = ~(layer0_outputs[8097]);
    assign outputs[383] = ~(layer0_outputs[6712]) | (layer0_outputs[6425]);
    assign outputs[384] = ~(layer0_outputs[3013]);
    assign outputs[385] = ~(layer0_outputs[9657]);
    assign outputs[386] = layer0_outputs[8894];
    assign outputs[387] = (layer0_outputs[6723]) & ~(layer0_outputs[1168]);
    assign outputs[388] = layer0_outputs[3130];
    assign outputs[389] = ~(layer0_outputs[2515]);
    assign outputs[390] = (layer0_outputs[2183]) & ~(layer0_outputs[7241]);
    assign outputs[391] = layer0_outputs[4068];
    assign outputs[392] = ~(layer0_outputs[10003]) | (layer0_outputs[1524]);
    assign outputs[393] = ~((layer0_outputs[9457]) | (layer0_outputs[7567]));
    assign outputs[394] = layer0_outputs[3795];
    assign outputs[395] = layer0_outputs[2759];
    assign outputs[396] = ~(layer0_outputs[227]);
    assign outputs[397] = ~((layer0_outputs[5599]) | (layer0_outputs[325]));
    assign outputs[398] = ~(layer0_outputs[6679]) | (layer0_outputs[8556]);
    assign outputs[399] = ~(layer0_outputs[3568]);
    assign outputs[400] = ~(layer0_outputs[6285]);
    assign outputs[401] = layer0_outputs[3405];
    assign outputs[402] = ~(layer0_outputs[8045]) | (layer0_outputs[7392]);
    assign outputs[403] = (layer0_outputs[1714]) & (layer0_outputs[6232]);
    assign outputs[404] = (layer0_outputs[2710]) ^ (layer0_outputs[4043]);
    assign outputs[405] = layer0_outputs[6786];
    assign outputs[406] = ~(layer0_outputs[1118]);
    assign outputs[407] = (layer0_outputs[2869]) & ~(layer0_outputs[5022]);
    assign outputs[408] = ~((layer0_outputs[2638]) & (layer0_outputs[7455]));
    assign outputs[409] = (layer0_outputs[1604]) & ~(layer0_outputs[7349]);
    assign outputs[410] = ~(layer0_outputs[4256]);
    assign outputs[411] = layer0_outputs[1426];
    assign outputs[412] = ~(layer0_outputs[3455]);
    assign outputs[413] = layer0_outputs[7283];
    assign outputs[414] = (layer0_outputs[3915]) ^ (layer0_outputs[9453]);
    assign outputs[415] = (layer0_outputs[3718]) | (layer0_outputs[9881]);
    assign outputs[416] = (layer0_outputs[7292]) ^ (layer0_outputs[2071]);
    assign outputs[417] = layer0_outputs[4487];
    assign outputs[418] = layer0_outputs[5627];
    assign outputs[419] = ~(layer0_outputs[7899]);
    assign outputs[420] = (layer0_outputs[1362]) ^ (layer0_outputs[1830]);
    assign outputs[421] = layer0_outputs[5459];
    assign outputs[422] = ~(layer0_outputs[1748]);
    assign outputs[423] = ~(layer0_outputs[8372]) | (layer0_outputs[8931]);
    assign outputs[424] = ~((layer0_outputs[2593]) ^ (layer0_outputs[9775]));
    assign outputs[425] = ~(layer0_outputs[5946]) | (layer0_outputs[518]);
    assign outputs[426] = ~((layer0_outputs[5399]) ^ (layer0_outputs[4607]));
    assign outputs[427] = layer0_outputs[2032];
    assign outputs[428] = ~((layer0_outputs[5921]) & (layer0_outputs[4887]));
    assign outputs[429] = ~(layer0_outputs[7650]);
    assign outputs[430] = (layer0_outputs[6862]) | (layer0_outputs[9725]);
    assign outputs[431] = ~(layer0_outputs[5352]);
    assign outputs[432] = layer0_outputs[3501];
    assign outputs[433] = ~((layer0_outputs[1658]) ^ (layer0_outputs[3655]));
    assign outputs[434] = ~(layer0_outputs[7433]);
    assign outputs[435] = ~(layer0_outputs[9347]);
    assign outputs[436] = ~(layer0_outputs[994]);
    assign outputs[437] = ~((layer0_outputs[167]) ^ (layer0_outputs[7483]));
    assign outputs[438] = ~((layer0_outputs[1519]) ^ (layer0_outputs[9701]));
    assign outputs[439] = (layer0_outputs[59]) ^ (layer0_outputs[1434]);
    assign outputs[440] = layer0_outputs[190];
    assign outputs[441] = layer0_outputs[775];
    assign outputs[442] = ~(layer0_outputs[1968]) | (layer0_outputs[853]);
    assign outputs[443] = ~(layer0_outputs[9245]);
    assign outputs[444] = ~(layer0_outputs[3265]);
    assign outputs[445] = ~(layer0_outputs[3474]);
    assign outputs[446] = ~((layer0_outputs[1582]) & (layer0_outputs[5296]));
    assign outputs[447] = (layer0_outputs[4750]) ^ (layer0_outputs[973]);
    assign outputs[448] = layer0_outputs[5931];
    assign outputs[449] = ~((layer0_outputs[7701]) ^ (layer0_outputs[7427]));
    assign outputs[450] = ~(layer0_outputs[4739]);
    assign outputs[451] = ~((layer0_outputs[4782]) | (layer0_outputs[8794]));
    assign outputs[452] = layer0_outputs[2829];
    assign outputs[453] = layer0_outputs[5066];
    assign outputs[454] = (layer0_outputs[7601]) ^ (layer0_outputs[3857]);
    assign outputs[455] = layer0_outputs[9146];
    assign outputs[456] = ~(layer0_outputs[8030]);
    assign outputs[457] = ~((layer0_outputs[3306]) & (layer0_outputs[2004]));
    assign outputs[458] = (layer0_outputs[1888]) ^ (layer0_outputs[549]);
    assign outputs[459] = layer0_outputs[4756];
    assign outputs[460] = layer0_outputs[9530];
    assign outputs[461] = ~((layer0_outputs[6721]) | (layer0_outputs[7970]));
    assign outputs[462] = ~(layer0_outputs[3167]) | (layer0_outputs[2172]);
    assign outputs[463] = layer0_outputs[2526];
    assign outputs[464] = ~(layer0_outputs[5895]);
    assign outputs[465] = ~(layer0_outputs[2244]);
    assign outputs[466] = (layer0_outputs[1039]) & ~(layer0_outputs[5767]);
    assign outputs[467] = (layer0_outputs[3466]) | (layer0_outputs[10184]);
    assign outputs[468] = ~(layer0_outputs[7417]);
    assign outputs[469] = ~((layer0_outputs[2651]) ^ (layer0_outputs[5578]));
    assign outputs[470] = (layer0_outputs[4354]) ^ (layer0_outputs[6687]);
    assign outputs[471] = ~((layer0_outputs[7091]) ^ (layer0_outputs[7167]));
    assign outputs[472] = (layer0_outputs[10009]) ^ (layer0_outputs[3724]);
    assign outputs[473] = ~(layer0_outputs[6496]) | (layer0_outputs[4059]);
    assign outputs[474] = (layer0_outputs[596]) & ~(layer0_outputs[8916]);
    assign outputs[475] = ~(layer0_outputs[9144]);
    assign outputs[476] = ~((layer0_outputs[4103]) & (layer0_outputs[7390]));
    assign outputs[477] = ~((layer0_outputs[4133]) | (layer0_outputs[1588]));
    assign outputs[478] = (layer0_outputs[7435]) | (layer0_outputs[5389]);
    assign outputs[479] = layer0_outputs[369];
    assign outputs[480] = (layer0_outputs[674]) & ~(layer0_outputs[903]);
    assign outputs[481] = layer0_outputs[6338];
    assign outputs[482] = ~(layer0_outputs[8869]) | (layer0_outputs[4001]);
    assign outputs[483] = (layer0_outputs[9129]) & ~(layer0_outputs[10027]);
    assign outputs[484] = (layer0_outputs[737]) & ~(layer0_outputs[946]);
    assign outputs[485] = layer0_outputs[4125];
    assign outputs[486] = layer0_outputs[8198];
    assign outputs[487] = (layer0_outputs[3919]) & ~(layer0_outputs[9573]);
    assign outputs[488] = layer0_outputs[6230];
    assign outputs[489] = ~(layer0_outputs[7947]) | (layer0_outputs[519]);
    assign outputs[490] = ~((layer0_outputs[7270]) ^ (layer0_outputs[7101]));
    assign outputs[491] = ~((layer0_outputs[8547]) ^ (layer0_outputs[3870]));
    assign outputs[492] = ~((layer0_outputs[9937]) ^ (layer0_outputs[7246]));
    assign outputs[493] = layer0_outputs[4098];
    assign outputs[494] = layer0_outputs[5093];
    assign outputs[495] = ~(layer0_outputs[4545]);
    assign outputs[496] = layer0_outputs[3186];
    assign outputs[497] = (layer0_outputs[1837]) & ~(layer0_outputs[6072]);
    assign outputs[498] = (layer0_outputs[1694]) ^ (layer0_outputs[7158]);
    assign outputs[499] = ~(layer0_outputs[88]);
    assign outputs[500] = (layer0_outputs[1531]) & ~(layer0_outputs[9115]);
    assign outputs[501] = layer0_outputs[615];
    assign outputs[502] = ~(layer0_outputs[1094]);
    assign outputs[503] = (layer0_outputs[9354]) | (layer0_outputs[4315]);
    assign outputs[504] = ~(layer0_outputs[5181]) | (layer0_outputs[969]);
    assign outputs[505] = layer0_outputs[4421];
    assign outputs[506] = ~((layer0_outputs[5323]) | (layer0_outputs[4616]));
    assign outputs[507] = layer0_outputs[3803];
    assign outputs[508] = ~(layer0_outputs[8399]) | (layer0_outputs[5211]);
    assign outputs[509] = ~(layer0_outputs[7319]) | (layer0_outputs[5317]);
    assign outputs[510] = ~(layer0_outputs[1685]);
    assign outputs[511] = ~((layer0_outputs[1855]) ^ (layer0_outputs[3732]));
    assign outputs[512] = ~(layer0_outputs[379]) | (layer0_outputs[1393]);
    assign outputs[513] = ~(layer0_outputs[3793]) | (layer0_outputs[9350]);
    assign outputs[514] = ~(layer0_outputs[3824]);
    assign outputs[515] = (layer0_outputs[1975]) & ~(layer0_outputs[6944]);
    assign outputs[516] = ~(layer0_outputs[2090]) | (layer0_outputs[6043]);
    assign outputs[517] = layer0_outputs[6839];
    assign outputs[518] = layer0_outputs[9077];
    assign outputs[519] = ~((layer0_outputs[6402]) ^ (layer0_outputs[9907]));
    assign outputs[520] = ~((layer0_outputs[2928]) & (layer0_outputs[8183]));
    assign outputs[521] = layer0_outputs[8950];
    assign outputs[522] = (layer0_outputs[4163]) & (layer0_outputs[5967]);
    assign outputs[523] = layer0_outputs[66];
    assign outputs[524] = (layer0_outputs[3697]) | (layer0_outputs[9154]);
    assign outputs[525] = ~((layer0_outputs[3573]) | (layer0_outputs[7766]));
    assign outputs[526] = ~(layer0_outputs[6115]);
    assign outputs[527] = layer0_outputs[2880];
    assign outputs[528] = ~(layer0_outputs[4990]) | (layer0_outputs[8211]);
    assign outputs[529] = ~(layer0_outputs[1690]);
    assign outputs[530] = ~(layer0_outputs[6175]);
    assign outputs[531] = ~(layer0_outputs[4481]) | (layer0_outputs[395]);
    assign outputs[532] = ~((layer0_outputs[2125]) & (layer0_outputs[8095]));
    assign outputs[533] = layer0_outputs[525];
    assign outputs[534] = ~((layer0_outputs[3541]) ^ (layer0_outputs[9034]));
    assign outputs[535] = layer0_outputs[7613];
    assign outputs[536] = (layer0_outputs[4578]) ^ (layer0_outputs[3700]);
    assign outputs[537] = layer0_outputs[3049];
    assign outputs[538] = ~((layer0_outputs[7335]) ^ (layer0_outputs[8697]));
    assign outputs[539] = (layer0_outputs[7554]) ^ (layer0_outputs[4709]);
    assign outputs[540] = layer0_outputs[4826];
    assign outputs[541] = ~(layer0_outputs[8798]);
    assign outputs[542] = ~(layer0_outputs[390]) | (layer0_outputs[9848]);
    assign outputs[543] = layer0_outputs[522];
    assign outputs[544] = ~(layer0_outputs[5109]) | (layer0_outputs[8770]);
    assign outputs[545] = ~(layer0_outputs[3169]) | (layer0_outputs[8842]);
    assign outputs[546] = (layer0_outputs[5211]) | (layer0_outputs[2212]);
    assign outputs[547] = ~((layer0_outputs[4807]) & (layer0_outputs[916]));
    assign outputs[548] = ~((layer0_outputs[8176]) & (layer0_outputs[7658]));
    assign outputs[549] = (layer0_outputs[6500]) ^ (layer0_outputs[6565]);
    assign outputs[550] = ~(layer0_outputs[965]);
    assign outputs[551] = ~(layer0_outputs[4403]);
    assign outputs[552] = ~(layer0_outputs[629]);
    assign outputs[553] = layer0_outputs[6073];
    assign outputs[554] = layer0_outputs[6227];
    assign outputs[555] = (layer0_outputs[6767]) ^ (layer0_outputs[5153]);
    assign outputs[556] = (layer0_outputs[2513]) ^ (layer0_outputs[8949]);
    assign outputs[557] = (layer0_outputs[10169]) ^ (layer0_outputs[9556]);
    assign outputs[558] = ~(layer0_outputs[10191]) | (layer0_outputs[4872]);
    assign outputs[559] = layer0_outputs[8460];
    assign outputs[560] = layer0_outputs[7155];
    assign outputs[561] = (layer0_outputs[6152]) & ~(layer0_outputs[8793]);
    assign outputs[562] = ~((layer0_outputs[3023]) & (layer0_outputs[7109]));
    assign outputs[563] = ~(layer0_outputs[7632]);
    assign outputs[564] = ~((layer0_outputs[3578]) ^ (layer0_outputs[1876]));
    assign outputs[565] = ~(layer0_outputs[1965]);
    assign outputs[566] = (layer0_outputs[734]) & ~(layer0_outputs[550]);
    assign outputs[567] = ~((layer0_outputs[1676]) ^ (layer0_outputs[9409]));
    assign outputs[568] = (layer0_outputs[1450]) | (layer0_outputs[9914]);
    assign outputs[569] = layer0_outputs[9363];
    assign outputs[570] = (layer0_outputs[2461]) | (layer0_outputs[1696]);
    assign outputs[571] = layer0_outputs[9067];
    assign outputs[572] = (layer0_outputs[4252]) | (layer0_outputs[2827]);
    assign outputs[573] = layer0_outputs[104];
    assign outputs[574] = ~(layer0_outputs[8389]);
    assign outputs[575] = ~((layer0_outputs[4192]) ^ (layer0_outputs[2654]));
    assign outputs[576] = layer0_outputs[7356];
    assign outputs[577] = ~(layer0_outputs[3765]);
    assign outputs[578] = layer0_outputs[3699];
    assign outputs[579] = ~(layer0_outputs[3461]);
    assign outputs[580] = (layer0_outputs[117]) ^ (layer0_outputs[1004]);
    assign outputs[581] = (layer0_outputs[1451]) & ~(layer0_outputs[2812]);
    assign outputs[582] = ~((layer0_outputs[4613]) | (layer0_outputs[4815]));
    assign outputs[583] = ~((layer0_outputs[3080]) & (layer0_outputs[556]));
    assign outputs[584] = (layer0_outputs[7424]) | (layer0_outputs[1711]);
    assign outputs[585] = ~(layer0_outputs[9306]);
    assign outputs[586] = layer0_outputs[9565];
    assign outputs[587] = (layer0_outputs[232]) & ~(layer0_outputs[4497]);
    assign outputs[588] = ~((layer0_outputs[9018]) & (layer0_outputs[2686]));
    assign outputs[589] = ~((layer0_outputs[6013]) | (layer0_outputs[7113]));
    assign outputs[590] = ~(layer0_outputs[587]);
    assign outputs[591] = ~((layer0_outputs[8841]) ^ (layer0_outputs[7122]));
    assign outputs[592] = layer0_outputs[7374];
    assign outputs[593] = (layer0_outputs[4645]) ^ (layer0_outputs[3030]);
    assign outputs[594] = ~(layer0_outputs[233]);
    assign outputs[595] = layer0_outputs[1235];
    assign outputs[596] = 1'b0;
    assign outputs[597] = ~((layer0_outputs[5873]) | (layer0_outputs[5049]));
    assign outputs[598] = ~((layer0_outputs[2300]) ^ (layer0_outputs[7061]));
    assign outputs[599] = ~((layer0_outputs[3321]) | (layer0_outputs[1168]));
    assign outputs[600] = ~(layer0_outputs[6872]);
    assign outputs[601] = ~(layer0_outputs[5736]);
    assign outputs[602] = ~(layer0_outputs[4688]);
    assign outputs[603] = layer0_outputs[605];
    assign outputs[604] = 1'b0;
    assign outputs[605] = ~(layer0_outputs[9326]);
    assign outputs[606] = layer0_outputs[9535];
    assign outputs[607] = ~(layer0_outputs[4350]);
    assign outputs[608] = (layer0_outputs[3269]) ^ (layer0_outputs[1026]);
    assign outputs[609] = layer0_outputs[9062];
    assign outputs[610] = (layer0_outputs[1990]) ^ (layer0_outputs[8408]);
    assign outputs[611] = layer0_outputs[7922];
    assign outputs[612] = ~(layer0_outputs[6485]);
    assign outputs[613] = ~((layer0_outputs[1593]) & (layer0_outputs[9815]));
    assign outputs[614] = ~((layer0_outputs[4856]) | (layer0_outputs[5438]));
    assign outputs[615] = ~(layer0_outputs[580]) | (layer0_outputs[4537]);
    assign outputs[616] = ~(layer0_outputs[9888]);
    assign outputs[617] = ~(layer0_outputs[2362]);
    assign outputs[618] = (layer0_outputs[5748]) & ~(layer0_outputs[6547]);
    assign outputs[619] = layer0_outputs[8083];
    assign outputs[620] = ~(layer0_outputs[5612]) | (layer0_outputs[1420]);
    assign outputs[621] = ~(layer0_outputs[6851]);
    assign outputs[622] = (layer0_outputs[4899]) & (layer0_outputs[9853]);
    assign outputs[623] = layer0_outputs[2368];
    assign outputs[624] = ~((layer0_outputs[3921]) | (layer0_outputs[9502]));
    assign outputs[625] = layer0_outputs[8571];
    assign outputs[626] = layer0_outputs[1350];
    assign outputs[627] = ~(layer0_outputs[799]);
    assign outputs[628] = (layer0_outputs[5060]) & ~(layer0_outputs[10134]);
    assign outputs[629] = (layer0_outputs[6715]) & (layer0_outputs[8395]);
    assign outputs[630] = (layer0_outputs[6220]) & ~(layer0_outputs[9215]);
    assign outputs[631] = ~((layer0_outputs[5758]) | (layer0_outputs[9750]));
    assign outputs[632] = ~(layer0_outputs[1394]);
    assign outputs[633] = layer0_outputs[6123];
    assign outputs[634] = ~((layer0_outputs[3148]) & (layer0_outputs[8833]));
    assign outputs[635] = (layer0_outputs[1334]) | (layer0_outputs[1009]);
    assign outputs[636] = ~(layer0_outputs[8364]);
    assign outputs[637] = (layer0_outputs[7470]) & ~(layer0_outputs[3416]);
    assign outputs[638] = (layer0_outputs[1501]) ^ (layer0_outputs[8192]);
    assign outputs[639] = ~(layer0_outputs[10176]);
    assign outputs[640] = (layer0_outputs[324]) | (layer0_outputs[1391]);
    assign outputs[641] = ~((layer0_outputs[252]) & (layer0_outputs[7187]));
    assign outputs[642] = (layer0_outputs[172]) ^ (layer0_outputs[443]);
    assign outputs[643] = (layer0_outputs[5971]) & (layer0_outputs[3293]);
    assign outputs[644] = (layer0_outputs[3704]) & (layer0_outputs[9942]);
    assign outputs[645] = layer0_outputs[5366];
    assign outputs[646] = ~(layer0_outputs[3611]) | (layer0_outputs[10224]);
    assign outputs[647] = (layer0_outputs[2377]) | (layer0_outputs[2457]);
    assign outputs[648] = ~(layer0_outputs[570]);
    assign outputs[649] = ~(layer0_outputs[7016]);
    assign outputs[650] = ~(layer0_outputs[7711]) | (layer0_outputs[5163]);
    assign outputs[651] = layer0_outputs[42];
    assign outputs[652] = layer0_outputs[5504];
    assign outputs[653] = (layer0_outputs[798]) ^ (layer0_outputs[5811]);
    assign outputs[654] = ~((layer0_outputs[1072]) & (layer0_outputs[5436]));
    assign outputs[655] = ~(layer0_outputs[7149]);
    assign outputs[656] = ~(layer0_outputs[2874]);
    assign outputs[657] = ~(layer0_outputs[3711]) | (layer0_outputs[4410]);
    assign outputs[658] = (layer0_outputs[9462]) ^ (layer0_outputs[10028]);
    assign outputs[659] = (layer0_outputs[5060]) & (layer0_outputs[7125]);
    assign outputs[660] = ~(layer0_outputs[9718]);
    assign outputs[661] = (layer0_outputs[5935]) & ~(layer0_outputs[6511]);
    assign outputs[662] = ~((layer0_outputs[1955]) ^ (layer0_outputs[1808]));
    assign outputs[663] = layer0_outputs[8280];
    assign outputs[664] = (layer0_outputs[4657]) & ~(layer0_outputs[9012]);
    assign outputs[665] = (layer0_outputs[10069]) | (layer0_outputs[2046]);
    assign outputs[666] = layer0_outputs[2247];
    assign outputs[667] = layer0_outputs[3483];
    assign outputs[668] = ~(layer0_outputs[7044]) | (layer0_outputs[6993]);
    assign outputs[669] = layer0_outputs[4101];
    assign outputs[670] = layer0_outputs[2748];
    assign outputs[671] = (layer0_outputs[1612]) ^ (layer0_outputs[9905]);
    assign outputs[672] = ~((layer0_outputs[711]) ^ (layer0_outputs[7703]));
    assign outputs[673] = layer0_outputs[6126];
    assign outputs[674] = ~(layer0_outputs[7001]);
    assign outputs[675] = (layer0_outputs[4970]) & (layer0_outputs[2299]);
    assign outputs[676] = layer0_outputs[905];
    assign outputs[677] = ~(layer0_outputs[2379]);
    assign outputs[678] = ~(layer0_outputs[9803]);
    assign outputs[679] = (layer0_outputs[2537]) & (layer0_outputs[3097]);
    assign outputs[680] = layer0_outputs[6917];
    assign outputs[681] = ~(layer0_outputs[46]) | (layer0_outputs[3632]);
    assign outputs[682] = ~((layer0_outputs[9356]) ^ (layer0_outputs[3935]));
    assign outputs[683] = 1'b1;
    assign outputs[684] = (layer0_outputs[7276]) ^ (layer0_outputs[8492]);
    assign outputs[685] = layer0_outputs[10105];
    assign outputs[686] = layer0_outputs[1727];
    assign outputs[687] = ~(layer0_outputs[9831]);
    assign outputs[688] = (layer0_outputs[6886]) & (layer0_outputs[2234]);
    assign outputs[689] = layer0_outputs[5086];
    assign outputs[690] = ~(layer0_outputs[1385]) | (layer0_outputs[2850]);
    assign outputs[691] = ~(layer0_outputs[4531]);
    assign outputs[692] = layer0_outputs[8989];
    assign outputs[693] = ~(layer0_outputs[3990]);
    assign outputs[694] = ~((layer0_outputs[7074]) & (layer0_outputs[4799]));
    assign outputs[695] = layer0_outputs[3930];
    assign outputs[696] = (layer0_outputs[2438]) ^ (layer0_outputs[4775]);
    assign outputs[697] = ~((layer0_outputs[8291]) ^ (layer0_outputs[6625]));
    assign outputs[698] = (layer0_outputs[9497]) ^ (layer0_outputs[1250]);
    assign outputs[699] = ~(layer0_outputs[8798]);
    assign outputs[700] = ~(layer0_outputs[8585]) | (layer0_outputs[8009]);
    assign outputs[701] = layer0_outputs[8904];
    assign outputs[702] = (layer0_outputs[5740]) & (layer0_outputs[1663]);
    assign outputs[703] = ~((layer0_outputs[9811]) & (layer0_outputs[10132]));
    assign outputs[704] = (layer0_outputs[5192]) ^ (layer0_outputs[2705]);
    assign outputs[705] = ~(layer0_outputs[1757]);
    assign outputs[706] = (layer0_outputs[5374]) & ~(layer0_outputs[5071]);
    assign outputs[707] = layer0_outputs[7470];
    assign outputs[708] = ~((layer0_outputs[3477]) & (layer0_outputs[2945]));
    assign outputs[709] = (layer0_outputs[7354]) & (layer0_outputs[5837]);
    assign outputs[710] = ~((layer0_outputs[3813]) ^ (layer0_outputs[4608]));
    assign outputs[711] = layer0_outputs[3488];
    assign outputs[712] = ~(layer0_outputs[7248]);
    assign outputs[713] = ~((layer0_outputs[2651]) | (layer0_outputs[9335]));
    assign outputs[714] = ~((layer0_outputs[1374]) ^ (layer0_outputs[390]));
    assign outputs[715] = layer0_outputs[5522];
    assign outputs[716] = layer0_outputs[7294];
    assign outputs[717] = ~(layer0_outputs[1520]);
    assign outputs[718] = layer0_outputs[3032];
    assign outputs[719] = ~(layer0_outputs[8042]);
    assign outputs[720] = layer0_outputs[3331];
    assign outputs[721] = ~(layer0_outputs[8332]);
    assign outputs[722] = (layer0_outputs[4473]) & ~(layer0_outputs[9255]);
    assign outputs[723] = layer0_outputs[6734];
    assign outputs[724] = 1'b1;
    assign outputs[725] = layer0_outputs[4806];
    assign outputs[726] = ~((layer0_outputs[5063]) & (layer0_outputs[1913]));
    assign outputs[727] = layer0_outputs[9553];
    assign outputs[728] = ~(layer0_outputs[2620]);
    assign outputs[729] = ~(layer0_outputs[7514]);
    assign outputs[730] = ~(layer0_outputs[9247]) | (layer0_outputs[5887]);
    assign outputs[731] = ~((layer0_outputs[4013]) & (layer0_outputs[10231]));
    assign outputs[732] = (layer0_outputs[5999]) & (layer0_outputs[3139]);
    assign outputs[733] = ~(layer0_outputs[6247]);
    assign outputs[734] = layer0_outputs[10129];
    assign outputs[735] = (layer0_outputs[8006]) ^ (layer0_outputs[504]);
    assign outputs[736] = ~((layer0_outputs[4273]) ^ (layer0_outputs[1556]));
    assign outputs[737] = (layer0_outputs[2055]) | (layer0_outputs[10175]);
    assign outputs[738] = layer0_outputs[7809];
    assign outputs[739] = ~((layer0_outputs[1531]) ^ (layer0_outputs[2347]));
    assign outputs[740] = ~((layer0_outputs[7816]) & (layer0_outputs[1602]));
    assign outputs[741] = (layer0_outputs[5712]) & ~(layer0_outputs[6299]);
    assign outputs[742] = ~(layer0_outputs[3004]);
    assign outputs[743] = ~(layer0_outputs[861]) | (layer0_outputs[2510]);
    assign outputs[744] = 1'b1;
    assign outputs[745] = (layer0_outputs[663]) ^ (layer0_outputs[4011]);
    assign outputs[746] = ~(layer0_outputs[7016]);
    assign outputs[747] = (layer0_outputs[5148]) & (layer0_outputs[5421]);
    assign outputs[748] = (layer0_outputs[1962]) ^ (layer0_outputs[7936]);
    assign outputs[749] = ~((layer0_outputs[1369]) ^ (layer0_outputs[10120]));
    assign outputs[750] = ~(layer0_outputs[981]);
    assign outputs[751] = ~((layer0_outputs[9825]) & (layer0_outputs[7960]));
    assign outputs[752] = ~((layer0_outputs[9257]) ^ (layer0_outputs[7926]));
    assign outputs[753] = (layer0_outputs[3783]) ^ (layer0_outputs[2098]);
    assign outputs[754] = layer0_outputs[8245];
    assign outputs[755] = ~(layer0_outputs[3419]);
    assign outputs[756] = ~(layer0_outputs[9388]);
    assign outputs[757] = ~(layer0_outputs[8228]) | (layer0_outputs[9038]);
    assign outputs[758] = ~(layer0_outputs[6974]);
    assign outputs[759] = ~((layer0_outputs[3816]) ^ (layer0_outputs[7607]));
    assign outputs[760] = (layer0_outputs[1078]) ^ (layer0_outputs[2412]);
    assign outputs[761] = layer0_outputs[5247];
    assign outputs[762] = ~(layer0_outputs[2407]);
    assign outputs[763] = ~(layer0_outputs[3962]);
    assign outputs[764] = ~((layer0_outputs[1061]) ^ (layer0_outputs[7615]));
    assign outputs[765] = ~(layer0_outputs[7693]);
    assign outputs[766] = layer0_outputs[8517];
    assign outputs[767] = ~(layer0_outputs[1242]);
    assign outputs[768] = (layer0_outputs[2518]) | (layer0_outputs[1477]);
    assign outputs[769] = ~((layer0_outputs[2835]) ^ (layer0_outputs[8713]));
    assign outputs[770] = ~(layer0_outputs[5676]);
    assign outputs[771] = (layer0_outputs[3126]) & ~(layer0_outputs[8269]);
    assign outputs[772] = ~(layer0_outputs[1386]);
    assign outputs[773] = ~((layer0_outputs[2506]) ^ (layer0_outputs[728]));
    assign outputs[774] = (layer0_outputs[8987]) | (layer0_outputs[6781]);
    assign outputs[775] = (layer0_outputs[3131]) | (layer0_outputs[920]);
    assign outputs[776] = ~(layer0_outputs[7930]);
    assign outputs[777] = ~((layer0_outputs[5108]) ^ (layer0_outputs[811]));
    assign outputs[778] = ~(layer0_outputs[4785]);
    assign outputs[779] = layer0_outputs[6234];
    assign outputs[780] = (layer0_outputs[1760]) ^ (layer0_outputs[9244]);
    assign outputs[781] = ~((layer0_outputs[10074]) & (layer0_outputs[685]));
    assign outputs[782] = layer0_outputs[8517];
    assign outputs[783] = ~(layer0_outputs[8338]);
    assign outputs[784] = ~((layer0_outputs[5604]) & (layer0_outputs[7462]));
    assign outputs[785] = layer0_outputs[9497];
    assign outputs[786] = ~(layer0_outputs[9601]);
    assign outputs[787] = ~(layer0_outputs[2332]);
    assign outputs[788] = 1'b1;
    assign outputs[789] = ~((layer0_outputs[9790]) & (layer0_outputs[3905]));
    assign outputs[790] = ~(layer0_outputs[7173]);
    assign outputs[791] = layer0_outputs[667];
    assign outputs[792] = (layer0_outputs[2604]) | (layer0_outputs[4933]);
    assign outputs[793] = 1'b0;
    assign outputs[794] = ~((layer0_outputs[9543]) | (layer0_outputs[3169]));
    assign outputs[795] = ~((layer0_outputs[8251]) ^ (layer0_outputs[6728]));
    assign outputs[796] = (layer0_outputs[5693]) ^ (layer0_outputs[7213]);
    assign outputs[797] = (layer0_outputs[7083]) ^ (layer0_outputs[4402]);
    assign outputs[798] = ~(layer0_outputs[4234]);
    assign outputs[799] = ~(layer0_outputs[5720]);
    assign outputs[800] = ~((layer0_outputs[2606]) | (layer0_outputs[9300]));
    assign outputs[801] = layer0_outputs[7488];
    assign outputs[802] = ~(layer0_outputs[9712]) | (layer0_outputs[1549]);
    assign outputs[803] = layer0_outputs[5461];
    assign outputs[804] = (layer0_outputs[8114]) ^ (layer0_outputs[7790]);
    assign outputs[805] = (layer0_outputs[5127]) | (layer0_outputs[6169]);
    assign outputs[806] = ~(layer0_outputs[67]);
    assign outputs[807] = ~(layer0_outputs[8941]);
    assign outputs[808] = layer0_outputs[9456];
    assign outputs[809] = ~(layer0_outputs[2245]) | (layer0_outputs[7721]);
    assign outputs[810] = ~(layer0_outputs[2915]);
    assign outputs[811] = layer0_outputs[3313];
    assign outputs[812] = layer0_outputs[3713];
    assign outputs[813] = ~(layer0_outputs[1703]);
    assign outputs[814] = ~(layer0_outputs[4480]);
    assign outputs[815] = ~(layer0_outputs[3976]);
    assign outputs[816] = (layer0_outputs[9741]) & (layer0_outputs[350]);
    assign outputs[817] = (layer0_outputs[499]) ^ (layer0_outputs[6449]);
    assign outputs[818] = (layer0_outputs[8786]) & ~(layer0_outputs[2261]);
    assign outputs[819] = ~((layer0_outputs[5626]) | (layer0_outputs[8075]));
    assign outputs[820] = ~((layer0_outputs[9958]) ^ (layer0_outputs[6995]));
    assign outputs[821] = layer0_outputs[174];
    assign outputs[822] = ~((layer0_outputs[10018]) ^ (layer0_outputs[3565]));
    assign outputs[823] = ~(layer0_outputs[9911]) | (layer0_outputs[2778]);
    assign outputs[824] = ~((layer0_outputs[8527]) ^ (layer0_outputs[2794]));
    assign outputs[825] = layer0_outputs[3839];
    assign outputs[826] = (layer0_outputs[10055]) | (layer0_outputs[9634]);
    assign outputs[827] = ~(layer0_outputs[9192]);
    assign outputs[828] = ~((layer0_outputs[2776]) ^ (layer0_outputs[5481]));
    assign outputs[829] = layer0_outputs[9427];
    assign outputs[830] = ~((layer0_outputs[6209]) ^ (layer0_outputs[6955]));
    assign outputs[831] = layer0_outputs[2154];
    assign outputs[832] = layer0_outputs[3847];
    assign outputs[833] = (layer0_outputs[5858]) ^ (layer0_outputs[194]);
    assign outputs[834] = (layer0_outputs[1745]) | (layer0_outputs[3387]);
    assign outputs[835] = (layer0_outputs[1880]) ^ (layer0_outputs[5366]);
    assign outputs[836] = ~((layer0_outputs[4601]) | (layer0_outputs[994]));
    assign outputs[837] = ~(layer0_outputs[7557]);
    assign outputs[838] = ~(layer0_outputs[9055]);
    assign outputs[839] = ~((layer0_outputs[4080]) ^ (layer0_outputs[2086]));
    assign outputs[840] = ~((layer0_outputs[9708]) ^ (layer0_outputs[2378]));
    assign outputs[841] = ~(layer0_outputs[2459]);
    assign outputs[842] = layer0_outputs[3841];
    assign outputs[843] = ~(layer0_outputs[916]) | (layer0_outputs[2826]);
    assign outputs[844] = (layer0_outputs[4546]) ^ (layer0_outputs[3061]);
    assign outputs[845] = layer0_outputs[1836];
    assign outputs[846] = ~((layer0_outputs[9022]) & (layer0_outputs[1076]));
    assign outputs[847] = ~(layer0_outputs[7762]);
    assign outputs[848] = layer0_outputs[666];
    assign outputs[849] = ~(layer0_outputs[9155]);
    assign outputs[850] = layer0_outputs[3298];
    assign outputs[851] = ~((layer0_outputs[2447]) ^ (layer0_outputs[6606]));
    assign outputs[852] = layer0_outputs[8140];
    assign outputs[853] = layer0_outputs[1660];
    assign outputs[854] = (layer0_outputs[5299]) ^ (layer0_outputs[4789]);
    assign outputs[855] = ~((layer0_outputs[4902]) ^ (layer0_outputs[6813]));
    assign outputs[856] = (layer0_outputs[5706]) & ~(layer0_outputs[10183]);
    assign outputs[857] = ~(layer0_outputs[1659]);
    assign outputs[858] = ~(layer0_outputs[5676]);
    assign outputs[859] = ~(layer0_outputs[237]) | (layer0_outputs[7824]);
    assign outputs[860] = ~(layer0_outputs[5390]);
    assign outputs[861] = ~(layer0_outputs[5049]);
    assign outputs[862] = ~((layer0_outputs[2888]) ^ (layer0_outputs[4550]));
    assign outputs[863] = layer0_outputs[8699];
    assign outputs[864] = ~(layer0_outputs[7415]) | (layer0_outputs[5236]);
    assign outputs[865] = ~(layer0_outputs[3107]) | (layer0_outputs[5263]);
    assign outputs[866] = ~(layer0_outputs[3295]) | (layer0_outputs[1651]);
    assign outputs[867] = (layer0_outputs[1732]) ^ (layer0_outputs[6213]);
    assign outputs[868] = ~(layer0_outputs[8046]);
    assign outputs[869] = (layer0_outputs[762]) | (layer0_outputs[4311]);
    assign outputs[870] = ~(layer0_outputs[2300]);
    assign outputs[871] = layer0_outputs[6228];
    assign outputs[872] = 1'b1;
    assign outputs[873] = (layer0_outputs[106]) & (layer0_outputs[6666]);
    assign outputs[874] = layer0_outputs[5643];
    assign outputs[875] = (layer0_outputs[2416]) & (layer0_outputs[3766]);
    assign outputs[876] = (layer0_outputs[2799]) & ~(layer0_outputs[1791]);
    assign outputs[877] = (layer0_outputs[6480]) | (layer0_outputs[2360]);
    assign outputs[878] = (layer0_outputs[4652]) ^ (layer0_outputs[9930]);
    assign outputs[879] = ~(layer0_outputs[4347]);
    assign outputs[880] = ~(layer0_outputs[4057]) | (layer0_outputs[511]);
    assign outputs[881] = ~(layer0_outputs[2332]);
    assign outputs[882] = ~(layer0_outputs[8368]);
    assign outputs[883] = ~((layer0_outputs[6756]) ^ (layer0_outputs[10048]));
    assign outputs[884] = layer0_outputs[7382];
    assign outputs[885] = ~((layer0_outputs[1614]) ^ (layer0_outputs[9474]));
    assign outputs[886] = (layer0_outputs[5766]) & ~(layer0_outputs[4599]);
    assign outputs[887] = layer0_outputs[1303];
    assign outputs[888] = (layer0_outputs[7361]) & ~(layer0_outputs[9672]);
    assign outputs[889] = ~(layer0_outputs[3676]);
    assign outputs[890] = ~(layer0_outputs[9653]);
    assign outputs[891] = layer0_outputs[1104];
    assign outputs[892] = (layer0_outputs[1272]) & ~(layer0_outputs[1373]);
    assign outputs[893] = ~(layer0_outputs[6364]) | (layer0_outputs[150]);
    assign outputs[894] = (layer0_outputs[1442]) | (layer0_outputs[8196]);
    assign outputs[895] = ~(layer0_outputs[7233]) | (layer0_outputs[7498]);
    assign outputs[896] = ~(layer0_outputs[5497]);
    assign outputs[897] = ~(layer0_outputs[1032]);
    assign outputs[898] = layer0_outputs[8805];
    assign outputs[899] = ~(layer0_outputs[5610]);
    assign outputs[900] = ~((layer0_outputs[6342]) & (layer0_outputs[4682]));
    assign outputs[901] = layer0_outputs[4319];
    assign outputs[902] = (layer0_outputs[7698]) & (layer0_outputs[10200]);
    assign outputs[903] = layer0_outputs[8259];
    assign outputs[904] = ~(layer0_outputs[4395]);
    assign outputs[905] = (layer0_outputs[3506]) ^ (layer0_outputs[9081]);
    assign outputs[906] = ~(layer0_outputs[7408]);
    assign outputs[907] = (layer0_outputs[6944]) | (layer0_outputs[10135]);
    assign outputs[908] = ~(layer0_outputs[7419]) | (layer0_outputs[4506]);
    assign outputs[909] = ~(layer0_outputs[8106]) | (layer0_outputs[3500]);
    assign outputs[910] = ~((layer0_outputs[10110]) & (layer0_outputs[8223]));
    assign outputs[911] = ~((layer0_outputs[6424]) ^ (layer0_outputs[1977]));
    assign outputs[912] = ~(layer0_outputs[8956]);
    assign outputs[913] = ~(layer0_outputs[396]);
    assign outputs[914] = layer0_outputs[1233];
    assign outputs[915] = layer0_outputs[6573];
    assign outputs[916] = ~(layer0_outputs[10048]);
    assign outputs[917] = ~(layer0_outputs[8324]) | (layer0_outputs[5556]);
    assign outputs[918] = ~(layer0_outputs[3194]);
    assign outputs[919] = ~(layer0_outputs[5781]);
    assign outputs[920] = (layer0_outputs[9068]) & (layer0_outputs[4258]);
    assign outputs[921] = layer0_outputs[3882];
    assign outputs[922] = layer0_outputs[1704];
    assign outputs[923] = ~(layer0_outputs[7810]);
    assign outputs[924] = layer0_outputs[8569];
    assign outputs[925] = ~(layer0_outputs[5962]);
    assign outputs[926] = ~(layer0_outputs[4764]);
    assign outputs[927] = ~(layer0_outputs[562]);
    assign outputs[928] = ~(layer0_outputs[5494]) | (layer0_outputs[2510]);
    assign outputs[929] = (layer0_outputs[2524]) ^ (layer0_outputs[8702]);
    assign outputs[930] = ~(layer0_outputs[9448]);
    assign outputs[931] = layer0_outputs[5362];
    assign outputs[932] = ~(layer0_outputs[6782]) | (layer0_outputs[5136]);
    assign outputs[933] = ~((layer0_outputs[5181]) & (layer0_outputs[5956]));
    assign outputs[934] = layer0_outputs[7943];
    assign outputs[935] = ~(layer0_outputs[9391]) | (layer0_outputs[3572]);
    assign outputs[936] = ~(layer0_outputs[4977]);
    assign outputs[937] = ~(layer0_outputs[3235]);
    assign outputs[938] = (layer0_outputs[10181]) ^ (layer0_outputs[3596]);
    assign outputs[939] = layer0_outputs[2158];
    assign outputs[940] = layer0_outputs[1722];
    assign outputs[941] = ~(layer0_outputs[6730]);
    assign outputs[942] = ~(layer0_outputs[7161]);
    assign outputs[943] = ~(layer0_outputs[1821]);
    assign outputs[944] = ~((layer0_outputs[2008]) ^ (layer0_outputs[6005]));
    assign outputs[945] = (layer0_outputs[8513]) & ~(layer0_outputs[1765]);
    assign outputs[946] = ~(layer0_outputs[7578]) | (layer0_outputs[3229]);
    assign outputs[947] = layer0_outputs[3617];
    assign outputs[948] = ~((layer0_outputs[992]) ^ (layer0_outputs[1293]));
    assign outputs[949] = ~((layer0_outputs[764]) ^ (layer0_outputs[2109]));
    assign outputs[950] = ~((layer0_outputs[4223]) & (layer0_outputs[9578]));
    assign outputs[951] = layer0_outputs[2489];
    assign outputs[952] = layer0_outputs[5914];
    assign outputs[953] = (layer0_outputs[7742]) & ~(layer0_outputs[10032]);
    assign outputs[954] = ~((layer0_outputs[6265]) | (layer0_outputs[3625]));
    assign outputs[955] = ~((layer0_outputs[9241]) | (layer0_outputs[2273]));
    assign outputs[956] = layer0_outputs[8556];
    assign outputs[957] = (layer0_outputs[9475]) ^ (layer0_outputs[2220]);
    assign outputs[958] = ~(layer0_outputs[4619]);
    assign outputs[959] = layer0_outputs[8985];
    assign outputs[960] = ~(layer0_outputs[8522]);
    assign outputs[961] = ~((layer0_outputs[4638]) | (layer0_outputs[9258]));
    assign outputs[962] = (layer0_outputs[4035]) & ~(layer0_outputs[8829]);
    assign outputs[963] = (layer0_outputs[1767]) ^ (layer0_outputs[10050]);
    assign outputs[964] = ~(layer0_outputs[268]);
    assign outputs[965] = 1'b1;
    assign outputs[966] = ~(layer0_outputs[9046]);
    assign outputs[967] = layer0_outputs[1509];
    assign outputs[968] = (layer0_outputs[10142]) ^ (layer0_outputs[4448]);
    assign outputs[969] = ~((layer0_outputs[10209]) ^ (layer0_outputs[8131]));
    assign outputs[970] = ~((layer0_outputs[5268]) | (layer0_outputs[968]));
    assign outputs[971] = (layer0_outputs[9181]) ^ (layer0_outputs[5322]);
    assign outputs[972] = layer0_outputs[8501];
    assign outputs[973] = layer0_outputs[2814];
    assign outputs[974] = ~((layer0_outputs[8647]) ^ (layer0_outputs[4027]));
    assign outputs[975] = layer0_outputs[4970];
    assign outputs[976] = layer0_outputs[5931];
    assign outputs[977] = 1'b1;
    assign outputs[978] = ~(layer0_outputs[5002]);
    assign outputs[979] = ~((layer0_outputs[3785]) ^ (layer0_outputs[1356]));
    assign outputs[980] = layer0_outputs[6688];
    assign outputs[981] = (layer0_outputs[840]) | (layer0_outputs[1370]);
    assign outputs[982] = ~(layer0_outputs[3970]);
    assign outputs[983] = ~(layer0_outputs[6591]);
    assign outputs[984] = ~((layer0_outputs[1675]) & (layer0_outputs[4452]));
    assign outputs[985] = ~(layer0_outputs[9851]) | (layer0_outputs[9409]);
    assign outputs[986] = ~(layer0_outputs[3302]);
    assign outputs[987] = ~(layer0_outputs[7844]);
    assign outputs[988] = ~(layer0_outputs[1916]);
    assign outputs[989] = ~(layer0_outputs[4985]);
    assign outputs[990] = ~((layer0_outputs[2281]) ^ (layer0_outputs[3401]));
    assign outputs[991] = (layer0_outputs[1657]) | (layer0_outputs[9583]);
    assign outputs[992] = ~((layer0_outputs[2548]) ^ (layer0_outputs[4138]));
    assign outputs[993] = layer0_outputs[3498];
    assign outputs[994] = layer0_outputs[3504];
    assign outputs[995] = ~((layer0_outputs[5496]) & (layer0_outputs[2002]));
    assign outputs[996] = ~(layer0_outputs[4603]) | (layer0_outputs[2278]);
    assign outputs[997] = ~((layer0_outputs[3992]) ^ (layer0_outputs[5950]));
    assign outputs[998] = ~((layer0_outputs[5273]) | (layer0_outputs[5387]));
    assign outputs[999] = ~(layer0_outputs[690]);
    assign outputs[1000] = ~(layer0_outputs[6770]);
    assign outputs[1001] = ~(layer0_outputs[1610]);
    assign outputs[1002] = layer0_outputs[3671];
    assign outputs[1003] = ~((layer0_outputs[8274]) ^ (layer0_outputs[4842]));
    assign outputs[1004] = layer0_outputs[1871];
    assign outputs[1005] = 1'b1;
    assign outputs[1006] = (layer0_outputs[2527]) & ~(layer0_outputs[3222]);
    assign outputs[1007] = ~(layer0_outputs[940]);
    assign outputs[1008] = (layer0_outputs[2741]) & (layer0_outputs[7689]);
    assign outputs[1009] = ~(layer0_outputs[5302]) | (layer0_outputs[6561]);
    assign outputs[1010] = ~(layer0_outputs[1463]) | (layer0_outputs[3212]);
    assign outputs[1011] = ~((layer0_outputs[7612]) | (layer0_outputs[8644]));
    assign outputs[1012] = ~((layer0_outputs[6124]) ^ (layer0_outputs[3481]));
    assign outputs[1013] = (layer0_outputs[5062]) ^ (layer0_outputs[2117]);
    assign outputs[1014] = layer0_outputs[9027];
    assign outputs[1015] = layer0_outputs[1313];
    assign outputs[1016] = ~(layer0_outputs[822]);
    assign outputs[1017] = (layer0_outputs[1693]) & ~(layer0_outputs[2971]);
    assign outputs[1018] = layer0_outputs[8738];
    assign outputs[1019] = ~(layer0_outputs[3099]);
    assign outputs[1020] = layer0_outputs[6200];
    assign outputs[1021] = ~((layer0_outputs[3326]) | (layer0_outputs[8979]));
    assign outputs[1022] = (layer0_outputs[9120]) ^ (layer0_outputs[7940]);
    assign outputs[1023] = ~(layer0_outputs[1523]) | (layer0_outputs[7576]);
    assign outputs[1024] = ~((layer0_outputs[1844]) ^ (layer0_outputs[2167]));
    assign outputs[1025] = (layer0_outputs[3898]) & ~(layer0_outputs[3190]);
    assign outputs[1026] = ~(layer0_outputs[454]);
    assign outputs[1027] = (layer0_outputs[4840]) & ~(layer0_outputs[4197]);
    assign outputs[1028] = (layer0_outputs[847]) & ~(layer0_outputs[6913]);
    assign outputs[1029] = ~(layer0_outputs[899]);
    assign outputs[1030] = (layer0_outputs[3126]) ^ (layer0_outputs[8849]);
    assign outputs[1031] = ~(layer0_outputs[5601]);
    assign outputs[1032] = (layer0_outputs[975]) ^ (layer0_outputs[3240]);
    assign outputs[1033] = ~(layer0_outputs[4548]);
    assign outputs[1034] = (layer0_outputs[5568]) ^ (layer0_outputs[4936]);
    assign outputs[1035] = (layer0_outputs[3216]) & ~(layer0_outputs[8680]);
    assign outputs[1036] = ~(layer0_outputs[3593]);
    assign outputs[1037] = (layer0_outputs[9981]) & ~(layer0_outputs[288]);
    assign outputs[1038] = (layer0_outputs[388]) & ~(layer0_outputs[9605]);
    assign outputs[1039] = (layer0_outputs[6860]) ^ (layer0_outputs[8859]);
    assign outputs[1040] = layer0_outputs[8757];
    assign outputs[1041] = (layer0_outputs[4598]) & ~(layer0_outputs[7170]);
    assign outputs[1042] = (layer0_outputs[10190]) & ~(layer0_outputs[3748]);
    assign outputs[1043] = (layer0_outputs[5140]) & ~(layer0_outputs[75]);
    assign outputs[1044] = ~(layer0_outputs[6718]);
    assign outputs[1045] = (layer0_outputs[10042]) ^ (layer0_outputs[7511]);
    assign outputs[1046] = ~(layer0_outputs[7670]);
    assign outputs[1047] = (layer0_outputs[3964]) & ~(layer0_outputs[9084]);
    assign outputs[1048] = (layer0_outputs[7389]) & ~(layer0_outputs[2080]);
    assign outputs[1049] = ~((layer0_outputs[5937]) | (layer0_outputs[2148]));
    assign outputs[1050] = layer0_outputs[9040];
    assign outputs[1051] = ~(layer0_outputs[9902]);
    assign outputs[1052] = layer0_outputs[4928];
    assign outputs[1053] = layer0_outputs[8520];
    assign outputs[1054] = (layer0_outputs[934]) & ~(layer0_outputs[6406]);
    assign outputs[1055] = ~(layer0_outputs[1917]);
    assign outputs[1056] = ~((layer0_outputs[9156]) ^ (layer0_outputs[9825]));
    assign outputs[1057] = ~(layer0_outputs[6426]);
    assign outputs[1058] = (layer0_outputs[2104]) & ~(layer0_outputs[5548]);
    assign outputs[1059] = (layer0_outputs[1064]) & ~(layer0_outputs[5352]);
    assign outputs[1060] = ~(layer0_outputs[1231]);
    assign outputs[1061] = ~(layer0_outputs[4804]);
    assign outputs[1062] = ~((layer0_outputs[9212]) | (layer0_outputs[2742]));
    assign outputs[1063] = ~((layer0_outputs[4226]) | (layer0_outputs[8184]));
    assign outputs[1064] = (layer0_outputs[8077]) & (layer0_outputs[10076]);
    assign outputs[1065] = ~((layer0_outputs[10171]) ^ (layer0_outputs[6401]));
    assign outputs[1066] = (layer0_outputs[5232]) ^ (layer0_outputs[482]);
    assign outputs[1067] = 1'b0;
    assign outputs[1068] = ~((layer0_outputs[348]) | (layer0_outputs[6548]));
    assign outputs[1069] = (layer0_outputs[3291]) & ~(layer0_outputs[4733]);
    assign outputs[1070] = ~((layer0_outputs[1]) | (layer0_outputs[4260]));
    assign outputs[1071] = layer0_outputs[9504];
    assign outputs[1072] = ~((layer0_outputs[3071]) | (layer0_outputs[8677]));
    assign outputs[1073] = (layer0_outputs[1554]) ^ (layer0_outputs[6379]);
    assign outputs[1074] = (layer0_outputs[9262]) & ~(layer0_outputs[4325]);
    assign outputs[1075] = ~(layer0_outputs[9459]);
    assign outputs[1076] = (layer0_outputs[10230]) & ~(layer0_outputs[1233]);
    assign outputs[1077] = (layer0_outputs[533]) & ~(layer0_outputs[8497]);
    assign outputs[1078] = (layer0_outputs[10172]) ^ (layer0_outputs[7153]);
    assign outputs[1079] = (layer0_outputs[3806]) & (layer0_outputs[1484]);
    assign outputs[1080] = (layer0_outputs[8439]) & ~(layer0_outputs[5161]);
    assign outputs[1081] = (layer0_outputs[8326]) & ~(layer0_outputs[5193]);
    assign outputs[1082] = (layer0_outputs[5812]) & ~(layer0_outputs[9261]);
    assign outputs[1083] = ~((layer0_outputs[3364]) | (layer0_outputs[8248]));
    assign outputs[1084] = layer0_outputs[478];
    assign outputs[1085] = ~(layer0_outputs[6880]);
    assign outputs[1086] = 1'b0;
    assign outputs[1087] = (layer0_outputs[5215]) & ~(layer0_outputs[4342]);
    assign outputs[1088] = layer0_outputs[1194];
    assign outputs[1089] = (layer0_outputs[0]) & ~(layer0_outputs[3750]);
    assign outputs[1090] = ~((layer0_outputs[5867]) ^ (layer0_outputs[4895]));
    assign outputs[1091] = (layer0_outputs[2251]) & ~(layer0_outputs[7917]);
    assign outputs[1092] = ~(layer0_outputs[9974]);
    assign outputs[1093] = ~((layer0_outputs[9569]) | (layer0_outputs[2116]));
    assign outputs[1094] = ~((layer0_outputs[380]) | (layer0_outputs[5096]));
    assign outputs[1095] = ~((layer0_outputs[5926]) & (layer0_outputs[5375]));
    assign outputs[1096] = ~((layer0_outputs[7965]) | (layer0_outputs[7140]));
    assign outputs[1097] = (layer0_outputs[9206]) & (layer0_outputs[7838]);
    assign outputs[1098] = (layer0_outputs[4721]) & ~(layer0_outputs[1767]);
    assign outputs[1099] = (layer0_outputs[742]) & ~(layer0_outputs[4688]);
    assign outputs[1100] = ~(layer0_outputs[5189]);
    assign outputs[1101] = layer0_outputs[3808];
    assign outputs[1102] = (layer0_outputs[1315]) ^ (layer0_outputs[6037]);
    assign outputs[1103] = (layer0_outputs[7038]) & (layer0_outputs[3653]);
    assign outputs[1104] = (layer0_outputs[4028]) & ~(layer0_outputs[3394]);
    assign outputs[1105] = (layer0_outputs[1226]) ^ (layer0_outputs[6930]);
    assign outputs[1106] = ~(layer0_outputs[9807]);
    assign outputs[1107] = ~(layer0_outputs[7652]);
    assign outputs[1108] = 1'b0;
    assign outputs[1109] = layer0_outputs[6267];
    assign outputs[1110] = (layer0_outputs[5533]) & ~(layer0_outputs[7518]);
    assign outputs[1111] = ~(layer0_outputs[1162]) | (layer0_outputs[183]);
    assign outputs[1112] = ~(layer0_outputs[3036]) | (layer0_outputs[5589]);
    assign outputs[1113] = (layer0_outputs[5262]) & ~(layer0_outputs[8683]);
    assign outputs[1114] = (layer0_outputs[5816]) & ~(layer0_outputs[4501]);
    assign outputs[1115] = layer0_outputs[9571];
    assign outputs[1116] = layer0_outputs[6090];
    assign outputs[1117] = (layer0_outputs[5215]) & (layer0_outputs[8593]);
    assign outputs[1118] = layer0_outputs[8866];
    assign outputs[1119] = layer0_outputs[2539];
    assign outputs[1120] = (layer0_outputs[2455]) & ~(layer0_outputs[7198]);
    assign outputs[1121] = layer0_outputs[4592];
    assign outputs[1122] = (layer0_outputs[533]) & ~(layer0_outputs[2044]);
    assign outputs[1123] = (layer0_outputs[9065]) & ~(layer0_outputs[6572]);
    assign outputs[1124] = layer0_outputs[2411];
    assign outputs[1125] = ~((layer0_outputs[5729]) ^ (layer0_outputs[6103]));
    assign outputs[1126] = (layer0_outputs[807]) ^ (layer0_outputs[8229]);
    assign outputs[1127] = layer0_outputs[6783];
    assign outputs[1128] = ~(layer0_outputs[1979]);
    assign outputs[1129] = (layer0_outputs[8283]) ^ (layer0_outputs[9386]);
    assign outputs[1130] = ~(layer0_outputs[7512]) | (layer0_outputs[2849]);
    assign outputs[1131] = ~(layer0_outputs[8123]);
    assign outputs[1132] = ~((layer0_outputs[737]) ^ (layer0_outputs[6293]));
    assign outputs[1133] = ~((layer0_outputs[314]) ^ (layer0_outputs[5754]));
    assign outputs[1134] = ~((layer0_outputs[513]) ^ (layer0_outputs[3371]));
    assign outputs[1135] = (layer0_outputs[5308]) & ~(layer0_outputs[7665]);
    assign outputs[1136] = (layer0_outputs[2763]) & (layer0_outputs[2943]);
    assign outputs[1137] = (layer0_outputs[9125]) ^ (layer0_outputs[7916]);
    assign outputs[1138] = ~((layer0_outputs[2276]) | (layer0_outputs[3948]));
    assign outputs[1139] = ~((layer0_outputs[9473]) ^ (layer0_outputs[7837]));
    assign outputs[1140] = ~((layer0_outputs[2587]) | (layer0_outputs[8033]));
    assign outputs[1141] = 1'b0;
    assign outputs[1142] = ~(layer0_outputs[886]);
    assign outputs[1143] = layer0_outputs[4000];
    assign outputs[1144] = layer0_outputs[3868];
    assign outputs[1145] = (layer0_outputs[9958]) & (layer0_outputs[809]);
    assign outputs[1146] = (layer0_outputs[7391]) & ~(layer0_outputs[5654]);
    assign outputs[1147] = ~((layer0_outputs[4971]) ^ (layer0_outputs[8567]));
    assign outputs[1148] = (layer0_outputs[9813]) & ~(layer0_outputs[4604]);
    assign outputs[1149] = (layer0_outputs[5958]) & ~(layer0_outputs[1640]);
    assign outputs[1150] = ~((layer0_outputs[7875]) | (layer0_outputs[622]));
    assign outputs[1151] = 1'b0;
    assign outputs[1152] = ~((layer0_outputs[9304]) | (layer0_outputs[7194]));
    assign outputs[1153] = (layer0_outputs[664]) ^ (layer0_outputs[8766]);
    assign outputs[1154] = ~(layer0_outputs[9999]);
    assign outputs[1155] = (layer0_outputs[8516]) & (layer0_outputs[3606]);
    assign outputs[1156] = (layer0_outputs[2541]) ^ (layer0_outputs[10008]);
    assign outputs[1157] = (layer0_outputs[8013]) & ~(layer0_outputs[5947]);
    assign outputs[1158] = (layer0_outputs[2519]) ^ (layer0_outputs[5351]);
    assign outputs[1159] = (layer0_outputs[1911]) & (layer0_outputs[1403]);
    assign outputs[1160] = layer0_outputs[103];
    assign outputs[1161] = layer0_outputs[7520];
    assign outputs[1162] = ~(layer0_outputs[8328]);
    assign outputs[1163] = ~((layer0_outputs[446]) ^ (layer0_outputs[98]));
    assign outputs[1164] = (layer0_outputs[2359]) ^ (layer0_outputs[2302]);
    assign outputs[1165] = ~((layer0_outputs[4174]) ^ (layer0_outputs[4173]));
    assign outputs[1166] = (layer0_outputs[6041]) ^ (layer0_outputs[2487]);
    assign outputs[1167] = (layer0_outputs[3184]) ^ (layer0_outputs[3188]);
    assign outputs[1168] = (layer0_outputs[1541]) ^ (layer0_outputs[1441]);
    assign outputs[1169] = (layer0_outputs[6587]) & (layer0_outputs[9978]);
    assign outputs[1170] = (layer0_outputs[8767]) ^ (layer0_outputs[9913]);
    assign outputs[1171] = layer0_outputs[5661];
    assign outputs[1172] = ~(layer0_outputs[883]);
    assign outputs[1173] = ~((layer0_outputs[5331]) | (layer0_outputs[2904]));
    assign outputs[1174] = layer0_outputs[6677];
    assign outputs[1175] = ~((layer0_outputs[2675]) | (layer0_outputs[2780]));
    assign outputs[1176] = (layer0_outputs[368]) & (layer0_outputs[4240]);
    assign outputs[1177] = (layer0_outputs[6663]) & (layer0_outputs[2462]);
    assign outputs[1178] = (layer0_outputs[7548]) | (layer0_outputs[3077]);
    assign outputs[1179] = (layer0_outputs[6991]) & ~(layer0_outputs[1646]);
    assign outputs[1180] = (layer0_outputs[9715]) & ~(layer0_outputs[9004]);
    assign outputs[1181] = layer0_outputs[1586];
    assign outputs[1182] = ~(layer0_outputs[4351]);
    assign outputs[1183] = (layer0_outputs[6267]) & (layer0_outputs[6468]);
    assign outputs[1184] = ~(layer0_outputs[7486]) | (layer0_outputs[9757]);
    assign outputs[1185] = (layer0_outputs[5395]) & (layer0_outputs[7041]);
    assign outputs[1186] = layer0_outputs[6689];
    assign outputs[1187] = (layer0_outputs[8401]) & ~(layer0_outputs[7757]);
    assign outputs[1188] = layer0_outputs[9661];
    assign outputs[1189] = (layer0_outputs[1799]) & (layer0_outputs[274]);
    assign outputs[1190] = 1'b0;
    assign outputs[1191] = ~((layer0_outputs[1853]) ^ (layer0_outputs[1319]));
    assign outputs[1192] = ~(layer0_outputs[7084]);
    assign outputs[1193] = ~(layer0_outputs[5838]) | (layer0_outputs[230]);
    assign outputs[1194] = (layer0_outputs[8144]) & ~(layer0_outputs[8265]);
    assign outputs[1195] = ~(layer0_outputs[1155]);
    assign outputs[1196] = 1'b0;
    assign outputs[1197] = layer0_outputs[9547];
    assign outputs[1198] = ~(layer0_outputs[8466]);
    assign outputs[1199] = ~(layer0_outputs[10065]);
    assign outputs[1200] = ~(layer0_outputs[8846]);
    assign outputs[1201] = ~(layer0_outputs[3568]);
    assign outputs[1202] = ~((layer0_outputs[860]) ^ (layer0_outputs[3908]));
    assign outputs[1203] = ~((layer0_outputs[3854]) | (layer0_outputs[8884]));
    assign outputs[1204] = (layer0_outputs[6199]) | (layer0_outputs[3626]);
    assign outputs[1205] = layer0_outputs[4460];
    assign outputs[1206] = (layer0_outputs[4257]) ^ (layer0_outputs[564]);
    assign outputs[1207] = (layer0_outputs[7818]) & (layer0_outputs[9868]);
    assign outputs[1208] = 1'b0;
    assign outputs[1209] = (layer0_outputs[9184]) & ~(layer0_outputs[3764]);
    assign outputs[1210] = ~(layer0_outputs[3389]);
    assign outputs[1211] = ~((layer0_outputs[10171]) | (layer0_outputs[1228]));
    assign outputs[1212] = ~((layer0_outputs[1812]) ^ (layer0_outputs[4772]));
    assign outputs[1213] = 1'b0;
    assign outputs[1214] = (layer0_outputs[4137]) & (layer0_outputs[2043]);
    assign outputs[1215] = (layer0_outputs[10191]) & ~(layer0_outputs[5619]);
    assign outputs[1216] = ~(layer0_outputs[7826]);
    assign outputs[1217] = (layer0_outputs[9379]) ^ (layer0_outputs[7927]);
    assign outputs[1218] = layer0_outputs[4203];
    assign outputs[1219] = layer0_outputs[1287];
    assign outputs[1220] = ~((layer0_outputs[909]) | (layer0_outputs[4907]));
    assign outputs[1221] = (layer0_outputs[5402]) & ~(layer0_outputs[7012]);
    assign outputs[1222] = (layer0_outputs[2018]) ^ (layer0_outputs[5037]);
    assign outputs[1223] = ~((layer0_outputs[1709]) ^ (layer0_outputs[4713]));
    assign outputs[1224] = (layer0_outputs[3688]) ^ (layer0_outputs[996]);
    assign outputs[1225] = (layer0_outputs[3353]) & ~(layer0_outputs[3551]);
    assign outputs[1226] = layer0_outputs[5205];
    assign outputs[1227] = ~(layer0_outputs[9487]);
    assign outputs[1228] = 1'b0;
    assign outputs[1229] = ~((layer0_outputs[4660]) | (layer0_outputs[6013]));
    assign outputs[1230] = ~((layer0_outputs[4085]) ^ (layer0_outputs[2776]));
    assign outputs[1231] = (layer0_outputs[1788]) ^ (layer0_outputs[596]);
    assign outputs[1232] = ~((layer0_outputs[251]) | (layer0_outputs[4697]));
    assign outputs[1233] = (layer0_outputs[1742]) ^ (layer0_outputs[951]);
    assign outputs[1234] = 1'b0;
    assign outputs[1235] = (layer0_outputs[7210]) & ~(layer0_outputs[6047]);
    assign outputs[1236] = ~((layer0_outputs[3112]) ^ (layer0_outputs[181]));
    assign outputs[1237] = ~((layer0_outputs[2059]) ^ (layer0_outputs[5055]));
    assign outputs[1238] = ~((layer0_outputs[6082]) | (layer0_outputs[2179]));
    assign outputs[1239] = ~(layer0_outputs[7397]);
    assign outputs[1240] = ~((layer0_outputs[4384]) ^ (layer0_outputs[3074]));
    assign outputs[1241] = (layer0_outputs[5965]) | (layer0_outputs[1827]);
    assign outputs[1242] = (layer0_outputs[1700]) & ~(layer0_outputs[5096]);
    assign outputs[1243] = layer0_outputs[8478];
    assign outputs[1244] = layer0_outputs[4099];
    assign outputs[1245] = ~(layer0_outputs[9167]);
    assign outputs[1246] = layer0_outputs[4966];
    assign outputs[1247] = ~((layer0_outputs[8585]) | (layer0_outputs[9137]));
    assign outputs[1248] = ~((layer0_outputs[6869]) ^ (layer0_outputs[9598]));
    assign outputs[1249] = ~((layer0_outputs[5316]) ^ (layer0_outputs[5303]));
    assign outputs[1250] = (layer0_outputs[8880]) & ~(layer0_outputs[1117]);
    assign outputs[1251] = (layer0_outputs[6908]) & ~(layer0_outputs[1175]);
    assign outputs[1252] = ~((layer0_outputs[4533]) | (layer0_outputs[464]));
    assign outputs[1253] = (layer0_outputs[8627]) & (layer0_outputs[7932]);
    assign outputs[1254] = (layer0_outputs[6638]) & ~(layer0_outputs[5972]);
    assign outputs[1255] = ~(layer0_outputs[1713]);
    assign outputs[1256] = ~(layer0_outputs[6735]);
    assign outputs[1257] = (layer0_outputs[8537]) & (layer0_outputs[6532]);
    assign outputs[1258] = ~(layer0_outputs[8569]);
    assign outputs[1259] = (layer0_outputs[8319]) ^ (layer0_outputs[5675]);
    assign outputs[1260] = ~(layer0_outputs[278]);
    assign outputs[1261] = layer0_outputs[3855];
    assign outputs[1262] = ~((layer0_outputs[7481]) | (layer0_outputs[2639]));
    assign outputs[1263] = ~((layer0_outputs[9682]) | (layer0_outputs[9204]));
    assign outputs[1264] = (layer0_outputs[5991]) & (layer0_outputs[2653]);
    assign outputs[1265] = ~(layer0_outputs[850]);
    assign outputs[1266] = (layer0_outputs[8573]) & ~(layer0_outputs[8476]);
    assign outputs[1267] = layer0_outputs[7625];
    assign outputs[1268] = (layer0_outputs[4007]) & ~(layer0_outputs[7731]);
    assign outputs[1269] = ~(layer0_outputs[8279]);
    assign outputs[1270] = ~((layer0_outputs[7707]) ^ (layer0_outputs[9051]));
    assign outputs[1271] = (layer0_outputs[3898]) & ~(layer0_outputs[1966]);
    assign outputs[1272] = layer0_outputs[5860];
    assign outputs[1273] = ~(layer0_outputs[7021]) | (layer0_outputs[331]);
    assign outputs[1274] = layer0_outputs[3159];
    assign outputs[1275] = (layer0_outputs[7218]) & ~(layer0_outputs[1980]);
    assign outputs[1276] = ~((layer0_outputs[8344]) ^ (layer0_outputs[3152]));
    assign outputs[1277] = ~(layer0_outputs[5601]);
    assign outputs[1278] = (layer0_outputs[6135]) & ~(layer0_outputs[1827]);
    assign outputs[1279] = ~((layer0_outputs[3266]) | (layer0_outputs[5624]));
    assign outputs[1280] = (layer0_outputs[9499]) & ~(layer0_outputs[9610]);
    assign outputs[1281] = layer0_outputs[5915];
    assign outputs[1282] = ~((layer0_outputs[5379]) ^ (layer0_outputs[6682]));
    assign outputs[1283] = ~((layer0_outputs[398]) | (layer0_outputs[1352]));
    assign outputs[1284] = layer0_outputs[1848];
    assign outputs[1285] = (layer0_outputs[10022]) & ~(layer0_outputs[7191]);
    assign outputs[1286] = ~(layer0_outputs[936]);
    assign outputs[1287] = ~(layer0_outputs[10201]);
    assign outputs[1288] = ~(layer0_outputs[936]);
    assign outputs[1289] = layer0_outputs[5741];
    assign outputs[1290] = ~((layer0_outputs[3248]) | (layer0_outputs[7226]));
    assign outputs[1291] = (layer0_outputs[4941]) & ~(layer0_outputs[2649]);
    assign outputs[1292] = layer0_outputs[1569];
    assign outputs[1293] = ~((layer0_outputs[2644]) ^ (layer0_outputs[5373]));
    assign outputs[1294] = ~(layer0_outputs[7197]);
    assign outputs[1295] = layer0_outputs[7212];
    assign outputs[1296] = layer0_outputs[3078];
    assign outputs[1297] = (layer0_outputs[1354]) ^ (layer0_outputs[2200]);
    assign outputs[1298] = 1'b0;
    assign outputs[1299] = (layer0_outputs[4886]) & ~(layer0_outputs[6190]);
    assign outputs[1300] = (layer0_outputs[9994]) & ~(layer0_outputs[5046]);
    assign outputs[1301] = (layer0_outputs[2676]) & ~(layer0_outputs[4052]);
    assign outputs[1302] = (layer0_outputs[9591]) & ~(layer0_outputs[2322]);
    assign outputs[1303] = layer0_outputs[2795];
    assign outputs[1304] = ~((layer0_outputs[4877]) ^ (layer0_outputs[6509]));
    assign outputs[1305] = ~(layer0_outputs[4647]);
    assign outputs[1306] = (layer0_outputs[9408]) & ~(layer0_outputs[978]);
    assign outputs[1307] = ~(layer0_outputs[2587]);
    assign outputs[1308] = layer0_outputs[224];
    assign outputs[1309] = ~((layer0_outputs[3525]) ^ (layer0_outputs[4047]));
    assign outputs[1310] = (layer0_outputs[3552]) ^ (layer0_outputs[1085]);
    assign outputs[1311] = (layer0_outputs[6580]) & ~(layer0_outputs[842]);
    assign outputs[1312] = (layer0_outputs[6893]) & (layer0_outputs[8990]);
    assign outputs[1313] = (layer0_outputs[9465]) & ~(layer0_outputs[9090]);
    assign outputs[1314] = ~(layer0_outputs[8122]) | (layer0_outputs[5040]);
    assign outputs[1315] = (layer0_outputs[1455]) & ~(layer0_outputs[773]);
    assign outputs[1316] = (layer0_outputs[2524]) | (layer0_outputs[8579]);
    assign outputs[1317] = ~(layer0_outputs[4055]);
    assign outputs[1318] = ~((layer0_outputs[3120]) ^ (layer0_outputs[7235]));
    assign outputs[1319] = (layer0_outputs[6532]) ^ (layer0_outputs[6068]);
    assign outputs[1320] = 1'b0;
    assign outputs[1321] = (layer0_outputs[4984]) & ~(layer0_outputs[8488]);
    assign outputs[1322] = layer0_outputs[797];
    assign outputs[1323] = ~((layer0_outputs[6093]) | (layer0_outputs[4499]));
    assign outputs[1324] = (layer0_outputs[1736]) & (layer0_outputs[3804]);
    assign outputs[1325] = (layer0_outputs[309]) & (layer0_outputs[5745]);
    assign outputs[1326] = (layer0_outputs[7499]) & (layer0_outputs[9896]);
    assign outputs[1327] = ~((layer0_outputs[2187]) ^ (layer0_outputs[3830]));
    assign outputs[1328] = (layer0_outputs[4230]) ^ (layer0_outputs[8064]);
    assign outputs[1329] = ~((layer0_outputs[3270]) ^ (layer0_outputs[5326]));
    assign outputs[1330] = (layer0_outputs[7082]) & ~(layer0_outputs[3377]);
    assign outputs[1331] = (layer0_outputs[6403]) & ~(layer0_outputs[4952]);
    assign outputs[1332] = (layer0_outputs[443]) & ~(layer0_outputs[8246]);
    assign outputs[1333] = ~((layer0_outputs[6399]) | (layer0_outputs[9431]));
    assign outputs[1334] = ~((layer0_outputs[2840]) ^ (layer0_outputs[3962]));
    assign outputs[1335] = (layer0_outputs[711]) & ~(layer0_outputs[7483]);
    assign outputs[1336] = (layer0_outputs[2295]) ^ (layer0_outputs[555]);
    assign outputs[1337] = ~((layer0_outputs[9944]) | (layer0_outputs[7090]));
    assign outputs[1338] = (layer0_outputs[6345]) & (layer0_outputs[3834]);
    assign outputs[1339] = ~((layer0_outputs[3421]) | (layer0_outputs[7211]));
    assign outputs[1340] = (layer0_outputs[5044]) & (layer0_outputs[6659]);
    assign outputs[1341] = (layer0_outputs[2125]) & ~(layer0_outputs[4634]);
    assign outputs[1342] = 1'b0;
    assign outputs[1343] = layer0_outputs[3302];
    assign outputs[1344] = (layer0_outputs[8143]) & ~(layer0_outputs[7967]);
    assign outputs[1345] = ~(layer0_outputs[5787]);
    assign outputs[1346] = (layer0_outputs[8222]) & ~(layer0_outputs[2634]);
    assign outputs[1347] = layer0_outputs[2358];
    assign outputs[1348] = (layer0_outputs[6506]) & ~(layer0_outputs[7830]);
    assign outputs[1349] = (layer0_outputs[4025]) & (layer0_outputs[3250]);
    assign outputs[1350] = layer0_outputs[8016];
    assign outputs[1351] = ~((layer0_outputs[4280]) ^ (layer0_outputs[5034]));
    assign outputs[1352] = (layer0_outputs[302]) ^ (layer0_outputs[1919]);
    assign outputs[1353] = layer0_outputs[8608];
    assign outputs[1354] = (layer0_outputs[7366]) & ~(layer0_outputs[8700]);
    assign outputs[1355] = ~(layer0_outputs[4962]);
    assign outputs[1356] = ~(layer0_outputs[9070]);
    assign outputs[1357] = ~((layer0_outputs[6924]) | (layer0_outputs[9297]));
    assign outputs[1358] = (layer0_outputs[9578]) ^ (layer0_outputs[7805]);
    assign outputs[1359] = (layer0_outputs[8738]) ^ (layer0_outputs[2851]);
    assign outputs[1360] = (layer0_outputs[3550]) & ~(layer0_outputs[7144]);
    assign outputs[1361] = (layer0_outputs[9913]) & (layer0_outputs[7310]);
    assign outputs[1362] = (layer0_outputs[7007]) & ~(layer0_outputs[1955]);
    assign outputs[1363] = (layer0_outputs[477]) & ~(layer0_outputs[602]);
    assign outputs[1364] = ~((layer0_outputs[7256]) | (layer0_outputs[4731]));
    assign outputs[1365] = layer0_outputs[2568];
    assign outputs[1366] = layer0_outputs[6533];
    assign outputs[1367] = 1'b0;
    assign outputs[1368] = (layer0_outputs[6742]) ^ (layer0_outputs[7254]);
    assign outputs[1369] = layer0_outputs[8626];
    assign outputs[1370] = layer0_outputs[5547];
    assign outputs[1371] = layer0_outputs[8375];
    assign outputs[1372] = layer0_outputs[4675];
    assign outputs[1373] = ~((layer0_outputs[9021]) ^ (layer0_outputs[5579]));
    assign outputs[1374] = (layer0_outputs[1479]) & ~(layer0_outputs[375]);
    assign outputs[1375] = ~((layer0_outputs[4744]) ^ (layer0_outputs[4244]));
    assign outputs[1376] = (layer0_outputs[3694]) & ~(layer0_outputs[1262]);
    assign outputs[1377] = (layer0_outputs[2304]) & ~(layer0_outputs[243]);
    assign outputs[1378] = (layer0_outputs[590]) | (layer0_outputs[1636]);
    assign outputs[1379] = (layer0_outputs[4625]) ^ (layer0_outputs[7995]);
    assign outputs[1380] = ~((layer0_outputs[2350]) | (layer0_outputs[6878]));
    assign outputs[1381] = (layer0_outputs[1081]) & (layer0_outputs[2688]);
    assign outputs[1382] = (layer0_outputs[8819]) ^ (layer0_outputs[7854]);
    assign outputs[1383] = (layer0_outputs[10020]) ^ (layer0_outputs[2622]);
    assign outputs[1384] = (layer0_outputs[3842]) & (layer0_outputs[6697]);
    assign outputs[1385] = (layer0_outputs[5770]) | (layer0_outputs[5462]);
    assign outputs[1386] = (layer0_outputs[1273]) & ~(layer0_outputs[10138]);
    assign outputs[1387] = (layer0_outputs[1387]) & ~(layer0_outputs[4243]);
    assign outputs[1388] = layer0_outputs[8218];
    assign outputs[1389] = ~(layer0_outputs[3141]);
    assign outputs[1390] = (layer0_outputs[2867]) ^ (layer0_outputs[2957]);
    assign outputs[1391] = (layer0_outputs[13]) & (layer0_outputs[9900]);
    assign outputs[1392] = (layer0_outputs[3785]) & ~(layer0_outputs[3189]);
    assign outputs[1393] = ~((layer0_outputs[2671]) | (layer0_outputs[7472]));
    assign outputs[1394] = (layer0_outputs[2106]) & ~(layer0_outputs[4349]);
    assign outputs[1395] = (layer0_outputs[5133]) & ~(layer0_outputs[5587]);
    assign outputs[1396] = (layer0_outputs[1435]) & ~(layer0_outputs[4041]);
    assign outputs[1397] = (layer0_outputs[4328]) | (layer0_outputs[8871]);
    assign outputs[1398] = (layer0_outputs[10179]) & (layer0_outputs[4478]);
    assign outputs[1399] = (layer0_outputs[9096]) & (layer0_outputs[5590]);
    assign outputs[1400] = layer0_outputs[5266];
    assign outputs[1401] = ~(layer0_outputs[7116]);
    assign outputs[1402] = ~((layer0_outputs[1877]) | (layer0_outputs[1887]));
    assign outputs[1403] = 1'b0;
    assign outputs[1404] = ~((layer0_outputs[4988]) ^ (layer0_outputs[2269]));
    assign outputs[1405] = (layer0_outputs[2844]) & ~(layer0_outputs[8572]);
    assign outputs[1406] = (layer0_outputs[2668]) & ~(layer0_outputs[8515]);
    assign outputs[1407] = ~(layer0_outputs[9778]);
    assign outputs[1408] = (layer0_outputs[6722]) & ~(layer0_outputs[1005]);
    assign outputs[1409] = (layer0_outputs[2049]) & ~(layer0_outputs[6731]);
    assign outputs[1410] = layer0_outputs[9703];
    assign outputs[1411] = ~((layer0_outputs[4878]) & (layer0_outputs[3549]));
    assign outputs[1412] = (layer0_outputs[6695]) & (layer0_outputs[2164]);
    assign outputs[1413] = ~((layer0_outputs[6387]) ^ (layer0_outputs[445]));
    assign outputs[1414] = ~((layer0_outputs[9250]) ^ (layer0_outputs[2145]));
    assign outputs[1415] = layer0_outputs[6953];
    assign outputs[1416] = ~((layer0_outputs[5443]) | (layer0_outputs[176]));
    assign outputs[1417] = (layer0_outputs[180]) & ~(layer0_outputs[4441]);
    assign outputs[1418] = (layer0_outputs[4178]) & ~(layer0_outputs[2648]);
    assign outputs[1419] = ~((layer0_outputs[4938]) | (layer0_outputs[5468]));
    assign outputs[1420] = 1'b0;
    assign outputs[1421] = ~(layer0_outputs[5597]) | (layer0_outputs[7646]);
    assign outputs[1422] = ~((layer0_outputs[2565]) & (layer0_outputs[3368]));
    assign outputs[1423] = 1'b0;
    assign outputs[1424] = layer0_outputs[1882];
    assign outputs[1425] = (layer0_outputs[5001]) & ~(layer0_outputs[6459]);
    assign outputs[1426] = ~((layer0_outputs[4377]) | (layer0_outputs[6241]));
    assign outputs[1427] = (layer0_outputs[7082]) & (layer0_outputs[4038]);
    assign outputs[1428] = layer0_outputs[3236];
    assign outputs[1429] = (layer0_outputs[3736]) & ~(layer0_outputs[1204]);
    assign outputs[1430] = (layer0_outputs[9922]) & (layer0_outputs[9122]);
    assign outputs[1431] = (layer0_outputs[6398]) & (layer0_outputs[8242]);
    assign outputs[1432] = ~((layer0_outputs[3774]) ^ (layer0_outputs[1378]));
    assign outputs[1433] = layer0_outputs[6895];
    assign outputs[1434] = ~(layer0_outputs[8914]);
    assign outputs[1435] = ~(layer0_outputs[3467]);
    assign outputs[1436] = ~(layer0_outputs[6426]);
    assign outputs[1437] = layer0_outputs[4661];
    assign outputs[1438] = (layer0_outputs[4219]) & (layer0_outputs[7426]);
    assign outputs[1439] = layer0_outputs[301];
    assign outputs[1440] = 1'b0;
    assign outputs[1441] = layer0_outputs[3168];
    assign outputs[1442] = layer0_outputs[9471];
    assign outputs[1443] = ~((layer0_outputs[6098]) & (layer0_outputs[4929]));
    assign outputs[1444] = ~((layer0_outputs[4247]) | (layer0_outputs[2442]));
    assign outputs[1445] = ~(layer0_outputs[340]);
    assign outputs[1446] = (layer0_outputs[6247]) ^ (layer0_outputs[4551]);
    assign outputs[1447] = layer0_outputs[7839];
    assign outputs[1448] = ~((layer0_outputs[8886]) ^ (layer0_outputs[4837]));
    assign outputs[1449] = layer0_outputs[3129];
    assign outputs[1450] = ~((layer0_outputs[7915]) | (layer0_outputs[10106]));
    assign outputs[1451] = layer0_outputs[1079];
    assign outputs[1452] = ~(layer0_outputs[3501]);
    assign outputs[1453] = (layer0_outputs[9143]) & ~(layer0_outputs[3689]);
    assign outputs[1454] = ~((layer0_outputs[1054]) | (layer0_outputs[3642]));
    assign outputs[1455] = ~((layer0_outputs[9983]) ^ (layer0_outputs[3867]));
    assign outputs[1456] = (layer0_outputs[7748]) & (layer0_outputs[31]);
    assign outputs[1457] = ~(layer0_outputs[4795]);
    assign outputs[1458] = (layer0_outputs[5876]) & (layer0_outputs[2326]);
    assign outputs[1459] = ~((layer0_outputs[1627]) | (layer0_outputs[677]));
    assign outputs[1460] = ~((layer0_outputs[7359]) ^ (layer0_outputs[8053]));
    assign outputs[1461] = ~(layer0_outputs[5474]);
    assign outputs[1462] = 1'b0;
    assign outputs[1463] = ~(layer0_outputs[2711]);
    assign outputs[1464] = ~((layer0_outputs[2190]) ^ (layer0_outputs[248]));
    assign outputs[1465] = ~(layer0_outputs[886]);
    assign outputs[1466] = ~(layer0_outputs[4344]);
    assign outputs[1467] = layer0_outputs[849];
    assign outputs[1468] = ~(layer0_outputs[597]);
    assign outputs[1469] = (layer0_outputs[2256]) & ~(layer0_outputs[2149]);
    assign outputs[1470] = ~((layer0_outputs[6688]) | (layer0_outputs[4108]));
    assign outputs[1471] = (layer0_outputs[816]) & ~(layer0_outputs[9555]);
    assign outputs[1472] = ~((layer0_outputs[8532]) ^ (layer0_outputs[9108]));
    assign outputs[1473] = (layer0_outputs[5246]) ^ (layer0_outputs[7739]);
    assign outputs[1474] = ~(layer0_outputs[8158]);
    assign outputs[1475] = ~(layer0_outputs[1502]);
    assign outputs[1476] = ~(layer0_outputs[169]);
    assign outputs[1477] = ~(layer0_outputs[5238]);
    assign outputs[1478] = ~((layer0_outputs[241]) | (layer0_outputs[3493]));
    assign outputs[1479] = (layer0_outputs[9642]) & (layer0_outputs[8182]);
    assign outputs[1480] = ~(layer0_outputs[1162]);
    assign outputs[1481] = ~(layer0_outputs[4677]);
    assign outputs[1482] = ~((layer0_outputs[7635]) | (layer0_outputs[7984]));
    assign outputs[1483] = ~(layer0_outputs[1252]);
    assign outputs[1484] = ~((layer0_outputs[6214]) | (layer0_outputs[7958]));
    assign outputs[1485] = ~((layer0_outputs[4684]) | (layer0_outputs[3664]));
    assign outputs[1486] = ~(layer0_outputs[10214]);
    assign outputs[1487] = ~((layer0_outputs[4068]) | (layer0_outputs[7789]));
    assign outputs[1488] = (layer0_outputs[1254]) ^ (layer0_outputs[2391]);
    assign outputs[1489] = ~(layer0_outputs[5953]);
    assign outputs[1490] = (layer0_outputs[5275]) & ~(layer0_outputs[3998]);
    assign outputs[1491] = (layer0_outputs[1757]) & ~(layer0_outputs[1266]);
    assign outputs[1492] = ~((layer0_outputs[5545]) | (layer0_outputs[240]));
    assign outputs[1493] = ~((layer0_outputs[3360]) ^ (layer0_outputs[8913]));
    assign outputs[1494] = 1'b0;
    assign outputs[1495] = ~((layer0_outputs[5147]) ^ (layer0_outputs[1659]));
    assign outputs[1496] = ~(layer0_outputs[9658]);
    assign outputs[1497] = ~(layer0_outputs[4962]);
    assign outputs[1498] = (layer0_outputs[8276]) ^ (layer0_outputs[1445]);
    assign outputs[1499] = ~((layer0_outputs[1083]) | (layer0_outputs[3906]));
    assign outputs[1500] = ~(layer0_outputs[2592]);
    assign outputs[1501] = ~(layer0_outputs[9184]);
    assign outputs[1502] = (layer0_outputs[302]) & (layer0_outputs[5483]);
    assign outputs[1503] = (layer0_outputs[7544]) ^ (layer0_outputs[3548]);
    assign outputs[1504] = (layer0_outputs[848]) ^ (layer0_outputs[372]);
    assign outputs[1505] = (layer0_outputs[1957]) ^ (layer0_outputs[6350]);
    assign outputs[1506] = (layer0_outputs[2103]) ^ (layer0_outputs[3454]);
    assign outputs[1507] = (layer0_outputs[5195]) & ~(layer0_outputs[9503]);
    assign outputs[1508] = layer0_outputs[836];
    assign outputs[1509] = (layer0_outputs[1467]) & (layer0_outputs[9635]);
    assign outputs[1510] = ~(layer0_outputs[984]);
    assign outputs[1511] = (layer0_outputs[1692]) & ~(layer0_outputs[8467]);
    assign outputs[1512] = ~((layer0_outputs[8027]) | (layer0_outputs[6493]));
    assign outputs[1513] = (layer0_outputs[1785]) ^ (layer0_outputs[8804]);
    assign outputs[1514] = 1'b0;
    assign outputs[1515] = layer0_outputs[5139];
    assign outputs[1516] = (layer0_outputs[5720]) & ~(layer0_outputs[6388]);
    assign outputs[1517] = ~(layer0_outputs[6727]);
    assign outputs[1518] = (layer0_outputs[9724]) ^ (layer0_outputs[10206]);
    assign outputs[1519] = ~((layer0_outputs[962]) ^ (layer0_outputs[8358]));
    assign outputs[1520] = ~(layer0_outputs[7918]);
    assign outputs[1521] = ~(layer0_outputs[10056]);
    assign outputs[1522] = (layer0_outputs[8994]) & (layer0_outputs[9491]);
    assign outputs[1523] = ~((layer0_outputs[4994]) | (layer0_outputs[4639]));
    assign outputs[1524] = ~(layer0_outputs[9328]);
    assign outputs[1525] = layer0_outputs[2632];
    assign outputs[1526] = (layer0_outputs[9236]) ^ (layer0_outputs[6975]);
    assign outputs[1527] = (layer0_outputs[3108]) & (layer0_outputs[4158]);
    assign outputs[1528] = ~(layer0_outputs[10078]);
    assign outputs[1529] = (layer0_outputs[4427]) & ~(layer0_outputs[1025]);
    assign outputs[1530] = ~(layer0_outputs[6451]);
    assign outputs[1531] = layer0_outputs[8716];
    assign outputs[1532] = (layer0_outputs[7187]) & ~(layer0_outputs[5224]);
    assign outputs[1533] = ~(layer0_outputs[4868]);
    assign outputs[1534] = (layer0_outputs[3345]) & ~(layer0_outputs[7859]);
    assign outputs[1535] = (layer0_outputs[7622]) & ~(layer0_outputs[195]);
    assign outputs[1536] = (layer0_outputs[2588]) & (layer0_outputs[9271]);
    assign outputs[1537] = ~((layer0_outputs[5214]) ^ (layer0_outputs[8329]));
    assign outputs[1538] = ~(layer0_outputs[1339]) | (layer0_outputs[7540]);
    assign outputs[1539] = ~(layer0_outputs[3941]);
    assign outputs[1540] = (layer0_outputs[2431]) & ~(layer0_outputs[2555]);
    assign outputs[1541] = ~((layer0_outputs[4658]) | (layer0_outputs[2311]));
    assign outputs[1542] = layer0_outputs[7178];
    assign outputs[1543] = ~(layer0_outputs[9022]);
    assign outputs[1544] = ~((layer0_outputs[2531]) | (layer0_outputs[3978]));
    assign outputs[1545] = layer0_outputs[2239];
    assign outputs[1546] = ~(layer0_outputs[6876]);
    assign outputs[1547] = (layer0_outputs[4540]) & ~(layer0_outputs[2331]);
    assign outputs[1548] = (layer0_outputs[1779]) & ~(layer0_outputs[4761]);
    assign outputs[1549] = ~(layer0_outputs[7052]);
    assign outputs[1550] = 1'b0;
    assign outputs[1551] = (layer0_outputs[3080]) & ~(layer0_outputs[3141]);
    assign outputs[1552] = (layer0_outputs[6289]) & (layer0_outputs[2273]);
    assign outputs[1553] = (layer0_outputs[8194]) & (layer0_outputs[2214]);
    assign outputs[1554] = layer0_outputs[4448];
    assign outputs[1555] = (layer0_outputs[2859]) & (layer0_outputs[5119]);
    assign outputs[1556] = (layer0_outputs[8924]) & ~(layer0_outputs[5013]);
    assign outputs[1557] = ~((layer0_outputs[884]) | (layer0_outputs[7205]));
    assign outputs[1558] = ~((layer0_outputs[2610]) | (layer0_outputs[687]));
    assign outputs[1559] = (layer0_outputs[7775]) & ~(layer0_outputs[5811]);
    assign outputs[1560] = ~(layer0_outputs[3813]);
    assign outputs[1561] = ~((layer0_outputs[4801]) & (layer0_outputs[5235]));
    assign outputs[1562] = (layer0_outputs[4155]) & ~(layer0_outputs[5782]);
    assign outputs[1563] = layer0_outputs[3076];
    assign outputs[1564] = layer0_outputs[396];
    assign outputs[1565] = (layer0_outputs[2194]) & ~(layer0_outputs[8824]);
    assign outputs[1566] = layer0_outputs[5018];
    assign outputs[1567] = ~((layer0_outputs[7010]) ^ (layer0_outputs[1847]));
    assign outputs[1568] = layer0_outputs[9097];
    assign outputs[1569] = ~(layer0_outputs[1252]);
    assign outputs[1570] = (layer0_outputs[4157]) & (layer0_outputs[4745]);
    assign outputs[1571] = ~(layer0_outputs[8180]);
    assign outputs[1572] = (layer0_outputs[8834]) ^ (layer0_outputs[10079]);
    assign outputs[1573] = (layer0_outputs[3396]) & ~(layer0_outputs[7132]);
    assign outputs[1574] = ~((layer0_outputs[6067]) ^ (layer0_outputs[616]));
    assign outputs[1575] = (layer0_outputs[5954]) & (layer0_outputs[6807]);
    assign outputs[1576] = ~((layer0_outputs[4513]) | (layer0_outputs[4302]));
    assign outputs[1577] = ~((layer0_outputs[3688]) | (layer0_outputs[7615]));
    assign outputs[1578] = (layer0_outputs[2967]) & (layer0_outputs[10124]);
    assign outputs[1579] = (layer0_outputs[3537]) & (layer0_outputs[8467]);
    assign outputs[1580] = (layer0_outputs[3547]) & ~(layer0_outputs[3027]);
    assign outputs[1581] = layer0_outputs[4549];
    assign outputs[1582] = (layer0_outputs[8800]) & ~(layer0_outputs[6521]);
    assign outputs[1583] = ~((layer0_outputs[4267]) | (layer0_outputs[4890]));
    assign outputs[1584] = (layer0_outputs[7877]) & ~(layer0_outputs[123]);
    assign outputs[1585] = ~(layer0_outputs[3445]);
    assign outputs[1586] = layer0_outputs[932];
    assign outputs[1587] = ~(layer0_outputs[2336]);
    assign outputs[1588] = ~((layer0_outputs[2021]) ^ (layer0_outputs[9520]));
    assign outputs[1589] = ~((layer0_outputs[5820]) ^ (layer0_outputs[3455]));
    assign outputs[1590] = (layer0_outputs[7238]) & (layer0_outputs[4676]);
    assign outputs[1591] = (layer0_outputs[2110]) ^ (layer0_outputs[9347]);
    assign outputs[1592] = ~(layer0_outputs[9973]);
    assign outputs[1593] = (layer0_outputs[8439]) ^ (layer0_outputs[2149]);
    assign outputs[1594] = layer0_outputs[4294];
    assign outputs[1595] = ~((layer0_outputs[988]) | (layer0_outputs[2659]));
    assign outputs[1596] = ~((layer0_outputs[8877]) | (layer0_outputs[7294]));
    assign outputs[1597] = (layer0_outputs[7348]) ^ (layer0_outputs[5444]);
    assign outputs[1598] = ~((layer0_outputs[3429]) ^ (layer0_outputs[7193]));
    assign outputs[1599] = ~(layer0_outputs[4926]);
    assign outputs[1600] = layer0_outputs[2833];
    assign outputs[1601] = layer0_outputs[6899];
    assign outputs[1602] = (layer0_outputs[3554]) & ~(layer0_outputs[4013]);
    assign outputs[1603] = ~(layer0_outputs[5356]);
    assign outputs[1604] = ~((layer0_outputs[966]) | (layer0_outputs[9550]));
    assign outputs[1605] = (layer0_outputs[5397]) | (layer0_outputs[9407]);
    assign outputs[1606] = ~((layer0_outputs[3477]) ^ (layer0_outputs[6790]));
    assign outputs[1607] = ~((layer0_outputs[9201]) ^ (layer0_outputs[7920]));
    assign outputs[1608] = ~(layer0_outputs[4756]);
    assign outputs[1609] = (layer0_outputs[9007]) ^ (layer0_outputs[2226]);
    assign outputs[1610] = (layer0_outputs[5184]) & ~(layer0_outputs[9952]);
    assign outputs[1611] = ~(layer0_outputs[96]);
    assign outputs[1612] = (layer0_outputs[4908]) & ~(layer0_outputs[68]);
    assign outputs[1613] = ~((layer0_outputs[2303]) | (layer0_outputs[10169]));
    assign outputs[1614] = ~(layer0_outputs[6508]);
    assign outputs[1615] = (layer0_outputs[3157]) & ~(layer0_outputs[5614]);
    assign outputs[1616] = (layer0_outputs[6816]) & ~(layer0_outputs[479]);
    assign outputs[1617] = ~(layer0_outputs[4717]);
    assign outputs[1618] = ~(layer0_outputs[7736]) | (layer0_outputs[7702]);
    assign outputs[1619] = (layer0_outputs[720]) & (layer0_outputs[3644]);
    assign outputs[1620] = (layer0_outputs[9553]) & ~(layer0_outputs[6750]);
    assign outputs[1621] = ~((layer0_outputs[8651]) ^ (layer0_outputs[2005]));
    assign outputs[1622] = layer0_outputs[2786];
    assign outputs[1623] = ~(layer0_outputs[5896]);
    assign outputs[1624] = ~((layer0_outputs[1477]) ^ (layer0_outputs[8570]));
    assign outputs[1625] = (layer0_outputs[8812]) & ~(layer0_outputs[8351]);
    assign outputs[1626] = ~((layer0_outputs[2390]) ^ (layer0_outputs[8244]));
    assign outputs[1627] = layer0_outputs[4249];
    assign outputs[1628] = ~((layer0_outputs[1670]) | (layer0_outputs[4313]));
    assign outputs[1629] = ~((layer0_outputs[5518]) ^ (layer0_outputs[9740]));
    assign outputs[1630] = ~(layer0_outputs[1325]);
    assign outputs[1631] = layer0_outputs[3696];
    assign outputs[1632] = layer0_outputs[1638];
    assign outputs[1633] = (layer0_outputs[9996]) ^ (layer0_outputs[5499]);
    assign outputs[1634] = layer0_outputs[7981];
    assign outputs[1635] = ~((layer0_outputs[4173]) ^ (layer0_outputs[4293]));
    assign outputs[1636] = (layer0_outputs[5496]) & (layer0_outputs[8971]);
    assign outputs[1637] = ~(layer0_outputs[5416]);
    assign outputs[1638] = layer0_outputs[7520];
    assign outputs[1639] = ~((layer0_outputs[4146]) | (layer0_outputs[3376]));
    assign outputs[1640] = (layer0_outputs[8475]) ^ (layer0_outputs[5551]);
    assign outputs[1641] = ~(layer0_outputs[7316]);
    assign outputs[1642] = ~((layer0_outputs[2394]) | (layer0_outputs[2012]));
    assign outputs[1643] = layer0_outputs[1710];
    assign outputs[1644] = ~((layer0_outputs[8813]) | (layer0_outputs[9066]));
    assign outputs[1645] = (layer0_outputs[7115]) & (layer0_outputs[4079]);
    assign outputs[1646] = (layer0_outputs[7215]) ^ (layer0_outputs[6634]);
    assign outputs[1647] = (layer0_outputs[1619]) ^ (layer0_outputs[8201]);
    assign outputs[1648] = (layer0_outputs[4079]) & ~(layer0_outputs[9346]);
    assign outputs[1649] = (layer0_outputs[3585]) & ~(layer0_outputs[3559]);
    assign outputs[1650] = (layer0_outputs[6491]) | (layer0_outputs[6348]);
    assign outputs[1651] = (layer0_outputs[1978]) & (layer0_outputs[8258]);
    assign outputs[1652] = ~((layer0_outputs[491]) | (layer0_outputs[1419]));
    assign outputs[1653] = layer0_outputs[2664];
    assign outputs[1654] = ~(layer0_outputs[4514]);
    assign outputs[1655] = layer0_outputs[10119];
    assign outputs[1656] = ~((layer0_outputs[9587]) | (layer0_outputs[9612]));
    assign outputs[1657] = layer0_outputs[5286];
    assign outputs[1658] = ~(layer0_outputs[8601]);
    assign outputs[1659] = ~((layer0_outputs[4644]) | (layer0_outputs[1718]));
    assign outputs[1660] = (layer0_outputs[8722]) & ~(layer0_outputs[7313]);
    assign outputs[1661] = (layer0_outputs[3493]) ^ (layer0_outputs[772]);
    assign outputs[1662] = ~(layer0_outputs[3428]);
    assign outputs[1663] = layer0_outputs[7309];
    assign outputs[1664] = ~((layer0_outputs[6181]) | (layer0_outputs[5426]));
    assign outputs[1665] = layer0_outputs[7695];
    assign outputs[1666] = (layer0_outputs[4687]) & (layer0_outputs[1557]);
    assign outputs[1667] = layer0_outputs[9540];
    assign outputs[1668] = (layer0_outputs[7929]) & (layer0_outputs[5217]);
    assign outputs[1669] = layer0_outputs[4896];
    assign outputs[1670] = ~((layer0_outputs[2703]) | (layer0_outputs[6025]));
    assign outputs[1671] = ~(layer0_outputs[7360]);
    assign outputs[1672] = (layer0_outputs[5374]) & ~(layer0_outputs[1137]);
    assign outputs[1673] = layer0_outputs[5673];
    assign outputs[1674] = (layer0_outputs[4526]) & ~(layer0_outputs[5453]);
    assign outputs[1675] = layer0_outputs[8204];
    assign outputs[1676] = (layer0_outputs[5281]) & ~(layer0_outputs[6607]);
    assign outputs[1677] = ~((layer0_outputs[8246]) | (layer0_outputs[1873]));
    assign outputs[1678] = ~((layer0_outputs[7437]) ^ (layer0_outputs[1567]));
    assign outputs[1679] = layer0_outputs[5579];
    assign outputs[1680] = ~((layer0_outputs[7429]) ^ (layer0_outputs[9284]));
    assign outputs[1681] = (layer0_outputs[10043]) & ~(layer0_outputs[3378]);
    assign outputs[1682] = ~((layer0_outputs[6286]) | (layer0_outputs[4438]));
    assign outputs[1683] = ~((layer0_outputs[7371]) ^ (layer0_outputs[7863]));
    assign outputs[1684] = (layer0_outputs[9309]) & ~(layer0_outputs[7206]);
    assign outputs[1685] = ~((layer0_outputs[6461]) ^ (layer0_outputs[10182]));
    assign outputs[1686] = ~((layer0_outputs[10211]) | (layer0_outputs[2826]));
    assign outputs[1687] = (layer0_outputs[9820]) & ~(layer0_outputs[9381]);
    assign outputs[1688] = ~((layer0_outputs[6589]) | (layer0_outputs[4226]));
    assign outputs[1689] = layer0_outputs[4396];
    assign outputs[1690] = ~((layer0_outputs[1740]) | (layer0_outputs[658]));
    assign outputs[1691] = (layer0_outputs[2686]) & ~(layer0_outputs[3234]);
    assign outputs[1692] = (layer0_outputs[5469]) & (layer0_outputs[2948]);
    assign outputs[1693] = (layer0_outputs[6020]) & ~(layer0_outputs[4393]);
    assign outputs[1694] = (layer0_outputs[1443]) ^ (layer0_outputs[6627]);
    assign outputs[1695] = (layer0_outputs[9462]) & (layer0_outputs[4456]);
    assign outputs[1696] = (layer0_outputs[3643]) & (layer0_outputs[8691]);
    assign outputs[1697] = (layer0_outputs[2182]) ^ (layer0_outputs[7717]);
    assign outputs[1698] = (layer0_outputs[2128]) & (layer0_outputs[4651]);
    assign outputs[1699] = ~(layer0_outputs[6941]);
    assign outputs[1700] = (layer0_outputs[4348]) & ~(layer0_outputs[2256]);
    assign outputs[1701] = layer0_outputs[4177];
    assign outputs[1702] = layer0_outputs[6304];
    assign outputs[1703] = layer0_outputs[9679];
    assign outputs[1704] = (layer0_outputs[4331]) & ~(layer0_outputs[1053]);
    assign outputs[1705] = ~(layer0_outputs[1481]);
    assign outputs[1706] = ~((layer0_outputs[9083]) | (layer0_outputs[5028]));
    assign outputs[1707] = (layer0_outputs[3273]) & (layer0_outputs[2118]);
    assign outputs[1708] = ~((layer0_outputs[6835]) ^ (layer0_outputs[8695]));
    assign outputs[1709] = (layer0_outputs[36]) & (layer0_outputs[808]);
    assign outputs[1710] = (layer0_outputs[5027]) ^ (layer0_outputs[5187]);
    assign outputs[1711] = (layer0_outputs[4212]) & (layer0_outputs[9631]);
    assign outputs[1712] = ~(layer0_outputs[5029]);
    assign outputs[1713] = ~((layer0_outputs[2126]) ^ (layer0_outputs[7443]));
    assign outputs[1714] = (layer0_outputs[292]) & (layer0_outputs[1000]);
    assign outputs[1715] = (layer0_outputs[3182]) & ~(layer0_outputs[5772]);
    assign outputs[1716] = ~((layer0_outputs[3436]) & (layer0_outputs[2159]));
    assign outputs[1717] = ~((layer0_outputs[5714]) ^ (layer0_outputs[1292]));
    assign outputs[1718] = ~(layer0_outputs[6337]);
    assign outputs[1719] = ~(layer0_outputs[2956]);
    assign outputs[1720] = ~(layer0_outputs[1366]);
    assign outputs[1721] = (layer0_outputs[7973]) & ~(layer0_outputs[2573]);
    assign outputs[1722] = (layer0_outputs[9240]) ^ (layer0_outputs[9441]);
    assign outputs[1723] = (layer0_outputs[3359]) & ~(layer0_outputs[7457]);
    assign outputs[1724] = ~((layer0_outputs[6976]) & (layer0_outputs[3008]));
    assign outputs[1725] = layer0_outputs[6933];
    assign outputs[1726] = (layer0_outputs[9053]) ^ (layer0_outputs[5563]);
    assign outputs[1727] = (layer0_outputs[7467]) & ~(layer0_outputs[6400]);
    assign outputs[1728] = ~(layer0_outputs[7387]);
    assign outputs[1729] = (layer0_outputs[6103]) & ~(layer0_outputs[411]);
    assign outputs[1730] = ~((layer0_outputs[2757]) | (layer0_outputs[9574]));
    assign outputs[1731] = (layer0_outputs[8250]) & ~(layer0_outputs[8503]);
    assign outputs[1732] = (layer0_outputs[8718]) & ~(layer0_outputs[3716]);
    assign outputs[1733] = layer0_outputs[2699];
    assign outputs[1734] = (layer0_outputs[9114]) ^ (layer0_outputs[5332]);
    assign outputs[1735] = (layer0_outputs[7383]) & ~(layer0_outputs[8686]);
    assign outputs[1736] = (layer0_outputs[7073]) & ~(layer0_outputs[4866]);
    assign outputs[1737] = ~((layer0_outputs[4152]) | (layer0_outputs[747]));
    assign outputs[1738] = (layer0_outputs[5075]) ^ (layer0_outputs[5728]);
    assign outputs[1739] = layer0_outputs[6596];
    assign outputs[1740] = (layer0_outputs[218]) & ~(layer0_outputs[7182]);
    assign outputs[1741] = ~((layer0_outputs[7039]) ^ (layer0_outputs[4010]));
    assign outputs[1742] = ~(layer0_outputs[6141]);
    assign outputs[1743] = (layer0_outputs[168]) & ~(layer0_outputs[2555]);
    assign outputs[1744] = ~((layer0_outputs[9977]) ^ (layer0_outputs[8420]));
    assign outputs[1745] = (layer0_outputs[3002]) ^ (layer0_outputs[9878]);
    assign outputs[1746] = ~(layer0_outputs[9638]);
    assign outputs[1747] = (layer0_outputs[6596]) & (layer0_outputs[3570]);
    assign outputs[1748] = ~((layer0_outputs[3937]) | (layer0_outputs[1945]));
    assign outputs[1749] = (layer0_outputs[3802]) & ~(layer0_outputs[7357]);
    assign outputs[1750] = ~((layer0_outputs[7540]) | (layer0_outputs[6347]));
    assign outputs[1751] = (layer0_outputs[3488]) & ~(layer0_outputs[4978]);
    assign outputs[1752] = layer0_outputs[8334];
    assign outputs[1753] = (layer0_outputs[6568]) & ~(layer0_outputs[5665]);
    assign outputs[1754] = ~(layer0_outputs[656]);
    assign outputs[1755] = ~((layer0_outputs[937]) | (layer0_outputs[531]));
    assign outputs[1756] = ~((layer0_outputs[5219]) | (layer0_outputs[5540]));
    assign outputs[1757] = ~((layer0_outputs[9101]) | (layer0_outputs[7305]));
    assign outputs[1758] = (layer0_outputs[5652]) & ~(layer0_outputs[7530]);
    assign outputs[1759] = ~((layer0_outputs[6255]) ^ (layer0_outputs[8241]));
    assign outputs[1760] = (layer0_outputs[9801]) & (layer0_outputs[2088]);
    assign outputs[1761] = layer0_outputs[1592];
    assign outputs[1762] = layer0_outputs[854];
    assign outputs[1763] = (layer0_outputs[220]) & ~(layer0_outputs[10]);
    assign outputs[1764] = ~(layer0_outputs[9269]);
    assign outputs[1765] = (layer0_outputs[3729]) & (layer0_outputs[1044]);
    assign outputs[1766] = ~((layer0_outputs[8436]) ^ (layer0_outputs[5970]));
    assign outputs[1767] = 1'b0;
    assign outputs[1768] = ~(layer0_outputs[8977]);
    assign outputs[1769] = (layer0_outputs[137]) & ~(layer0_outputs[8792]);
    assign outputs[1770] = ~(layer0_outputs[4927]);
    assign outputs[1771] = (layer0_outputs[10101]) ^ (layer0_outputs[8675]);
    assign outputs[1772] = (layer0_outputs[2691]) & (layer0_outputs[2972]);
    assign outputs[1773] = layer0_outputs[8419];
    assign outputs[1774] = (layer0_outputs[205]) ^ (layer0_outputs[5828]);
    assign outputs[1775] = (layer0_outputs[5337]) & ~(layer0_outputs[1964]);
    assign outputs[1776] = ~((layer0_outputs[9000]) | (layer0_outputs[7571]));
    assign outputs[1777] = ~((layer0_outputs[682]) | (layer0_outputs[9431]));
    assign outputs[1778] = ~(layer0_outputs[6436]);
    assign outputs[1779] = (layer0_outputs[4450]) & ~(layer0_outputs[5988]);
    assign outputs[1780] = (layer0_outputs[6943]) & ~(layer0_outputs[8559]);
    assign outputs[1781] = layer0_outputs[3241];
    assign outputs[1782] = ~((layer0_outputs[1453]) ^ (layer0_outputs[9884]));
    assign outputs[1783] = ~((layer0_outputs[7080]) ^ (layer0_outputs[8486]));
    assign outputs[1784] = 1'b0;
    assign outputs[1785] = (layer0_outputs[505]) ^ (layer0_outputs[2201]);
    assign outputs[1786] = ~((layer0_outputs[7562]) | (layer0_outputs[6451]));
    assign outputs[1787] = ~((layer0_outputs[154]) | (layer0_outputs[9361]));
    assign outputs[1788] = (layer0_outputs[529]) & ~(layer0_outputs[7729]);
    assign outputs[1789] = (layer0_outputs[689]) ^ (layer0_outputs[9529]);
    assign outputs[1790] = (layer0_outputs[6485]) & ~(layer0_outputs[687]);
    assign outputs[1791] = (layer0_outputs[8253]) & (layer0_outputs[5620]);
    assign outputs[1792] = ~((layer0_outputs[2736]) | (layer0_outputs[9884]));
    assign outputs[1793] = ~(layer0_outputs[1949]);
    assign outputs[1794] = layer0_outputs[9164];
    assign outputs[1795] = layer0_outputs[7788];
    assign outputs[1796] = ~((layer0_outputs[1529]) ^ (layer0_outputs[2181]));
    assign outputs[1797] = ~(layer0_outputs[4631]);
    assign outputs[1798] = layer0_outputs[9471];
    assign outputs[1799] = layer0_outputs[30];
    assign outputs[1800] = layer0_outputs[5133];
    assign outputs[1801] = (layer0_outputs[64]) ^ (layer0_outputs[5116]);
    assign outputs[1802] = ~(layer0_outputs[8043]);
    assign outputs[1803] = ~(layer0_outputs[6800]);
    assign outputs[1804] = (layer0_outputs[1164]) ^ (layer0_outputs[2622]);
    assign outputs[1805] = (layer0_outputs[5955]) & ~(layer0_outputs[8526]);
    assign outputs[1806] = ~(layer0_outputs[3457]);
    assign outputs[1807] = ~((layer0_outputs[733]) ^ (layer0_outputs[7176]));
    assign outputs[1808] = (layer0_outputs[5919]) & ~(layer0_outputs[1938]);
    assign outputs[1809] = ~((layer0_outputs[5859]) ^ (layer0_outputs[6782]));
    assign outputs[1810] = layer0_outputs[9401];
    assign outputs[1811] = (layer0_outputs[6461]) & ~(layer0_outputs[4342]);
    assign outputs[1812] = layer0_outputs[181];
    assign outputs[1813] = ~(layer0_outputs[8457]);
    assign outputs[1814] = (layer0_outputs[676]) ^ (layer0_outputs[2734]);
    assign outputs[1815] = layer0_outputs[8298];
    assign outputs[1816] = (layer0_outputs[9650]) & (layer0_outputs[7101]);
    assign outputs[1817] = (layer0_outputs[3215]) & (layer0_outputs[6361]);
    assign outputs[1818] = (layer0_outputs[2861]) & ~(layer0_outputs[5861]);
    assign outputs[1819] = ~((layer0_outputs[1281]) | (layer0_outputs[8677]));
    assign outputs[1820] = layer0_outputs[9102];
    assign outputs[1821] = (layer0_outputs[8179]) & ~(layer0_outputs[6182]);
    assign outputs[1822] = (layer0_outputs[950]) & (layer0_outputs[6812]);
    assign outputs[1823] = (layer0_outputs[3460]) & ~(layer0_outputs[8604]);
    assign outputs[1824] = layer0_outputs[6124];
    assign outputs[1825] = ~((layer0_outputs[3576]) | (layer0_outputs[2791]));
    assign outputs[1826] = 1'b0;
    assign outputs[1827] = (layer0_outputs[4809]) & ~(layer0_outputs[463]);
    assign outputs[1828] = layer0_outputs[8565];
    assign outputs[1829] = (layer0_outputs[3777]) & ~(layer0_outputs[10039]);
    assign outputs[1830] = layer0_outputs[8586];
    assign outputs[1831] = (layer0_outputs[7701]) ^ (layer0_outputs[1114]);
    assign outputs[1832] = ~((layer0_outputs[7918]) | (layer0_outputs[1009]));
    assign outputs[1833] = (layer0_outputs[5297]) & ~(layer0_outputs[1329]);
    assign outputs[1834] = ~((layer0_outputs[7576]) | (layer0_outputs[5226]));
    assign outputs[1835] = ~(layer0_outputs[5971]);
    assign outputs[1836] = layer0_outputs[849];
    assign outputs[1837] = (layer0_outputs[1754]) & ~(layer0_outputs[4600]);
    assign outputs[1838] = ~(layer0_outputs[6323]);
    assign outputs[1839] = (layer0_outputs[1546]) & (layer0_outputs[5707]);
    assign outputs[1840] = (layer0_outputs[7070]) & ~(layer0_outputs[5742]);
    assign outputs[1841] = (layer0_outputs[9612]) & ~(layer0_outputs[9939]);
    assign outputs[1842] = (layer0_outputs[5746]) & ~(layer0_outputs[9677]);
    assign outputs[1843] = ~(layer0_outputs[8959]);
    assign outputs[1844] = layer0_outputs[9241];
    assign outputs[1845] = 1'b0;
    assign outputs[1846] = ~((layer0_outputs[8117]) ^ (layer0_outputs[3273]));
    assign outputs[1847] = (layer0_outputs[5735]) & ~(layer0_outputs[9400]);
    assign outputs[1848] = ~(layer0_outputs[9515]);
    assign outputs[1849] = (layer0_outputs[1976]) ^ (layer0_outputs[9200]);
    assign outputs[1850] = (layer0_outputs[1720]) ^ (layer0_outputs[8821]);
    assign outputs[1851] = (layer0_outputs[3365]) & ~(layer0_outputs[7087]);
    assign outputs[1852] = 1'b0;
    assign outputs[1853] = ~((layer0_outputs[7113]) | (layer0_outputs[7801]));
    assign outputs[1854] = ~((layer0_outputs[9277]) | (layer0_outputs[9249]));
    assign outputs[1855] = layer0_outputs[2589];
    assign outputs[1856] = (layer0_outputs[1585]) & ~(layer0_outputs[3750]);
    assign outputs[1857] = layer0_outputs[1019];
    assign outputs[1858] = ~((layer0_outputs[7352]) ^ (layer0_outputs[1155]));
    assign outputs[1859] = (layer0_outputs[3139]) & ~(layer0_outputs[8715]);
    assign outputs[1860] = layer0_outputs[5743];
    assign outputs[1861] = (layer0_outputs[2470]) ^ (layer0_outputs[9200]);
    assign outputs[1862] = (layer0_outputs[8366]) & (layer0_outputs[5757]);
    assign outputs[1863] = (layer0_outputs[8550]) ^ (layer0_outputs[8864]);
    assign outputs[1864] = (layer0_outputs[767]) & ~(layer0_outputs[1154]);
    assign outputs[1865] = ~((layer0_outputs[3966]) ^ (layer0_outputs[8025]));
    assign outputs[1866] = (layer0_outputs[4231]) & ~(layer0_outputs[6444]);
    assign outputs[1867] = layer0_outputs[4956];
    assign outputs[1868] = ~(layer0_outputs[3602]);
    assign outputs[1869] = ~(layer0_outputs[1795]);
    assign outputs[1870] = 1'b0;
    assign outputs[1871] = (layer0_outputs[6287]) ^ (layer0_outputs[2704]);
    assign outputs[1872] = ~(layer0_outputs[4449]);
    assign outputs[1873] = (layer0_outputs[2106]) ^ (layer0_outputs[8425]);
    assign outputs[1874] = ~((layer0_outputs[8003]) | (layer0_outputs[10207]));
    assign outputs[1875] = (layer0_outputs[10002]) & ~(layer0_outputs[8214]);
    assign outputs[1876] = ~((layer0_outputs[3588]) | (layer0_outputs[6096]));
    assign outputs[1877] = ~(layer0_outputs[79]);
    assign outputs[1878] = ~(layer0_outputs[7910]) | (layer0_outputs[6308]);
    assign outputs[1879] = ~((layer0_outputs[744]) ^ (layer0_outputs[369]));
    assign outputs[1880] = ~(layer0_outputs[597]);
    assign outputs[1881] = (layer0_outputs[9635]) & ~(layer0_outputs[9218]);
    assign outputs[1882] = ~((layer0_outputs[1981]) | (layer0_outputs[188]));
    assign outputs[1883] = layer0_outputs[4282];
    assign outputs[1884] = ~(layer0_outputs[8020]);
    assign outputs[1885] = ~((layer0_outputs[2911]) | (layer0_outputs[9166]));
    assign outputs[1886] = layer0_outputs[2230];
    assign outputs[1887] = (layer0_outputs[6076]) & (layer0_outputs[9511]);
    assign outputs[1888] = ~(layer0_outputs[7360]);
    assign outputs[1889] = (layer0_outputs[1496]) & ~(layer0_outputs[2877]);
    assign outputs[1890] = (layer0_outputs[7109]) & ~(layer0_outputs[565]);
    assign outputs[1891] = (layer0_outputs[6760]) & ~(layer0_outputs[2580]);
    assign outputs[1892] = (layer0_outputs[2333]) & ~(layer0_outputs[3458]);
    assign outputs[1893] = layer0_outputs[9583];
    assign outputs[1894] = (layer0_outputs[2695]) & ~(layer0_outputs[363]);
    assign outputs[1895] = (layer0_outputs[7526]) ^ (layer0_outputs[3544]);
    assign outputs[1896] = ~((layer0_outputs[715]) ^ (layer0_outputs[6667]));
    assign outputs[1897] = (layer0_outputs[5403]) & (layer0_outputs[6440]);
    assign outputs[1898] = (layer0_outputs[7955]) & (layer0_outputs[2854]);
    assign outputs[1899] = ~(layer0_outputs[6752]);
    assign outputs[1900] = ~(layer0_outputs[4985]);
    assign outputs[1901] = (layer0_outputs[10179]) & (layer0_outputs[8584]);
    assign outputs[1902] = (layer0_outputs[1719]) & ~(layer0_outputs[6236]);
    assign outputs[1903] = (layer0_outputs[8050]) & ~(layer0_outputs[7281]);
    assign outputs[1904] = (layer0_outputs[345]) & ~(layer0_outputs[7924]);
    assign outputs[1905] = ~(layer0_outputs[1069]);
    assign outputs[1906] = (layer0_outputs[3426]) & ~(layer0_outputs[8750]);
    assign outputs[1907] = (layer0_outputs[2087]) ^ (layer0_outputs[2768]);
    assign outputs[1908] = ~((layer0_outputs[5034]) ^ (layer0_outputs[4207]));
    assign outputs[1909] = (layer0_outputs[2028]) & ~(layer0_outputs[8350]);
    assign outputs[1910] = layer0_outputs[2053];
    assign outputs[1911] = ~(layer0_outputs[5858]);
    assign outputs[1912] = layer0_outputs[638];
    assign outputs[1913] = 1'b0;
    assign outputs[1914] = layer0_outputs[89];
    assign outputs[1915] = (layer0_outputs[7763]) & (layer0_outputs[9834]);
    assign outputs[1916] = (layer0_outputs[4099]) & ~(layer0_outputs[9717]);
    assign outputs[1917] = (layer0_outputs[111]) & ~(layer0_outputs[2726]);
    assign outputs[1918] = ~(layer0_outputs[2497]);
    assign outputs[1919] = (layer0_outputs[1165]) & ~(layer0_outputs[567]);
    assign outputs[1920] = (layer0_outputs[5042]) & ~(layer0_outputs[6324]);
    assign outputs[1921] = ~((layer0_outputs[1734]) ^ (layer0_outputs[1670]));
    assign outputs[1922] = layer0_outputs[8593];
    assign outputs[1923] = layer0_outputs[7531];
    assign outputs[1924] = layer0_outputs[6787];
    assign outputs[1925] = ~((layer0_outputs[1918]) | (layer0_outputs[1758]));
    assign outputs[1926] = (layer0_outputs[1774]) & ~(layer0_outputs[5067]);
    assign outputs[1927] = (layer0_outputs[1933]) ^ (layer0_outputs[5481]);
    assign outputs[1928] = (layer0_outputs[592]) ^ (layer0_outputs[5473]);
    assign outputs[1929] = ~(layer0_outputs[8590]);
    assign outputs[1930] = ~(layer0_outputs[9748]);
    assign outputs[1931] = layer0_outputs[6350];
    assign outputs[1932] = ~((layer0_outputs[9964]) ^ (layer0_outputs[5719]));
    assign outputs[1933] = layer0_outputs[9374];
    assign outputs[1934] = (layer0_outputs[10212]) ^ (layer0_outputs[6437]);
    assign outputs[1935] = (layer0_outputs[2741]) & (layer0_outputs[6687]);
    assign outputs[1936] = ~(layer0_outputs[1254]) | (layer0_outputs[5821]);
    assign outputs[1937] = (layer0_outputs[1701]) & (layer0_outputs[4754]);
    assign outputs[1938] = layer0_outputs[3286];
    assign outputs[1939] = layer0_outputs[1971];
    assign outputs[1940] = ~((layer0_outputs[2376]) | (layer0_outputs[6889]));
    assign outputs[1941] = layer0_outputs[2086];
    assign outputs[1942] = (layer0_outputs[1159]) & ~(layer0_outputs[1232]);
    assign outputs[1943] = ~(layer0_outputs[8951]);
    assign outputs[1944] = ~((layer0_outputs[9586]) | (layer0_outputs[5408]));
    assign outputs[1945] = (layer0_outputs[2594]) ^ (layer0_outputs[6509]);
    assign outputs[1946] = (layer0_outputs[2625]) & (layer0_outputs[5379]);
    assign outputs[1947] = 1'b0;
    assign outputs[1948] = ~(layer0_outputs[2895]);
    assign outputs[1949] = (layer0_outputs[4596]) & ~(layer0_outputs[2959]);
    assign outputs[1950] = (layer0_outputs[7897]) ^ (layer0_outputs[1169]);
    assign outputs[1951] = (layer0_outputs[3057]) ^ (layer0_outputs[5383]);
    assign outputs[1952] = (layer0_outputs[7860]) & ~(layer0_outputs[8624]);
    assign outputs[1953] = (layer0_outputs[2307]) ^ (layer0_outputs[10125]);
    assign outputs[1954] = ~(layer0_outputs[9912]);
    assign outputs[1955] = ~((layer0_outputs[8156]) | (layer0_outputs[1089]));
    assign outputs[1956] = (layer0_outputs[7630]) & (layer0_outputs[1220]);
    assign outputs[1957] = ~(layer0_outputs[10129]);
    assign outputs[1958] = ~((layer0_outputs[6455]) ^ (layer0_outputs[6923]));
    assign outputs[1959] = (layer0_outputs[5721]) & ~(layer0_outputs[1895]);
    assign outputs[1960] = (layer0_outputs[7503]) & ~(layer0_outputs[1115]);
    assign outputs[1961] = layer0_outputs[7207];
    assign outputs[1962] = layer0_outputs[1867];
    assign outputs[1963] = (layer0_outputs[3933]) ^ (layer0_outputs[8186]);
    assign outputs[1964] = layer0_outputs[3634];
    assign outputs[1965] = ~((layer0_outputs[2561]) ^ (layer0_outputs[8444]));
    assign outputs[1966] = (layer0_outputs[4157]) & (layer0_outputs[3365]);
    assign outputs[1967] = (layer0_outputs[5418]) & ~(layer0_outputs[5691]);
    assign outputs[1968] = ~((layer0_outputs[9772]) | (layer0_outputs[527]));
    assign outputs[1969] = (layer0_outputs[963]) & ~(layer0_outputs[7641]);
    assign outputs[1970] = (layer0_outputs[4867]) & (layer0_outputs[4335]);
    assign outputs[1971] = (layer0_outputs[2190]) & (layer0_outputs[9067]);
    assign outputs[1972] = (layer0_outputs[9444]) & ~(layer0_outputs[6192]);
    assign outputs[1973] = (layer0_outputs[3517]) & ~(layer0_outputs[4429]);
    assign outputs[1974] = layer0_outputs[5292];
    assign outputs[1975] = layer0_outputs[3600];
    assign outputs[1976] = ~(layer0_outputs[2907]) | (layer0_outputs[7234]);
    assign outputs[1977] = ~(layer0_outputs[7303]);
    assign outputs[1978] = layer0_outputs[6966];
    assign outputs[1979] = ~(layer0_outputs[6330]);
    assign outputs[1980] = (layer0_outputs[9072]) & (layer0_outputs[6154]);
    assign outputs[1981] = ~((layer0_outputs[9625]) ^ (layer0_outputs[6086]));
    assign outputs[1982] = (layer0_outputs[5666]) ^ (layer0_outputs[8086]);
    assign outputs[1983] = ~((layer0_outputs[8832]) | (layer0_outputs[2783]));
    assign outputs[1984] = layer0_outputs[4723];
    assign outputs[1985] = (layer0_outputs[1291]) & ~(layer0_outputs[7869]);
    assign outputs[1986] = (layer0_outputs[4519]) & ~(layer0_outputs[3144]);
    assign outputs[1987] = ~(layer0_outputs[10131]);
    assign outputs[1988] = (layer0_outputs[1111]) ^ (layer0_outputs[5909]);
    assign outputs[1989] = ~((layer0_outputs[9613]) & (layer0_outputs[3341]));
    assign outputs[1990] = ~((layer0_outputs[1539]) | (layer0_outputs[5521]));
    assign outputs[1991] = (layer0_outputs[8962]) & (layer0_outputs[3285]);
    assign outputs[1992] = ~((layer0_outputs[7266]) ^ (layer0_outputs[2788]));
    assign outputs[1993] = ~((layer0_outputs[6370]) ^ (layer0_outputs[1280]));
    assign outputs[1994] = (layer0_outputs[3733]) & (layer0_outputs[7182]);
    assign outputs[1995] = 1'b0;
    assign outputs[1996] = ~((layer0_outputs[2846]) ^ (layer0_outputs[1677]));
    assign outputs[1997] = ~((layer0_outputs[6645]) | (layer0_outputs[559]));
    assign outputs[1998] = (layer0_outputs[5878]) & (layer0_outputs[2473]);
    assign outputs[1999] = layer0_outputs[1296];
    assign outputs[2000] = (layer0_outputs[4981]) & ~(layer0_outputs[4333]);
    assign outputs[2001] = layer0_outputs[7452];
    assign outputs[2002] = (layer0_outputs[3335]) & (layer0_outputs[7277]);
    assign outputs[2003] = ~((layer0_outputs[9529]) ^ (layer0_outputs[3146]));
    assign outputs[2004] = ~(layer0_outputs[3841]);
    assign outputs[2005] = (layer0_outputs[5847]) ^ (layer0_outputs[2931]);
    assign outputs[2006] = (layer0_outputs[871]) ^ (layer0_outputs[1008]);
    assign outputs[2007] = 1'b0;
    assign outputs[2008] = (layer0_outputs[8720]) & (layer0_outputs[3111]);
    assign outputs[2009] = 1'b0;
    assign outputs[2010] = (layer0_outputs[2174]) & (layer0_outputs[2433]);
    assign outputs[2011] = ~((layer0_outputs[10187]) ^ (layer0_outputs[2504]));
    assign outputs[2012] = (layer0_outputs[6268]) & ~(layer0_outputs[3174]);
    assign outputs[2013] = layer0_outputs[4986];
    assign outputs[2014] = ~(layer0_outputs[3430]);
    assign outputs[2015] = ~(layer0_outputs[3530]);
    assign outputs[2016] = ~((layer0_outputs[10205]) ^ (layer0_outputs[3556]));
    assign outputs[2017] = layer0_outputs[9988];
    assign outputs[2018] = ~(layer0_outputs[193]);
    assign outputs[2019] = ~((layer0_outputs[8469]) ^ (layer0_outputs[7463]));
    assign outputs[2020] = layer0_outputs[9947];
    assign outputs[2021] = ~((layer0_outputs[872]) ^ (layer0_outputs[1208]));
    assign outputs[2022] = layer0_outputs[416];
    assign outputs[2023] = ~((layer0_outputs[6511]) | (layer0_outputs[9384]));
    assign outputs[2024] = (layer0_outputs[5757]) & ~(layer0_outputs[2284]);
    assign outputs[2025] = ~(layer0_outputs[3883]);
    assign outputs[2026] = ~((layer0_outputs[528]) ^ (layer0_outputs[354]));
    assign outputs[2027] = (layer0_outputs[1681]) & ~(layer0_outputs[771]);
    assign outputs[2028] = ~((layer0_outputs[8054]) ^ (layer0_outputs[9883]));
    assign outputs[2029] = (layer0_outputs[270]) & ~(layer0_outputs[6747]);
    assign outputs[2030] = layer0_outputs[3711];
    assign outputs[2031] = (layer0_outputs[9327]) & ~(layer0_outputs[6129]);
    assign outputs[2032] = layer0_outputs[2051];
    assign outputs[2033] = layer0_outputs[7572];
    assign outputs[2034] = ~(layer0_outputs[4281]);
    assign outputs[2035] = (layer0_outputs[1447]) & (layer0_outputs[326]);
    assign outputs[2036] = (layer0_outputs[5347]) & ~(layer0_outputs[622]);
    assign outputs[2037] = ~((layer0_outputs[6576]) | (layer0_outputs[4744]));
    assign outputs[2038] = ~(layer0_outputs[202]);
    assign outputs[2039] = ~(layer0_outputs[1959]);
    assign outputs[2040] = ~((layer0_outputs[60]) & (layer0_outputs[5863]));
    assign outputs[2041] = ~(layer0_outputs[5247]);
    assign outputs[2042] = (layer0_outputs[6812]) & ~(layer0_outputs[3225]);
    assign outputs[2043] = ~((layer0_outputs[6148]) & (layer0_outputs[684]));
    assign outputs[2044] = (layer0_outputs[5801]) & ~(layer0_outputs[6641]);
    assign outputs[2045] = (layer0_outputs[9413]) | (layer0_outputs[5180]);
    assign outputs[2046] = layer0_outputs[8101];
    assign outputs[2047] = ~(layer0_outputs[6306]);
    assign outputs[2048] = ~(layer0_outputs[8791]);
    assign outputs[2049] = ~((layer0_outputs[3219]) & (layer0_outputs[2263]));
    assign outputs[2050] = (layer0_outputs[9765]) | (layer0_outputs[347]);
    assign outputs[2051] = ~(layer0_outputs[8445]);
    assign outputs[2052] = ~((layer0_outputs[8642]) & (layer0_outputs[10178]));
    assign outputs[2053] = (layer0_outputs[1309]) ^ (layer0_outputs[7977]);
    assign outputs[2054] = layer0_outputs[296];
    assign outputs[2055] = layer0_outputs[2368];
    assign outputs[2056] = ~((layer0_outputs[4780]) & (layer0_outputs[101]));
    assign outputs[2057] = ~((layer0_outputs[7322]) ^ (layer0_outputs[2655]));
    assign outputs[2058] = ~((layer0_outputs[3977]) ^ (layer0_outputs[38]));
    assign outputs[2059] = ~((layer0_outputs[876]) | (layer0_outputs[238]));
    assign outputs[2060] = ~((layer0_outputs[5692]) | (layer0_outputs[6044]));
    assign outputs[2061] = ~(layer0_outputs[702]);
    assign outputs[2062] = ~(layer0_outputs[3839]);
    assign outputs[2063] = layer0_outputs[2361];
    assign outputs[2064] = ~(layer0_outputs[7031]);
    assign outputs[2065] = ~(layer0_outputs[1150]);
    assign outputs[2066] = layer0_outputs[7547];
    assign outputs[2067] = (layer0_outputs[1566]) ^ (layer0_outputs[6492]);
    assign outputs[2068] = ~((layer0_outputs[1773]) ^ (layer0_outputs[8697]));
    assign outputs[2069] = ~(layer0_outputs[6095]);
    assign outputs[2070] = layer0_outputs[841];
    assign outputs[2071] = (layer0_outputs[8897]) & ~(layer0_outputs[4230]);
    assign outputs[2072] = ~((layer0_outputs[9709]) ^ (layer0_outputs[7878]));
    assign outputs[2073] = ~((layer0_outputs[1695]) ^ (layer0_outputs[10008]));
    assign outputs[2074] = ~((layer0_outputs[801]) ^ (layer0_outputs[4836]));
    assign outputs[2075] = ~((layer0_outputs[3887]) ^ (layer0_outputs[6452]));
    assign outputs[2076] = (layer0_outputs[5348]) & ~(layer0_outputs[9352]);
    assign outputs[2077] = 1'b1;
    assign outputs[2078] = ~((layer0_outputs[5820]) ^ (layer0_outputs[1433]));
    assign outputs[2079] = layer0_outputs[9321];
    assign outputs[2080] = ~((layer0_outputs[3238]) ^ (layer0_outputs[1099]));
    assign outputs[2081] = ~((layer0_outputs[3843]) & (layer0_outputs[1001]));
    assign outputs[2082] = (layer0_outputs[6559]) & ~(layer0_outputs[8243]);
    assign outputs[2083] = layer0_outputs[5716];
    assign outputs[2084] = layer0_outputs[649];
    assign outputs[2085] = ~(layer0_outputs[3050]);
    assign outputs[2086] = ~(layer0_outputs[4466]);
    assign outputs[2087] = ~((layer0_outputs[5950]) ^ (layer0_outputs[8067]));
    assign outputs[2088] = ~(layer0_outputs[5151]) | (layer0_outputs[5864]);
    assign outputs[2089] = ~(layer0_outputs[5368]) | (layer0_outputs[2937]);
    assign outputs[2090] = layer0_outputs[7065];
    assign outputs[2091] = layer0_outputs[4134];
    assign outputs[2092] = ~((layer0_outputs[9449]) ^ (layer0_outputs[3842]));
    assign outputs[2093] = ~(layer0_outputs[1777]);
    assign outputs[2094] = layer0_outputs[7441];
    assign outputs[2095] = ~(layer0_outputs[7592]) | (layer0_outputs[258]);
    assign outputs[2096] = ~(layer0_outputs[4365]);
    assign outputs[2097] = (layer0_outputs[8954]) & ~(layer0_outputs[6143]);
    assign outputs[2098] = layer0_outputs[516];
    assign outputs[2099] = layer0_outputs[4217];
    assign outputs[2100] = ~((layer0_outputs[5890]) ^ (layer0_outputs[1834]));
    assign outputs[2101] = ~((layer0_outputs[4054]) ^ (layer0_outputs[7501]));
    assign outputs[2102] = layer0_outputs[8813];
    assign outputs[2103] = ~((layer0_outputs[6015]) ^ (layer0_outputs[9247]));
    assign outputs[2104] = layer0_outputs[2995];
    assign outputs[2105] = layer0_outputs[10117];
    assign outputs[2106] = (layer0_outputs[6994]) & ~(layer0_outputs[3943]);
    assign outputs[2107] = ~((layer0_outputs[1188]) & (layer0_outputs[457]));
    assign outputs[2108] = layer0_outputs[4092];
    assign outputs[2109] = layer0_outputs[5595];
    assign outputs[2110] = layer0_outputs[7272];
    assign outputs[2111] = ~((layer0_outputs[7296]) & (layer0_outputs[7336]));
    assign outputs[2112] = layer0_outputs[1116];
    assign outputs[2113] = ~((layer0_outputs[8254]) | (layer0_outputs[1626]));
    assign outputs[2114] = ~((layer0_outputs[2019]) ^ (layer0_outputs[9944]));
    assign outputs[2115] = ~(layer0_outputs[2100]) | (layer0_outputs[1138]);
    assign outputs[2116] = (layer0_outputs[9965]) ^ (layer0_outputs[48]);
    assign outputs[2117] = (layer0_outputs[7981]) ^ (layer0_outputs[6548]);
    assign outputs[2118] = (layer0_outputs[6975]) | (layer0_outputs[3757]);
    assign outputs[2119] = layer0_outputs[7136];
    assign outputs[2120] = ~((layer0_outputs[5334]) ^ (layer0_outputs[6057]));
    assign outputs[2121] = layer0_outputs[7893];
    assign outputs[2122] = (layer0_outputs[4119]) ^ (layer0_outputs[569]);
    assign outputs[2123] = ~(layer0_outputs[1100]) | (layer0_outputs[9480]);
    assign outputs[2124] = ~((layer0_outputs[2888]) ^ (layer0_outputs[5863]));
    assign outputs[2125] = ~(layer0_outputs[307]) | (layer0_outputs[8882]);
    assign outputs[2126] = ~((layer0_outputs[3683]) ^ (layer0_outputs[380]));
    assign outputs[2127] = ~(layer0_outputs[9252]);
    assign outputs[2128] = ~(layer0_outputs[1096]);
    assign outputs[2129] = ~(layer0_outputs[2737]) | (layer0_outputs[3595]);
    assign outputs[2130] = ~((layer0_outputs[304]) & (layer0_outputs[7948]));
    assign outputs[2131] = layer0_outputs[9230];
    assign outputs[2132] = ~(layer0_outputs[3244]);
    assign outputs[2133] = ~((layer0_outputs[2224]) ^ (layer0_outputs[9071]));
    assign outputs[2134] = ~(layer0_outputs[49]);
    assign outputs[2135] = layer0_outputs[7307];
    assign outputs[2136] = (layer0_outputs[536]) & ~(layer0_outputs[7841]);
    assign outputs[2137] = layer0_outputs[9254];
    assign outputs[2138] = (layer0_outputs[5183]) ^ (layer0_outputs[1668]);
    assign outputs[2139] = ~(layer0_outputs[8774]);
    assign outputs[2140] = ~(layer0_outputs[9633]);
    assign outputs[2141] = ~((layer0_outputs[37]) | (layer0_outputs[4395]));
    assign outputs[2142] = (layer0_outputs[7480]) ^ (layer0_outputs[6008]);
    assign outputs[2143] = ~(layer0_outputs[6628]) | (layer0_outputs[7803]);
    assign outputs[2144] = ~(layer0_outputs[1584]) | (layer0_outputs[8215]);
    assign outputs[2145] = ~(layer0_outputs[8387]);
    assign outputs[2146] = (layer0_outputs[255]) & ~(layer0_outputs[5381]);
    assign outputs[2147] = (layer0_outputs[312]) ^ (layer0_outputs[400]);
    assign outputs[2148] = (layer0_outputs[5852]) & (layer0_outputs[512]);
    assign outputs[2149] = ~(layer0_outputs[4713]) | (layer0_outputs[6078]);
    assign outputs[2150] = ~(layer0_outputs[9319]);
    assign outputs[2151] = (layer0_outputs[3958]) | (layer0_outputs[7263]);
    assign outputs[2152] = ~((layer0_outputs[5930]) ^ (layer0_outputs[2177]));
    assign outputs[2153] = ~(layer0_outputs[9124]);
    assign outputs[2154] = ~(layer0_outputs[4109]);
    assign outputs[2155] = ~((layer0_outputs[5489]) ^ (layer0_outputs[6231]));
    assign outputs[2156] = ~((layer0_outputs[7248]) ^ (layer0_outputs[269]));
    assign outputs[2157] = layer0_outputs[4442];
    assign outputs[2158] = (layer0_outputs[3778]) ^ (layer0_outputs[6635]);
    assign outputs[2159] = layer0_outputs[4458];
    assign outputs[2160] = ~((layer0_outputs[3667]) & (layer0_outputs[3820]));
    assign outputs[2161] = ~((layer0_outputs[1637]) ^ (layer0_outputs[4710]));
    assign outputs[2162] = ~((layer0_outputs[153]) ^ (layer0_outputs[6534]));
    assign outputs[2163] = ~((layer0_outputs[9629]) & (layer0_outputs[194]));
    assign outputs[2164] = (layer0_outputs[5264]) | (layer0_outputs[6942]);
    assign outputs[2165] = ~((layer0_outputs[6738]) ^ (layer0_outputs[5510]));
    assign outputs[2166] = ~((layer0_outputs[1368]) & (layer0_outputs[4739]));
    assign outputs[2167] = layer0_outputs[8720];
    assign outputs[2168] = (layer0_outputs[1831]) ^ (layer0_outputs[7842]);
    assign outputs[2169] = ~(layer0_outputs[8730]);
    assign outputs[2170] = ~((layer0_outputs[519]) & (layer0_outputs[10096]));
    assign outputs[2171] = ~(layer0_outputs[915]) | (layer0_outputs[10208]);
    assign outputs[2172] = ~(layer0_outputs[2255]) | (layer0_outputs[5769]);
    assign outputs[2173] = ~((layer0_outputs[6849]) ^ (layer0_outputs[6165]));
    assign outputs[2174] = ~((layer0_outputs[9420]) & (layer0_outputs[2402]));
    assign outputs[2175] = ~(layer0_outputs[5951]);
    assign outputs[2176] = ~((layer0_outputs[7994]) ^ (layer0_outputs[8615]));
    assign outputs[2177] = ~(layer0_outputs[6172]);
    assign outputs[2178] = layer0_outputs[9120];
    assign outputs[2179] = (layer0_outputs[2196]) | (layer0_outputs[8453]);
    assign outputs[2180] = ~((layer0_outputs[7050]) & (layer0_outputs[7806]));
    assign outputs[2181] = ~((layer0_outputs[4918]) ^ (layer0_outputs[283]));
    assign outputs[2182] = ~(layer0_outputs[2452]);
    assign outputs[2183] = layer0_outputs[9853];
    assign outputs[2184] = (layer0_outputs[6034]) ^ (layer0_outputs[5231]);
    assign outputs[2185] = ~(layer0_outputs[8515]) | (layer0_outputs[3744]);
    assign outputs[2186] = (layer0_outputs[2479]) ^ (layer0_outputs[1112]);
    assign outputs[2187] = layer0_outputs[5535];
    assign outputs[2188] = (layer0_outputs[5032]) | (layer0_outputs[583]);
    assign outputs[2189] = (layer0_outputs[7223]) ^ (layer0_outputs[5665]);
    assign outputs[2190] = layer0_outputs[6741];
    assign outputs[2191] = ~(layer0_outputs[6084]);
    assign outputs[2192] = ~(layer0_outputs[1029]);
    assign outputs[2193] = ~(layer0_outputs[8157]);
    assign outputs[2194] = layer0_outputs[2966];
    assign outputs[2195] = (layer0_outputs[1341]) ^ (layer0_outputs[5859]);
    assign outputs[2196] = ~((layer0_outputs[10082]) | (layer0_outputs[7528]));
    assign outputs[2197] = (layer0_outputs[7460]) & ~(layer0_outputs[2026]);
    assign outputs[2198] = ~(layer0_outputs[8672]);
    assign outputs[2199] = ~(layer0_outputs[3327]) | (layer0_outputs[5087]);
    assign outputs[2200] = ~(layer0_outputs[7336]) | (layer0_outputs[3323]);
    assign outputs[2201] = ~((layer0_outputs[2659]) & (layer0_outputs[5817]));
    assign outputs[2202] = layer0_outputs[1680];
    assign outputs[2203] = ~(layer0_outputs[84]);
    assign outputs[2204] = ~(layer0_outputs[9617]) | (layer0_outputs[5398]);
    assign outputs[2205] = ~((layer0_outputs[874]) & (layer0_outputs[655]));
    assign outputs[2206] = (layer0_outputs[3149]) & ~(layer0_outputs[8081]);
    assign outputs[2207] = ~(layer0_outputs[2797]);
    assign outputs[2208] = ~(layer0_outputs[7558]);
    assign outputs[2209] = ~((layer0_outputs[2523]) ^ (layer0_outputs[8644]));
    assign outputs[2210] = ~(layer0_outputs[7413]) | (layer0_outputs[4583]);
    assign outputs[2211] = layer0_outputs[8224];
    assign outputs[2212] = ~(layer0_outputs[7507]);
    assign outputs[2213] = ~(layer0_outputs[754]) | (layer0_outputs[6421]);
    assign outputs[2214] = ~((layer0_outputs[3796]) ^ (layer0_outputs[612]));
    assign outputs[2215] = ~(layer0_outputs[6915]);
    assign outputs[2216] = ~((layer0_outputs[7761]) & (layer0_outputs[8753]));
    assign outputs[2217] = ~(layer0_outputs[9370]) | (layer0_outputs[5453]);
    assign outputs[2218] = ~(layer0_outputs[6604]);
    assign outputs[2219] = (layer0_outputs[8029]) ^ (layer0_outputs[5628]);
    assign outputs[2220] = ~((layer0_outputs[2462]) & (layer0_outputs[468]));
    assign outputs[2221] = (layer0_outputs[7974]) | (layer0_outputs[2960]);
    assign outputs[2222] = ~(layer0_outputs[4310]);
    assign outputs[2223] = (layer0_outputs[9484]) ^ (layer0_outputs[1178]);
    assign outputs[2224] = ~(layer0_outputs[9352]);
    assign outputs[2225] = ~(layer0_outputs[7720]) | (layer0_outputs[6647]);
    assign outputs[2226] = 1'b0;
    assign outputs[2227] = ~((layer0_outputs[133]) ^ (layer0_outputs[1398]));
    assign outputs[2228] = (layer0_outputs[1267]) & ~(layer0_outputs[7912]);
    assign outputs[2229] = ~((layer0_outputs[9516]) ^ (layer0_outputs[3468]));
    assign outputs[2230] = ~(layer0_outputs[3797]);
    assign outputs[2231] = (layer0_outputs[1487]) | (layer0_outputs[3027]);
    assign outputs[2232] = ~(layer0_outputs[2829]);
    assign outputs[2233] = ~(layer0_outputs[8939]) | (layer0_outputs[2666]);
    assign outputs[2234] = layer0_outputs[6710];
    assign outputs[2235] = ~(layer0_outputs[5237]);
    assign outputs[2236] = ~(layer0_outputs[7298]);
    assign outputs[2237] = layer0_outputs[1879];
    assign outputs[2238] = ~(layer0_outputs[7841]);
    assign outputs[2239] = (layer0_outputs[5004]) ^ (layer0_outputs[7114]);
    assign outputs[2240] = layer0_outputs[1401];
    assign outputs[2241] = ~((layer0_outputs[7888]) ^ (layer0_outputs[6883]));
    assign outputs[2242] = (layer0_outputs[1201]) | (layer0_outputs[4252]);
    assign outputs[2243] = (layer0_outputs[8779]) & (layer0_outputs[1755]);
    assign outputs[2244] = ~((layer0_outputs[2397]) | (layer0_outputs[7582]));
    assign outputs[2245] = ~(layer0_outputs[5923]) | (layer0_outputs[795]);
    assign outputs[2246] = layer0_outputs[7673];
    assign outputs[2247] = ~(layer0_outputs[7354]);
    assign outputs[2248] = (layer0_outputs[6969]) & ~(layer0_outputs[267]);
    assign outputs[2249] = ~(layer0_outputs[2011]);
    assign outputs[2250] = ~(layer0_outputs[6764]);
    assign outputs[2251] = ~(layer0_outputs[3064]);
    assign outputs[2252] = (layer0_outputs[3819]) & (layer0_outputs[1570]);
    assign outputs[2253] = (layer0_outputs[6342]) & (layer0_outputs[3659]);
    assign outputs[2254] = ~(layer0_outputs[8874]);
    assign outputs[2255] = ~((layer0_outputs[461]) ^ (layer0_outputs[7713]));
    assign outputs[2256] = (layer0_outputs[7401]) ^ (layer0_outputs[9356]);
    assign outputs[2257] = ~(layer0_outputs[7660]);
    assign outputs[2258] = ~(layer0_outputs[3102]);
    assign outputs[2259] = layer0_outputs[5266];
    assign outputs[2260] = layer0_outputs[4737];
    assign outputs[2261] = layer0_outputs[10000];
    assign outputs[2262] = ~((layer0_outputs[4463]) ^ (layer0_outputs[1047]));
    assign outputs[2263] = ~((layer0_outputs[6006]) & (layer0_outputs[4144]));
    assign outputs[2264] = 1'b1;
    assign outputs[2265] = 1'b1;
    assign outputs[2266] = ~((layer0_outputs[929]) ^ (layer0_outputs[2160]));
    assign outputs[2267] = ~(layer0_outputs[2801]) | (layer0_outputs[2538]);
    assign outputs[2268] = ~(layer0_outputs[10093]);
    assign outputs[2269] = ~(layer0_outputs[940]);
    assign outputs[2270] = ~(layer0_outputs[7835]);
    assign outputs[2271] = ~(layer0_outputs[9028]);
    assign outputs[2272] = ~(layer0_outputs[1257]);
    assign outputs[2273] = layer0_outputs[431];
    assign outputs[2274] = ~(layer0_outputs[510]);
    assign outputs[2275] = layer0_outputs[6012];
    assign outputs[2276] = (layer0_outputs[9174]) | (layer0_outputs[2285]);
    assign outputs[2277] = layer0_outputs[5538];
    assign outputs[2278] = ~((layer0_outputs[956]) ^ (layer0_outputs[4581]));
    assign outputs[2279] = layer0_outputs[7252];
    assign outputs[2280] = 1'b1;
    assign outputs[2281] = ~(layer0_outputs[2488]) | (layer0_outputs[6276]);
    assign outputs[2282] = ~(layer0_outputs[529]);
    assign outputs[2283] = (layer0_outputs[4167]) ^ (layer0_outputs[7169]);
    assign outputs[2284] = (layer0_outputs[4434]) & ~(layer0_outputs[2957]);
    assign outputs[2285] = ~(layer0_outputs[4770]) | (layer0_outputs[7156]);
    assign outputs[2286] = layer0_outputs[8739];
    assign outputs[2287] = layer0_outputs[8105];
    assign outputs[2288] = (layer0_outputs[576]) ^ (layer0_outputs[165]);
    assign outputs[2289] = layer0_outputs[7800];
    assign outputs[2290] = ~(layer0_outputs[5633]) | (layer0_outputs[8689]);
    assign outputs[2291] = (layer0_outputs[4171]) & ~(layer0_outputs[993]);
    assign outputs[2292] = ~(layer0_outputs[5874]);
    assign outputs[2293] = (layer0_outputs[304]) & ~(layer0_outputs[5723]);
    assign outputs[2294] = ~(layer0_outputs[9706]) | (layer0_outputs[8472]);
    assign outputs[2295] = ~(layer0_outputs[7696]);
    assign outputs[2296] = layer0_outputs[2949];
    assign outputs[2297] = ~((layer0_outputs[5877]) & (layer0_outputs[4922]));
    assign outputs[2298] = ~(layer0_outputs[1219]);
    assign outputs[2299] = ~((layer0_outputs[44]) ^ (layer0_outputs[955]));
    assign outputs[2300] = (layer0_outputs[1566]) & ~(layer0_outputs[7680]);
    assign outputs[2301] = ~((layer0_outputs[8446]) ^ (layer0_outputs[1537]));
    assign outputs[2302] = ~(layer0_outputs[5679]) | (layer0_outputs[5796]);
    assign outputs[2303] = ~(layer0_outputs[5024]);
    assign outputs[2304] = ~(layer0_outputs[6435]);
    assign outputs[2305] = (layer0_outputs[488]) & (layer0_outputs[7599]);
    assign outputs[2306] = (layer0_outputs[3199]) ^ (layer0_outputs[295]);
    assign outputs[2307] = ~(layer0_outputs[4958]);
    assign outputs[2308] = ~((layer0_outputs[821]) ^ (layer0_outputs[9311]));
    assign outputs[2309] = ~(layer0_outputs[1847]) | (layer0_outputs[5870]);
    assign outputs[2310] = ~((layer0_outputs[265]) ^ (layer0_outputs[7560]));
    assign outputs[2311] = ~(layer0_outputs[4943]) | (layer0_outputs[4290]);
    assign outputs[2312] = ~(layer0_outputs[3826]);
    assign outputs[2313] = layer0_outputs[649];
    assign outputs[2314] = ~(layer0_outputs[6520]) | (layer0_outputs[3180]);
    assign outputs[2315] = ~(layer0_outputs[4880]) | (layer0_outputs[2031]);
    assign outputs[2316] = ~(layer0_outputs[5884]);
    assign outputs[2317] = layer0_outputs[4465];
    assign outputs[2318] = ~((layer0_outputs[9294]) ^ (layer0_outputs[432]));
    assign outputs[2319] = ~(layer0_outputs[3902]) | (layer0_outputs[9454]);
    assign outputs[2320] = layer0_outputs[3307];
    assign outputs[2321] = ~((layer0_outputs[124]) ^ (layer0_outputs[4166]));
    assign outputs[2322] = ~((layer0_outputs[4429]) ^ (layer0_outputs[7506]));
    assign outputs[2323] = ~(layer0_outputs[702]);
    assign outputs[2324] = (layer0_outputs[1915]) & (layer0_outputs[5161]);
    assign outputs[2325] = layer0_outputs[6138];
    assign outputs[2326] = 1'b1;
    assign outputs[2327] = ~(layer0_outputs[7631]);
    assign outputs[2328] = ~(layer0_outputs[4184]);
    assign outputs[2329] = ~(layer0_outputs[899]);
    assign outputs[2330] = (layer0_outputs[5907]) & (layer0_outputs[9614]);
    assign outputs[2331] = ~((layer0_outputs[6957]) ^ (layer0_outputs[6653]));
    assign outputs[2332] = (layer0_outputs[361]) | (layer0_outputs[1786]);
    assign outputs[2333] = ~(layer0_outputs[3438]);
    assign outputs[2334] = ~(layer0_outputs[7892]);
    assign outputs[2335] = layer0_outputs[890];
    assign outputs[2336] = ~(layer0_outputs[905]);
    assign outputs[2337] = (layer0_outputs[8572]) | (layer0_outputs[6875]);
    assign outputs[2338] = layer0_outputs[8943];
    assign outputs[2339] = (layer0_outputs[7297]) ^ (layer0_outputs[6085]);
    assign outputs[2340] = (layer0_outputs[6567]) ^ (layer0_outputs[1868]);
    assign outputs[2341] = ~((layer0_outputs[4150]) & (layer0_outputs[2232]));
    assign outputs[2342] = layer0_outputs[7380];
    assign outputs[2343] = ~((layer0_outputs[7935]) | (layer0_outputs[2309]));
    assign outputs[2344] = ~((layer0_outputs[2746]) ^ (layer0_outputs[3956]));
    assign outputs[2345] = ~(layer0_outputs[9168]);
    assign outputs[2346] = ~(layer0_outputs[4833]) | (layer0_outputs[9893]);
    assign outputs[2347] = ~(layer0_outputs[8849]);
    assign outputs[2348] = ~(layer0_outputs[7405]) | (layer0_outputs[5979]);
    assign outputs[2349] = layer0_outputs[8153];
    assign outputs[2350] = 1'b1;
    assign outputs[2351] = (layer0_outputs[9274]) & (layer0_outputs[6692]);
    assign outputs[2352] = ~((layer0_outputs[9762]) & (layer0_outputs[3559]));
    assign outputs[2353] = ~(layer0_outputs[3236]);
    assign outputs[2354] = ~(layer0_outputs[9793]);
    assign outputs[2355] = layer0_outputs[9029];
    assign outputs[2356] = ~((layer0_outputs[8860]) ^ (layer0_outputs[7902]));
    assign outputs[2357] = ~(layer0_outputs[715]);
    assign outputs[2358] = ~(layer0_outputs[7966]);
    assign outputs[2359] = (layer0_outputs[2725]) | (layer0_outputs[2752]);
    assign outputs[2360] = 1'b1;
    assign outputs[2361] = ~((layer0_outputs[1536]) ^ (layer0_outputs[1645]));
    assign outputs[2362] = ~((layer0_outputs[9272]) ^ (layer0_outputs[6190]));
    assign outputs[2363] = ~(layer0_outputs[1381]);
    assign outputs[2364] = layer0_outputs[4752];
    assign outputs[2365] = layer0_outputs[1331];
    assign outputs[2366] = ~(layer0_outputs[5943]);
    assign outputs[2367] = ~(layer0_outputs[4884]);
    assign outputs[2368] = layer0_outputs[9760];
    assign outputs[2369] = (layer0_outputs[3278]) & ~(layer0_outputs[3884]);
    assign outputs[2370] = layer0_outputs[7462];
    assign outputs[2371] = (layer0_outputs[2852]) | (layer0_outputs[2858]);
    assign outputs[2372] = (layer0_outputs[2795]) ^ (layer0_outputs[7977]);
    assign outputs[2373] = layer0_outputs[3659];
    assign outputs[2374] = ~((layer0_outputs[8743]) ^ (layer0_outputs[5031]));
    assign outputs[2375] = (layer0_outputs[4033]) & ~(layer0_outputs[1642]);
    assign outputs[2376] = layer0_outputs[4464];
    assign outputs[2377] = layer0_outputs[3059];
    assign outputs[2378] = layer0_outputs[7141];
    assign outputs[2379] = ~((layer0_outputs[9722]) & (layer0_outputs[1259]));
    assign outputs[2380] = ~((layer0_outputs[9768]) & (layer0_outputs[6931]));
    assign outputs[2381] = ~(layer0_outputs[8898]) | (layer0_outputs[8247]);
    assign outputs[2382] = ~((layer0_outputs[438]) ^ (layer0_outputs[6368]));
    assign outputs[2383] = ~((layer0_outputs[8735]) & (layer0_outputs[1617]));
    assign outputs[2384] = ~(layer0_outputs[9087]) | (layer0_outputs[1809]);
    assign outputs[2385] = (layer0_outputs[3882]) & (layer0_outputs[3691]);
    assign outputs[2386] = ~(layer0_outputs[9901]) | (layer0_outputs[5119]);
    assign outputs[2387] = layer0_outputs[6215];
    assign outputs[2388] = ~((layer0_outputs[517]) ^ (layer0_outputs[6413]));
    assign outputs[2389] = layer0_outputs[10232];
    assign outputs[2390] = ~(layer0_outputs[8449]);
    assign outputs[2391] = ~((layer0_outputs[4071]) ^ (layer0_outputs[1393]));
    assign outputs[2392] = ~(layer0_outputs[6182]);
    assign outputs[2393] = ~((layer0_outputs[10235]) & (layer0_outputs[5779]));
    assign outputs[2394] = (layer0_outputs[2223]) & (layer0_outputs[9969]);
    assign outputs[2395] = ~(layer0_outputs[3011]);
    assign outputs[2396] = layer0_outputs[4902];
    assign outputs[2397] = (layer0_outputs[3381]) | (layer0_outputs[5734]);
    assign outputs[2398] = ~((layer0_outputs[2962]) ^ (layer0_outputs[6083]));
    assign outputs[2399] = layer0_outputs[5305];
    assign outputs[2400] = ~((layer0_outputs[5137]) ^ (layer0_outputs[8645]));
    assign outputs[2401] = ~(layer0_outputs[4372]);
    assign outputs[2402] = ~(layer0_outputs[8801]) | (layer0_outputs[9703]);
    assign outputs[2403] = (layer0_outputs[7764]) & ~(layer0_outputs[1408]);
    assign outputs[2404] = (layer0_outputs[4495]) ^ (layer0_outputs[231]);
    assign outputs[2405] = layer0_outputs[7024];
    assign outputs[2406] = ~(layer0_outputs[5755]);
    assign outputs[2407] = (layer0_outputs[8253]) ^ (layer0_outputs[1021]);
    assign outputs[2408] = (layer0_outputs[8505]) | (layer0_outputs[5365]);
    assign outputs[2409] = ~(layer0_outputs[1687]);
    assign outputs[2410] = layer0_outputs[3601];
    assign outputs[2411] = ~(layer0_outputs[9468]);
    assign outputs[2412] = layer0_outputs[334];
    assign outputs[2413] = (layer0_outputs[4557]) ^ (layer0_outputs[4084]);
    assign outputs[2414] = layer0_outputs[10070];
    assign outputs[2415] = ~(layer0_outputs[2969]);
    assign outputs[2416] = ~((layer0_outputs[1420]) ^ (layer0_outputs[3942]));
    assign outputs[2417] = ~(layer0_outputs[3350]);
    assign outputs[2418] = ~((layer0_outputs[3610]) ^ (layer0_outputs[4508]));
    assign outputs[2419] = ~(layer0_outputs[1050]) | (layer0_outputs[10059]);
    assign outputs[2420] = (layer0_outputs[7771]) & (layer0_outputs[3059]);
    assign outputs[2421] = ~(layer0_outputs[1290]) | (layer0_outputs[5332]);
    assign outputs[2422] = ~((layer0_outputs[4439]) | (layer0_outputs[8532]));
    assign outputs[2423] = ~(layer0_outputs[6250]);
    assign outputs[2424] = ~(layer0_outputs[7135]);
    assign outputs[2425] = layer0_outputs[8540];
    assign outputs[2426] = (layer0_outputs[1511]) & ~(layer0_outputs[1572]);
    assign outputs[2427] = ~(layer0_outputs[8656]);
    assign outputs[2428] = ~(layer0_outputs[8634]) | (layer0_outputs[6649]);
    assign outputs[2429] = ~(layer0_outputs[4892]) | (layer0_outputs[4185]);
    assign outputs[2430] = ~(layer0_outputs[4501]);
    assign outputs[2431] = (layer0_outputs[8451]) ^ (layer0_outputs[2803]);
    assign outputs[2432] = 1'b1;
    assign outputs[2433] = ~((layer0_outputs[1236]) & (layer0_outputs[6719]));
    assign outputs[2434] = (layer0_outputs[5125]) & ~(layer0_outputs[825]);
    assign outputs[2435] = ~(layer0_outputs[6291]);
    assign outputs[2436] = ~(layer0_outputs[4852]);
    assign outputs[2437] = ~((layer0_outputs[9375]) ^ (layer0_outputs[5798]));
    assign outputs[2438] = ~(layer0_outputs[4309]);
    assign outputs[2439] = ~(layer0_outputs[5410]);
    assign outputs[2440] = ~(layer0_outputs[69]);
    assign outputs[2441] = ~(layer0_outputs[3829]);
    assign outputs[2442] = ~(layer0_outputs[4005]);
    assign outputs[2443] = ~(layer0_outputs[8139]);
    assign outputs[2444] = (layer0_outputs[1768]) & ~(layer0_outputs[8452]);
    assign outputs[2445] = ~(layer0_outputs[5522]) | (layer0_outputs[8419]);
    assign outputs[2446] = ~((layer0_outputs[8141]) ^ (layer0_outputs[2366]));
    assign outputs[2447] = ~((layer0_outputs[4070]) ^ (layer0_outputs[6868]));
    assign outputs[2448] = layer0_outputs[5610];
    assign outputs[2449] = ~(layer0_outputs[4272]);
    assign outputs[2450] = ~((layer0_outputs[9408]) & (layer0_outputs[2444]));
    assign outputs[2451] = layer0_outputs[10010];
    assign outputs[2452] = ~(layer0_outputs[4298]);
    assign outputs[2453] = ~(layer0_outputs[1157]);
    assign outputs[2454] = ~(layer0_outputs[5198]);
    assign outputs[2455] = (layer0_outputs[675]) ^ (layer0_outputs[136]);
    assign outputs[2456] = ~(layer0_outputs[8314]) | (layer0_outputs[7683]);
    assign outputs[2457] = layer0_outputs[3798];
    assign outputs[2458] = ~(layer0_outputs[418]) | (layer0_outputs[9432]);
    assign outputs[2459] = layer0_outputs[97];
    assign outputs[2460] = ~(layer0_outputs[641]);
    assign outputs[2461] = ~((layer0_outputs[2799]) & (layer0_outputs[789]));
    assign outputs[2462] = ~(layer0_outputs[9049]) | (layer0_outputs[7021]);
    assign outputs[2463] = ~(layer0_outputs[3651]);
    assign outputs[2464] = (layer0_outputs[7722]) ^ (layer0_outputs[4304]);
    assign outputs[2465] = (layer0_outputs[36]) & ~(layer0_outputs[446]);
    assign outputs[2466] = ~(layer0_outputs[5433]) | (layer0_outputs[9443]);
    assign outputs[2467] = ~((layer0_outputs[881]) | (layer0_outputs[5923]));
    assign outputs[2468] = layer0_outputs[2962];
    assign outputs[2469] = ~((layer0_outputs[7399]) ^ (layer0_outputs[8928]));
    assign outputs[2470] = ~((layer0_outputs[5071]) ^ (layer0_outputs[5543]));
    assign outputs[2471] = ~((layer0_outputs[6301]) ^ (layer0_outputs[9126]));
    assign outputs[2472] = layer0_outputs[8495];
    assign outputs[2473] = layer0_outputs[4928];
    assign outputs[2474] = ~((layer0_outputs[2979]) & (layer0_outputs[9554]));
    assign outputs[2475] = ~(layer0_outputs[3622]) | (layer0_outputs[6332]);
    assign outputs[2476] = ~((layer0_outputs[4345]) | (layer0_outputs[8613]));
    assign outputs[2477] = ~((layer0_outputs[5367]) ^ (layer0_outputs[8506]));
    assign outputs[2478] = ~(layer0_outputs[9775]);
    assign outputs[2479] = ~(layer0_outputs[3037]);
    assign outputs[2480] = ~((layer0_outputs[1505]) ^ (layer0_outputs[6793]));
    assign outputs[2481] = (layer0_outputs[195]) ^ (layer0_outputs[3626]);
    assign outputs[2482] = layer0_outputs[55];
    assign outputs[2483] = ~(layer0_outputs[8147]);
    assign outputs[2484] = layer0_outputs[5949];
    assign outputs[2485] = ~((layer0_outputs[7608]) ^ (layer0_outputs[4484]));
    assign outputs[2486] = ~(layer0_outputs[7241]) | (layer0_outputs[1947]);
    assign outputs[2487] = layer0_outputs[5434];
    assign outputs[2488] = (layer0_outputs[5528]) & (layer0_outputs[5993]);
    assign outputs[2489] = ~((layer0_outputs[7260]) ^ (layer0_outputs[5333]));
    assign outputs[2490] = (layer0_outputs[4055]) | (layer0_outputs[7963]);
    assign outputs[2491] = (layer0_outputs[5821]) ^ (layer0_outputs[2767]);
    assign outputs[2492] = ~(layer0_outputs[3102]);
    assign outputs[2493] = ~(layer0_outputs[5304]);
    assign outputs[2494] = ~(layer0_outputs[4046]) | (layer0_outputs[2887]);
    assign outputs[2495] = layer0_outputs[1681];
    assign outputs[2496] = (layer0_outputs[8620]) ^ (layer0_outputs[1579]);
    assign outputs[2497] = (layer0_outputs[4236]) | (layer0_outputs[7839]);
    assign outputs[2498] = ~(layer0_outputs[10142]) | (layer0_outputs[3483]);
    assign outputs[2499] = layer0_outputs[6157];
    assign outputs[2500] = ~(layer0_outputs[9351]);
    assign outputs[2501] = (layer0_outputs[5117]) | (layer0_outputs[4344]);
    assign outputs[2502] = layer0_outputs[9525];
    assign outputs[2503] = ~(layer0_outputs[5364]);
    assign outputs[2504] = (layer0_outputs[9941]) | (layer0_outputs[3838]);
    assign outputs[2505] = layer0_outputs[9039];
    assign outputs[2506] = (layer0_outputs[6669]) ^ (layer0_outputs[3621]);
    assign outputs[2507] = ~((layer0_outputs[4178]) ^ (layer0_outputs[1802]));
    assign outputs[2508] = ~(layer0_outputs[6717]) | (layer0_outputs[1356]);
    assign outputs[2509] = layer0_outputs[3706];
    assign outputs[2510] = ~(layer0_outputs[4794]) | (layer0_outputs[7491]);
    assign outputs[2511] = ~(layer0_outputs[10067]) | (layer0_outputs[6686]);
    assign outputs[2512] = ~(layer0_outputs[7300]);
    assign outputs[2513] = layer0_outputs[8450];
    assign outputs[2514] = (layer0_outputs[9007]) & ~(layer0_outputs[5406]);
    assign outputs[2515] = ~((layer0_outputs[828]) & (layer0_outputs[6151]));
    assign outputs[2516] = (layer0_outputs[6998]) | (layer0_outputs[4797]);
    assign outputs[2517] = ~((layer0_outputs[9782]) & (layer0_outputs[7343]));
    assign outputs[2518] = (layer0_outputs[6605]) & ~(layer0_outputs[783]);
    assign outputs[2519] = (layer0_outputs[4788]) & (layer0_outputs[2130]);
    assign outputs[2520] = ~(layer0_outputs[1358]);
    assign outputs[2521] = (layer0_outputs[2100]) ^ (layer0_outputs[5055]);
    assign outputs[2522] = layer0_outputs[9230];
    assign outputs[2523] = ~(layer0_outputs[595]);
    assign outputs[2524] = ~(layer0_outputs[4590]) | (layer0_outputs[9434]);
    assign outputs[2525] = layer0_outputs[5973];
    assign outputs[2526] = ~(layer0_outputs[6880]);
    assign outputs[2527] = ~(layer0_outputs[7319]);
    assign outputs[2528] = layer0_outputs[2951];
    assign outputs[2529] = ~(layer0_outputs[5048]);
    assign outputs[2530] = ~(layer0_outputs[5433]);
    assign outputs[2531] = (layer0_outputs[3957]) & ~(layer0_outputs[2670]);
    assign outputs[2532] = layer0_outputs[2215];
    assign outputs[2533] = layer0_outputs[6520];
    assign outputs[2534] = ~((layer0_outputs[122]) & (layer0_outputs[2077]));
    assign outputs[2535] = ~((layer0_outputs[7475]) ^ (layer0_outputs[1746]));
    assign outputs[2536] = (layer0_outputs[9041]) & (layer0_outputs[8748]);
    assign outputs[2537] = layer0_outputs[9219];
    assign outputs[2538] = (layer0_outputs[4844]) & ~(layer0_outputs[8519]);
    assign outputs[2539] = layer0_outputs[5668];
    assign outputs[2540] = ~(layer0_outputs[10224]) | (layer0_outputs[8019]);
    assign outputs[2541] = ~((layer0_outputs[1535]) | (layer0_outputs[9820]));
    assign outputs[2542] = layer0_outputs[5979];
    assign outputs[2543] = layer0_outputs[9795];
    assign outputs[2544] = ~((layer0_outputs[9141]) & (layer0_outputs[6139]));
    assign outputs[2545] = ~(layer0_outputs[7257]);
    assign outputs[2546] = layer0_outputs[7794];
    assign outputs[2547] = (layer0_outputs[8320]) & (layer0_outputs[704]);
    assign outputs[2548] = ~(layer0_outputs[7832]);
    assign outputs[2549] = (layer0_outputs[8927]) | (layer0_outputs[9954]);
    assign outputs[2550] = layer0_outputs[3772];
    assign outputs[2551] = ~((layer0_outputs[7894]) | (layer0_outputs[8248]));
    assign outputs[2552] = ~(layer0_outputs[7422]) | (layer0_outputs[8047]);
    assign outputs[2553] = ~((layer0_outputs[7484]) & (layer0_outputs[3707]));
    assign outputs[2554] = layer0_outputs[3079];
    assign outputs[2555] = layer0_outputs[9029];
    assign outputs[2556] = ~(layer0_outputs[8481]);
    assign outputs[2557] = layer0_outputs[8512];
    assign outputs[2558] = layer0_outputs[8159];
    assign outputs[2559] = (layer0_outputs[2787]) ^ (layer0_outputs[9546]);
    assign outputs[2560] = (layer0_outputs[1758]) ^ (layer0_outputs[2831]);
    assign outputs[2561] = ~(layer0_outputs[4453]);
    assign outputs[2562] = layer0_outputs[1031];
    assign outputs[2563] = layer0_outputs[5472];
    assign outputs[2564] = ~(layer0_outputs[3282]);
    assign outputs[2565] = layer0_outputs[606];
    assign outputs[2566] = ~(layer0_outputs[5480]);
    assign outputs[2567] = ~(layer0_outputs[8840]);
    assign outputs[2568] = ~((layer0_outputs[3689]) ^ (layer0_outputs[2339]));
    assign outputs[2569] = ~(layer0_outputs[1092]);
    assign outputs[2570] = layer0_outputs[9506];
    assign outputs[2571] = (layer0_outputs[9915]) & (layer0_outputs[4605]);
    assign outputs[2572] = (layer0_outputs[3545]) ^ (layer0_outputs[3127]);
    assign outputs[2573] = ~((layer0_outputs[1231]) ^ (layer0_outputs[1609]));
    assign outputs[2574] = (layer0_outputs[8994]) & ~(layer0_outputs[5325]);
    assign outputs[2575] = ~(layer0_outputs[7449]);
    assign outputs[2576] = layer0_outputs[2083];
    assign outputs[2577] = ~((layer0_outputs[7887]) & (layer0_outputs[3181]));
    assign outputs[2578] = ~((layer0_outputs[7026]) ^ (layer0_outputs[6177]));
    assign outputs[2579] = (layer0_outputs[237]) ^ (layer0_outputs[1985]);
    assign outputs[2580] = (layer0_outputs[2296]) ^ (layer0_outputs[1074]);
    assign outputs[2581] = ~(layer0_outputs[5761]);
    assign outputs[2582] = (layer0_outputs[2980]) | (layer0_outputs[455]);
    assign outputs[2583] = ~((layer0_outputs[5485]) ^ (layer0_outputs[10131]));
    assign outputs[2584] = ~((layer0_outputs[3413]) | (layer0_outputs[3242]));
    assign outputs[2585] = layer0_outputs[5593];
    assign outputs[2586] = ~(layer0_outputs[7363]) | (layer0_outputs[6]);
    assign outputs[2587] = ~((layer0_outputs[5514]) | (layer0_outputs[8729]));
    assign outputs[2588] = ~(layer0_outputs[9324]);
    assign outputs[2589] = layer0_outputs[6775];
    assign outputs[2590] = (layer0_outputs[4352]) ^ (layer0_outputs[3368]);
    assign outputs[2591] = ~(layer0_outputs[6344]);
    assign outputs[2592] = layer0_outputs[5249];
    assign outputs[2593] = layer0_outputs[4716];
    assign outputs[2594] = ~(layer0_outputs[3739]);
    assign outputs[2595] = (layer0_outputs[2707]) | (layer0_outputs[9602]);
    assign outputs[2596] = ~((layer0_outputs[4495]) & (layer0_outputs[10225]));
    assign outputs[2597] = (layer0_outputs[8115]) | (layer0_outputs[9282]);
    assign outputs[2598] = ~(layer0_outputs[1010]) | (layer0_outputs[2069]);
    assign outputs[2599] = ~(layer0_outputs[5836]);
    assign outputs[2600] = (layer0_outputs[9990]) ^ (layer0_outputs[8523]);
    assign outputs[2601] = ~(layer0_outputs[4781]) | (layer0_outputs[4180]);
    assign outputs[2602] = (layer0_outputs[2542]) ^ (layer0_outputs[4326]);
    assign outputs[2603] = ~(layer0_outputs[9333]);
    assign outputs[2604] = ~((layer0_outputs[7225]) ^ (layer0_outputs[9264]));
    assign outputs[2605] = layer0_outputs[5190];
    assign outputs[2606] = layer0_outputs[9428];
    assign outputs[2607] = (layer0_outputs[2884]) ^ (layer0_outputs[9004]);
    assign outputs[2608] = layer0_outputs[9984];
    assign outputs[2609] = (layer0_outputs[1277]) ^ (layer0_outputs[2975]);
    assign outputs[2610] = ~(layer0_outputs[9936]) | (layer0_outputs[2963]);
    assign outputs[2611] = (layer0_outputs[4382]) & (layer0_outputs[10086]);
    assign outputs[2612] = ~((layer0_outputs[6302]) & (layer0_outputs[7030]));
    assign outputs[2613] = ~(layer0_outputs[10061]) | (layer0_outputs[4868]);
    assign outputs[2614] = (layer0_outputs[1365]) ^ (layer0_outputs[9590]);
    assign outputs[2615] = layer0_outputs[9343];
    assign outputs[2616] = ~(layer0_outputs[2065]) | (layer0_outputs[8832]);
    assign outputs[2617] = (layer0_outputs[1592]) & ~(layer0_outputs[1502]);
    assign outputs[2618] = (layer0_outputs[5105]) & ~(layer0_outputs[653]);
    assign outputs[2619] = layer0_outputs[834];
    assign outputs[2620] = ~(layer0_outputs[3773]);
    assign outputs[2621] = layer0_outputs[5573];
    assign outputs[2622] = layer0_outputs[6298];
    assign outputs[2623] = ~((layer0_outputs[8920]) & (layer0_outputs[2805]));
    assign outputs[2624] = ~((layer0_outputs[5646]) ^ (layer0_outputs[3440]));
    assign outputs[2625] = ~(layer0_outputs[7896]);
    assign outputs[2626] = (layer0_outputs[1087]) & ~(layer0_outputs[2618]);
    assign outputs[2627] = (layer0_outputs[790]) & (layer0_outputs[1172]);
    assign outputs[2628] = layer0_outputs[5488];
    assign outputs[2629] = ~((layer0_outputs[33]) & (layer0_outputs[9778]));
    assign outputs[2630] = layer0_outputs[9466];
    assign outputs[2631] = ~((layer0_outputs[6428]) & (layer0_outputs[8146]));
    assign outputs[2632] = (layer0_outputs[9590]) ^ (layer0_outputs[6695]);
    assign outputs[2633] = ~(layer0_outputs[3064]);
    assign outputs[2634] = ~(layer0_outputs[9291]);
    assign outputs[2635] = ~(layer0_outputs[3947]);
    assign outputs[2636] = layer0_outputs[3958];
    assign outputs[2637] = ~(layer0_outputs[5448]);
    assign outputs[2638] = layer0_outputs[921];
    assign outputs[2639] = ~(layer0_outputs[6488]);
    assign outputs[2640] = layer0_outputs[3783];
    assign outputs[2641] = ~(layer0_outputs[1394]);
    assign outputs[2642] = layer0_outputs[7671];
    assign outputs[2643] = ~(layer0_outputs[4030]);
    assign outputs[2644] = ~(layer0_outputs[9946]);
    assign outputs[2645] = layer0_outputs[6904];
    assign outputs[2646] = layer0_outputs[5197];
    assign outputs[2647] = ~(layer0_outputs[4973]);
    assign outputs[2648] = layer0_outputs[10094];
    assign outputs[2649] = ~(layer0_outputs[520]);
    assign outputs[2650] = ~(layer0_outputs[6719]);
    assign outputs[2651] = (layer0_outputs[7744]) ^ (layer0_outputs[7872]);
    assign outputs[2652] = ~((layer0_outputs[4451]) | (layer0_outputs[6111]));
    assign outputs[2653] = (layer0_outputs[9872]) ^ (layer0_outputs[4170]);
    assign outputs[2654] = ~((layer0_outputs[8942]) ^ (layer0_outputs[6527]));
    assign outputs[2655] = ~(layer0_outputs[6346]);
    assign outputs[2656] = ~(layer0_outputs[3423]) | (layer0_outputs[3742]);
    assign outputs[2657] = (layer0_outputs[8526]) ^ (layer0_outputs[6703]);
    assign outputs[2658] = ~((layer0_outputs[5603]) & (layer0_outputs[6592]));
    assign outputs[2659] = ~(layer0_outputs[611]);
    assign outputs[2660] = ~(layer0_outputs[8401]);
    assign outputs[2661] = ~((layer0_outputs[10188]) ^ (layer0_outputs[4186]));
    assign outputs[2662] = ~(layer0_outputs[6970]);
    assign outputs[2663] = layer0_outputs[933];
    assign outputs[2664] = ~((layer0_outputs[8305]) ^ (layer0_outputs[2784]));
    assign outputs[2665] = ~(layer0_outputs[1983]) | (layer0_outputs[3865]);
    assign outputs[2666] = (layer0_outputs[9447]) ^ (layer0_outputs[8258]);
    assign outputs[2667] = (layer0_outputs[1543]) ^ (layer0_outputs[570]);
    assign outputs[2668] = ~(layer0_outputs[2062]);
    assign outputs[2669] = ~((layer0_outputs[5910]) & (layer0_outputs[5465]));
    assign outputs[2670] = layer0_outputs[3440];
    assign outputs[2671] = layer0_outputs[7024];
    assign outputs[2672] = layer0_outputs[1951];
    assign outputs[2673] = ~((layer0_outputs[9541]) & (layer0_outputs[3002]));
    assign outputs[2674] = ~(layer0_outputs[6772]);
    assign outputs[2675] = layer0_outputs[2895];
    assign outputs[2676] = layer0_outputs[7905];
    assign outputs[2677] = (layer0_outputs[8434]) & ~(layer0_outputs[10108]);
    assign outputs[2678] = ~((layer0_outputs[6665]) ^ (layer0_outputs[7949]));
    assign outputs[2679] = ~(layer0_outputs[7574]);
    assign outputs[2680] = (layer0_outputs[859]) ^ (layer0_outputs[2779]);
    assign outputs[2681] = layer0_outputs[4663];
    assign outputs[2682] = (layer0_outputs[8244]) ^ (layer0_outputs[9882]);
    assign outputs[2683] = layer0_outputs[824];
    assign outputs[2684] = ~(layer0_outputs[3790]);
    assign outputs[2685] = layer0_outputs[4725];
    assign outputs[2686] = (layer0_outputs[3113]) & ~(layer0_outputs[2769]);
    assign outputs[2687] = ~((layer0_outputs[3926]) & (layer0_outputs[6858]));
    assign outputs[2688] = ~(layer0_outputs[1986]);
    assign outputs[2689] = layer0_outputs[9880];
    assign outputs[2690] = ~(layer0_outputs[6160]);
    assign outputs[2691] = ~((layer0_outputs[7504]) ^ (layer0_outputs[3717]));
    assign outputs[2692] = layer0_outputs[3282];
    assign outputs[2693] = ~(layer0_outputs[6446]);
    assign outputs[2694] = ~(layer0_outputs[1771]);
    assign outputs[2695] = layer0_outputs[4221];
    assign outputs[2696] = ~((layer0_outputs[3817]) | (layer0_outputs[6827]));
    assign outputs[2697] = ~(layer0_outputs[6778]) | (layer0_outputs[3425]);
    assign outputs[2698] = ~((layer0_outputs[4302]) ^ (layer0_outputs[3304]));
    assign outputs[2699] = (layer0_outputs[3647]) ^ (layer0_outputs[4830]);
    assign outputs[2700] = ~((layer0_outputs[327]) ^ (layer0_outputs[4086]));
    assign outputs[2701] = layer0_outputs[3045];
    assign outputs[2702] = layer0_outputs[6766];
    assign outputs[2703] = ~((layer0_outputs[152]) | (layer0_outputs[2062]));
    assign outputs[2704] = (layer0_outputs[9585]) & (layer0_outputs[7755]);
    assign outputs[2705] = (layer0_outputs[2210]) ^ (layer0_outputs[2601]);
    assign outputs[2706] = (layer0_outputs[5570]) ^ (layer0_outputs[6843]);
    assign outputs[2707] = ~(layer0_outputs[2773]);
    assign outputs[2708] = ~(layer0_outputs[8562]);
    assign outputs[2709] = ~(layer0_outputs[8724]) | (layer0_outputs[7386]);
    assign outputs[2710] = ~((layer0_outputs[3532]) ^ (layer0_outputs[10053]));
    assign outputs[2711] = (layer0_outputs[5574]) | (layer0_outputs[10210]);
    assign outputs[2712] = ~(layer0_outputs[7517]);
    assign outputs[2713] = ~(layer0_outputs[573]);
    assign outputs[2714] = layer0_outputs[2217];
    assign outputs[2715] = ~(layer0_outputs[8380]) | (layer0_outputs[10122]);
    assign outputs[2716] = ~((layer0_outputs[1006]) ^ (layer0_outputs[7450]));
    assign outputs[2717] = ~(layer0_outputs[8095]) | (layer0_outputs[4772]);
    assign outputs[2718] = (layer0_outputs[8746]) | (layer0_outputs[7474]);
    assign outputs[2719] = ~(layer0_outputs[5794]) | (layer0_outputs[3000]);
    assign outputs[2720] = layer0_outputs[5815];
    assign outputs[2721] = ~((layer0_outputs[9390]) ^ (layer0_outputs[2843]));
    assign outputs[2722] = (layer0_outputs[4337]) & (layer0_outputs[8736]);
    assign outputs[2723] = layer0_outputs[8805];
    assign outputs[2724] = ~((layer0_outputs[7105]) ^ (layer0_outputs[1884]));
    assign outputs[2725] = ~(layer0_outputs[1644]);
    assign outputs[2726] = ~(layer0_outputs[7033]);
    assign outputs[2727] = (layer0_outputs[480]) | (layer0_outputs[9616]);
    assign outputs[2728] = layer0_outputs[3028];
    assign outputs[2729] = ~(layer0_outputs[9639]) | (layer0_outputs[1469]);
    assign outputs[2730] = ~(layer0_outputs[3178]);
    assign outputs[2731] = layer0_outputs[507];
    assign outputs[2732] = ~(layer0_outputs[1983]) | (layer0_outputs[6499]);
    assign outputs[2733] = ~(layer0_outputs[4802]);
    assign outputs[2734] = ~(layer0_outputs[8213]);
    assign outputs[2735] = ~((layer0_outputs[636]) & (layer0_outputs[1020]));
    assign outputs[2736] = ~(layer0_outputs[5804]);
    assign outputs[2737] = (layer0_outputs[2317]) ^ (layer0_outputs[1212]);
    assign outputs[2738] = (layer0_outputs[3799]) & ~(layer0_outputs[576]);
    assign outputs[2739] = ~(layer0_outputs[8107]);
    assign outputs[2740] = layer0_outputs[9837];
    assign outputs[2741] = (layer0_outputs[309]) | (layer0_outputs[5795]);
    assign outputs[2742] = (layer0_outputs[8461]) & ~(layer0_outputs[4532]);
    assign outputs[2743] = ~(layer0_outputs[3862]);
    assign outputs[2744] = ~((layer0_outputs[5253]) & (layer0_outputs[5861]));
    assign outputs[2745] = ~(layer0_outputs[5440]);
    assign outputs[2746] = (layer0_outputs[9058]) ^ (layer0_outputs[875]);
    assign outputs[2747] = ~(layer0_outputs[2257]);
    assign outputs[2748] = layer0_outputs[1683];
    assign outputs[2749] = (layer0_outputs[1440]) ^ (layer0_outputs[4916]);
    assign outputs[2750] = ~(layer0_outputs[4563]) | (layer0_outputs[763]);
    assign outputs[2751] = ~((layer0_outputs[4337]) & (layer0_outputs[1596]));
    assign outputs[2752] = ~(layer0_outputs[6132]);
    assign outputs[2753] = ~(layer0_outputs[2483]);
    assign outputs[2754] = ~(layer0_outputs[8207]) | (layer0_outputs[5529]);
    assign outputs[2755] = (layer0_outputs[3388]) ^ (layer0_outputs[1317]);
    assign outputs[2756] = ~((layer0_outputs[2912]) | (layer0_outputs[4848]));
    assign outputs[2757] = ~(layer0_outputs[7573]);
    assign outputs[2758] = (layer0_outputs[10225]) ^ (layer0_outputs[4196]);
    assign outputs[2759] = (layer0_outputs[3502]) ^ (layer0_outputs[5250]);
    assign outputs[2760] = (layer0_outputs[8340]) ^ (layer0_outputs[6979]);
    assign outputs[2761] = ~((layer0_outputs[7946]) & (layer0_outputs[1452]));
    assign outputs[2762] = ~((layer0_outputs[7616]) ^ (layer0_outputs[9365]));
    assign outputs[2763] = layer0_outputs[5789];
    assign outputs[2764] = layer0_outputs[7677];
    assign outputs[2765] = layer0_outputs[2732];
    assign outputs[2766] = ~(layer0_outputs[2938]);
    assign outputs[2767] = ~(layer0_outputs[4633]) | (layer0_outputs[335]);
    assign outputs[2768] = ~(layer0_outputs[8243]);
    assign outputs[2769] = ~((layer0_outputs[1307]) & (layer0_outputs[2629]));
    assign outputs[2770] = ~(layer0_outputs[4196]);
    assign outputs[2771] = ~((layer0_outputs[5725]) ^ (layer0_outputs[6153]));
    assign outputs[2772] = ~(layer0_outputs[6815]) | (layer0_outputs[6234]);
    assign outputs[2773] = (layer0_outputs[6551]) & (layer0_outputs[7651]);
    assign outputs[2774] = (layer0_outputs[4373]) & ~(layer0_outputs[2998]);
    assign outputs[2775] = (layer0_outputs[337]) & ~(layer0_outputs[8818]);
    assign outputs[2776] = 1'b1;
    assign outputs[2777] = layer0_outputs[2089];
    assign outputs[2778] = layer0_outputs[5641];
    assign outputs[2779] = ~(layer0_outputs[4321]);
    assign outputs[2780] = (layer0_outputs[5748]) ^ (layer0_outputs[9015]);
    assign outputs[2781] = ~(layer0_outputs[9847]);
    assign outputs[2782] = (layer0_outputs[2324]) & (layer0_outputs[3861]);
    assign outputs[2783] = ~(layer0_outputs[8059]) | (layer0_outputs[6696]);
    assign outputs[2784] = (layer0_outputs[7630]) ^ (layer0_outputs[6176]);
    assign outputs[2785] = ~((layer0_outputs[815]) ^ (layer0_outputs[7752]));
    assign outputs[2786] = ~(layer0_outputs[3762]) | (layer0_outputs[2385]);
    assign outputs[2787] = ~(layer0_outputs[8774]) | (layer0_outputs[9253]);
    assign outputs[2788] = ~((layer0_outputs[2796]) ^ (layer0_outputs[5749]));
    assign outputs[2789] = ~(layer0_outputs[4762]);
    assign outputs[2790] = layer0_outputs[358];
    assign outputs[2791] = layer0_outputs[8189];
    assign outputs[2792] = ~(layer0_outputs[7385]);
    assign outputs[2793] = (layer0_outputs[7261]) ^ (layer0_outputs[115]);
    assign outputs[2794] = ~(layer0_outputs[3341]);
    assign outputs[2795] = (layer0_outputs[6630]) & (layer0_outputs[3531]);
    assign outputs[2796] = ~((layer0_outputs[7909]) & (layer0_outputs[7696]));
    assign outputs[2797] = ~(layer0_outputs[6139]);
    assign outputs[2798] = layer0_outputs[6494];
    assign outputs[2799] = ~(layer0_outputs[6837]);
    assign outputs[2800] = layer0_outputs[8708];
    assign outputs[2801] = layer0_outputs[9923];
    assign outputs[2802] = (layer0_outputs[4595]) & ~(layer0_outputs[2660]);
    assign outputs[2803] = ~(layer0_outputs[4847]) | (layer0_outputs[6018]);
    assign outputs[2804] = (layer0_outputs[5499]) ^ (layer0_outputs[939]);
    assign outputs[2805] = ~(layer0_outputs[10077]);
    assign outputs[2806] = (layer0_outputs[2794]) & (layer0_outputs[7711]);
    assign outputs[2807] = (layer0_outputs[9674]) ^ (layer0_outputs[6310]);
    assign outputs[2808] = layer0_outputs[8521];
    assign outputs[2809] = (layer0_outputs[4167]) & ~(layer0_outputs[6111]);
    assign outputs[2810] = ~(layer0_outputs[6390]);
    assign outputs[2811] = ~(layer0_outputs[5482]) | (layer0_outputs[950]);
    assign outputs[2812] = ~((layer0_outputs[2896]) ^ (layer0_outputs[4255]));
    assign outputs[2813] = ~(layer0_outputs[6011]);
    assign outputs[2814] = ~((layer0_outputs[6653]) ^ (layer0_outputs[6093]));
    assign outputs[2815] = ~(layer0_outputs[4799]) | (layer0_outputs[9180]);
    assign outputs[2816] = (layer0_outputs[3450]) & ~(layer0_outputs[2716]);
    assign outputs[2817] = ~(layer0_outputs[6652]);
    assign outputs[2818] = layer0_outputs[7637];
    assign outputs[2819] = ~((layer0_outputs[7913]) ^ (layer0_outputs[4040]));
    assign outputs[2820] = layer0_outputs[3357];
    assign outputs[2821] = (layer0_outputs[6343]) ^ (layer0_outputs[8367]);
    assign outputs[2822] = (layer0_outputs[2396]) ^ (layer0_outputs[9442]);
    assign outputs[2823] = (layer0_outputs[2022]) & ~(layer0_outputs[3094]);
    assign outputs[2824] = ~(layer0_outputs[6845]);
    assign outputs[2825] = ~(layer0_outputs[6709]);
    assign outputs[2826] = layer0_outputs[4435];
    assign outputs[2827] = (layer0_outputs[3925]) ^ (layer0_outputs[5942]);
    assign outputs[2828] = layer0_outputs[6824];
    assign outputs[2829] = ~(layer0_outputs[5025]) | (layer0_outputs[1943]);
    assign outputs[2830] = (layer0_outputs[2696]) & ~(layer0_outputs[6612]);
    assign outputs[2831] = (layer0_outputs[2202]) & ~(layer0_outputs[3354]);
    assign outputs[2832] = layer0_outputs[1843];
    assign outputs[2833] = ~((layer0_outputs[6061]) & (layer0_outputs[271]));
    assign outputs[2834] = (layer0_outputs[5594]) ^ (layer0_outputs[6382]);
    assign outputs[2835] = (layer0_outputs[9696]) & ~(layer0_outputs[2313]);
    assign outputs[2836] = layer0_outputs[4060];
    assign outputs[2837] = ~(layer0_outputs[4938]);
    assign outputs[2838] = ~((layer0_outputs[2211]) ^ (layer0_outputs[5786]));
    assign outputs[2839] = ~(layer0_outputs[6562]);
    assign outputs[2840] = ~((layer0_outputs[1377]) ^ (layer0_outputs[7291]));
    assign outputs[2841] = ~((layer0_outputs[7668]) | (layer0_outputs[5594]));
    assign outputs[2842] = ~(layer0_outputs[9033]);
    assign outputs[2843] = layer0_outputs[824];
    assign outputs[2844] = (layer0_outputs[1282]) & ~(layer0_outputs[2693]);
    assign outputs[2845] = ~(layer0_outputs[9879]);
    assign outputs[2846] = (layer0_outputs[3573]) | (layer0_outputs[6016]);
    assign outputs[2847] = layer0_outputs[5418];
    assign outputs[2848] = ~(layer0_outputs[5710]) | (layer0_outputs[7456]);
    assign outputs[2849] = ~(layer0_outputs[1158]);
    assign outputs[2850] = ~((layer0_outputs[5471]) ^ (layer0_outputs[9507]));
    assign outputs[2851] = layer0_outputs[9870];
    assign outputs[2852] = (layer0_outputs[2879]) ^ (layer0_outputs[6154]);
    assign outputs[2853] = 1'b1;
    assign outputs[2854] = ~(layer0_outputs[9157]);
    assign outputs[2855] = ~(layer0_outputs[10197]);
    assign outputs[2856] = layer0_outputs[1414];
    assign outputs[2857] = ~((layer0_outputs[394]) ^ (layer0_outputs[1066]));
    assign outputs[2858] = layer0_outputs[10052];
    assign outputs[2859] = ~((layer0_outputs[6384]) ^ (layer0_outputs[1866]));
    assign outputs[2860] = ~((layer0_outputs[0]) & (layer0_outputs[2756]));
    assign outputs[2861] = ~(layer0_outputs[9060]);
    assign outputs[2862] = layer0_outputs[5503];
    assign outputs[2863] = ~((layer0_outputs[2560]) | (layer0_outputs[8020]));
    assign outputs[2864] = ~((layer0_outputs[1807]) ^ (layer0_outputs[5186]));
    assign outputs[2865] = layer0_outputs[4441];
    assign outputs[2866] = layer0_outputs[2471];
    assign outputs[2867] = ~(layer0_outputs[9797]) | (layer0_outputs[10107]);
    assign outputs[2868] = (layer0_outputs[6409]) & (layer0_outputs[3770]);
    assign outputs[2869] = layer0_outputs[8930];
    assign outputs[2870] = ~(layer0_outputs[1001]);
    assign outputs[2871] = (layer0_outputs[7111]) | (layer0_outputs[991]);
    assign outputs[2872] = ~((layer0_outputs[3479]) & (layer0_outputs[2400]));
    assign outputs[2873] = ~(layer0_outputs[1013]) | (layer0_outputs[6037]);
    assign outputs[2874] = (layer0_outputs[588]) ^ (layer0_outputs[4120]);
    assign outputs[2875] = (layer0_outputs[8863]) | (layer0_outputs[979]);
    assign outputs[2876] = ~(layer0_outputs[9292]) | (layer0_outputs[9683]);
    assign outputs[2877] = ~((layer0_outputs[3404]) ^ (layer0_outputs[6784]));
    assign outputs[2878] = layer0_outputs[6473];
    assign outputs[2879] = ~((layer0_outputs[7719]) ^ (layer0_outputs[4301]));
    assign outputs[2880] = ~(layer0_outputs[2575]) | (layer0_outputs[1820]);
    assign outputs[2881] = (layer0_outputs[4056]) & ~(layer0_outputs[2058]);
    assign outputs[2882] = ~((layer0_outputs[6609]) & (layer0_outputs[180]));
    assign outputs[2883] = ~(layer0_outputs[10227]);
    assign outputs[2884] = ~((layer0_outputs[6978]) ^ (layer0_outputs[7047]));
    assign outputs[2885] = layer0_outputs[1683];
    assign outputs[2886] = ~(layer0_outputs[149]);
    assign outputs[2887] = ~(layer0_outputs[1552]);
    assign outputs[2888] = layer0_outputs[4584];
    assign outputs[2889] = ~((layer0_outputs[5373]) ^ (layer0_outputs[6893]));
    assign outputs[2890] = (layer0_outputs[1779]) | (layer0_outputs[5894]);
    assign outputs[2891] = (layer0_outputs[6275]) ^ (layer0_outputs[5412]);
    assign outputs[2892] = ~((layer0_outputs[2139]) ^ (layer0_outputs[8357]));
    assign outputs[2893] = ~(layer0_outputs[3181]) | (layer0_outputs[2538]);
    assign outputs[2894] = (layer0_outputs[7004]) ^ (layer0_outputs[2533]);
    assign outputs[2895] = layer0_outputs[3448];
    assign outputs[2896] = ~(layer0_outputs[4678]);
    assign outputs[2897] = ~((layer0_outputs[564]) ^ (layer0_outputs[8771]));
    assign outputs[2898] = (layer0_outputs[119]) ^ (layer0_outputs[4941]);
    assign outputs[2899] = layer0_outputs[3806];
    assign outputs[2900] = ~(layer0_outputs[8489]);
    assign outputs[2901] = (layer0_outputs[5790]) & ~(layer0_outputs[6574]);
    assign outputs[2902] = layer0_outputs[402];
    assign outputs[2903] = layer0_outputs[6467];
    assign outputs[2904] = (layer0_outputs[9304]) | (layer0_outputs[3123]);
    assign outputs[2905] = ~(layer0_outputs[273]) | (layer0_outputs[3735]);
    assign outputs[2906] = (layer0_outputs[469]) & ~(layer0_outputs[9821]);
    assign outputs[2907] = (layer0_outputs[2963]) | (layer0_outputs[1263]);
    assign outputs[2908] = (layer0_outputs[8485]) & ~(layer0_outputs[9319]);
    assign outputs[2909] = ~((layer0_outputs[10109]) ^ (layer0_outputs[7014]));
    assign outputs[2910] = (layer0_outputs[1514]) | (layer0_outputs[7399]);
    assign outputs[2911] = ~(layer0_outputs[6770]) | (layer0_outputs[574]);
    assign outputs[2912] = layer0_outputs[5331];
    assign outputs[2913] = ~(layer0_outputs[7943]) | (layer0_outputs[10202]);
    assign outputs[2914] = layer0_outputs[7914];
    assign outputs[2915] = layer0_outputs[2447];
    assign outputs[2916] = (layer0_outputs[869]) ^ (layer0_outputs[1813]);
    assign outputs[2917] = ~(layer0_outputs[1797]) | (layer0_outputs[1808]);
    assign outputs[2918] = ~((layer0_outputs[9476]) | (layer0_outputs[5393]));
    assign outputs[2919] = ~(layer0_outputs[5169]);
    assign outputs[2920] = (layer0_outputs[7980]) ^ (layer0_outputs[508]);
    assign outputs[2921] = ~(layer0_outputs[338]) | (layer0_outputs[1405]);
    assign outputs[2922] = ~(layer0_outputs[8107]);
    assign outputs[2923] = (layer0_outputs[2074]) ^ (layer0_outputs[7658]);
    assign outputs[2924] = (layer0_outputs[8876]) ^ (layer0_outputs[6078]);
    assign outputs[2925] = ~(layer0_outputs[3485]) | (layer0_outputs[1775]);
    assign outputs[2926] = layer0_outputs[10010];
    assign outputs[2927] = ~((layer0_outputs[6219]) ^ (layer0_outputs[219]));
    assign outputs[2928] = ~(layer0_outputs[174]);
    assign outputs[2929] = ~(layer0_outputs[5905]);
    assign outputs[2930] = ~((layer0_outputs[8541]) | (layer0_outputs[1099]));
    assign outputs[2931] = (layer0_outputs[538]) & ~(layer0_outputs[7262]);
    assign outputs[2932] = ~(layer0_outputs[6704]);
    assign outputs[2933] = layer0_outputs[8099];
    assign outputs[2934] = layer0_outputs[8984];
    assign outputs[2935] = ~((layer0_outputs[129]) | (layer0_outputs[697]));
    assign outputs[2936] = ~(layer0_outputs[6642]);
    assign outputs[2937] = layer0_outputs[2722];
    assign outputs[2938] = ~((layer0_outputs[1554]) | (layer0_outputs[5261]));
    assign outputs[2939] = (layer0_outputs[2209]) ^ (layer0_outputs[125]);
    assign outputs[2940] = (layer0_outputs[4258]) & (layer0_outputs[6171]);
    assign outputs[2941] = (layer0_outputs[8339]) ^ (layer0_outputs[3516]);
    assign outputs[2942] = ~((layer0_outputs[4710]) ^ (layer0_outputs[2472]));
    assign outputs[2943] = (layer0_outputs[10239]) ^ (layer0_outputs[8170]);
    assign outputs[2944] = (layer0_outputs[8215]) | (layer0_outputs[3147]);
    assign outputs[2945] = ~(layer0_outputs[4277]);
    assign outputs[2946] = (layer0_outputs[734]) & (layer0_outputs[8855]);
    assign outputs[2947] = (layer0_outputs[10044]) & ~(layer0_outputs[1494]);
    assign outputs[2948] = ~(layer0_outputs[2291]) | (layer0_outputs[2822]);
    assign outputs[2949] = (layer0_outputs[8440]) & (layer0_outputs[7813]);
    assign outputs[2950] = (layer0_outputs[2399]) & ~(layer0_outputs[2605]);
    assign outputs[2951] = (layer0_outputs[3669]) & (layer0_outputs[2530]);
    assign outputs[2952] = ~((layer0_outputs[4668]) & (layer0_outputs[6683]));
    assign outputs[2953] = layer0_outputs[6090];
    assign outputs[2954] = layer0_outputs[91];
    assign outputs[2955] = ~(layer0_outputs[793]);
    assign outputs[2956] = ~(layer0_outputs[582]);
    assign outputs[2957] = (layer0_outputs[4303]) ^ (layer0_outputs[6296]);
    assign outputs[2958] = ~(layer0_outputs[7878]);
    assign outputs[2959] = ~((layer0_outputs[6981]) & (layer0_outputs[4917]));
    assign outputs[2960] = ~((layer0_outputs[974]) ^ (layer0_outputs[6628]));
    assign outputs[2961] = (layer0_outputs[3257]) & ~(layer0_outputs[4508]);
    assign outputs[2962] = 1'b1;
    assign outputs[2963] = layer0_outputs[6423];
    assign outputs[2964] = (layer0_outputs[6408]) & ~(layer0_outputs[7959]);
    assign outputs[2965] = ~(layer0_outputs[5078]) | (layer0_outputs[9789]);
    assign outputs[2966] = layer0_outputs[7120];
    assign outputs[2967] = ~(layer0_outputs[3610]);
    assign outputs[2968] = ~(layer0_outputs[7888]);
    assign outputs[2969] = layer0_outputs[4242];
    assign outputs[2970] = layer0_outputs[8462];
    assign outputs[2971] = ~(layer0_outputs[4944]);
    assign outputs[2972] = (layer0_outputs[7759]) & ~(layer0_outputs[9043]);
    assign outputs[2973] = ~(layer0_outputs[8055]);
    assign outputs[2974] = ~(layer0_outputs[3879]) | (layer0_outputs[3990]);
    assign outputs[2975] = ~((layer0_outputs[5463]) ^ (layer0_outputs[8879]));
    assign outputs[2976] = (layer0_outputs[628]) ^ (layer0_outputs[1468]);
    assign outputs[2977] = layer0_outputs[5914];
    assign outputs[2978] = ~(layer0_outputs[696]);
    assign outputs[2979] = ~(layer0_outputs[2647]);
    assign outputs[2980] = ~((layer0_outputs[7693]) & (layer0_outputs[8628]));
    assign outputs[2981] = ~((layer0_outputs[3263]) & (layer0_outputs[5419]));
    assign outputs[2982] = layer0_outputs[530];
    assign outputs[2983] = (layer0_outputs[2070]) | (layer0_outputs[2978]);
    assign outputs[2984] = ~(layer0_outputs[9673]);
    assign outputs[2985] = ~(layer0_outputs[7678]) | (layer0_outputs[10213]);
    assign outputs[2986] = (layer0_outputs[3836]) | (layer0_outputs[6924]);
    assign outputs[2987] = ~((layer0_outputs[5708]) | (layer0_outputs[8480]));
    assign outputs[2988] = ~(layer0_outputs[8385]);
    assign outputs[2989] = (layer0_outputs[4521]) | (layer0_outputs[3406]);
    assign outputs[2990] = (layer0_outputs[10221]) & ~(layer0_outputs[9117]);
    assign outputs[2991] = ~((layer0_outputs[8251]) | (layer0_outputs[4874]));
    assign outputs[2992] = ~((layer0_outputs[2318]) | (layer0_outputs[7107]));
    assign outputs[2993] = layer0_outputs[7546];
    assign outputs[2994] = ~(layer0_outputs[9764]) | (layer0_outputs[3115]);
    assign outputs[2995] = (layer0_outputs[8171]) & ~(layer0_outputs[2917]);
    assign outputs[2996] = ~((layer0_outputs[1110]) ^ (layer0_outputs[9577]));
    assign outputs[2997] = ~((layer0_outputs[425]) | (layer0_outputs[983]));
    assign outputs[2998] = layer0_outputs[6502];
    assign outputs[2999] = (layer0_outputs[1092]) ^ (layer0_outputs[5705]);
    assign outputs[3000] = (layer0_outputs[9602]) & (layer0_outputs[2981]);
    assign outputs[3001] = layer0_outputs[5519];
    assign outputs[3002] = layer0_outputs[4031];
    assign outputs[3003] = layer0_outputs[1481];
    assign outputs[3004] = ~(layer0_outputs[145]);
    assign outputs[3005] = layer0_outputs[2310];
    assign outputs[3006] = ~((layer0_outputs[1324]) ^ (layer0_outputs[9645]));
    assign outputs[3007] = (layer0_outputs[3924]) & ~(layer0_outputs[6180]);
    assign outputs[3008] = (layer0_outputs[3636]) ^ (layer0_outputs[6632]);
    assign outputs[3009] = (layer0_outputs[5916]) & ~(layer0_outputs[10132]);
    assign outputs[3010] = (layer0_outputs[8076]) ^ (layer0_outputs[10113]);
    assign outputs[3011] = layer0_outputs[5337];
    assign outputs[3012] = ~((layer0_outputs[3358]) & (layer0_outputs[3166]));
    assign outputs[3013] = (layer0_outputs[2303]) | (layer0_outputs[3156]);
    assign outputs[3014] = (layer0_outputs[885]) | (layer0_outputs[1678]);
    assign outputs[3015] = (layer0_outputs[927]) & ~(layer0_outputs[4327]);
    assign outputs[3016] = layer0_outputs[5561];
    assign outputs[3017] = ~(layer0_outputs[4592]);
    assign outputs[3018] = (layer0_outputs[8346]) ^ (layer0_outputs[5250]);
    assign outputs[3019] = (layer0_outputs[8128]) & ~(layer0_outputs[6950]);
    assign outputs[3020] = ~((layer0_outputs[2474]) ^ (layer0_outputs[8881]));
    assign outputs[3021] = ~((layer0_outputs[1944]) | (layer0_outputs[3497]));
    assign outputs[3022] = (layer0_outputs[4727]) ^ (layer0_outputs[4346]);
    assign outputs[3023] = ~(layer0_outputs[386]);
    assign outputs[3024] = ~(layer0_outputs[4278]);
    assign outputs[3025] = layer0_outputs[1667];
    assign outputs[3026] = layer0_outputs[5365];
    assign outputs[3027] = (layer0_outputs[7996]) ^ (layer0_outputs[1052]);
    assign outputs[3028] = (layer0_outputs[6689]) | (layer0_outputs[6185]);
    assign outputs[3029] = ~((layer0_outputs[6385]) ^ (layer0_outputs[2684]));
    assign outputs[3030] = ~(layer0_outputs[1147]) | (layer0_outputs[779]);
    assign outputs[3031] = ~((layer0_outputs[3579]) ^ (layer0_outputs[8970]));
    assign outputs[3032] = (layer0_outputs[356]) ^ (layer0_outputs[3395]);
    assign outputs[3033] = (layer0_outputs[4004]) ^ (layer0_outputs[1763]);
    assign outputs[3034] = (layer0_outputs[1509]) ^ (layer0_outputs[9089]);
    assign outputs[3035] = ~(layer0_outputs[8776]) | (layer0_outputs[9747]);
    assign outputs[3036] = (layer0_outputs[4354]) ^ (layer0_outputs[1942]);
    assign outputs[3037] = ~((layer0_outputs[2448]) | (layer0_outputs[9441]));
    assign outputs[3038] = ~((layer0_outputs[7325]) & (layer0_outputs[3243]));
    assign outputs[3039] = ~(layer0_outputs[9528]) | (layer0_outputs[6009]);
    assign outputs[3040] = ~((layer0_outputs[6715]) & (layer0_outputs[8747]));
    assign outputs[3041] = ~((layer0_outputs[9464]) & (layer0_outputs[4590]));
    assign outputs[3042] = ~(layer0_outputs[6057]);
    assign outputs[3043] = ~(layer0_outputs[3096]) | (layer0_outputs[3576]);
    assign outputs[3044] = layer0_outputs[1320];
    assign outputs[3045] = 1'b1;
    assign outputs[3046] = layer0_outputs[1720];
    assign outputs[3047] = layer0_outputs[7638];
    assign outputs[3048] = ~(layer0_outputs[8894]);
    assign outputs[3049] = layer0_outputs[4061];
    assign outputs[3050] = (layer0_outputs[6583]) & ~(layer0_outputs[370]);
    assign outputs[3051] = layer0_outputs[1187];
    assign outputs[3052] = ~((layer0_outputs[6955]) | (layer0_outputs[3721]));
    assign outputs[3053] = ~((layer0_outputs[8554]) ^ (layer0_outputs[9115]));
    assign outputs[3054] = ~(layer0_outputs[9872]);
    assign outputs[3055] = ~(layer0_outputs[4837]);
    assign outputs[3056] = ~(layer0_outputs[53]);
    assign outputs[3057] = ~(layer0_outputs[7596]) | (layer0_outputs[9424]);
    assign outputs[3058] = ~((layer0_outputs[9752]) | (layer0_outputs[7135]));
    assign outputs[3059] = ~(layer0_outputs[5629]);
    assign outputs[3060] = ~((layer0_outputs[2629]) & (layer0_outputs[8957]));
    assign outputs[3061] = (layer0_outputs[9776]) ^ (layer0_outputs[1209]);
    assign outputs[3062] = ~((layer0_outputs[4796]) ^ (layer0_outputs[9806]));
    assign outputs[3063] = layer0_outputs[3928];
    assign outputs[3064] = (layer0_outputs[1017]) ^ (layer0_outputs[1174]);
    assign outputs[3065] = ~(layer0_outputs[9360]);
    assign outputs[3066] = ~((layer0_outputs[9989]) ^ (layer0_outputs[2898]));
    assign outputs[3067] = ~(layer0_outputs[3030]);
    assign outputs[3068] = ~((layer0_outputs[652]) & (layer0_outputs[9543]));
    assign outputs[3069] = (layer0_outputs[4625]) ^ (layer0_outputs[8564]);
    assign outputs[3070] = ~((layer0_outputs[1828]) & (layer0_outputs[10146]));
    assign outputs[3071] = ~((layer0_outputs[10066]) ^ (layer0_outputs[8909]));
    assign outputs[3072] = ~((layer0_outputs[633]) ^ (layer0_outputs[6644]));
    assign outputs[3073] = ~((layer0_outputs[6946]) & (layer0_outputs[10217]));
    assign outputs[3074] = ~(layer0_outputs[4622]);
    assign outputs[3075] = ~((layer0_outputs[7952]) | (layer0_outputs[3759]));
    assign outputs[3076] = (layer0_outputs[9546]) | (layer0_outputs[9163]);
    assign outputs[3077] = ~((layer0_outputs[6798]) & (layer0_outputs[6736]));
    assign outputs[3078] = ~(layer0_outputs[9743]);
    assign outputs[3079] = layer0_outputs[997];
    assign outputs[3080] = ~((layer0_outputs[6268]) ^ (layer0_outputs[4193]));
    assign outputs[3081] = ~(layer0_outputs[1903]) | (layer0_outputs[5667]);
    assign outputs[3082] = ~(layer0_outputs[2412]) | (layer0_outputs[9365]);
    assign outputs[3083] = layer0_outputs[9468];
    assign outputs[3084] = (layer0_outputs[8058]) & ~(layer0_outputs[6463]);
    assign outputs[3085] = ~((layer0_outputs[7032]) ^ (layer0_outputs[2219]));
    assign outputs[3086] = ~((layer0_outputs[9134]) ^ (layer0_outputs[5290]));
    assign outputs[3087] = layer0_outputs[5977];
    assign outputs[3088] = ~(layer0_outputs[5653]) | (layer0_outputs[653]);
    assign outputs[3089] = ~(layer0_outputs[8731]) | (layer0_outputs[3190]);
    assign outputs[3090] = ~(layer0_outputs[3794]);
    assign outputs[3091] = (layer0_outputs[2473]) ^ (layer0_outputs[2670]);
    assign outputs[3092] = ~(layer0_outputs[1361]);
    assign outputs[3093] = (layer0_outputs[6948]) ^ (layer0_outputs[8029]);
    assign outputs[3094] = ~(layer0_outputs[9835]);
    assign outputs[3095] = ~(layer0_outputs[1907]);
    assign outputs[3096] = ~(layer0_outputs[3490]);
    assign outputs[3097] = layer0_outputs[2441];
    assign outputs[3098] = ~((layer0_outputs[8116]) & (layer0_outputs[8709]));
    assign outputs[3099] = layer0_outputs[5149];
    assign outputs[3100] = ~(layer0_outputs[2947]);
    assign outputs[3101] = layer0_outputs[5829];
    assign outputs[3102] = ~((layer0_outputs[7013]) | (layer0_outputs[2331]));
    assign outputs[3103] = (layer0_outputs[1485]) ^ (layer0_outputs[5590]);
    assign outputs[3104] = layer0_outputs[2014];
    assign outputs[3105] = ~((layer0_outputs[7012]) ^ (layer0_outputs[4206]));
    assign outputs[3106] = layer0_outputs[3315];
    assign outputs[3107] = layer0_outputs[4693];
    assign outputs[3108] = ~(layer0_outputs[6550]);
    assign outputs[3109] = ~((layer0_outputs[2834]) ^ (layer0_outputs[5898]));
    assign outputs[3110] = layer0_outputs[6011];
    assign outputs[3111] = ~(layer0_outputs[8432]);
    assign outputs[3112] = (layer0_outputs[7181]) ^ (layer0_outputs[316]);
    assign outputs[3113] = layer0_outputs[9822];
    assign outputs[3114] = layer0_outputs[8538];
    assign outputs[3115] = ~(layer0_outputs[2195]);
    assign outputs[3116] = ~(layer0_outputs[901]);
    assign outputs[3117] = layer0_outputs[9871];
    assign outputs[3118] = (layer0_outputs[413]) ^ (layer0_outputs[6224]);
    assign outputs[3119] = ~(layer0_outputs[3136]);
    assign outputs[3120] = ~((layer0_outputs[261]) ^ (layer0_outputs[56]));
    assign outputs[3121] = layer0_outputs[9861];
    assign outputs[3122] = (layer0_outputs[3309]) ^ (layer0_outputs[6018]);
    assign outputs[3123] = (layer0_outputs[5328]) | (layer0_outputs[3015]);
    assign outputs[3124] = ~((layer0_outputs[7003]) ^ (layer0_outputs[2926]));
    assign outputs[3125] = ~(layer0_outputs[3434]) | (layer0_outputs[3704]);
    assign outputs[3126] = layer0_outputs[6091];
    assign outputs[3127] = (layer0_outputs[4869]) & (layer0_outputs[7955]);
    assign outputs[3128] = ~(layer0_outputs[1450]);
    assign outputs[3129] = ~((layer0_outputs[5885]) & (layer0_outputs[7525]));
    assign outputs[3130] = ~(layer0_outputs[8347]);
    assign outputs[3131] = ~(layer0_outputs[1318]);
    assign outputs[3132] = (layer0_outputs[4814]) ^ (layer0_outputs[9287]);
    assign outputs[3133] = ~((layer0_outputs[9809]) ^ (layer0_outputs[1105]));
    assign outputs[3134] = ~((layer0_outputs[7453]) ^ (layer0_outputs[518]));
    assign outputs[3135] = ~((layer0_outputs[4979]) ^ (layer0_outputs[5725]));
    assign outputs[3136] = ~(layer0_outputs[543]);
    assign outputs[3137] = (layer0_outputs[9011]) & (layer0_outputs[8031]);
    assign outputs[3138] = layer0_outputs[5047];
    assign outputs[3139] = ~((layer0_outputs[10002]) ^ (layer0_outputs[10080]));
    assign outputs[3140] = (layer0_outputs[7802]) | (layer0_outputs[3715]);
    assign outputs[3141] = ~(layer0_outputs[4712]);
    assign outputs[3142] = (layer0_outputs[2490]) ^ (layer0_outputs[4078]);
    assign outputs[3143] = ~(layer0_outputs[9651]);
    assign outputs[3144] = (layer0_outputs[6626]) & ~(layer0_outputs[9392]);
    assign outputs[3145] = ~(layer0_outputs[9876]) | (layer0_outputs[9117]);
    assign outputs[3146] = layer0_outputs[2113];
    assign outputs[3147] = layer0_outputs[900];
    assign outputs[3148] = ~(layer0_outputs[8130]);
    assign outputs[3149] = ~(layer0_outputs[4522]);
    assign outputs[3150] = layer0_outputs[9732];
    assign outputs[3151] = (layer0_outputs[2386]) ^ (layer0_outputs[1082]);
    assign outputs[3152] = (layer0_outputs[5938]) ^ (layer0_outputs[10200]);
    assign outputs[3153] = ~((layer0_outputs[9245]) | (layer0_outputs[6433]));
    assign outputs[3154] = ~((layer0_outputs[9755]) ^ (layer0_outputs[10149]));
    assign outputs[3155] = (layer0_outputs[8231]) ^ (layer0_outputs[5194]);
    assign outputs[3156] = layer0_outputs[6245];
    assign outputs[3157] = ~(layer0_outputs[8947]) | (layer0_outputs[6064]);
    assign outputs[3158] = ~(layer0_outputs[7301]);
    assign outputs[3159] = (layer0_outputs[7344]) ^ (layer0_outputs[2410]);
    assign outputs[3160] = ~(layer0_outputs[6465]);
    assign outputs[3161] = ~(layer0_outputs[7006]);
    assign outputs[3162] = layer0_outputs[4907];
    assign outputs[3163] = ~(layer0_outputs[4390]);
    assign outputs[3164] = ~(layer0_outputs[7366]) | (layer0_outputs[8088]);
    assign outputs[3165] = ~(layer0_outputs[4843]) | (layer0_outputs[725]);
    assign outputs[3166] = layer0_outputs[7976];
    assign outputs[3167] = (layer0_outputs[9577]) ^ (layer0_outputs[4181]);
    assign outputs[3168] = ~((layer0_outputs[3122]) ^ (layer0_outputs[4254]));
    assign outputs[3169] = (layer0_outputs[6315]) & (layer0_outputs[9581]);
    assign outputs[3170] = layer0_outputs[2150];
    assign outputs[3171] = ~(layer0_outputs[8420]);
    assign outputs[3172] = ~((layer0_outputs[4800]) ^ (layer0_outputs[6575]));
    assign outputs[3173] = ~(layer0_outputs[9394]) | (layer0_outputs[9052]);
    assign outputs[3174] = ~((layer0_outputs[8289]) | (layer0_outputs[8955]));
    assign outputs[3175] = ~(layer0_outputs[1190]) | (layer0_outputs[2857]);
    assign outputs[3176] = (layer0_outputs[8778]) & ~(layer0_outputs[4813]);
    assign outputs[3177] = layer0_outputs[4670];
    assign outputs[3178] = ~(layer0_outputs[4539]);
    assign outputs[3179] = (layer0_outputs[4394]) ^ (layer0_outputs[2673]);
    assign outputs[3180] = ~(layer0_outputs[1265]);
    assign outputs[3181] = (layer0_outputs[4955]) | (layer0_outputs[9790]);
    assign outputs[3182] = ~((layer0_outputs[3276]) & (layer0_outputs[5737]));
    assign outputs[3183] = ~(layer0_outputs[1028]) | (layer0_outputs[9990]);
    assign outputs[3184] = ~(layer0_outputs[545]);
    assign outputs[3185] = ~(layer0_outputs[7431]);
    assign outputs[3186] = layer0_outputs[2747];
    assign outputs[3187] = ~((layer0_outputs[5222]) ^ (layer0_outputs[3678]));
    assign outputs[3188] = ~(layer0_outputs[1114]);
    assign outputs[3189] = ~((layer0_outputs[4159]) & (layer0_outputs[81]));
    assign outputs[3190] = ~(layer0_outputs[4002]);
    assign outputs[3191] = ~((layer0_outputs[2162]) ^ (layer0_outputs[6780]));
    assign outputs[3192] = (layer0_outputs[7521]) ^ (layer0_outputs[261]);
    assign outputs[3193] = ~((layer0_outputs[7131]) | (layer0_outputs[6329]));
    assign outputs[3194] = layer0_outputs[8882];
    assign outputs[3195] = ~(layer0_outputs[1330]) | (layer0_outputs[1476]);
    assign outputs[3196] = layer0_outputs[9011];
    assign outputs[3197] = ~(layer0_outputs[2278]) | (layer0_outputs[3200]);
    assign outputs[3198] = ~(layer0_outputs[5052]);
    assign outputs[3199] = ~((layer0_outputs[3915]) ^ (layer0_outputs[8974]));
    assign outputs[3200] = layer0_outputs[6140];
    assign outputs[3201] = ~((layer0_outputs[2647]) | (layer0_outputs[7782]));
    assign outputs[3202] = ~(layer0_outputs[2560]);
    assign outputs[3203] = ~(layer0_outputs[5074]);
    assign outputs[3204] = ~((layer0_outputs[2448]) ^ (layer0_outputs[6900]));
    assign outputs[3205] = ~(layer0_outputs[9325]);
    assign outputs[3206] = layer0_outputs[1106];
    assign outputs[3207] = (layer0_outputs[1937]) & ~(layer0_outputs[8704]);
    assign outputs[3208] = ~((layer0_outputs[5880]) & (layer0_outputs[7051]));
    assign outputs[3209] = ~(layer0_outputs[7078]) | (layer0_outputs[1517]);
    assign outputs[3210] = ~(layer0_outputs[8525]);
    assign outputs[3211] = (layer0_outputs[2840]) & ~(layer0_outputs[5052]);
    assign outputs[3212] = ~(layer0_outputs[2720]) | (layer0_outputs[5562]);
    assign outputs[3213] = layer0_outputs[3092];
    assign outputs[3214] = ~(layer0_outputs[2921]);
    assign outputs[3215] = ~((layer0_outputs[3619]) ^ (layer0_outputs[9303]));
    assign outputs[3216] = (layer0_outputs[4134]) & ~(layer0_outputs[3362]);
    assign outputs[3217] = layer0_outputs[7033];
    assign outputs[3218] = ~(layer0_outputs[9340]);
    assign outputs[3219] = ~((layer0_outputs[6909]) ^ (layer0_outputs[4399]));
    assign outputs[3220] = ~(layer0_outputs[8102]);
    assign outputs[3221] = layer0_outputs[1321];
    assign outputs[3222] = (layer0_outputs[8549]) ^ (layer0_outputs[6416]);
    assign outputs[3223] = (layer0_outputs[4726]) | (layer0_outputs[6560]);
    assign outputs[3224] = (layer0_outputs[5494]) ^ (layer0_outputs[1104]);
    assign outputs[3225] = layer0_outputs[3569];
    assign outputs[3226] = ~((layer0_outputs[3642]) | (layer0_outputs[7633]));
    assign outputs[3227] = ~(layer0_outputs[5056]);
    assign outputs[3228] = ~((layer0_outputs[9909]) ^ (layer0_outputs[4517]));
    assign outputs[3229] = ~(layer0_outputs[639]);
    assign outputs[3230] = ~((layer0_outputs[5484]) & (layer0_outputs[1534]));
    assign outputs[3231] = ~(layer0_outputs[4883]) | (layer0_outputs[955]);
    assign outputs[3232] = layer0_outputs[1226];
    assign outputs[3233] = ~((layer0_outputs[7378]) ^ (layer0_outputs[1634]));
    assign outputs[3234] = ~(layer0_outputs[3759]);
    assign outputs[3235] = (layer0_outputs[1029]) ^ (layer0_outputs[1829]);
    assign outputs[3236] = (layer0_outputs[9041]) & ~(layer0_outputs[5527]);
    assign outputs[3237] = ~(layer0_outputs[3405]) | (layer0_outputs[4484]);
    assign outputs[3238] = (layer0_outputs[6106]) ^ (layer0_outputs[3025]);
    assign outputs[3239] = layer0_outputs[7104];
    assign outputs[3240] = ~((layer0_outputs[1974]) & (layer0_outputs[8139]));
    assign outputs[3241] = layer0_outputs[4463];
    assign outputs[3242] = ~(layer0_outputs[4825]) | (layer0_outputs[2631]);
    assign outputs[3243] = layer0_outputs[9998];
    assign outputs[3244] = ~((layer0_outputs[1804]) & (layer0_outputs[7190]));
    assign outputs[3245] = (layer0_outputs[1259]) ^ (layer0_outputs[4122]);
    assign outputs[3246] = (layer0_outputs[4145]) ^ (layer0_outputs[2559]);
    assign outputs[3247] = ~((layer0_outputs[9632]) ^ (layer0_outputs[949]));
    assign outputs[3248] = ~(layer0_outputs[3808]);
    assign outputs[3249] = (layer0_outputs[9631]) & ~(layer0_outputs[3123]);
    assign outputs[3250] = (layer0_outputs[4583]) | (layer0_outputs[9128]);
    assign outputs[3251] = layer0_outputs[5333];
    assign outputs[3252] = layer0_outputs[5605];
    assign outputs[3253] = ~((layer0_outputs[3495]) ^ (layer0_outputs[5227]));
    assign outputs[3254] = layer0_outputs[5182];
    assign outputs[3255] = ~(layer0_outputs[2096]) | (layer0_outputs[4217]);
    assign outputs[3256] = ~(layer0_outputs[5532]);
    assign outputs[3257] = (layer0_outputs[8891]) | (layer0_outputs[6386]);
    assign outputs[3258] = (layer0_outputs[113]) & (layer0_outputs[2979]);
    assign outputs[3259] = (layer0_outputs[3001]) | (layer0_outputs[3792]);
    assign outputs[3260] = (layer0_outputs[2203]) & ~(layer0_outputs[4336]);
    assign outputs[3261] = ~(layer0_outputs[6716]);
    assign outputs[3262] = ~(layer0_outputs[3119]) | (layer0_outputs[9560]);
    assign outputs[3263] = (layer0_outputs[4582]) ^ (layer0_outputs[5842]);
    assign outputs[3264] = layer0_outputs[3435];
    assign outputs[3265] = ~(layer0_outputs[5080]);
    assign outputs[3266] = layer0_outputs[9987];
    assign outputs[3267] = (layer0_outputs[1669]) & ~(layer0_outputs[5924]);
    assign outputs[3268] = layer0_outputs[7054];
    assign outputs[3269] = (layer0_outputs[39]) & (layer0_outputs[4721]);
    assign outputs[3270] = ~(layer0_outputs[10209]);
    assign outputs[3271] = ~(layer0_outputs[2268]);
    assign outputs[3272] = layer0_outputs[1833];
    assign outputs[3273] = layer0_outputs[5771];
    assign outputs[3274] = (layer0_outputs[8056]) ^ (layer0_outputs[6866]);
    assign outputs[3275] = (layer0_outputs[2315]) ^ (layer0_outputs[7442]);
    assign outputs[3276] = ~((layer0_outputs[2068]) ^ (layer0_outputs[1988]));
    assign outputs[3277] = ~(layer0_outputs[2531]) | (layer0_outputs[6817]);
    assign outputs[3278] = 1'b1;
    assign outputs[3279] = layer0_outputs[4604];
    assign outputs[3280] = ~(layer0_outputs[8795]);
    assign outputs[3281] = ~((layer0_outputs[2305]) & (layer0_outputs[1454]));
    assign outputs[3282] = layer0_outputs[1349];
    assign outputs[3283] = layer0_outputs[1340];
    assign outputs[3284] = (layer0_outputs[8991]) | (layer0_outputs[3727]);
    assign outputs[3285] = layer0_outputs[5358];
    assign outputs[3286] = ~(layer0_outputs[5976]);
    assign outputs[3287] = (layer0_outputs[6144]) | (layer0_outputs[7270]);
    assign outputs[3288] = ~((layer0_outputs[1094]) ^ (layer0_outputs[5213]));
    assign outputs[3289] = layer0_outputs[89];
    assign outputs[3290] = ~(layer0_outputs[8609]) | (layer0_outputs[9849]);
    assign outputs[3291] = layer0_outputs[5479];
    assign outputs[3292] = layer0_outputs[6792];
    assign outputs[3293] = (layer0_outputs[1277]) & ~(layer0_outputs[5893]);
    assign outputs[3294] = layer0_outputs[2674];
    assign outputs[3295] = ~((layer0_outputs[6740]) & (layer0_outputs[4431]));
    assign outputs[3296] = ~((layer0_outputs[5854]) & (layer0_outputs[226]));
    assign outputs[3297] = layer0_outputs[2033];
    assign outputs[3298] = layer0_outputs[4216];
    assign outputs[3299] = (layer0_outputs[9411]) & ~(layer0_outputs[8454]);
    assign outputs[3300] = ~((layer0_outputs[7944]) ^ (layer0_outputs[9489]));
    assign outputs[3301] = ~((layer0_outputs[7195]) | (layer0_outputs[1424]));
    assign outputs[3302] = (layer0_outputs[9170]) | (layer0_outputs[1651]);
    assign outputs[3303] = layer0_outputs[4088];
    assign outputs[3304] = layer0_outputs[9256];
    assign outputs[3305] = ~(layer0_outputs[5411]);
    assign outputs[3306] = layer0_outputs[2392];
    assign outputs[3307] = ~(layer0_outputs[4403]);
    assign outputs[3308] = ~((layer0_outputs[8940]) ^ (layer0_outputs[5545]));
    assign outputs[3309] = layer0_outputs[153];
    assign outputs[3310] = ~(layer0_outputs[8715]) | (layer0_outputs[5416]);
    assign outputs[3311] = (layer0_outputs[3645]) | (layer0_outputs[957]);
    assign outputs[3312] = ~(layer0_outputs[8433]) | (layer0_outputs[1733]);
    assign outputs[3313] = (layer0_outputs[467]) & ~(layer0_outputs[4972]);
    assign outputs[3314] = layer0_outputs[3757];
    assign outputs[3315] = ~((layer0_outputs[383]) ^ (layer0_outputs[145]));
    assign outputs[3316] = ~(layer0_outputs[2379]);
    assign outputs[3317] = layer0_outputs[7476];
    assign outputs[3318] = ~(layer0_outputs[2603]) | (layer0_outputs[8872]);
    assign outputs[3319] = layer0_outputs[8199];
    assign outputs[3320] = ~(layer0_outputs[3893]) | (layer0_outputs[588]);
    assign outputs[3321] = (layer0_outputs[215]) ^ (layer0_outputs[2713]);
    assign outputs[3322] = ~(layer0_outputs[4671]);
    assign outputs[3323] = ~(layer0_outputs[10117]);
    assign outputs[3324] = layer0_outputs[7548];
    assign outputs[3325] = ~(layer0_outputs[7356]);
    assign outputs[3326] = ~(layer0_outputs[1782]);
    assign outputs[3327] = (layer0_outputs[3876]) & ~(layer0_outputs[3183]);
    assign outputs[3328] = ~(layer0_outputs[5775]);
    assign outputs[3329] = (layer0_outputs[6435]) & ~(layer0_outputs[5225]);
    assign outputs[3330] = ~(layer0_outputs[1710]);
    assign outputs[3331] = ~((layer0_outputs[5074]) & (layer0_outputs[9848]));
    assign outputs[3332] = (layer0_outputs[1206]) & ~(layer0_outputs[1879]);
    assign outputs[3333] = ~(layer0_outputs[982]);
    assign outputs[3334] = ~(layer0_outputs[8167]);
    assign outputs[3335] = (layer0_outputs[9406]) & ~(layer0_outputs[182]);
    assign outputs[3336] = ~((layer0_outputs[3520]) & (layer0_outputs[4665]));
    assign outputs[3337] = ~((layer0_outputs[1351]) ^ (layer0_outputs[541]));
    assign outputs[3338] = layer0_outputs[5826];
    assign outputs[3339] = 1'b1;
    assign outputs[3340] = layer0_outputs[8888];
    assign outputs[3341] = ~(layer0_outputs[10015]);
    assign outputs[3342] = (layer0_outputs[4163]) ^ (layer0_outputs[917]);
    assign outputs[3343] = ~(layer0_outputs[8418]);
    assign outputs[3344] = ~((layer0_outputs[3847]) ^ (layer0_outputs[1007]));
    assign outputs[3345] = layer0_outputs[6765];
    assign outputs[3346] = ~(layer0_outputs[9300]) | (layer0_outputs[1723]);
    assign outputs[3347] = ~(layer0_outputs[5120]);
    assign outputs[3348] = layer0_outputs[4123];
    assign outputs[3349] = ~((layer0_outputs[7377]) & (layer0_outputs[9715]));
    assign outputs[3350] = layer0_outputs[6556];
    assign outputs[3351] = ~(layer0_outputs[5404]);
    assign outputs[3352] = ~(layer0_outputs[9401]) | (layer0_outputs[2727]);
    assign outputs[3353] = ~((layer0_outputs[5812]) ^ (layer0_outputs[1770]));
    assign outputs[3354] = ~(layer0_outputs[2792]) | (layer0_outputs[6155]);
    assign outputs[3355] = ~(layer0_outputs[3446]);
    assign outputs[3356] = (layer0_outputs[6161]) & ~(layer0_outputs[2564]);
    assign outputs[3357] = (layer0_outputs[4132]) ^ (layer0_outputs[3145]);
    assign outputs[3358] = (layer0_outputs[8557]) | (layer0_outputs[78]);
    assign outputs[3359] = (layer0_outputs[4468]) & ~(layer0_outputs[1130]);
    assign outputs[3360] = ~(layer0_outputs[1217]) | (layer0_outputs[6767]);
    assign outputs[3361] = ~(layer0_outputs[1843]);
    assign outputs[3362] = layer0_outputs[5806];
    assign outputs[3363] = (layer0_outputs[6338]) & ~(layer0_outputs[2015]);
    assign outputs[3364] = (layer0_outputs[1439]) ^ (layer0_outputs[362]);
    assign outputs[3365] = ~(layer0_outputs[6896]);
    assign outputs[3366] = ~(layer0_outputs[4641]);
    assign outputs[3367] = (layer0_outputs[4324]) ^ (layer0_outputs[4316]);
    assign outputs[3368] = (layer0_outputs[7931]) ^ (layer0_outputs[3802]);
    assign outputs[3369] = layer0_outputs[7692];
    assign outputs[3370] = layer0_outputs[4904];
    assign outputs[3371] = ~((layer0_outputs[7035]) ^ (layer0_outputs[4093]));
    assign outputs[3372] = ~((layer0_outputs[6805]) ^ (layer0_outputs[10106]));
    assign outputs[3373] = ~(layer0_outputs[1326]) | (layer0_outputs[8673]);
    assign outputs[3374] = (layer0_outputs[7088]) ^ (layer0_outputs[1941]);
    assign outputs[3375] = ~(layer0_outputs[235]);
    assign outputs[3376] = ~((layer0_outputs[8722]) ^ (layer0_outputs[9301]));
    assign outputs[3377] = (layer0_outputs[76]) ^ (layer0_outputs[4085]);
    assign outputs[3378] = layer0_outputs[5635];
    assign outputs[3379] = ~((layer0_outputs[451]) ^ (layer0_outputs[1817]));
    assign outputs[3380] = ~(layer0_outputs[9091]);
    assign outputs[3381] = (layer0_outputs[10107]) | (layer0_outputs[3186]);
    assign outputs[3382] = ~(layer0_outputs[1215]) | (layer0_outputs[2679]);
    assign outputs[3383] = (layer0_outputs[3266]) ^ (layer0_outputs[3746]);
    assign outputs[3384] = ~((layer0_outputs[1969]) & (layer0_outputs[1956]));
    assign outputs[3385] = (layer0_outputs[4631]) & ~(layer0_outputs[8412]);
    assign outputs[3386] = (layer0_outputs[2090]) & (layer0_outputs[7865]);
    assign outputs[3387] = ~(layer0_outputs[9647]);
    assign outputs[3388] = ~((layer0_outputs[6569]) ^ (layer0_outputs[5882]));
    assign outputs[3389] = ~(layer0_outputs[7822]) | (layer0_outputs[5962]);
    assign outputs[3390] = (layer0_outputs[8619]) & (layer0_outputs[5905]);
    assign outputs[3391] = layer0_outputs[303];
    assign outputs[3392] = ~((layer0_outputs[2906]) | (layer0_outputs[6835]));
    assign outputs[3393] = (layer0_outputs[3555]) ^ (layer0_outputs[6365]);
    assign outputs[3394] = ~(layer0_outputs[2824]) | (layer0_outputs[4451]);
    assign outputs[3395] = ~((layer0_outputs[8711]) & (layer0_outputs[254]));
    assign outputs[3396] = ~(layer0_outputs[2735]) | (layer0_outputs[8867]);
    assign outputs[3397] = ~((layer0_outputs[10038]) & (layer0_outputs[6207]));
    assign outputs[3398] = (layer0_outputs[2013]) & ~(layer0_outputs[1329]);
    assign outputs[3399] = (layer0_outputs[2286]) ^ (layer0_outputs[7392]);
    assign outputs[3400] = ~((layer0_outputs[3347]) ^ (layer0_outputs[9272]));
    assign outputs[3401] = (layer0_outputs[417]) & ~(layer0_outputs[2785]);
    assign outputs[3402] = ~((layer0_outputs[384]) ^ (layer0_outputs[2066]));
    assign outputs[3403] = ~(layer0_outputs[645]);
    assign outputs[3404] = (layer0_outputs[4137]) & (layer0_outputs[4988]);
    assign outputs[3405] = (layer0_outputs[158]) ^ (layer0_outputs[6110]);
    assign outputs[3406] = layer0_outputs[6972];
    assign outputs[3407] = (layer0_outputs[6118]) & ~(layer0_outputs[6210]);
    assign outputs[3408] = ~((layer0_outputs[6599]) ^ (layer0_outputs[8533]));
    assign outputs[3409] = ~(layer0_outputs[3480]) | (layer0_outputs[9105]);
    assign outputs[3410] = 1'b1;
    assign outputs[3411] = ~(layer0_outputs[496]);
    assign outputs[3412] = layer0_outputs[4854];
    assign outputs[3413] = layer0_outputs[6049];
    assign outputs[3414] = ~((layer0_outputs[9458]) ^ (layer0_outputs[1448]));
    assign outputs[3415] = (layer0_outputs[3403]) | (layer0_outputs[679]);
    assign outputs[3416] = (layer0_outputs[9098]) ^ (layer0_outputs[8630]);
    assign outputs[3417] = (layer0_outputs[2241]) ^ (layer0_outputs[1181]);
    assign outputs[3418] = (layer0_outputs[7618]) & ~(layer0_outputs[8129]);
    assign outputs[3419] = (layer0_outputs[8633]) | (layer0_outputs[3605]);
    assign outputs[3420] = ~((layer0_outputs[9101]) ^ (layer0_outputs[1635]));
    assign outputs[3421] = (layer0_outputs[1002]) ^ (layer0_outputs[9720]);
    assign outputs[3422] = layer0_outputs[1682];
    assign outputs[3423] = ~(layer0_outputs[7890]);
    assign outputs[3424] = ~((layer0_outputs[8535]) | (layer0_outputs[3482]));
    assign outputs[3425] = (layer0_outputs[5322]) & ~(layer0_outputs[2649]);
    assign outputs[3426] = ~((layer0_outputs[9094]) | (layer0_outputs[1790]));
    assign outputs[3427] = layer0_outputs[9748];
    assign outputs[3428] = ~(layer0_outputs[8694]);
    assign outputs[3429] = ~(layer0_outputs[986]);
    assign outputs[3430] = ~(layer0_outputs[4509]) | (layer0_outputs[9580]);
    assign outputs[3431] = ~(layer0_outputs[7338]) | (layer0_outputs[5162]);
    assign outputs[3432] = (layer0_outputs[286]) ^ (layer0_outputs[1016]);
    assign outputs[3433] = ~(layer0_outputs[7890]);
    assign outputs[3434] = ~((layer0_outputs[250]) ^ (layer0_outputs[200]));
    assign outputs[3435] = ~(layer0_outputs[6926]);
    assign outputs[3436] = layer0_outputs[5230];
    assign outputs[3437] = layer0_outputs[6918];
    assign outputs[3438] = (layer0_outputs[6525]) & (layer0_outputs[4312]);
    assign outputs[3439] = layer0_outputs[8052];
    assign outputs[3440] = (layer0_outputs[8560]) ^ (layer0_outputs[2254]);
    assign outputs[3441] = ~((layer0_outputs[9526]) & (layer0_outputs[8731]));
    assign outputs[3442] = layer0_outputs[7745];
    assign outputs[3443] = (layer0_outputs[6807]) & ~(layer0_outputs[6339]);
    assign outputs[3444] = (layer0_outputs[8058]) ^ (layer0_outputs[7715]);
    assign outputs[3445] = (layer0_outputs[7134]) ^ (layer0_outputs[6899]);
    assign outputs[3446] = ~(layer0_outputs[4379]);
    assign outputs[3447] = ~(layer0_outputs[5265]);
    assign outputs[3448] = ~(layer0_outputs[5196]);
    assign outputs[3449] = ~(layer0_outputs[8149]);
    assign outputs[3450] = ~(layer0_outputs[8172]);
    assign outputs[3451] = (layer0_outputs[1506]) ^ (layer0_outputs[4109]);
    assign outputs[3452] = layer0_outputs[5762];
    assign outputs[3453] = ~(layer0_outputs[1221]);
    assign outputs[3454] = ~(layer0_outputs[3244]);
    assign outputs[3455] = (layer0_outputs[10079]) ^ (layer0_outputs[2410]);
    assign outputs[3456] = ~(layer0_outputs[5432]);
    assign outputs[3457] = (layer0_outputs[127]) ^ (layer0_outputs[5284]);
    assign outputs[3458] = layer0_outputs[2764];
    assign outputs[3459] = layer0_outputs[5954];
    assign outputs[3460] = ~(layer0_outputs[8893]);
    assign outputs[3461] = ~(layer0_outputs[3237]);
    assign outputs[3462] = layer0_outputs[3932];
    assign outputs[3463] = ~((layer0_outputs[3392]) ^ (layer0_outputs[2863]));
    assign outputs[3464] = ~(layer0_outputs[5485]);
    assign outputs[3465] = ~((layer0_outputs[2097]) ^ (layer0_outputs[9259]));
    assign outputs[3466] = (layer0_outputs[6137]) & ~(layer0_outputs[8016]);
    assign outputs[3467] = ~(layer0_outputs[722]);
    assign outputs[3468] = (layer0_outputs[7147]) & ~(layer0_outputs[4233]);
    assign outputs[3469] = ~(layer0_outputs[2458]) | (layer0_outputs[2350]);
    assign outputs[3470] = layer0_outputs[5788];
    assign outputs[3471] = layer0_outputs[1305];
    assign outputs[3472] = (layer0_outputs[5454]) ^ (layer0_outputs[7285]);
    assign outputs[3473] = ~(layer0_outputs[8862]) | (layer0_outputs[3886]);
    assign outputs[3474] = ~((layer0_outputs[1617]) ^ (layer0_outputs[10217]));
    assign outputs[3475] = (layer0_outputs[5714]) & (layer0_outputs[8257]);
    assign outputs[3476] = (layer0_outputs[8617]) & (layer0_outputs[1898]);
    assign outputs[3477] = ~((layer0_outputs[4366]) ^ (layer0_outputs[2930]));
    assign outputs[3478] = ~((layer0_outputs[6166]) | (layer0_outputs[5344]));
    assign outputs[3479] = (layer0_outputs[4010]) | (layer0_outputs[887]);
    assign outputs[3480] = layer0_outputs[1884];
    assign outputs[3481] = ~(layer0_outputs[4445]);
    assign outputs[3482] = (layer0_outputs[7917]) ^ (layer0_outputs[8256]);
    assign outputs[3483] = layer0_outputs[4915];
    assign outputs[3484] = layer0_outputs[6590];
    assign outputs[3485] = ~((layer0_outputs[6178]) ^ (layer0_outputs[8103]));
    assign outputs[3486] = (layer0_outputs[1426]) ^ (layer0_outputs[3710]);
    assign outputs[3487] = layer0_outputs[9887];
    assign outputs[3488] = ~((layer0_outputs[4320]) & (layer0_outputs[3155]));
    assign outputs[3489] = (layer0_outputs[9660]) ^ (layer0_outputs[2940]);
    assign outputs[3490] = ~((layer0_outputs[8848]) | (layer0_outputs[9755]));
    assign outputs[3491] = ~(layer0_outputs[5175]) | (layer0_outputs[5662]);
    assign outputs[3492] = ~(layer0_outputs[3465]);
    assign outputs[3493] = ~((layer0_outputs[2265]) ^ (layer0_outputs[7431]));
    assign outputs[3494] = layer0_outputs[3814];
    assign outputs[3495] = ~(layer0_outputs[7466]);
    assign outputs[3496] = (layer0_outputs[3132]) ^ (layer0_outputs[6643]);
    assign outputs[3497] = ~(layer0_outputs[7084]) | (layer0_outputs[6673]);
    assign outputs[3498] = (layer0_outputs[1248]) | (layer0_outputs[5305]);
    assign outputs[3499] = layer0_outputs[1355];
    assign outputs[3500] = layer0_outputs[1997];
    assign outputs[3501] = (layer0_outputs[7009]) | (layer0_outputs[7718]);
    assign outputs[3502] = layer0_outputs[3285];
    assign outputs[3503] = layer0_outputs[4730];
    assign outputs[3504] = (layer0_outputs[9588]) ^ (layer0_outputs[5212]);
    assign outputs[3505] = (layer0_outputs[5903]) & ~(layer0_outputs[3832]);
    assign outputs[3506] = (layer0_outputs[6098]) & ~(layer0_outputs[4093]);
    assign outputs[3507] = ~(layer0_outputs[3871]);
    assign outputs[3508] = ~(layer0_outputs[5487]);
    assign outputs[3509] = layer0_outputs[1963];
    assign outputs[3510] = layer0_outputs[3699];
    assign outputs[3511] = ~(layer0_outputs[2395]);
    assign outputs[3512] = ~((layer0_outputs[891]) & (layer0_outputs[6833]));
    assign outputs[3513] = (layer0_outputs[6619]) & ~(layer0_outputs[1953]);
    assign outputs[3514] = (layer0_outputs[8816]) ^ (layer0_outputs[7048]);
    assign outputs[3515] = layer0_outputs[4987];
    assign outputs[3516] = layer0_outputs[10239];
    assign outputs[3517] = ~(layer0_outputs[196]) | (layer0_outputs[3980]);
    assign outputs[3518] = ~((layer0_outputs[1437]) ^ (layer0_outputs[6656]));
    assign outputs[3519] = layer0_outputs[5427];
    assign outputs[3520] = (layer0_outputs[5835]) ^ (layer0_outputs[3195]);
    assign outputs[3521] = ~((layer0_outputs[829]) & (layer0_outputs[1577]));
    assign outputs[3522] = layer0_outputs[3262];
    assign outputs[3523] = ~(layer0_outputs[9842]) | (layer0_outputs[2374]);
    assign outputs[3524] = ~(layer0_outputs[724]);
    assign outputs[3525] = ~(layer0_outputs[524]);
    assign outputs[3526] = ~(layer0_outputs[8691]) | (layer0_outputs[7617]);
    assign outputs[3527] = ~(layer0_outputs[3762]) | (layer0_outputs[254]);
    assign outputs[3528] = ~((layer0_outputs[2194]) ^ (layer0_outputs[3072]));
    assign outputs[3529] = (layer0_outputs[6038]) ^ (layer0_outputs[894]);
    assign outputs[3530] = ~((layer0_outputs[4974]) | (layer0_outputs[2268]));
    assign outputs[3531] = layer0_outputs[8782];
    assign outputs[3532] = ~(layer0_outputs[1976]);
    assign outputs[3533] = 1'b1;
    assign outputs[3534] = layer0_outputs[8188];
    assign outputs[3535] = ~((layer0_outputs[8119]) ^ (layer0_outputs[91]));
    assign outputs[3536] = ~((layer0_outputs[1613]) ^ (layer0_outputs[893]));
    assign outputs[3537] = (layer0_outputs[6357]) | (layer0_outputs[5061]);
    assign outputs[3538] = layer0_outputs[3215];
    assign outputs[3539] = layer0_outputs[2326];
    assign outputs[3540] = layer0_outputs[5600];
    assign outputs[3541] = (layer0_outputs[6121]) & (layer0_outputs[2952]);
    assign outputs[3542] = ~(layer0_outputs[8167]) | (layer0_outputs[9253]);
    assign outputs[3543] = (layer0_outputs[1470]) & ~(layer0_outputs[9682]);
    assign outputs[3544] = layer0_outputs[290];
    assign outputs[3545] = ~(layer0_outputs[415]);
    assign outputs[3546] = layer0_outputs[5909];
    assign outputs[3547] = (layer0_outputs[586]) ^ (layer0_outputs[1932]);
    assign outputs[3548] = ~(layer0_outputs[7647]);
    assign outputs[3549] = layer0_outputs[5090];
    assign outputs[3550] = ~(layer0_outputs[7624]);
    assign outputs[3551] = ~((layer0_outputs[7064]) ^ (layer0_outputs[6598]));
    assign outputs[3552] = layer0_outputs[4187];
    assign outputs[3553] = layer0_outputs[8688];
    assign outputs[3554] = 1'b0;
    assign outputs[3555] = ~((layer0_outputs[7782]) ^ (layer0_outputs[2738]));
    assign outputs[3556] = (layer0_outputs[9364]) ^ (layer0_outputs[5753]);
    assign outputs[3557] = 1'b1;
    assign outputs[3558] = layer0_outputs[1520];
    assign outputs[3559] = (layer0_outputs[7461]) & (layer0_outputs[1747]);
    assign outputs[3560] = (layer0_outputs[9674]) | (layer0_outputs[2405]);
    assign outputs[3561] = layer0_outputs[5602];
    assign outputs[3562] = (layer0_outputs[648]) & ~(layer0_outputs[4711]);
    assign outputs[3563] = (layer0_outputs[7205]) ^ (layer0_outputs[2242]);
    assign outputs[3564] = layer0_outputs[8285];
    assign outputs[3565] = ~((layer0_outputs[3972]) ^ (layer0_outputs[9926]));
    assign outputs[3566] = layer0_outputs[8085];
    assign outputs[3567] = ~(layer0_outputs[661]);
    assign outputs[3568] = (layer0_outputs[7626]) | (layer0_outputs[7883]);
    assign outputs[3569] = ~(layer0_outputs[4748]);
    assign outputs[3570] = ~((layer0_outputs[5371]) | (layer0_outputs[3945]));
    assign outputs[3571] = layer0_outputs[2639];
    assign outputs[3572] = ~((layer0_outputs[9209]) | (layer0_outputs[7420]));
    assign outputs[3573] = ~((layer0_outputs[5067]) ^ (layer0_outputs[2864]));
    assign outputs[3574] = layer0_outputs[4094];
    assign outputs[3575] = (layer0_outputs[3743]) & ~(layer0_outputs[2748]);
    assign outputs[3576] = (layer0_outputs[5713]) ^ (layer0_outputs[9204]);
    assign outputs[3577] = (layer0_outputs[2235]) & ~(layer0_outputs[461]);
    assign outputs[3578] = layer0_outputs[8822];
    assign outputs[3579] = ~((layer0_outputs[7812]) ^ (layer0_outputs[9176]));
    assign outputs[3580] = layer0_outputs[2120];
    assign outputs[3581] = (layer0_outputs[7828]) | (layer0_outputs[9148]);
    assign outputs[3582] = ~(layer0_outputs[5146]) | (layer0_outputs[9600]);
    assign outputs[3583] = layer0_outputs[4602];
    assign outputs[3584] = layer0_outputs[8614];
    assign outputs[3585] = ~(layer0_outputs[4285]);
    assign outputs[3586] = ~(layer0_outputs[2571]);
    assign outputs[3587] = layer0_outputs[1491];
    assign outputs[3588] = (layer0_outputs[6765]) | (layer0_outputs[9505]);
    assign outputs[3589] = ~((layer0_outputs[7575]) ^ (layer0_outputs[3047]));
    assign outputs[3590] = ~(layer0_outputs[448]) | (layer0_outputs[9759]);
    assign outputs[3591] = ~((layer0_outputs[3106]) ^ (layer0_outputs[8584]));
    assign outputs[3592] = ~(layer0_outputs[719]);
    assign outputs[3593] = ~(layer0_outputs[2185]);
    assign outputs[3594] = (layer0_outputs[3377]) | (layer0_outputs[8079]);
    assign outputs[3595] = ~(layer0_outputs[5793]);
    assign outputs[3596] = layer0_outputs[7801];
    assign outputs[3597] = layer0_outputs[2147];
    assign outputs[3598] = (layer0_outputs[246]) ^ (layer0_outputs[8835]);
    assign outputs[3599] = ~(layer0_outputs[27]) | (layer0_outputs[1381]);
    assign outputs[3600] = ~(layer0_outputs[2817]);
    assign outputs[3601] = ~(layer0_outputs[5519]);
    assign outputs[3602] = (layer0_outputs[8165]) & ~(layer0_outputs[3811]);
    assign outputs[3603] = ~((layer0_outputs[414]) ^ (layer0_outputs[6612]));
    assign outputs[3604] = (layer0_outputs[6217]) & (layer0_outputs[7246]);
    assign outputs[3605] = ~(layer0_outputs[543]) | (layer0_outputs[2566]);
    assign outputs[3606] = ~(layer0_outputs[5578]);
    assign outputs[3607] = layer0_outputs[6757];
    assign outputs[3608] = layer0_outputs[7677];
    assign outputs[3609] = (layer0_outputs[25]) ^ (layer0_outputs[3939]);
    assign outputs[3610] = ~(layer0_outputs[6877]);
    assign outputs[3611] = ~((layer0_outputs[3741]) ^ (layer0_outputs[4333]));
    assign outputs[3612] = ~(layer0_outputs[1449]) | (layer0_outputs[9830]);
    assign outputs[3613] = ~(layer0_outputs[2293]) | (layer0_outputs[726]);
    assign outputs[3614] = ~(layer0_outputs[422]);
    assign outputs[3615] = ~((layer0_outputs[6418]) ^ (layer0_outputs[7689]));
    assign outputs[3616] = ~((layer0_outputs[9868]) & (layer0_outputs[8230]));
    assign outputs[3617] = (layer0_outputs[6100]) & ~(layer0_outputs[8110]);
    assign outputs[3618] = ~((layer0_outputs[4689]) ^ (layer0_outputs[1153]));
    assign outputs[3619] = ~(layer0_outputs[1546]);
    assign outputs[3620] = layer0_outputs[10045];
    assign outputs[3621] = layer0_outputs[7938];
    assign outputs[3622] = layer0_outputs[6970];
    assign outputs[3623] = layer0_outputs[6294];
    assign outputs[3624] = ~(layer0_outputs[5629]);
    assign outputs[3625] = ~(layer0_outputs[7587]);
    assign outputs[3626] = ~((layer0_outputs[2521]) & (layer0_outputs[7973]));
    assign outputs[3627] = ~(layer0_outputs[1709]);
    assign outputs[3628] = layer0_outputs[4982];
    assign outputs[3629] = (layer0_outputs[2261]) | (layer0_outputs[432]);
    assign outputs[3630] = layer0_outputs[6841];
    assign outputs[3631] = ~(layer0_outputs[3363]);
    assign outputs[3632] = (layer0_outputs[9413]) & (layer0_outputs[3863]);
    assign outputs[3633] = ~(layer0_outputs[8667]);
    assign outputs[3634] = layer0_outputs[6056];
    assign outputs[3635] = ~(layer0_outputs[6444]);
    assign outputs[3636] = layer0_outputs[6052];
    assign outputs[3637] = ~(layer0_outputs[5152]);
    assign outputs[3638] = (layer0_outputs[8651]) ^ (layer0_outputs[7202]);
    assign outputs[3639] = ~(layer0_outputs[5441]);
    assign outputs[3640] = ~(layer0_outputs[3997]);
    assign outputs[3641] = layer0_outputs[8019];
    assign outputs[3642] = ~(layer0_outputs[9579]) | (layer0_outputs[2736]);
    assign outputs[3643] = ~(layer0_outputs[3836]);
    assign outputs[3644] = (layer0_outputs[5267]) ^ (layer0_outputs[297]);
    assign outputs[3645] = layer0_outputs[8219];
    assign outputs[3646] = ~((layer0_outputs[1650]) | (layer0_outputs[5926]));
    assign outputs[3647] = layer0_outputs[259];
    assign outputs[3648] = ~(layer0_outputs[2195]);
    assign outputs[3649] = ~(layer0_outputs[9179]) | (layer0_outputs[4159]);
    assign outputs[3650] = ~(layer0_outputs[970]);
    assign outputs[3651] = layer0_outputs[2266];
    assign outputs[3652] = layer0_outputs[6202];
    assign outputs[3653] = ~(layer0_outputs[6341]);
    assign outputs[3654] = ~((layer0_outputs[691]) ^ (layer0_outputs[5498]));
    assign outputs[3655] = ~((layer0_outputs[4279]) ^ (layer0_outputs[5]));
    assign outputs[3656] = layer0_outputs[2227];
    assign outputs[3657] = (layer0_outputs[2322]) ^ (layer0_outputs[4488]);
    assign outputs[3658] = (layer0_outputs[1400]) ^ (layer0_outputs[1337]);
    assign outputs[3659] = (layer0_outputs[3745]) & ~(layer0_outputs[1246]);
    assign outputs[3660] = ~(layer0_outputs[9962]);
    assign outputs[3661] = ~(layer0_outputs[9038]) | (layer0_outputs[2316]);
    assign outputs[3662] = layer0_outputs[3732];
    assign outputs[3663] = ~(layer0_outputs[9302]) | (layer0_outputs[2914]);
    assign outputs[3664] = (layer0_outputs[3154]) | (layer0_outputs[6982]);
    assign outputs[3665] = ~(layer0_outputs[999]) | (layer0_outputs[6637]);
    assign outputs[3666] = ~(layer0_outputs[1781]);
    assign outputs[3667] = (layer0_outputs[4763]) ^ (layer0_outputs[1384]);
    assign outputs[3668] = ~(layer0_outputs[6134]) | (layer0_outputs[1577]);
    assign outputs[3669] = ~(layer0_outputs[8295]);
    assign outputs[3670] = layer0_outputs[8082];
    assign outputs[3671] = ~((layer0_outputs[8591]) ^ (layer0_outputs[3101]));
    assign outputs[3672] = (layer0_outputs[9721]) ^ (layer0_outputs[2526]);
    assign outputs[3673] = ~((layer0_outputs[101]) & (layer0_outputs[9023]));
    assign outputs[3674] = ~(layer0_outputs[6681]);
    assign outputs[3675] = ~(layer0_outputs[7308]);
    assign outputs[3676] = ~(layer0_outputs[2348]);
    assign outputs[3677] = ~(layer0_outputs[7469]);
    assign outputs[3678] = ~(layer0_outputs[7174]) | (layer0_outputs[6541]);
    assign outputs[3679] = ~((layer0_outputs[6119]) ^ (layer0_outputs[4307]));
    assign outputs[3680] = 1'b0;
    assign outputs[3681] = ~((layer0_outputs[7347]) ^ (layer0_outputs[8568]));
    assign outputs[3682] = ~((layer0_outputs[775]) ^ (layer0_outputs[8410]));
    assign outputs[3683] = ~((layer0_outputs[8153]) & (layer0_outputs[4641]));
    assign outputs[3684] = (layer0_outputs[3325]) | (layer0_outputs[5107]);
    assign outputs[3685] = ~(layer0_outputs[3039]);
    assign outputs[3686] = ~(layer0_outputs[2236]) | (layer0_outputs[4733]);
    assign outputs[3687] = layer0_outputs[7138];
    assign outputs[3688] = ~((layer0_outputs[1525]) ^ (layer0_outputs[1730]));
    assign outputs[3689] = ~(layer0_outputs[8785]);
    assign outputs[3690] = layer0_outputs[7286];
    assign outputs[3691] = (layer0_outputs[2657]) & ~(layer0_outputs[4090]);
    assign outputs[3692] = layer0_outputs[6196];
    assign outputs[3693] = (layer0_outputs[2956]) | (layer0_outputs[1371]);
    assign outputs[3694] = (layer0_outputs[9645]) | (layer0_outputs[58]);
    assign outputs[3695] = layer0_outputs[9822];
    assign outputs[3696] = ~(layer0_outputs[6533]);
    assign outputs[3697] = ~(layer0_outputs[6071]) | (layer0_outputs[10005]);
    assign outputs[3698] = ~(layer0_outputs[8438]);
    assign outputs[3699] = ~(layer0_outputs[838]);
    assign outputs[3700] = (layer0_outputs[2951]) ^ (layer0_outputs[4924]);
    assign outputs[3701] = ~(layer0_outputs[10165]);
    assign outputs[3702] = (layer0_outputs[964]) & (layer0_outputs[8491]);
    assign outputs[3703] = (layer0_outputs[3385]) ^ (layer0_outputs[861]);
    assign outputs[3704] = ~((layer0_outputs[4737]) ^ (layer0_outputs[8026]));
    assign outputs[3705] = layer0_outputs[120];
    assign outputs[3706] = (layer0_outputs[5930]) ^ (layer0_outputs[8561]);
    assign outputs[3707] = layer0_outputs[3017];
    assign outputs[3708] = ~(layer0_outputs[6130]);
    assign outputs[3709] = ~(layer0_outputs[4921]);
    assign outputs[3710] = ~(layer0_outputs[5877]);
    assign outputs[3711] = ~(layer0_outputs[6550]);
    assign outputs[3712] = layer0_outputs[9684];
    assign outputs[3713] = ~((layer0_outputs[3420]) & (layer0_outputs[3525]));
    assign outputs[3714] = ~((layer0_outputs[8905]) & (layer0_outputs[5809]));
    assign outputs[3715] = (layer0_outputs[6510]) & (layer0_outputs[5275]);
    assign outputs[3716] = (layer0_outputs[7797]) | (layer0_outputs[10211]);
    assign outputs[3717] = ~((layer0_outputs[2872]) ^ (layer0_outputs[7960]));
    assign outputs[3718] = layer0_outputs[4153];
    assign outputs[3719] = ~((layer0_outputs[3016]) ^ (layer0_outputs[5719]));
    assign outputs[3720] = (layer0_outputs[5290]) ^ (layer0_outputs[4004]);
    assign outputs[3721] = ~(layer0_outputs[2816]);
    assign outputs[3722] = ~((layer0_outputs[3765]) ^ (layer0_outputs[786]));
    assign outputs[3723] = ~(layer0_outputs[9298]) | (layer0_outputs[4694]);
    assign outputs[3724] = ~(layer0_outputs[3571]);
    assign outputs[3725] = (layer0_outputs[8266]) ^ (layer0_outputs[9086]);
    assign outputs[3726] = ~((layer0_outputs[4589]) & (layer0_outputs[2742]));
    assign outputs[3727] = (layer0_outputs[9073]) ^ (layer0_outputs[6136]);
    assign outputs[3728] = layer0_outputs[7974];
    assign outputs[3729] = ~(layer0_outputs[8861]);
    assign outputs[3730] = ~((layer0_outputs[1401]) ^ (layer0_outputs[3165]));
    assign outputs[3731] = layer0_outputs[9424];
    assign outputs[3732] = ~(layer0_outputs[9758]);
    assign outputs[3733] = ~((layer0_outputs[9223]) | (layer0_outputs[1948]));
    assign outputs[3734] = ~(layer0_outputs[5384]) | (layer0_outputs[5526]);
    assign outputs[3735] = ~(layer0_outputs[1431]);
    assign outputs[3736] = (layer0_outputs[8581]) & (layer0_outputs[6935]);
    assign outputs[3737] = ~(layer0_outputs[6419]);
    assign outputs[3738] = layer0_outputs[3846];
    assign outputs[3739] = (layer0_outputs[5734]) | (layer0_outputs[2076]);
    assign outputs[3740] = (layer0_outputs[6884]) ^ (layer0_outputs[9141]);
    assign outputs[3741] = 1'b1;
    assign outputs[3742] = ~((layer0_outputs[6229]) ^ (layer0_outputs[7275]));
    assign outputs[3743] = (layer0_outputs[10031]) | (layer0_outputs[5141]);
    assign outputs[3744] = (layer0_outputs[5561]) & ~(layer0_outputs[6952]);
    assign outputs[3745] = ~(layer0_outputs[9035]) | (layer0_outputs[4459]);
    assign outputs[3746] = layer0_outputs[4935];
    assign outputs[3747] = ~(layer0_outputs[4]);
    assign outputs[3748] = (layer0_outputs[2771]) & ~(layer0_outputs[424]);
    assign outputs[3749] = ~((layer0_outputs[9199]) ^ (layer0_outputs[1630]));
    assign outputs[3750] = ~((layer0_outputs[5335]) | (layer0_outputs[4857]));
    assign outputs[3751] = (layer0_outputs[7375]) ^ (layer0_outputs[3909]);
    assign outputs[3752] = layer0_outputs[7231];
    assign outputs[3753] = (layer0_outputs[9693]) ^ (layer0_outputs[3330]);
    assign outputs[3754] = (layer0_outputs[2270]) & ~(layer0_outputs[7895]);
    assign outputs[3755] = ~(layer0_outputs[4106]);
    assign outputs[3756] = ~((layer0_outputs[9800]) ^ (layer0_outputs[3983]));
    assign outputs[3757] = layer0_outputs[4189];
    assign outputs[3758] = (layer0_outputs[2527]) ^ (layer0_outputs[9867]);
    assign outputs[3759] = ~((layer0_outputs[6303]) ^ (layer0_outputs[9267]));
    assign outputs[3760] = ~(layer0_outputs[3664]);
    assign outputs[3761] = layer0_outputs[8235];
    assign outputs[3762] = layer0_outputs[5398];
    assign outputs[3763] = layer0_outputs[3441];
    assign outputs[3764] = ~(layer0_outputs[2401]);
    assign outputs[3765] = ~(layer0_outputs[5360]);
    assign outputs[3766] = (layer0_outputs[4241]) | (layer0_outputs[5422]);
    assign outputs[3767] = ~(layer0_outputs[5793]);
    assign outputs[3768] = (layer0_outputs[2899]) ^ (layer0_outputs[1440]);
    assign outputs[3769] = (layer0_outputs[706]) ^ (layer0_outputs[1889]);
    assign outputs[3770] = ~((layer0_outputs[9668]) ^ (layer0_outputs[6384]));
    assign outputs[3771] = ~(layer0_outputs[2815]);
    assign outputs[3772] = ~(layer0_outputs[5058]);
    assign outputs[3773] = layer0_outputs[3233];
    assign outputs[3774] = (layer0_outputs[8333]) ^ (layer0_outputs[4367]);
    assign outputs[3775] = (layer0_outputs[2242]) ^ (layer0_outputs[5994]);
    assign outputs[3776] = ~(layer0_outputs[10015]) | (layer0_outputs[8815]);
    assign outputs[3777] = ~((layer0_outputs[3120]) ^ (layer0_outputs[6257]));
    assign outputs[3778] = ~(layer0_outputs[1789]);
    assign outputs[3779] = ~((layer0_outputs[3103]) & (layer0_outputs[6004]));
    assign outputs[3780] = ~(layer0_outputs[5957]);
    assign outputs[3781] = (layer0_outputs[8460]) ^ (layer0_outputs[6445]);
    assign outputs[3782] = layer0_outputs[8769];
    assign outputs[3783] = (layer0_outputs[7990]) ^ (layer0_outputs[9513]);
    assign outputs[3784] = ~(layer0_outputs[5165]);
    assign outputs[3785] = (layer0_outputs[4866]) & (layer0_outputs[2421]);
    assign outputs[3786] = layer0_outputs[4240];
    assign outputs[3787] = ~(layer0_outputs[2456]) | (layer0_outputs[5689]);
    assign outputs[3788] = ~((layer0_outputs[24]) ^ (layer0_outputs[5495]));
    assign outputs[3789] = layer0_outputs[7545];
    assign outputs[3790] = layer0_outputs[1607];
    assign outputs[3791] = ~(layer0_outputs[7117]);
    assign outputs[3792] = ~(layer0_outputs[6887]);
    assign outputs[3793] = ~(layer0_outputs[6934]) | (layer0_outputs[1923]);
    assign outputs[3794] = (layer0_outputs[4322]) | (layer0_outputs[5560]);
    assign outputs[3795] = ~((layer0_outputs[6855]) ^ (layer0_outputs[5106]));
    assign outputs[3796] = ~((layer0_outputs[717]) ^ (layer0_outputs[1333]));
    assign outputs[3797] = ~(layer0_outputs[4210]);
    assign outputs[3798] = (layer0_outputs[6840]) & ~(layer0_outputs[6690]);
    assign outputs[3799] = ~((layer0_outputs[7954]) ^ (layer0_outputs[2837]));
    assign outputs[3800] = layer0_outputs[1214];
    assign outputs[3801] = ~(layer0_outputs[3944]);
    assign outputs[3802] = ~(layer0_outputs[7675]);
    assign outputs[3803] = (layer0_outputs[930]) & ~(layer0_outputs[7643]);
    assign outputs[3804] = ~((layer0_outputs[979]) ^ (layer0_outputs[973]));
    assign outputs[3805] = (layer0_outputs[7393]) & (layer0_outputs[2355]);
    assign outputs[3806] = layer0_outputs[6476];
    assign outputs[3807] = ~((layer0_outputs[7020]) | (layer0_outputs[9119]));
    assign outputs[3808] = ~(layer0_outputs[1707]) | (layer0_outputs[8504]);
    assign outputs[3809] = ~((layer0_outputs[417]) ^ (layer0_outputs[523]));
    assign outputs[3810] = ~((layer0_outputs[9024]) & (layer0_outputs[5751]));
    assign outputs[3811] = ~(layer0_outputs[3335]) | (layer0_outputs[8133]);
    assign outputs[3812] = ~(layer0_outputs[4411]);
    assign outputs[3813] = (layer0_outputs[139]) ^ (layer0_outputs[6642]);
    assign outputs[3814] = ~(layer0_outputs[5410]);
    assign outputs[3815] = ~((layer0_outputs[3198]) ^ (layer0_outputs[5634]));
    assign outputs[3816] = (layer0_outputs[1863]) & ~(layer0_outputs[6973]);
    assign outputs[3817] = ~(layer0_outputs[8221]);
    assign outputs[3818] = layer0_outputs[3115];
    assign outputs[3819] = ~((layer0_outputs[5000]) ^ (layer0_outputs[8365]));
    assign outputs[3820] = ~((layer0_outputs[10019]) ^ (layer0_outputs[2207]));
    assign outputs[3821] = ~((layer0_outputs[6708]) ^ (layer0_outputs[476]));
    assign outputs[3822] = layer0_outputs[7073];
    assign outputs[3823] = (layer0_outputs[2781]) & ~(layer0_outputs[9844]);
    assign outputs[3824] = ~((layer0_outputs[2913]) ^ (layer0_outputs[4340]));
    assign outputs[3825] = ~(layer0_outputs[1066]) | (layer0_outputs[4175]);
    assign outputs[3826] = (layer0_outputs[1525]) & ~(layer0_outputs[8993]);
    assign outputs[3827] = (layer0_outputs[7499]) ^ (layer0_outputs[7644]);
    assign outputs[3828] = (layer0_outputs[1674]) ^ (layer0_outputs[6173]);
    assign outputs[3829] = layer0_outputs[5707];
    assign outputs[3830] = (layer0_outputs[4539]) ^ (layer0_outputs[8534]);
    assign outputs[3831] = (layer0_outputs[938]) & ~(layer0_outputs[7364]);
    assign outputs[3832] = layer0_outputs[4575];
    assign outputs[3833] = layer0_outputs[7992];
    assign outputs[3834] = 1'b1;
    assign outputs[3835] = ~(layer0_outputs[7185]) | (layer0_outputs[6457]);
    assign outputs[3836] = ~(layer0_outputs[6036]);
    assign outputs[3837] = (layer0_outputs[2640]) ^ (layer0_outputs[9979]);
    assign outputs[3838] = ~(layer0_outputs[2851]);
    assign outputs[3839] = (layer0_outputs[5933]) | (layer0_outputs[6960]);
    assign outputs[3840] = (layer0_outputs[9104]) & ~(layer0_outputs[9766]);
    assign outputs[3841] = (layer0_outputs[8325]) & ~(layer0_outputs[716]);
    assign outputs[3842] = ~(layer0_outputs[9439]);
    assign outputs[3843] = ~(layer0_outputs[4050]);
    assign outputs[3844] = (layer0_outputs[1878]) ^ (layer0_outputs[5145]);
    assign outputs[3845] = ~((layer0_outputs[620]) ^ (layer0_outputs[9376]));
    assign outputs[3846] = ~(layer0_outputs[10181]) | (layer0_outputs[7151]);
    assign outputs[3847] = layer0_outputs[4021];
    assign outputs[3848] = layer0_outputs[5099];
    assign outputs[3849] = layer0_outputs[5288];
    assign outputs[3850] = (layer0_outputs[4244]) & ~(layer0_outputs[3584]);
    assign outputs[3851] = (layer0_outputs[9811]) & (layer0_outputs[5104]);
    assign outputs[3852] = ~(layer0_outputs[6739]);
    assign outputs[3853] = ~(layer0_outputs[4867]);
    assign outputs[3854] = (layer0_outputs[3428]) ^ (layer0_outputs[4810]);
    assign outputs[3855] = ~(layer0_outputs[5647]) | (layer0_outputs[3969]);
    assign outputs[3856] = layer0_outputs[8292];
    assign outputs[3857] = ~(layer0_outputs[7251]) | (layer0_outputs[3523]);
    assign outputs[3858] = (layer0_outputs[1801]) ^ (layer0_outputs[3070]);
    assign outputs[3859] = (layer0_outputs[7031]) | (layer0_outputs[7979]);
    assign outputs[3860] = layer0_outputs[10099];
    assign outputs[3861] = layer0_outputs[3539];
    assign outputs[3862] = ~(layer0_outputs[5173]);
    assign outputs[3863] = layer0_outputs[5311];
    assign outputs[3864] = ~((layer0_outputs[3993]) & (layer0_outputs[8931]));
    assign outputs[3865] = ~(layer0_outputs[6383]);
    assign outputs[3866] = ~(layer0_outputs[3980]);
    assign outputs[3867] = ~(layer0_outputs[5137]) | (layer0_outputs[910]);
    assign outputs[3868] = layer0_outputs[8961];
    assign outputs[3869] = (layer0_outputs[1319]) ^ (layer0_outputs[5070]);
    assign outputs[3870] = ~((layer0_outputs[6381]) ^ (layer0_outputs[483]));
    assign outputs[3871] = layer0_outputs[3623];
    assign outputs[3872] = (layer0_outputs[685]) ^ (layer0_outputs[9533]);
    assign outputs[3873] = layer0_outputs[3505];
    assign outputs[3874] = (layer0_outputs[9460]) & ~(layer0_outputs[2437]);
    assign outputs[3875] = (layer0_outputs[397]) ^ (layer0_outputs[305]);
    assign outputs[3876] = layer0_outputs[7224];
    assign outputs[3877] = (layer0_outputs[5105]) & ~(layer0_outputs[3068]);
    assign outputs[3878] = (layer0_outputs[2183]) & (layer0_outputs[7394]);
    assign outputs[3879] = ~(layer0_outputs[4335]);
    assign outputs[3880] = (layer0_outputs[9696]) & (layer0_outputs[7542]);
    assign outputs[3881] = layer0_outputs[2001];
    assign outputs[3882] = (layer0_outputs[6031]) | (layer0_outputs[2684]);
    assign outputs[3883] = (layer0_outputs[1496]) ^ (layer0_outputs[5261]);
    assign outputs[3884] = ~(layer0_outputs[4309]);
    assign outputs[3885] = (layer0_outputs[833]) | (layer0_outputs[1348]);
    assign outputs[3886] = ~((layer0_outputs[7999]) ^ (layer0_outputs[4790]));
    assign outputs[3887] = layer0_outputs[1364];
    assign outputs[3888] = (layer0_outputs[9832]) ^ (layer0_outputs[9084]);
    assign outputs[3889] = layer0_outputs[5788];
    assign outputs[3890] = ~(layer0_outputs[10013]);
    assign outputs[3891] = (layer0_outputs[6129]) ^ (layer0_outputs[3205]);
    assign outputs[3892] = (layer0_outputs[4007]) & (layer0_outputs[8116]);
    assign outputs[3893] = ~(layer0_outputs[6919]);
    assign outputs[3894] = ~(layer0_outputs[826]) | (layer0_outputs[5357]);
    assign outputs[3895] = ~(layer0_outputs[6570]) | (layer0_outputs[1766]);
    assign outputs[3896] = ~(layer0_outputs[8322]);
    assign outputs[3897] = ~(layer0_outputs[6483]);
    assign outputs[3898] = ~((layer0_outputs[8169]) | (layer0_outputs[344]));
    assign outputs[3899] = layer0_outputs[4922];
    assign outputs[3900] = ~((layer0_outputs[6574]) & (layer0_outputs[826]));
    assign outputs[3901] = layer0_outputs[9461];
    assign outputs[3902] = ~((layer0_outputs[5041]) ^ (layer0_outputs[8150]));
    assign outputs[3903] = layer0_outputs[28];
    assign outputs[3904] = ~((layer0_outputs[4996]) & (layer0_outputs[10163]));
    assign outputs[3905] = 1'b1;
    assign outputs[3906] = ~((layer0_outputs[8179]) & (layer0_outputs[6766]));
    assign outputs[3907] = ~((layer0_outputs[1048]) & (layer0_outputs[107]));
    assign outputs[3908] = (layer0_outputs[2501]) | (layer0_outputs[2553]);
    assign outputs[3909] = ~(layer0_outputs[4692]);
    assign outputs[3910] = ~(layer0_outputs[8135]);
    assign outputs[3911] = (layer0_outputs[5394]) & (layer0_outputs[2142]);
    assign outputs[3912] = layer0_outputs[1113];
    assign outputs[3913] = ~(layer0_outputs[86]);
    assign outputs[3914] = ~(layer0_outputs[4446]);
    assign outputs[3915] = ~(layer0_outputs[4212]);
    assign outputs[3916] = ~(layer0_outputs[1850]) | (layer0_outputs[9702]);
    assign outputs[3917] = layer0_outputs[5483];
    assign outputs[3918] = ~(layer0_outputs[9208]) | (layer0_outputs[9881]);
    assign outputs[3919] = layer0_outputs[785];
    assign outputs[3920] = ~(layer0_outputs[159]);
    assign outputs[3921] = ~(layer0_outputs[6512]) | (layer0_outputs[9513]);
    assign outputs[3922] = layer0_outputs[4559];
    assign outputs[3923] = ~(layer0_outputs[7629]);
    assign outputs[3924] = ~(layer0_outputs[3726]);
    assign outputs[3925] = layer0_outputs[3713];
    assign outputs[3926] = (layer0_outputs[5188]) ^ (layer0_outputs[8355]);
    assign outputs[3927] = layer0_outputs[8919];
    assign outputs[3928] = ~((layer0_outputs[6804]) ^ (layer0_outputs[4380]));
    assign outputs[3929] = (layer0_outputs[6997]) & (layer0_outputs[5541]);
    assign outputs[3930] = ~(layer0_outputs[5409]) | (layer0_outputs[8857]);
    assign outputs[3931] = (layer0_outputs[8771]) & ~(layer0_outputs[2477]);
    assign outputs[3932] = (layer0_outputs[10160]) | (layer0_outputs[5336]);
    assign outputs[3933] = ~(layer0_outputs[5033]);
    assign outputs[3934] = ~(layer0_outputs[4180]) | (layer0_outputs[9841]);
    assign outputs[3935] = (layer0_outputs[6735]) ^ (layer0_outputs[6441]);
    assign outputs[3936] = ~(layer0_outputs[3217]);
    assign outputs[3937] = (layer0_outputs[4798]) ^ (layer0_outputs[365]);
    assign outputs[3938] = ~((layer0_outputs[3502]) ^ (layer0_outputs[1876]));
    assign outputs[3939] = ~(layer0_outputs[6786]);
    assign outputs[3940] = ~(layer0_outputs[1454]) | (layer0_outputs[3045]);
    assign outputs[3941] = (layer0_outputs[7363]) & ~(layer0_outputs[6783]);
    assign outputs[3942] = ~(layer0_outputs[3359]) | (layer0_outputs[4724]);
    assign outputs[3943] = layer0_outputs[9601];
    assign outputs[3944] = ~((layer0_outputs[5164]) & (layer0_outputs[2216]));
    assign outputs[3945] = ~(layer0_outputs[9879]);
    assign outputs[3946] = layer0_outputs[1867];
    assign outputs[3947] = layer0_outputs[117];
    assign outputs[3948] = layer0_outputs[3218];
    assign outputs[3949] = ~(layer0_outputs[8457]);
    assign outputs[3950] = layer0_outputs[3437];
    assign outputs[3951] = layer0_outputs[3978];
    assign outputs[3952] = ~(layer0_outputs[8618]);
    assign outputs[3953] = ~(layer0_outputs[9992]) | (layer0_outputs[7582]);
    assign outputs[3954] = ~((layer0_outputs[10157]) ^ (layer0_outputs[3880]));
    assign outputs[3955] = (layer0_outputs[9619]) ^ (layer0_outputs[10153]);
    assign outputs[3956] = ~((layer0_outputs[5869]) | (layer0_outputs[2020]));
    assign outputs[3957] = ~(layer0_outputs[6521]);
    assign outputs[3958] = (layer0_outputs[1851]) ^ (layer0_outputs[9095]);
    assign outputs[3959] = ~((layer0_outputs[8966]) & (layer0_outputs[9517]));
    assign outputs[3960] = ~(layer0_outputs[8225]);
    assign outputs[3961] = ~((layer0_outputs[3062]) ^ (layer0_outputs[9556]));
    assign outputs[3962] = ~((layer0_outputs[2516]) ^ (layer0_outputs[47]));
    assign outputs[3963] = (layer0_outputs[4407]) & ~(layer0_outputs[1293]);
    assign outputs[3964] = (layer0_outputs[2723]) & (layer0_outputs[5291]);
    assign outputs[3965] = ~(layer0_outputs[6014]);
    assign outputs[3966] = (layer0_outputs[8855]) ^ (layer0_outputs[3101]);
    assign outputs[3967] = ~(layer0_outputs[3734]);
    assign outputs[3968] = ~(layer0_outputs[8379]);
    assign outputs[3969] = (layer0_outputs[796]) | (layer0_outputs[4209]);
    assign outputs[3970] = ~((layer0_outputs[4995]) | (layer0_outputs[878]));
    assign outputs[3971] = layer0_outputs[9997];
    assign outputs[3972] = (layer0_outputs[4943]) ^ (layer0_outputs[4204]);
    assign outputs[3973] = ~(layer0_outputs[8578]);
    assign outputs[3974] = ~(layer0_outputs[5789]);
    assign outputs[3975] = layer0_outputs[7914];
    assign outputs[3976] = (layer0_outputs[7326]) ^ (layer0_outputs[4761]);
    assign outputs[3977] = ~(layer0_outputs[341]) | (layer0_outputs[3305]);
    assign outputs[3978] = (layer0_outputs[759]) ^ (layer0_outputs[6588]);
    assign outputs[3979] = (layer0_outputs[7666]) ^ (layer0_outputs[9688]);
    assign outputs[3980] = ~(layer0_outputs[7444]);
    assign outputs[3981] = (layer0_outputs[5448]) ^ (layer0_outputs[7713]);
    assign outputs[3982] = (layer0_outputs[9514]) & ~(layer0_outputs[352]);
    assign outputs[3983] = layer0_outputs[8831];
    assign outputs[3984] = ~((layer0_outputs[2428]) ^ (layer0_outputs[10085]));
    assign outputs[3985] = ~(layer0_outputs[8803]) | (layer0_outputs[9151]);
    assign outputs[3986] = layer0_outputs[2138];
    assign outputs[3987] = layer0_outputs[9519];
    assign outputs[3988] = (layer0_outputs[923]) & (layer0_outputs[6015]);
    assign outputs[3989] = ~(layer0_outputs[4426]);
    assign outputs[3990] = layer0_outputs[603];
    assign outputs[3991] = (layer0_outputs[310]) | (layer0_outputs[6617]);
    assign outputs[3992] = ~(layer0_outputs[5147]);
    assign outputs[3993] = ~((layer0_outputs[3778]) ^ (layer0_outputs[5875]));
    assign outputs[3994] = ~((layer0_outputs[6526]) ^ (layer0_outputs[2713]));
    assign outputs[3995] = ~((layer0_outputs[6059]) & (layer0_outputs[382]));
    assign outputs[3996] = ~(layer0_outputs[444]);
    assign outputs[3997] = (layer0_outputs[4175]) | (layer0_outputs[7798]);
    assign outputs[3998] = ~(layer0_outputs[3229]);
    assign outputs[3999] = ~((layer0_outputs[6142]) ^ (layer0_outputs[3208]));
    assign outputs[4000] = ~(layer0_outputs[498]);
    assign outputs[4001] = (layer0_outputs[1517]) ^ (layer0_outputs[5839]);
    assign outputs[4002] = (layer0_outputs[4114]) ^ (layer0_outputs[3246]);
    assign outputs[4003] = layer0_outputs[6801];
    assign outputs[4004] = ~((layer0_outputs[3478]) & (layer0_outputs[3391]));
    assign outputs[4005] = (layer0_outputs[9582]) ^ (layer0_outputs[9951]);
    assign outputs[4006] = ~(layer0_outputs[2078]);
    assign outputs[4007] = ~((layer0_outputs[2652]) ^ (layer0_outputs[7153]));
    assign outputs[4008] = ~(layer0_outputs[6906]);
    assign outputs[4009] = (layer0_outputs[8566]) ^ (layer0_outputs[3581]);
    assign outputs[4010] = (layer0_outputs[2946]) & (layer0_outputs[3020]);
    assign outputs[4011] = (layer0_outputs[4071]) ^ (layer0_outputs[7145]);
    assign outputs[4012] = ~((layer0_outputs[3213]) ^ (layer0_outputs[7773]));
    assign outputs[4013] = layer0_outputs[7060];
    assign outputs[4014] = ~(layer0_outputs[5956]);
    assign outputs[4015] = ~((layer0_outputs[141]) & (layer0_outputs[490]));
    assign outputs[4016] = ~(layer0_outputs[1296]);
    assign outputs[4017] = 1'b1;
    assign outputs[4018] = (layer0_outputs[6197]) | (layer0_outputs[7697]);
    assign outputs[4019] = layer0_outputs[7217];
    assign outputs[4020] = (layer0_outputs[7295]) ^ (layer0_outputs[609]);
    assign outputs[4021] = layer0_outputs[3662];
    assign outputs[4022] = layer0_outputs[4215];
    assign outputs[4023] = ~(layer0_outputs[6170]);
    assign outputs[4024] = ~((layer0_outputs[6680]) & (layer0_outputs[1387]));
    assign outputs[4025] = ~(layer0_outputs[659]);
    assign outputs[4026] = (layer0_outputs[8880]) & (layer0_outputs[6885]);
    assign outputs[4027] = ~(layer0_outputs[10228]);
    assign outputs[4028] = ~((layer0_outputs[3399]) ^ (layer0_outputs[9030]));
    assign outputs[4029] = ~(layer0_outputs[6248]);
    assign outputs[4030] = (layer0_outputs[3231]) | (layer0_outputs[7115]);
    assign outputs[4031] = ~(layer0_outputs[8494]);
    assign outputs[4032] = layer0_outputs[3192];
    assign outputs[4033] = ~(layer0_outputs[6722]) | (layer0_outputs[2422]);
    assign outputs[4034] = ~(layer0_outputs[3413]);
    assign outputs[4035] = layer0_outputs[4220];
    assign outputs[4036] = layer0_outputs[8061];
    assign outputs[4037] = (layer0_outputs[536]) & (layer0_outputs[3597]);
    assign outputs[4038] = ~((layer0_outputs[4045]) ^ (layer0_outputs[9752]));
    assign outputs[4039] = ~(layer0_outputs[9774]);
    assign outputs[4040] = (layer0_outputs[7177]) ^ (layer0_outputs[4686]);
    assign outputs[4041] = layer0_outputs[6639];
    assign outputs[4042] = layer0_outputs[178];
    assign outputs[4043] = ~((layer0_outputs[6667]) ^ (layer0_outputs[9949]));
    assign outputs[4044] = ~(layer0_outputs[617]);
    assign outputs[4045] = ~(layer0_outputs[1131]);
    assign outputs[4046] = ~(layer0_outputs[839]) | (layer0_outputs[2641]);
    assign outputs[4047] = ~((layer0_outputs[258]) ^ (layer0_outputs[3251]));
    assign outputs[4048] = ~(layer0_outputs[756]);
    assign outputs[4049] = ~((layer0_outputs[4257]) ^ (layer0_outputs[7772]));
    assign outputs[4050] = ~(layer0_outputs[3906]);
    assign outputs[4051] = layer0_outputs[1638];
    assign outputs[4052] = layer0_outputs[421];
    assign outputs[4053] = layer0_outputs[3315];
    assign outputs[4054] = ~(layer0_outputs[5075]);
    assign outputs[4055] = ~(layer0_outputs[8030]);
    assign outputs[4056] = layer0_outputs[6477];
    assign outputs[4057] = layer0_outputs[9798];
    assign outputs[4058] = ~(layer0_outputs[5862]) | (layer0_outputs[151]);
    assign outputs[4059] = ~(layer0_outputs[2180]);
    assign outputs[4060] = ~(layer0_outputs[2141]);
    assign outputs[4061] = ~((layer0_outputs[8675]) & (layer0_outputs[4957]));
    assign outputs[4062] = ~((layer0_outputs[10009]) ^ (layer0_outputs[6167]));
    assign outputs[4063] = (layer0_outputs[3628]) | (layer0_outputs[6501]);
    assign outputs[4064] = ~(layer0_outputs[4691]) | (layer0_outputs[2936]);
    assign outputs[4065] = layer0_outputs[70];
    assign outputs[4066] = ~((layer0_outputs[1480]) ^ (layer0_outputs[7146]));
    assign outputs[4067] = ~((layer0_outputs[9476]) | (layer0_outputs[4148]));
    assign outputs[4068] = (layer0_outputs[9142]) ^ (layer0_outputs[3226]);
    assign outputs[4069] = (layer0_outputs[9677]) | (layer0_outputs[4536]);
    assign outputs[4070] = ~((layer0_outputs[9710]) ^ (layer0_outputs[2325]));
    assign outputs[4071] = (layer0_outputs[7614]) & ~(layer0_outputs[8296]);
    assign outputs[4072] = ~((layer0_outputs[8102]) & (layer0_outputs[9828]));
    assign outputs[4073] = layer0_outputs[2515];
    assign outputs[4074] = ~(layer0_outputs[8338]) | (layer0_outputs[1146]);
    assign outputs[4075] = layer0_outputs[7087];
    assign outputs[4076] = ~(layer0_outputs[8089]);
    assign outputs[4077] = (layer0_outputs[8514]) ^ (layer0_outputs[383]);
    assign outputs[4078] = layer0_outputs[6660];
    assign outputs[4079] = layer0_outputs[7586];
    assign outputs[4080] = layer0_outputs[2722];
    assign outputs[4081] = (layer0_outputs[1504]) ^ (layer0_outputs[2759]);
    assign outputs[4082] = (layer0_outputs[8598]) ^ (layer0_outputs[7891]);
    assign outputs[4083] = (layer0_outputs[4722]) & (layer0_outputs[18]);
    assign outputs[4084] = layer0_outputs[806];
    assign outputs[4085] = layer0_outputs[6788];
    assign outputs[4086] = layer0_outputs[4386];
    assign outputs[4087] = ~(layer0_outputs[10120]);
    assign outputs[4088] = ~(layer0_outputs[8289]);
    assign outputs[4089] = (layer0_outputs[2461]) & (layer0_outputs[1425]);
    assign outputs[4090] = ~(layer0_outputs[3746]);
    assign outputs[4091] = (layer0_outputs[5585]) ^ (layer0_outputs[5925]);
    assign outputs[4092] = ~(layer0_outputs[2961]);
    assign outputs[4093] = ~(layer0_outputs[1049]) | (layer0_outputs[2724]);
    assign outputs[4094] = ~((layer0_outputs[8988]) ^ (layer0_outputs[1508]));
    assign outputs[4095] = (layer0_outputs[6708]) ^ (layer0_outputs[4601]);
    assign outputs[4096] = layer0_outputs[5703];
    assign outputs[4097] = ~((layer0_outputs[6075]) | (layer0_outputs[6686]));
    assign outputs[4098] = (layer0_outputs[5438]) ^ (layer0_outputs[2783]);
    assign outputs[4099] = (layer0_outputs[4179]) ^ (layer0_outputs[668]);
    assign outputs[4100] = ~(layer0_outputs[5098]);
    assign outputs[4101] = ~(layer0_outputs[4605]);
    assign outputs[4102] = (layer0_outputs[7965]) ^ (layer0_outputs[2254]);
    assign outputs[4103] = ~((layer0_outputs[7618]) ^ (layer0_outputs[3394]));
    assign outputs[4104] = (layer0_outputs[10084]) ^ (layer0_outputs[1266]);
    assign outputs[4105] = (layer0_outputs[1316]) | (layer0_outputs[863]);
    assign outputs[4106] = (layer0_outputs[4762]) ^ (layer0_outputs[1848]);
    assign outputs[4107] = (layer0_outputs[4603]) ^ (layer0_outputs[2578]);
    assign outputs[4108] = ~((layer0_outputs[7342]) ^ (layer0_outputs[2750]));
    assign outputs[4109] = (layer0_outputs[5077]) & (layer0_outputs[8750]);
    assign outputs[4110] = layer0_outputs[4720];
    assign outputs[4111] = (layer0_outputs[5229]) ^ (layer0_outputs[8088]);
    assign outputs[4112] = (layer0_outputs[5945]) & ~(layer0_outputs[3752]);
    assign outputs[4113] = ~((layer0_outputs[7497]) & (layer0_outputs[4530]));
    assign outputs[4114] = ~(layer0_outputs[9845]);
    assign outputs[4115] = ~(layer0_outputs[3969]);
    assign outputs[4116] = (layer0_outputs[8232]) & ~(layer0_outputs[7096]);
    assign outputs[4117] = (layer0_outputs[8924]) & ~(layer0_outputs[1707]);
    assign outputs[4118] = ~(layer0_outputs[257]);
    assign outputs[4119] = ~((layer0_outputs[2142]) ^ (layer0_outputs[606]));
    assign outputs[4120] = layer0_outputs[10231];
    assign outputs[4121] = (layer0_outputs[5560]) & ~(layer0_outputs[574]);
    assign outputs[4122] = ~(layer0_outputs[4003]);
    assign outputs[4123] = ~(layer0_outputs[1284]);
    assign outputs[4124] = ~((layer0_outputs[5700]) ^ (layer0_outputs[8514]));
    assign outputs[4125] = (layer0_outputs[7847]) & ~(layer0_outputs[6501]);
    assign outputs[4126] = (layer0_outputs[761]) & ~(layer0_outputs[6280]);
    assign outputs[4127] = ~((layer0_outputs[4835]) | (layer0_outputs[5339]));
    assign outputs[4128] = ~((layer0_outputs[8408]) ^ (layer0_outputs[4026]));
    assign outputs[4129] = layer0_outputs[5450];
    assign outputs[4130] = (layer0_outputs[4073]) ^ (layer0_outputs[4005]);
    assign outputs[4131] = layer0_outputs[1942];
    assign outputs[4132] = ~((layer0_outputs[1472]) ^ (layer0_outputs[4325]));
    assign outputs[4133] = layer0_outputs[8944];
    assign outputs[4134] = (layer0_outputs[2822]) ^ (layer0_outputs[1211]);
    assign outputs[4135] = ~(layer0_outputs[7583]);
    assign outputs[4136] = (layer0_outputs[6389]) & ~(layer0_outputs[8009]);
    assign outputs[4137] = ~(layer0_outputs[495]) | (layer0_outputs[5445]);
    assign outputs[4138] = layer0_outputs[9856];
    assign outputs[4139] = (layer0_outputs[680]) & ~(layer0_outputs[5983]);
    assign outputs[4140] = layer0_outputs[4925];
    assign outputs[4141] = layer0_outputs[5165];
    assign outputs[4142] = (layer0_outputs[7168]) & ~(layer0_outputs[7578]);
    assign outputs[4143] = ~((layer0_outputs[8985]) | (layer0_outputs[4945]));
    assign outputs[4144] = (layer0_outputs[6886]) & ~(layer0_outputs[4142]);
    assign outputs[4145] = (layer0_outputs[5380]) & ~(layer0_outputs[2349]);
    assign outputs[4146] = layer0_outputs[7791];
    assign outputs[4147] = ~(layer0_outputs[9219]) | (layer0_outputs[5747]);
    assign outputs[4148] = ~((layer0_outputs[9739]) ^ (layer0_outputs[1874]));
    assign outputs[4149] = ~((layer0_outputs[3318]) | (layer0_outputs[7906]));
    assign outputs[4150] = (layer0_outputs[5231]) & (layer0_outputs[1891]);
    assign outputs[4151] = layer0_outputs[3322];
    assign outputs[4152] = layer0_outputs[8843];
    assign outputs[4153] = ~((layer0_outputs[2016]) ^ (layer0_outputs[4939]));
    assign outputs[4154] = ~(layer0_outputs[1996]);
    assign outputs[4155] = ~(layer0_outputs[9173]);
    assign outputs[4156] = ~(layer0_outputs[6610]);
    assign outputs[4157] = (layer0_outputs[8177]) & (layer0_outputs[19]);
    assign outputs[4158] = (layer0_outputs[9175]) | (layer0_outputs[774]);
    assign outputs[4159] = ~(layer0_outputs[7359]);
    assign outputs[4160] = layer0_outputs[6396];
    assign outputs[4161] = ~((layer0_outputs[5403]) ^ (layer0_outputs[7850]));
    assign outputs[4162] = ~(layer0_outputs[4373]);
    assign outputs[4163] = layer0_outputs[2919];
    assign outputs[4164] = (layer0_outputs[10114]) & ~(layer0_outputs[175]);
    assign outputs[4165] = (layer0_outputs[1014]) & ~(layer0_outputs[6598]);
    assign outputs[4166] = ~((layer0_outputs[4829]) & (layer0_outputs[8084]));
    assign outputs[4167] = ~((layer0_outputs[4064]) ^ (layer0_outputs[5062]));
    assign outputs[4168] = layer0_outputs[6496];
    assign outputs[4169] = layer0_outputs[967];
    assign outputs[4170] = (layer0_outputs[8546]) ^ (layer0_outputs[4920]);
    assign outputs[4171] = (layer0_outputs[7796]) & ~(layer0_outputs[4438]);
    assign outputs[4172] = (layer0_outputs[1782]) & ~(layer0_outputs[6478]);
    assign outputs[4173] = ~((layer0_outputs[5204]) ^ (layer0_outputs[3577]));
    assign outputs[4174] = ~(layer0_outputs[45]);
    assign outputs[4175] = layer0_outputs[6007];
    assign outputs[4176] = ~(layer0_outputs[4200]) | (layer0_outputs[2844]);
    assign outputs[4177] = (layer0_outputs[2314]) ^ (layer0_outputs[5167]);
    assign outputs[4178] = ~((layer0_outputs[5244]) ^ (layer0_outputs[51]));
    assign outputs[4179] = (layer0_outputs[954]) & ~(layer0_outputs[7705]);
    assign outputs[4180] = (layer0_outputs[8794]) & ~(layer0_outputs[7718]);
    assign outputs[4181] = (layer0_outputs[9970]) ^ (layer0_outputs[486]);
    assign outputs[4182] = ~(layer0_outputs[1078]) | (layer0_outputs[9903]);
    assign outputs[4183] = ~(layer0_outputs[6265]);
    assign outputs[4184] = (layer0_outputs[3582]) ^ (layer0_outputs[9485]);
    assign outputs[4185] = (layer0_outputs[3191]) ^ (layer0_outputs[260]);
    assign outputs[4186] = layer0_outputs[1871];
    assign outputs[4187] = (layer0_outputs[610]) & (layer0_outputs[10189]);
    assign outputs[4188] = layer0_outputs[5030];
    assign outputs[4189] = (layer0_outputs[4006]) ^ (layer0_outputs[947]);
    assign outputs[4190] = ~(layer0_outputs[4584]);
    assign outputs[4191] = ~((layer0_outputs[7277]) ^ (layer0_outputs[5456]));
    assign outputs[4192] = ~((layer0_outputs[7144]) | (layer0_outputs[6620]));
    assign outputs[4193] = (layer0_outputs[7050]) & ~(layer0_outputs[7289]);
    assign outputs[4194] = (layer0_outputs[9383]) ^ (layer0_outputs[3256]);
    assign outputs[4195] = layer0_outputs[4531];
    assign outputs[4196] = (layer0_outputs[961]) ^ (layer0_outputs[4127]);
    assign outputs[4197] = ~(layer0_outputs[8942]);
    assign outputs[4198] = (layer0_outputs[4091]) & ~(layer0_outputs[6959]);
    assign outputs[4199] = ~((layer0_outputs[294]) | (layer0_outputs[9950]));
    assign outputs[4200] = layer0_outputs[7254];
    assign outputs[4201] = ~(layer0_outputs[8856]);
    assign outputs[4202] = (layer0_outputs[8868]) & ~(layer0_outputs[8692]);
    assign outputs[4203] = (layer0_outputs[2710]) & (layer0_outputs[4949]);
    assign outputs[4204] = ~(layer0_outputs[2903]) | (layer0_outputs[3519]);
    assign outputs[4205] = (layer0_outputs[2590]) | (layer0_outputs[7493]);
    assign outputs[4206] = (layer0_outputs[5902]) & ~(layer0_outputs[851]);
    assign outputs[4207] = (layer0_outputs[4898]) ^ (layer0_outputs[7315]);
    assign outputs[4208] = (layer0_outputs[8035]) | (layer0_outputs[2627]);
    assign outputs[4209] = ~((layer0_outputs[860]) ^ (layer0_outputs[8624]));
    assign outputs[4210] = ~(layer0_outputs[7418]);
    assign outputs[4211] = 1'b0;
    assign outputs[4212] = ~(layer0_outputs[2252]);
    assign outputs[4213] = layer0_outputs[9489];
    assign outputs[4214] = ~(layer0_outputs[2417]);
    assign outputs[4215] = (layer0_outputs[1583]) & ~(layer0_outputs[4696]);
    assign outputs[4216] = ~(layer0_outputs[9206]);
    assign outputs[4217] = ~(layer0_outputs[7419]);
    assign outputs[4218] = (layer0_outputs[772]) & (layer0_outputs[1922]);
    assign outputs[4219] = (layer0_outputs[9368]) & ~(layer0_outputs[255]);
    assign outputs[4220] = ~(layer0_outputs[5656]);
    assign outputs[4221] = 1'b0;
    assign outputs[4222] = layer0_outputs[3185];
    assign outputs[4223] = (layer0_outputs[9773]) & ~(layer0_outputs[4515]);
    assign outputs[4224] = (layer0_outputs[1202]) & ~(layer0_outputs[2701]);
    assign outputs[4225] = ~((layer0_outputs[2415]) ^ (layer0_outputs[3861]));
    assign outputs[4226] = (layer0_outputs[2705]) ^ (layer0_outputs[3971]);
    assign outputs[4227] = (layer0_outputs[6563]) ^ (layer0_outputs[6100]);
    assign outputs[4228] = (layer0_outputs[3349]) & ~(layer0_outputs[6713]);
    assign outputs[4229] = ~(layer0_outputs[3901]);
    assign outputs[4230] = ~((layer0_outputs[8950]) & (layer0_outputs[10016]));
    assign outputs[4231] = ~((layer0_outputs[3777]) & (layer0_outputs[104]));
    assign outputs[4232] = ~(layer0_outputs[6483]);
    assign outputs[4233] = ~(layer0_outputs[4475]);
    assign outputs[4234] = ~((layer0_outputs[3040]) & (layer0_outputs[5904]));
    assign outputs[4235] = ~((layer0_outputs[3261]) ^ (layer0_outputs[3267]));
    assign outputs[4236] = (layer0_outputs[285]) ^ (layer0_outputs[2146]);
    assign outputs[4237] = 1'b0;
    assign outputs[4238] = layer0_outputs[3433];
    assign outputs[4239] = (layer0_outputs[411]) & ~(layer0_outputs[5446]);
    assign outputs[4240] = ~(layer0_outputs[2189]);
    assign outputs[4241] = ~((layer0_outputs[2678]) ^ (layer0_outputs[2334]));
    assign outputs[4242] = ~(layer0_outputs[9403]);
    assign outputs[4243] = layer0_outputs[2229];
    assign outputs[4244] = ~((layer0_outputs[7675]) ^ (layer0_outputs[5350]));
    assign outputs[4245] = ~((layer0_outputs[6971]) & (layer0_outputs[8500]));
    assign outputs[4246] = (layer0_outputs[6187]) & (layer0_outputs[2897]);
    assign outputs[4247] = ~((layer0_outputs[9975]) | (layer0_outputs[5766]));
    assign outputs[4248] = (layer0_outputs[1979]) & ~(layer0_outputs[1354]);
    assign outputs[4249] = (layer0_outputs[216]) ^ (layer0_outputs[5753]);
    assign outputs[4250] = (layer0_outputs[8598]) | (layer0_outputs[3124]);
    assign outputs[4251] = (layer0_outputs[4222]) ^ (layer0_outputs[1064]);
    assign outputs[4252] = (layer0_outputs[5006]) | (layer0_outputs[672]);
    assign outputs[4253] = (layer0_outputs[8024]) & ~(layer0_outputs[3819]);
    assign outputs[4254] = 1'b0;
    assign outputs[4255] = layer0_outputs[5196];
    assign outputs[4256] = ~((layer0_outputs[9307]) | (layer0_outputs[5011]));
    assign outputs[4257] = (layer0_outputs[7683]) ^ (layer0_outputs[5726]);
    assign outputs[4258] = (layer0_outputs[527]) & ~(layer0_outputs[5214]);
    assign outputs[4259] = ~(layer0_outputs[2734]);
    assign outputs[4260] = ~(layer0_outputs[6355]);
    assign outputs[4261] = (layer0_outputs[9131]) ^ (layer0_outputs[2906]);
    assign outputs[4262] = ~(layer0_outputs[2328]);
    assign outputs[4263] = ~(layer0_outputs[3595]);
    assign outputs[4264] = (layer0_outputs[3707]) & ~(layer0_outputs[4284]);
    assign outputs[4265] = (layer0_outputs[8648]) & ~(layer0_outputs[4678]);
    assign outputs[4266] = ~(layer0_outputs[8193]);
    assign outputs[4267] = ~(layer0_outputs[9537]);
    assign outputs[4268] = (layer0_outputs[7446]) | (layer0_outputs[7455]);
    assign outputs[4269] = ~(layer0_outputs[7673]) | (layer0_outputs[8837]);
    assign outputs[4270] = 1'b0;
    assign outputs[4271] = layer0_outputs[5990];
    assign outputs[4272] = ~(layer0_outputs[2488]);
    assign outputs[4273] = (layer0_outputs[155]) ^ (layer0_outputs[5694]);
    assign outputs[4274] = (layer0_outputs[211]) & (layer0_outputs[9816]);
    assign outputs[4275] = (layer0_outputs[7089]) & (layer0_outputs[7716]);
    assign outputs[4276] = ~(layer0_outputs[7007]);
    assign outputs[4277] = ~((layer0_outputs[842]) ^ (layer0_outputs[7222]));
    assign outputs[4278] = layer0_outputs[7362];
    assign outputs[4279] = ~((layer0_outputs[3091]) ^ (layer0_outputs[7862]));
    assign outputs[4280] = ~(layer0_outputs[1787]);
    assign outputs[4281] = ~(layer0_outputs[3192]);
    assign outputs[4282] = (layer0_outputs[1688]) & (layer0_outputs[6133]);
    assign outputs[4283] = ~(layer0_outputs[6107]) | (layer0_outputs[6443]);
    assign outputs[4284] = ~(layer0_outputs[9838]) | (layer0_outputs[7971]);
    assign outputs[4285] = layer0_outputs[6543];
    assign outputs[4286] = ~(layer0_outputs[5635]);
    assign outputs[4287] = (layer0_outputs[7166]) & ~(layer0_outputs[4556]);
    assign outputs[4288] = layer0_outputs[2458];
    assign outputs[4289] = ~(layer0_outputs[7505]);
    assign outputs[4290] = (layer0_outputs[8172]) & ~(layer0_outputs[695]);
    assign outputs[4291] = (layer0_outputs[691]) ^ (layer0_outputs[6513]);
    assign outputs[4292] = ~(layer0_outputs[6081]) | (layer0_outputs[4803]);
    assign outputs[4293] = ~((layer0_outputs[3326]) ^ (layer0_outputs[2566]));
    assign outputs[4294] = (layer0_outputs[6080]) & (layer0_outputs[1513]);
    assign outputs[4295] = ~(layer0_outputs[4053]);
    assign outputs[4296] = (layer0_outputs[1190]) & (layer0_outputs[2529]);
    assign outputs[4297] = layer0_outputs[8643];
    assign outputs[4298] = layer0_outputs[7250];
    assign outputs[4299] = layer0_outputs[7826];
    assign outputs[4300] = (layer0_outputs[62]) & ~(layer0_outputs[8865]);
    assign outputs[4301] = (layer0_outputs[8732]) & (layer0_outputs[1583]);
    assign outputs[4302] = (layer0_outputs[5319]) & ~(layer0_outputs[177]);
    assign outputs[4303] = (layer0_outputs[5738]) & (layer0_outputs[7523]);
    assign outputs[4304] = (layer0_outputs[5657]) & ~(layer0_outputs[6243]);
    assign outputs[4305] = layer0_outputs[5739];
    assign outputs[4306] = (layer0_outputs[6262]) & (layer0_outputs[1999]);
    assign outputs[4307] = ~(layer0_outputs[1365]);
    assign outputs[4308] = (layer0_outputs[9050]) & ~(layer0_outputs[926]);
    assign outputs[4309] = layer0_outputs[4552];
    assign outputs[4310] = (layer0_outputs[7899]) & (layer0_outputs[8155]);
    assign outputs[4311] = (layer0_outputs[7641]) ^ (layer0_outputs[4360]);
    assign outputs[4312] = layer0_outputs[2413];
    assign outputs[4313] = ~((layer0_outputs[2365]) ^ (layer0_outputs[3292]));
    assign outputs[4314] = ~((layer0_outputs[7228]) ^ (layer0_outputs[1035]));
    assign outputs[4315] = (layer0_outputs[6963]) ^ (layer0_outputs[1062]);
    assign outputs[4316] = (layer0_outputs[3797]) & ~(layer0_outputs[9228]);
    assign outputs[4317] = ~((layer0_outputs[6677]) | (layer0_outputs[8424]));
    assign outputs[4318] = ~((layer0_outputs[5759]) ^ (layer0_outputs[7908]));
    assign outputs[4319] = layer0_outputs[6264];
    assign outputs[4320] = (layer0_outputs[6512]) & ~(layer0_outputs[744]);
    assign outputs[4321] = ~((layer0_outputs[4810]) | (layer0_outputs[4003]));
    assign outputs[4322] = ~((layer0_outputs[7127]) & (layer0_outputs[5128]));
    assign outputs[4323] = ~((layer0_outputs[2077]) | (layer0_outputs[9255]));
    assign outputs[4324] = ~((layer0_outputs[729]) ^ (layer0_outputs[2186]));
    assign outputs[4325] = layer0_outputs[6358];
    assign outputs[4326] = layer0_outputs[4796];
    assign outputs[4327] = (layer0_outputs[4544]) ^ (layer0_outputs[4620]);
    assign outputs[4328] = ~((layer0_outputs[9924]) | (layer0_outputs[1073]));
    assign outputs[4329] = ~((layer0_outputs[6122]) ^ (layer0_outputs[1958]));
    assign outputs[4330] = layer0_outputs[644];
    assign outputs[4331] = ~((layer0_outputs[6362]) | (layer0_outputs[2934]));
    assign outputs[4332] = ~((layer0_outputs[817]) ^ (layer0_outputs[7177]));
    assign outputs[4333] = ~((layer0_outputs[6327]) | (layer0_outputs[6608]));
    assign outputs[4334] = layer0_outputs[7005];
    assign outputs[4335] = ~(layer0_outputs[1878]);
    assign outputs[4336] = (layer0_outputs[9740]) & ~(layer0_outputs[3286]);
    assign outputs[4337] = ~((layer0_outputs[999]) | (layer0_outputs[1054]));
    assign outputs[4338] = ~((layer0_outputs[7097]) ^ (layer0_outputs[9463]));
    assign outputs[4339] = (layer0_outputs[7118]) ^ (layer0_outputs[4696]);
    assign outputs[4340] = layer0_outputs[3773];
    assign outputs[4341] = layer0_outputs[9953];
    assign outputs[4342] = (layer0_outputs[2124]) ^ (layer0_outputs[6606]);
    assign outputs[4343] = ~(layer0_outputs[7799]);
    assign outputs[4344] = (layer0_outputs[5632]) ^ (layer0_outputs[7585]);
    assign outputs[4345] = ~((layer0_outputs[6321]) | (layer0_outputs[8313]));
    assign outputs[4346] = ~(layer0_outputs[1556]);
    assign outputs[4347] = (layer0_outputs[6271]) ^ (layer0_outputs[2820]);
    assign outputs[4348] = (layer0_outputs[5464]) & ~(layer0_outputs[2079]);
    assign outputs[4349] = ~((layer0_outputs[9327]) ^ (layer0_outputs[1263]));
    assign outputs[4350] = ~((layer0_outputs[3492]) ^ (layer0_outputs[3609]));
    assign outputs[4351] = ~((layer0_outputs[6054]) ^ (layer0_outputs[9193]));
    assign outputs[4352] = layer0_outputs[6321];
    assign outputs[4353] = layer0_outputs[5179];
    assign outputs[4354] = (layer0_outputs[3818]) & (layer0_outputs[2423]);
    assign outputs[4355] = ~(layer0_outputs[8861]);
    assign outputs[4356] = ~(layer0_outputs[9579]);
    assign outputs[4357] = ~(layer0_outputs[5059]);
    assign outputs[4358] = ~(layer0_outputs[6064]);
    assign outputs[4359] = ~((layer0_outputs[3650]) ^ (layer0_outputs[403]));
    assign outputs[4360] = ~(layer0_outputs[7057]);
    assign outputs[4361] = layer0_outputs[2370];
    assign outputs[4362] = ~((layer0_outputs[671]) | (layer0_outputs[5227]));
    assign outputs[4363] = (layer0_outputs[5516]) ^ (layer0_outputs[9242]);
    assign outputs[4364] = (layer0_outputs[4927]) & (layer0_outputs[328]);
    assign outputs[4365] = layer0_outputs[3670];
    assign outputs[4366] = (layer0_outputs[4769]) & ~(layer0_outputs[6248]);
    assign outputs[4367] = layer0_outputs[1396];
    assign outputs[4368] = ~(layer0_outputs[5270]);
    assign outputs[4369] = ~((layer0_outputs[7586]) ^ (layer0_outputs[3728]));
    assign outputs[4370] = layer0_outputs[4687];
    assign outputs[4371] = (layer0_outputs[9839]) ^ (layer0_outputs[6958]);
    assign outputs[4372] = ~((layer0_outputs[5028]) ^ (layer0_outputs[798]));
    assign outputs[4373] = (layer0_outputs[8078]) & ~(layer0_outputs[2115]);
    assign outputs[4374] = ~(layer0_outputs[3789]);
    assign outputs[4375] = (layer0_outputs[2069]) ^ (layer0_outputs[3324]);
    assign outputs[4376] = ~((layer0_outputs[8547]) ^ (layer0_outputs[9544]));
    assign outputs[4377] = ~((layer0_outputs[2970]) ^ (layer0_outputs[5887]));
    assign outputs[4378] = ~(layer0_outputs[1341]);
    assign outputs[4379] = ~((layer0_outputs[9650]) ^ (layer0_outputs[3981]));
    assign outputs[4380] = ~((layer0_outputs[1581]) ^ (layer0_outputs[5955]));
    assign outputs[4381] = layer0_outputs[9277];
    assign outputs[4382] = (layer0_outputs[3749]) ^ (layer0_outputs[6216]);
    assign outputs[4383] = ~((layer0_outputs[970]) ^ (layer0_outputs[9713]));
    assign outputs[4384] = ~(layer0_outputs[1268]);
    assign outputs[4385] = ~(layer0_outputs[4817]);
    assign outputs[4386] = ~(layer0_outputs[6622]);
    assign outputs[4387] = ~((layer0_outputs[3603]) | (layer0_outputs[782]));
    assign outputs[4388] = 1'b0;
    assign outputs[4389] = (layer0_outputs[1082]) & ~(layer0_outputs[6433]);
    assign outputs[4390] = ~((layer0_outputs[4408]) ^ (layer0_outputs[5763]));
    assign outputs[4391] = (layer0_outputs[3828]) & ~(layer0_outputs[29]);
    assign outputs[4392] = ~((layer0_outputs[1690]) | (layer0_outputs[9147]));
    assign outputs[4393] = ~(layer0_outputs[9736]);
    assign outputs[4394] = ~((layer0_outputs[7904]) ^ (layer0_outputs[6130]));
    assign outputs[4395] = ~(layer0_outputs[2683]) | (layer0_outputs[4410]);
    assign outputs[4396] = (layer0_outputs[4747]) ^ (layer0_outputs[8035]);
    assign outputs[4397] = (layer0_outputs[2901]) ^ (layer0_outputs[6290]);
    assign outputs[4398] = layer0_outputs[3807];
    assign outputs[4399] = layer0_outputs[6380];
    assign outputs[4400] = layer0_outputs[2351];
    assign outputs[4401] = (layer0_outputs[8160]) & (layer0_outputs[5449]);
    assign outputs[4402] = (layer0_outputs[7628]) ^ (layer0_outputs[8531]);
    assign outputs[4403] = layer0_outputs[10139];
    assign outputs[4404] = ~(layer0_outputs[9747]);
    assign outputs[4405] = (layer0_outputs[2468]) ^ (layer0_outputs[1413]);
    assign outputs[4406] = ~((layer0_outputs[6615]) ^ (layer0_outputs[5129]));
    assign outputs[4407] = ~((layer0_outputs[4092]) | (layer0_outputs[9681]));
    assign outputs[4408] = layer0_outputs[1518];
    assign outputs[4409] = (layer0_outputs[5596]) & (layer0_outputs[5531]);
    assign outputs[4410] = ~(layer0_outputs[8042]);
    assign outputs[4411] = ~((layer0_outputs[9256]) ^ (layer0_outputs[1207]));
    assign outputs[4412] = ~(layer0_outputs[8306]);
    assign outputs[4413] = ~(layer0_outputs[1654]);
    assign outputs[4414] = ~((layer0_outputs[315]) ^ (layer0_outputs[7426]));
    assign outputs[4415] = (layer0_outputs[1826]) & ~(layer0_outputs[4975]);
    assign outputs[4416] = (layer0_outputs[9453]) & ~(layer0_outputs[1085]);
    assign outputs[4417] = ~(layer0_outputs[9166]);
    assign outputs[4418] = layer0_outputs[2921];
    assign outputs[4419] = (layer0_outputs[1752]) & ~(layer0_outputs[6031]);
    assign outputs[4420] = ~(layer0_outputs[9297]) | (layer0_outputs[6986]);
    assign outputs[4421] = (layer0_outputs[10084]) & (layer0_outputs[1302]);
    assign outputs[4422] = ~(layer0_outputs[3552]);
    assign outputs[4423] = (layer0_outputs[9107]) ^ (layer0_outputs[9145]);
    assign outputs[4424] = ~(layer0_outputs[5670]);
    assign outputs[4425] = ~((layer0_outputs[9430]) ^ (layer0_outputs[132]));
    assign outputs[4426] = ~((layer0_outputs[6956]) ^ (layer0_outputs[4358]));
    assign outputs[4427] = ~(layer0_outputs[4078]);
    assign outputs[4428] = ~(layer0_outputs[402]);
    assign outputs[4429] = (layer0_outputs[9163]) ^ (layer0_outputs[4371]);
    assign outputs[4430] = ~(layer0_outputs[5093]);
    assign outputs[4431] = ~(layer0_outputs[3320]);
    assign outputs[4432] = ~((layer0_outputs[9473]) ^ (layer0_outputs[5003]));
    assign outputs[4433] = (layer0_outputs[4747]) & (layer0_outputs[7642]);
    assign outputs[4434] = ~(layer0_outputs[9609]);
    assign outputs[4435] = (layer0_outputs[9727]) & ~(layer0_outputs[1621]);
    assign outputs[4436] = (layer0_outputs[2801]) ^ (layer0_outputs[2617]);
    assign outputs[4437] = (layer0_outputs[1461]) ^ (layer0_outputs[6852]);
    assign outputs[4438] = ~(layer0_outputs[873]) | (layer0_outputs[9521]);
    assign outputs[4439] = layer0_outputs[2944];
    assign outputs[4440] = ~(layer0_outputs[2431]);
    assign outputs[4441] = (layer0_outputs[455]) ^ (layer0_outputs[5467]);
    assign outputs[4442] = ~((layer0_outputs[554]) & (layer0_outputs[3339]));
    assign outputs[4443] = ~(layer0_outputs[1362]);
    assign outputs[4444] = ~(layer0_outputs[6089]);
    assign outputs[4445] = (layer0_outputs[2623]) ^ (layer0_outputs[2756]);
    assign outputs[4446] = ~((layer0_outputs[2314]) ^ (layer0_outputs[678]));
    assign outputs[4447] = layer0_outputs[3871];
    assign outputs[4448] = (layer0_outputs[4108]) ^ (layer0_outputs[1763]);
    assign outputs[4449] = ~(layer0_outputs[8321]);
    assign outputs[4450] = (layer0_outputs[6907]) & ~(layer0_outputs[4054]);
    assign outputs[4451] = ~((layer0_outputs[7416]) ^ (layer0_outputs[9228]));
    assign outputs[4452] = ~(layer0_outputs[9818]);
    assign outputs[4453] = ~((layer0_outputs[9686]) ^ (layer0_outputs[1505]));
    assign outputs[4454] = (layer0_outputs[7854]) & (layer0_outputs[3907]);
    assign outputs[4455] = layer0_outputs[2824];
    assign outputs[4456] = ~((layer0_outputs[6377]) ^ (layer0_outputs[5385]));
    assign outputs[4457] = (layer0_outputs[2833]) ^ (layer0_outputs[9185]);
    assign outputs[4458] = (layer0_outputs[1530]) ^ (layer0_outputs[4268]);
    assign outputs[4459] = layer0_outputs[1389];
    assign outputs[4460] = layer0_outputs[173];
    assign outputs[4461] = ~((layer0_outputs[2079]) | (layer0_outputs[243]));
    assign outputs[4462] = (layer0_outputs[1091]) ^ (layer0_outputs[2744]);
    assign outputs[4463] = layer0_outputs[6841];
    assign outputs[4464] = ~(layer0_outputs[9160]);
    assign outputs[4465] = ~(layer0_outputs[1545]);
    assign outputs[4466] = ~(layer0_outputs[2845]);
    assign outputs[4467] = layer0_outputs[9132];
    assign outputs[4468] = (layer0_outputs[6079]) & ~(layer0_outputs[8545]);
    assign outputs[4469] = (layer0_outputs[4931]) & ~(layer0_outputs[7379]);
    assign outputs[4470] = ~((layer0_outputs[7723]) | (layer0_outputs[7666]));
    assign outputs[4471] = (layer0_outputs[503]) | (layer0_outputs[2607]);
    assign outputs[4472] = (layer0_outputs[5308]) ^ (layer0_outputs[2176]);
    assign outputs[4473] = layer0_outputs[3532];
    assign outputs[4474] = ~(layer0_outputs[7000]);
    assign outputs[4475] = (layer0_outputs[1249]) & ~(layer0_outputs[4513]);
    assign outputs[4476] = layer0_outputs[8146];
    assign outputs[4477] = (layer0_outputs[8468]) & (layer0_outputs[8760]);
    assign outputs[4478] = ~(layer0_outputs[9148]);
    assign outputs[4479] = layer0_outputs[4628];
    assign outputs[4480] = (layer0_outputs[10074]) & ~(layer0_outputs[1679]);
    assign outputs[4481] = ~((layer0_outputs[6943]) ^ (layer0_outputs[5908]));
    assign outputs[4482] = layer0_outputs[4718];
    assign outputs[4483] = ~((layer0_outputs[8999]) | (layer0_outputs[8468]));
    assign outputs[4484] = (layer0_outputs[3274]) & ~(layer0_outputs[1200]);
    assign outputs[4485] = ~(layer0_outputs[4483]) | (layer0_outputs[1796]);
    assign outputs[4486] = (layer0_outputs[4306]) & (layer0_outputs[1167]);
    assign outputs[4487] = layer0_outputs[1904];
    assign outputs[4488] = (layer0_outputs[4228]) & (layer0_outputs[8839]);
    assign outputs[4489] = layer0_outputs[5883];
    assign outputs[4490] = ~(layer0_outputs[2682]) | (layer0_outputs[7983]);
    assign outputs[4491] = ~(layer0_outputs[5870]);
    assign outputs[4492] = layer0_outputs[5773];
    assign outputs[4493] = ~((layer0_outputs[2239]) | (layer0_outputs[8586]));
    assign outputs[4494] = (layer0_outputs[2056]) ^ (layer0_outputs[6288]);
    assign outputs[4495] = ~((layer0_outputs[6984]) | (layer0_outputs[76]));
    assign outputs[4496] = layer0_outputs[1212];
    assign outputs[4497] = (layer0_outputs[9312]) & ~(layer0_outputs[2747]);
    assign outputs[4498] = (layer0_outputs[94]) | (layer0_outputs[5345]);
    assign outputs[4499] = (layer0_outputs[3526]) ^ (layer0_outputs[2109]);
    assign outputs[4500] = ~((layer0_outputs[9391]) ^ (layer0_outputs[8992]));
    assign outputs[4501] = ~((layer0_outputs[2860]) ^ (layer0_outputs[2983]));
    assign outputs[4502] = layer0_outputs[10007];
    assign outputs[4503] = ~((layer0_outputs[4211]) ^ (layer0_outputs[5758]));
    assign outputs[4504] = ~((layer0_outputs[4930]) ^ (layer0_outputs[1671]));
    assign outputs[4505] = ~((layer0_outputs[531]) ^ (layer0_outputs[6634]));
    assign outputs[4506] = ~(layer0_outputs[8706]);
    assign outputs[4507] = ~(layer0_outputs[7396]) | (layer0_outputs[3517]);
    assign outputs[4508] = (layer0_outputs[731]) ^ (layer0_outputs[5702]);
    assign outputs[4509] = ~((layer0_outputs[8727]) ^ (layer0_outputs[5841]));
    assign outputs[4510] = (layer0_outputs[7131]) ^ (layer0_outputs[7619]);
    assign outputs[4511] = (layer0_outputs[9593]) & ~(layer0_outputs[6734]);
    assign outputs[4512] = ~(layer0_outputs[2764]) | (layer0_outputs[2390]);
    assign outputs[4513] = ~(layer0_outputs[5891]);
    assign outputs[4514] = layer0_outputs[4204];
    assign outputs[4515] = ~((layer0_outputs[8178]) | (layer0_outputs[1555]));
    assign outputs[4516] = ~(layer0_outputs[6295]) | (layer0_outputs[6585]);
    assign outputs[4517] = ~(layer0_outputs[6597]);
    assign outputs[4518] = layer0_outputs[7377];
    assign outputs[4519] = layer0_outputs[5450];
    assign outputs[4520] = ~(layer0_outputs[1214]);
    assign outputs[4521] = ~(layer0_outputs[9697]) | (layer0_outputs[4626]);
    assign outputs[4522] = layer0_outputs[1281];
    assign outputs[4523] = ~(layer0_outputs[7593]);
    assign outputs[4524] = layer0_outputs[8668];
    assign outputs[4525] = ~((layer0_outputs[10148]) ^ (layer0_outputs[4663]));
    assign outputs[4526] = ~(layer0_outputs[7895]);
    assign outputs[4527] = (layer0_outputs[6578]) & ~(layer0_outputs[4523]);
    assign outputs[4528] = layer0_outputs[2805];
    assign outputs[4529] = ~(layer0_outputs[8564]);
    assign outputs[4530] = (layer0_outputs[9095]) ^ (layer0_outputs[87]);
    assign outputs[4531] = layer0_outputs[7477];
    assign outputs[4532] = (layer0_outputs[9336]) ^ (layer0_outputs[7535]);
    assign outputs[4533] = layer0_outputs[7649];
    assign outputs[4534] = (layer0_outputs[2012]) | (layer0_outputs[3833]);
    assign outputs[4535] = (layer0_outputs[7883]) ^ (layer0_outputs[6010]);
    assign outputs[4536] = ~((layer0_outputs[3136]) ^ (layer0_outputs[6989]));
    assign outputs[4537] = (layer0_outputs[3903]) ^ (layer0_outputs[4]);
    assign outputs[4538] = ~(layer0_outputs[3187]);
    assign outputs[4539] = ~((layer0_outputs[10024]) ^ (layer0_outputs[6476]));
    assign outputs[4540] = layer0_outputs[1823];
    assign outputs[4541] = ~(layer0_outputs[3187]);
    assign outputs[4542] = layer0_outputs[9299];
    assign outputs[4543] = layer0_outputs[3296];
    assign outputs[4544] = ~((layer0_outputs[8913]) & (layer0_outputs[8166]));
    assign outputs[4545] = (layer0_outputs[144]) ^ (layer0_outputs[971]);
    assign outputs[4546] = ~((layer0_outputs[8643]) ^ (layer0_outputs[7780]));
    assign outputs[4547] = ~(layer0_outputs[4383]);
    assign outputs[4548] = (layer0_outputs[8843]) ^ (layer0_outputs[9684]);
    assign outputs[4549] = ~(layer0_outputs[5455]);
    assign outputs[4550] = ~(layer0_outputs[8946]);
    assign outputs[4551] = ~((layer0_outputs[1482]) ^ (layer0_outputs[6297]));
    assign outputs[4552] = layer0_outputs[8456];
    assign outputs[4553] = ~((layer0_outputs[1177]) ^ (layer0_outputs[9213]));
    assign outputs[4554] = (layer0_outputs[5486]) & (layer0_outputs[6524]);
    assign outputs[4555] = layer0_outputs[1974];
    assign outputs[4556] = ~(layer0_outputs[9395]);
    assign outputs[4557] = ~(layer0_outputs[3853]);
    assign outputs[4558] = ~(layer0_outputs[8334]);
    assign outputs[4559] = layer0_outputs[6465];
    assign outputs[4560] = ~(layer0_outputs[2424]);
    assign outputs[4561] = layer0_outputs[245];
    assign outputs[4562] = layer0_outputs[235];
    assign outputs[4563] = ~(layer0_outputs[4291]);
    assign outputs[4564] = (layer0_outputs[4566]) | (layer0_outputs[3514]);
    assign outputs[4565] = ~(layer0_outputs[3835]);
    assign outputs[4566] = ~(layer0_outputs[2714]) | (layer0_outputs[5400]);
    assign outputs[4567] = ~(layer0_outputs[5192]);
    assign outputs[4568] = (layer0_outputs[2499]) ^ (layer0_outputs[1882]);
    assign outputs[4569] = (layer0_outputs[9905]) ^ (layer0_outputs[9800]);
    assign outputs[4570] = ~((layer0_outputs[1068]) | (layer0_outputs[9449]));
    assign outputs[4571] = ~((layer0_outputs[5402]) ^ (layer0_outputs[10140]));
    assign outputs[4572] = ~(layer0_outputs[1171]);
    assign outputs[4573] = (layer0_outputs[1444]) & (layer0_outputs[7991]);
    assign outputs[4574] = (layer0_outputs[2231]) ^ (layer0_outputs[10199]);
    assign outputs[4575] = ~(layer0_outputs[451]) | (layer0_outputs[6936]);
    assign outputs[4576] = ~(layer0_outputs[9348]);
    assign outputs[4577] = (layer0_outputs[5226]) ^ (layer0_outputs[1013]);
    assign outputs[4578] = ~((layer0_outputs[9609]) | (layer0_outputs[6505]));
    assign outputs[4579] = ~(layer0_outputs[5169]);
    assign outputs[4580] = (layer0_outputs[3138]) ^ (layer0_outputs[4661]);
    assign outputs[4581] = ~(layer0_outputs[10147]);
    assign outputs[4582] = ~(layer0_outputs[7515]);
    assign outputs[4583] = layer0_outputs[8652];
    assign outputs[4584] = (layer0_outputs[4414]) ^ (layer0_outputs[5644]);
    assign outputs[4585] = (layer0_outputs[9816]) & ~(layer0_outputs[572]);
    assign outputs[4586] = ~(layer0_outputs[9863]);
    assign outputs[4587] = ~(layer0_outputs[5457]);
    assign outputs[4588] = layer0_outputs[8433];
    assign outputs[4589] = (layer0_outputs[7860]) ^ (layer0_outputs[1548]);
    assign outputs[4590] = ~((layer0_outputs[1862]) ^ (layer0_outputs[686]));
    assign outputs[4591] = (layer0_outputs[830]) ^ (layer0_outputs[2049]);
    assign outputs[4592] = (layer0_outputs[6743]) ^ (layer0_outputs[9946]);
    assign outputs[4593] = ~(layer0_outputs[468]) | (layer0_outputs[792]);
    assign outputs[4594] = layer0_outputs[2558];
    assign outputs[4595] = layer0_outputs[3222];
    assign outputs[4596] = layer0_outputs[6738];
    assign outputs[4597] = ~(layer0_outputs[4963]);
    assign outputs[4598] = ~(layer0_outputs[9287]);
    assign outputs[4599] = ~(layer0_outputs[4832]);
    assign outputs[4600] = ~((layer0_outputs[6092]) ^ (layer0_outputs[3213]));
    assign outputs[4601] = (layer0_outputs[5359]) ^ (layer0_outputs[10219]);
    assign outputs[4602] = ~(layer0_outputs[8022]);
    assign outputs[4603] = (layer0_outputs[4862]) & ~(layer0_outputs[9171]);
    assign outputs[4604] = layer0_outputs[673];
    assign outputs[4605] = ~((layer0_outputs[646]) ^ (layer0_outputs[6654]));
    assign outputs[4606] = layer0_outputs[1160];
    assign outputs[4607] = (layer0_outputs[4640]) | (layer0_outputs[3947]);
    assign outputs[4608] = (layer0_outputs[2708]) & (layer0_outputs[500]);
    assign outputs[4609] = (layer0_outputs[1280]) ^ (layer0_outputs[8250]);
    assign outputs[4610] = layer0_outputs[701];
    assign outputs[4611] = ~((layer0_outputs[4667]) ^ (layer0_outputs[8875]));
    assign outputs[4612] = (layer0_outputs[3845]) & ~(layer0_outputs[8412]);
    assign outputs[4613] = ~(layer0_outputs[3151]);
    assign outputs[4614] = ~((layer0_outputs[4872]) | (layer0_outputs[2275]));
    assign outputs[4615] = layer0_outputs[2558];
    assign outputs[4616] = ~(layer0_outputs[6935]);
    assign outputs[4617] = (layer0_outputs[8639]) ^ (layer0_outputs[9096]);
    assign outputs[4618] = ~(layer0_outputs[2196]);
    assign outputs[4619] = ~(layer0_outputs[6603]);
    assign outputs[4620] = ~(layer0_outputs[9006]);
    assign outputs[4621] = ~((layer0_outputs[9423]) ^ (layer0_outputs[8132]));
    assign outputs[4622] = layer0_outputs[3056];
    assign outputs[4623] = ~(layer0_outputs[5567]) | (layer0_outputs[5493]);
    assign outputs[4624] = ~((layer0_outputs[7029]) | (layer0_outputs[8090]));
    assign outputs[4625] = (layer0_outputs[766]) & ~(layer0_outputs[8138]);
    assign outputs[4626] = ~(layer0_outputs[4091]) | (layer0_outputs[5685]);
    assign outputs[4627] = layer0_outputs[4541];
    assign outputs[4628] = (layer0_outputs[6651]) ^ (layer0_outputs[3263]);
    assign outputs[4629] = ~((layer0_outputs[6417]) ^ (layer0_outputs[8563]));
    assign outputs[4630] = layer0_outputs[3459];
    assign outputs[4631] = layer0_outputs[5708];
    assign outputs[4632] = (layer0_outputs[2028]) ^ (layer0_outputs[3844]);
    assign outputs[4633] = layer0_outputs[10109];
    assign outputs[4634] = (layer0_outputs[8780]) ^ (layer0_outputs[3952]);
    assign outputs[4635] = (layer0_outputs[9009]) ^ (layer0_outputs[1993]);
    assign outputs[4636] = (layer0_outputs[3183]) ^ (layer0_outputs[3865]);
    assign outputs[4637] = ~(layer0_outputs[7321]);
    assign outputs[4638] = ~((layer0_outputs[109]) | (layer0_outputs[9998]));
    assign outputs[4639] = (layer0_outputs[9730]) & ~(layer0_outputs[9621]);
    assign outputs[4640] = ~(layer0_outputs[1071]);
    assign outputs[4641] = layer0_outputs[9175];
    assign outputs[4642] = (layer0_outputs[3069]) ^ (layer0_outputs[5108]);
    assign outputs[4643] = (layer0_outputs[4223]) ^ (layer0_outputs[4694]);
    assign outputs[4644] = layer0_outputs[8106];
    assign outputs[4645] = (layer0_outputs[1762]) | (layer0_outputs[3243]);
    assign outputs[4646] = (layer0_outputs[7570]) & ~(layer0_outputs[5784]);
    assign outputs[4647] = layer0_outputs[1873];
    assign outputs[4648] = (layer0_outputs[6825]) & (layer0_outputs[5631]);
    assign outputs[4649] = ~((layer0_outputs[4881]) | (layer0_outputs[2934]));
    assign outputs[4650] = ~(layer0_outputs[9025]);
    assign outputs[4651] = (layer0_outputs[2923]) & (layer0_outputs[2484]);
    assign outputs[4652] = layer0_outputs[5729];
    assign outputs[4653] = (layer0_outputs[6322]) ^ (layer0_outputs[5506]);
    assign outputs[4654] = ~(layer0_outputs[410]);
    assign outputs[4655] = ~((layer0_outputs[3313]) | (layer0_outputs[8953]));
    assign outputs[4656] = ~(layer0_outputs[10043]);
    assign outputs[4657] = ~(layer0_outputs[5313]);
    assign outputs[4658] = (layer0_outputs[4066]) & (layer0_outputs[9972]);
    assign outputs[4659] = (layer0_outputs[5653]) ^ (layer0_outputs[5934]);
    assign outputs[4660] = ~(layer0_outputs[2552]);
    assign outputs[4661] = ~(layer0_outputs[10073]) | (layer0_outputs[217]);
    assign outputs[4662] = ~(layer0_outputs[6568]);
    assign outputs[4663] = 1'b0;
    assign outputs[4664] = ~(layer0_outputs[10159]);
    assign outputs[4665] = ~(layer0_outputs[4021]);
    assign outputs[4666] = (layer0_outputs[4726]) ^ (layer0_outputs[242]);
    assign outputs[4667] = ~((layer0_outputs[4665]) ^ (layer0_outputs[3444]));
    assign outputs[4668] = layer0_outputs[2868];
    assign outputs[4669] = ~(layer0_outputs[5051]);
    assign outputs[4670] = (layer0_outputs[6897]) ^ (layer0_outputs[5490]);
    assign outputs[4671] = (layer0_outputs[236]) ^ (layer0_outputs[3905]);
    assign outputs[4672] = ~(layer0_outputs[7301]);
    assign outputs[4673] = ~(layer0_outputs[10187]);
    assign outputs[4674] = 1'b0;
    assign outputs[4675] = layer0_outputs[9911];
    assign outputs[4676] = (layer0_outputs[6698]) & ~(layer0_outputs[1115]);
    assign outputs[4677] = (layer0_outputs[5171]) ^ (layer0_outputs[188]);
    assign outputs[4678] = (layer0_outputs[5683]) & ~(layer0_outputs[2241]);
    assign outputs[4679] = layer0_outputs[4498];
    assign outputs[4680] = (layer0_outputs[6806]) & ~(layer0_outputs[1237]);
    assign outputs[4681] = ~(layer0_outputs[6755]);
    assign outputs[4682] = (layer0_outputs[9130]) & ~(layer0_outputs[837]);
    assign outputs[4683] = (layer0_outputs[1132]) & (layer0_outputs[7733]);
    assign outputs[4684] = layer0_outputs[4270];
    assign outputs[4685] = ~(layer0_outputs[8954]);
    assign outputs[4686] = ~(layer0_outputs[6228]);
    assign outputs[4687] = ~(layer0_outputs[3630]) | (layer0_outputs[5010]);
    assign outputs[4688] = (layer0_outputs[6536]) | (layer0_outputs[4209]);
    assign outputs[4689] = ~(layer0_outputs[5184]);
    assign outputs[4690] = ~(layer0_outputs[5740]);
    assign outputs[4691] = (layer0_outputs[5554]) & (layer0_outputs[9344]);
    assign outputs[4692] = ~(layer0_outputs[1464]);
    assign outputs[4693] = layer0_outputs[2589];
    assign outputs[4694] = ~((layer0_outputs[5641]) ^ (layer0_outputs[3696]));
    assign outputs[4695] = ~(layer0_outputs[5040]);
    assign outputs[4696] = ~(layer0_outputs[458]);
    assign outputs[4697] = (layer0_outputs[3872]) & ~(layer0_outputs[7090]);
    assign outputs[4698] = ~((layer0_outputs[9897]) | (layer0_outputs[8396]));
    assign outputs[4699] = ~((layer0_outputs[5160]) ^ (layer0_outputs[7957]));
    assign outputs[4700] = ~((layer0_outputs[8177]) ^ (layer0_outputs[9679]));
    assign outputs[4701] = ~(layer0_outputs[4808]);
    assign outputs[4702] = (layer0_outputs[4386]) & ~(layer0_outputs[294]);
    assign outputs[4703] = ~((layer0_outputs[9988]) ^ (layer0_outputs[2199]));
    assign outputs[4704] = ~((layer0_outputs[9567]) | (layer0_outputs[3331]));
    assign outputs[4705] = layer0_outputs[1014];
    assign outputs[4706] = (layer0_outputs[6224]) | (layer0_outputs[5650]);
    assign outputs[4707] = ~((layer0_outputs[4549]) | (layer0_outputs[9293]));
    assign outputs[4708] = layer0_outputs[7229];
    assign outputs[4709] = ~((layer0_outputs[4656]) ^ (layer0_outputs[2529]));
    assign outputs[4710] = ~(layer0_outputs[2068]);
    assign outputs[4711] = ~(layer0_outputs[8661]);
    assign outputs[4712] = layer0_outputs[5173];
    assign outputs[4713] = ~((layer0_outputs[1427]) | (layer0_outputs[8185]));
    assign outputs[4714] = ~(layer0_outputs[3094]);
    assign outputs[4715] = ~(layer0_outputs[5894]);
    assign outputs[4716] = (layer0_outputs[701]) & ~(layer0_outputs[5511]);
    assign outputs[4717] = (layer0_outputs[6042]) ^ (layer0_outputs[9227]);
    assign outputs[4718] = (layer0_outputs[3548]) & ~(layer0_outputs[2532]);
    assign outputs[4719] = ~(layer0_outputs[678]);
    assign outputs[4720] = ~(layer0_outputs[5867]) | (layer0_outputs[2569]);
    assign outputs[4721] = (layer0_outputs[1734]) | (layer0_outputs[9608]);
    assign outputs[4722] = layer0_outputs[6881];
    assign outputs[4723] = layer0_outputs[5324];
    assign outputs[4724] = ~((layer0_outputs[1921]) | (layer0_outputs[8291]));
    assign outputs[4725] = layer0_outputs[4627];
    assign outputs[4726] = ~(layer0_outputs[3531]) | (layer0_outputs[7660]);
    assign outputs[4727] = ~((layer0_outputs[4476]) & (layer0_outputs[6328]));
    assign outputs[4728] = (layer0_outputs[2265]) | (layer0_outputs[6463]);
    assign outputs[4729] = (layer0_outputs[9842]) & (layer0_outputs[697]);
    assign outputs[4730] = (layer0_outputs[6257]) & (layer0_outputs[4446]);
    assign outputs[4731] = (layer0_outputs[5827]) ^ (layer0_outputs[5718]);
    assign outputs[4732] = ~((layer0_outputs[8796]) ^ (layer0_outputs[8531]));
    assign outputs[4733] = ~(layer0_outputs[1451]);
    assign outputs[4734] = ~((layer0_outputs[6164]) & (layer0_outputs[8765]));
    assign outputs[4735] = (layer0_outputs[4514]) & ~(layer0_outputs[1735]);
    assign outputs[4736] = ~(layer0_outputs[924]) | (layer0_outputs[464]);
    assign outputs[4737] = ~((layer0_outputs[9850]) ^ (layer0_outputs[3763]));
    assign outputs[4738] = (layer0_outputs[7489]) & ~(layer0_outputs[2221]);
    assign outputs[4739] = ~((layer0_outputs[3146]) ^ (layer0_outputs[3356]));
    assign outputs[4740] = layer0_outputs[4052];
    assign outputs[4741] = ~((layer0_outputs[699]) ^ (layer0_outputs[6289]));
    assign outputs[4742] = (layer0_outputs[8233]) ^ (layer0_outputs[7]);
    assign outputs[4743] = (layer0_outputs[7567]) & ~(layer0_outputs[7037]);
    assign outputs[4744] = layer0_outputs[863];
    assign outputs[4745] = ~(layer0_outputs[5271]);
    assign outputs[4746] = ~((layer0_outputs[6379]) ^ (layer0_outputs[4388]));
    assign outputs[4747] = ~((layer0_outputs[738]) ^ (layer0_outputs[4393]));
    assign outputs[4748] = ~((layer0_outputs[8670]) | (layer0_outputs[1588]));
    assign outputs[4749] = layer0_outputs[5848];
    assign outputs[4750] = layer0_outputs[3013];
    assign outputs[4751] = (layer0_outputs[5780]) | (layer0_outputs[4977]);
    assign outputs[4752] = ~((layer0_outputs[1044]) | (layer0_outputs[8284]));
    assign outputs[4753] = (layer0_outputs[8962]) & ~(layer0_outputs[1601]);
    assign outputs[4754] = layer0_outputs[8878];
    assign outputs[4755] = ~(layer0_outputs[7987]);
    assign outputs[4756] = ~(layer0_outputs[2405]);
    assign outputs[4757] = (layer0_outputs[9604]) ^ (layer0_outputs[4612]);
    assign outputs[4758] = ~((layer0_outputs[5168]) ^ (layer0_outputs[2992]));
    assign outputs[4759] = layer0_outputs[4376];
    assign outputs[4760] = ~((layer0_outputs[1800]) ^ (layer0_outputs[7962]));
    assign outputs[4761] = ~(layer0_outputs[280]);
    assign outputs[4762] = ~(layer0_outputs[9569]) | (layer0_outputs[8713]);
    assign outputs[4763] = layer0_outputs[9866];
    assign outputs[4764] = (layer0_outputs[5076]) & (layer0_outputs[5619]);
    assign outputs[4765] = (layer0_outputs[457]) & (layer0_outputs[8311]);
    assign outputs[4766] = ~((layer0_outputs[8521]) & (layer0_outputs[1192]));
    assign outputs[4767] = (layer0_outputs[5482]) | (layer0_outputs[5780]);
    assign outputs[4768] = (layer0_outputs[6873]) ^ (layer0_outputs[7978]);
    assign outputs[4769] = (layer0_outputs[8403]) | (layer0_outputs[12]);
    assign outputs[4770] = (layer0_outputs[1421]) ^ (layer0_outputs[2841]);
    assign outputs[4771] = ~(layer0_outputs[3782]);
    assign outputs[4772] = ~((layer0_outputs[1609]) ^ (layer0_outputs[3153]));
    assign outputs[4773] = layer0_outputs[4552];
    assign outputs[4774] = (layer0_outputs[4849]) ^ (layer0_outputs[7634]);
    assign outputs[4775] = layer0_outputs[1858];
    assign outputs[4776] = (layer0_outputs[1723]) ^ (layer0_outputs[8483]);
    assign outputs[4777] = ~(layer0_outputs[8330]);
    assign outputs[4778] = (layer0_outputs[7793]) & ~(layer0_outputs[9951]);
    assign outputs[4779] = ~((layer0_outputs[9565]) ^ (layer0_outputs[1590]));
    assign outputs[4780] = layer0_outputs[1804];
    assign outputs[4781] = layer0_outputs[4983];
    assign outputs[4782] = layer0_outputs[6927];
    assign outputs[4783] = (layer0_outputs[3068]) & ~(layer0_outputs[5045]);
    assign outputs[4784] = (layer0_outputs[9549]) & ~(layer0_outputs[480]);
    assign outputs[4785] = ~(layer0_outputs[5270]);
    assign outputs[4786] = ~((layer0_outputs[1693]) | (layer0_outputs[3384]));
    assign outputs[4787] = ~((layer0_outputs[7825]) ^ (layer0_outputs[9351]));
    assign outputs[4788] = layer0_outputs[3430];
    assign outputs[4789] = layer0_outputs[2961];
    assign outputs[4790] = ~((layer0_outputs[10064]) ^ (layer0_outputs[1022]));
    assign outputs[4791] = ~((layer0_outputs[2346]) ^ (layer0_outputs[7346]));
    assign outputs[4792] = ~((layer0_outputs[9079]) | (layer0_outputs[1008]));
    assign outputs[4793] = layer0_outputs[8772];
    assign outputs[4794] = ~(layer0_outputs[2600]);
    assign outputs[4795] = (layer0_outputs[3386]) & (layer0_outputs[3540]);
    assign outputs[4796] = ~(layer0_outputs[2213]);
    assign outputs[4797] = ~((layer0_outputs[2487]) | (layer0_outputs[5113]));
    assign outputs[4798] = ~(layer0_outputs[6194]) | (layer0_outputs[7855]);
    assign outputs[4799] = (layer0_outputs[1513]) & ~(layer0_outputs[1328]);
    assign outputs[4800] = ~(layer0_outputs[3340]);
    assign outputs[4801] = ~(layer0_outputs[7792]);
    assign outputs[4802] = ~(layer0_outputs[4468]);
    assign outputs[4803] = (layer0_outputs[8336]) ^ (layer0_outputs[10083]);
    assign outputs[4804] = layer0_outputs[4697];
    assign outputs[4805] = (layer0_outputs[6344]) & (layer0_outputs[5637]);
    assign outputs[4806] = ~((layer0_outputs[991]) & (layer0_outputs[741]));
    assign outputs[4807] = (layer0_outputs[425]) ^ (layer0_outputs[178]);
    assign outputs[4808] = ~((layer0_outputs[5421]) ^ (layer0_outputs[4804]));
    assign outputs[4809] = ~((layer0_outputs[6074]) ^ (layer0_outputs[6046]));
    assign outputs[4810] = ~((layer0_outputs[4058]) ^ (layer0_outputs[4892]));
    assign outputs[4811] = (layer0_outputs[9929]) & ~(layer0_outputs[4891]);
    assign outputs[4812] = layer0_outputs[7738];
    assign outputs[4813] = ~((layer0_outputs[4077]) ^ (layer0_outputs[3037]));
    assign outputs[4814] = (layer0_outputs[10023]) ^ (layer0_outputs[4644]);
    assign outputs[4815] = ~(layer0_outputs[2385]);
    assign outputs[4816] = (layer0_outputs[5613]) & (layer0_outputs[4525]);
    assign outputs[4817] = ~((layer0_outputs[65]) ^ (layer0_outputs[2517]));
    assign outputs[4818] = layer0_outputs[8263];
    assign outputs[4819] = ~(layer0_outputs[2612]);
    assign outputs[4820] = ~(layer0_outputs[3264]);
    assign outputs[4821] = layer0_outputs[6540];
    assign outputs[4822] = (layer0_outputs[3875]) & ~(layer0_outputs[2503]);
    assign outputs[4823] = (layer0_outputs[8227]) ^ (layer0_outputs[9804]);
    assign outputs[4824] = ~(layer0_outputs[712]);
    assign outputs[4825] = 1'b0;
    assign outputs[4826] = (layer0_outputs[5683]) & ~(layer0_outputs[9239]);
    assign outputs[4827] = ~(layer0_outputs[8723]) | (layer0_outputs[9106]);
    assign outputs[4828] = ~(layer0_outputs[6938]);
    assign outputs[4829] = (layer0_outputs[6967]) ^ (layer0_outputs[5085]);
    assign outputs[4830] = ~(layer0_outputs[4361]);
    assign outputs[4831] = (layer0_outputs[2435]) ^ (layer0_outputs[4066]);
    assign outputs[4832] = layer0_outputs[10137];
    assign outputs[4833] = (layer0_outputs[9]) & (layer0_outputs[6229]);
    assign outputs[4834] = layer0_outputs[5675];
    assign outputs[4835] = ~(layer0_outputs[3951]);
    assign outputs[4836] = ~(layer0_outputs[2512]);
    assign outputs[4837] = layer0_outputs[4924];
    assign outputs[4838] = (layer0_outputs[1548]) & ~(layer0_outputs[3933]);
    assign outputs[4839] = layer0_outputs[8828];
    assign outputs[4840] = ~(layer0_outputs[1343]);
    assign outputs[4841] = ~((layer0_outputs[6325]) ^ (layer0_outputs[6732]));
    assign outputs[4842] = layer0_outputs[9656];
    assign outputs[4843] = (layer0_outputs[5329]) & (layer0_outputs[2882]);
    assign outputs[4844] = layer0_outputs[6270];
    assign outputs[4845] = ~(layer0_outputs[972]) | (layer0_outputs[436]);
    assign outputs[4846] = (layer0_outputs[9281]) | (layer0_outputs[7235]);
    assign outputs[4847] = layer0_outputs[4381];
    assign outputs[4848] = ~(layer0_outputs[1491]);
    assign outputs[4849] = ~((layer0_outputs[8361]) ^ (layer0_outputs[4840]));
    assign outputs[4850] = layer0_outputs[2277];
    assign outputs[4851] = ~((layer0_outputs[5466]) | (layer0_outputs[2608]));
    assign outputs[4852] = (layer0_outputs[5194]) ^ (layer0_outputs[6019]);
    assign outputs[4853] = layer0_outputs[4824];
    assign outputs[4854] = layer0_outputs[9700];
    assign outputs[4855] = ~(layer0_outputs[5414]) | (layer0_outputs[1376]);
    assign outputs[4856] = ~((layer0_outputs[9380]) | (layer0_outputs[6544]));
    assign outputs[4857] = layer0_outputs[8559];
    assign outputs[4858] = layer0_outputs[6726];
    assign outputs[4859] = ~((layer0_outputs[651]) | (layer0_outputs[5815]));
    assign outputs[4860] = layer0_outputs[2633];
    assign outputs[4861] = ~((layer0_outputs[7222]) ^ (layer0_outputs[4376]));
    assign outputs[4862] = ~((layer0_outputs[10160]) | (layer0_outputs[4894]));
    assign outputs[4863] = ~((layer0_outputs[1558]) ^ (layer0_outputs[3633]));
    assign outputs[4864] = ~(layer0_outputs[9371]);
    assign outputs[4865] = layer0_outputs[9231];
    assign outputs[4866] = layer0_outputs[5779];
    assign outputs[4867] = ~((layer0_outputs[4154]) ^ (layer0_outputs[6251]));
    assign outputs[4868] = layer0_outputs[2790];
    assign outputs[4869] = (layer0_outputs[3034]) & (layer0_outputs[10144]);
    assign outputs[4870] = layer0_outputs[9810];
    assign outputs[4871] = ~(layer0_outputs[1801]) | (layer0_outputs[5340]);
    assign outputs[4872] = layer0_outputs[9346];
    assign outputs[4873] = ~((layer0_outputs[1090]) ^ (layer0_outputs[4049]));
    assign outputs[4874] = ~((layer0_outputs[5880]) ^ (layer0_outputs[4701]));
    assign outputs[4875] = (layer0_outputs[376]) ^ (layer0_outputs[8187]);
    assign outputs[4876] = layer0_outputs[3734];
    assign outputs[4877] = layer0_outputs[3052];
    assign outputs[4878] = ~((layer0_outputs[439]) ^ (layer0_outputs[6298]));
    assign outputs[4879] = layer0_outputs[6113];
    assign outputs[4880] = ~(layer0_outputs[8402]);
    assign outputs[4881] = layer0_outputs[2977];
    assign outputs[4882] = layer0_outputs[5823];
    assign outputs[4883] = ~((layer0_outputs[1666]) ^ (layer0_outputs[353]));
    assign outputs[4884] = ~(layer0_outputs[6157]) | (layer0_outputs[6855]);
    assign outputs[4885] = layer0_outputs[6250];
    assign outputs[4886] = ~(layer0_outputs[1134]);
    assign outputs[4887] = ~(layer0_outputs[2137]) | (layer0_outputs[3505]);
    assign outputs[4888] = ~((layer0_outputs[3339]) & (layer0_outputs[1490]));
    assign outputs[4889] = ~(layer0_outputs[3233]);
    assign outputs[4890] = layer0_outputs[696];
    assign outputs[4891] = ~((layer0_outputs[6475]) ^ (layer0_outputs[7998]));
    assign outputs[4892] = ~((layer0_outputs[4757]) | (layer0_outputs[7169]));
    assign outputs[4893] = ~((layer0_outputs[6552]) | (layer0_outputs[7704]));
    assign outputs[4894] = layer0_outputs[2480];
    assign outputs[4895] = (layer0_outputs[2053]) & ~(layer0_outputs[4227]);
    assign outputs[4896] = layer0_outputs[3720];
    assign outputs[4897] = (layer0_outputs[3461]) ^ (layer0_outputs[9846]);
    assign outputs[4898] = ~(layer0_outputs[5474]);
    assign outputs[4899] = layer0_outputs[3063];
    assign outputs[4900] = layer0_outputs[6334];
    assign outputs[4901] = layer0_outputs[4352];
    assign outputs[4902] = ~(layer0_outputs[1784]) | (layer0_outputs[6123]);
    assign outputs[4903] = ~((layer0_outputs[9197]) | (layer0_outputs[4908]));
    assign outputs[4904] = ~((layer0_outputs[5007]) ^ (layer0_outputs[9542]));
    assign outputs[4905] = (layer0_outputs[6398]) ^ (layer0_outputs[3319]);
    assign outputs[4906] = ~(layer0_outputs[102]);
    assign outputs[4907] = ~((layer0_outputs[8512]) ^ (layer0_outputs[9678]));
    assign outputs[4908] = ~((layer0_outputs[365]) ^ (layer0_outputs[7640]));
    assign outputs[4909] = layer0_outputs[804];
    assign outputs[4910] = ~(layer0_outputs[4297]) | (layer0_outputs[3179]);
    assign outputs[4911] = (layer0_outputs[7412]) ^ (layer0_outputs[2034]);
    assign outputs[4912] = layer0_outputs[1202];
    assign outputs[4913] = layer0_outputs[4505];
    assign outputs[4914] = (layer0_outputs[1093]) & ~(layer0_outputs[6699]);
    assign outputs[4915] = ~((layer0_outputs[6531]) ^ (layer0_outputs[4065]));
    assign outputs[4916] = ~((layer0_outputs[2787]) & (layer0_outputs[9877]));
    assign outputs[4917] = ~((layer0_outputs[1899]) ^ (layer0_outputs[4650]));
    assign outputs[4918] = ~(layer0_outputs[1550]) | (layer0_outputs[7023]);
    assign outputs[4919] = (layer0_outputs[7002]) ^ (layer0_outputs[3035]);
    assign outputs[4920] = ~(layer0_outputs[9378]);
    assign outputs[4921] = (layer0_outputs[3733]) & ~(layer0_outputs[9561]);
    assign outputs[4922] = layer0_outputs[8422];
    assign outputs[4923] = ~(layer0_outputs[5792]);
    assign outputs[4924] = ~((layer0_outputs[6144]) ^ (layer0_outputs[8185]));
    assign outputs[4925] = layer0_outputs[5886];
    assign outputs[4926] = ~((layer0_outputs[8545]) | (layer0_outputs[1611]));
    assign outputs[4927] = (layer0_outputs[3009]) & ~(layer0_outputs[9123]);
    assign outputs[4928] = ~(layer0_outputs[458]);
    assign outputs[4929] = ~(layer0_outputs[8012]);
    assign outputs[4930] = ~(layer0_outputs[2574]) | (layer0_outputs[644]);
    assign outputs[4931] = ~((layer0_outputs[4104]) ^ (layer0_outputs[9339]));
    assign outputs[4932] = ~(layer0_outputs[4274]);
    assign outputs[4933] = layer0_outputs[1643];
    assign outputs[4934] = ~(layer0_outputs[6736]) | (layer0_outputs[3670]);
    assign outputs[4935] = (layer0_outputs[1538]) & ~(layer0_outputs[5825]);
    assign outputs[4936] = (layer0_outputs[6238]) & (layer0_outputs[5969]);
    assign outputs[4937] = ~(layer0_outputs[8463]);
    assign outputs[4938] = layer0_outputs[5330];
    assign outputs[4939] = (layer0_outputs[7588]) ^ (layer0_outputs[2892]);
    assign outputs[4940] = ~(layer0_outputs[9021]);
    assign outputs[4941] = (layer0_outputs[4440]) & ~(layer0_outputs[1201]);
    assign outputs[4942] = ~(layer0_outputs[2482]);
    assign outputs[4943] = layer0_outputs[8119];
    assign outputs[4944] = (layer0_outputs[4860]) & ~(layer0_outputs[3538]);
    assign outputs[4945] = (layer0_outputs[7712]) ^ (layer0_outputs[3976]);
    assign outputs[4946] = layer0_outputs[8963];
    assign outputs[4947] = 1'b1;
    assign outputs[4948] = (layer0_outputs[7690]) ^ (layer0_outputs[1096]);
    assign outputs[4949] = ~(layer0_outputs[935]);
    assign outputs[4950] = layer0_outputs[9281];
    assign outputs[4951] = (layer0_outputs[9063]) ^ (layer0_outputs[1877]);
    assign outputs[4952] = layer0_outputs[5778];
    assign outputs[4953] = (layer0_outputs[827]) & (layer0_outputs[2662]);
    assign outputs[4954] = ~((layer0_outputs[6960]) ^ (layer0_outputs[1713]));
    assign outputs[4955] = layer0_outputs[9479];
    assign outputs[4956] = (layer0_outputs[5513]) & ~(layer0_outputs[2712]);
    assign outputs[4957] = (layer0_outputs[5251]) & (layer0_outputs[2953]);
    assign outputs[4958] = ~((layer0_outputs[2567]) ^ (layer0_outputs[1737]));
    assign outputs[4959] = ~(layer0_outputs[3874]) | (layer0_outputs[9270]);
    assign outputs[4960] = (layer0_outputs[6599]) & (layer0_outputs[4008]);
    assign outputs[4961] = ~((layer0_outputs[5996]) ^ (layer0_outputs[7546]));
    assign outputs[4962] = ~(layer0_outputs[6555]);
    assign outputs[4963] = (layer0_outputs[1729]) & ~(layer0_outputs[5172]);
    assign outputs[4964] = (layer0_outputs[2998]) ^ (layer0_outputs[7937]);
    assign outputs[4965] = (layer0_outputs[2954]) & ~(layer0_outputs[8664]);
    assign outputs[4966] = (layer0_outputs[8932]) & ~(layer0_outputs[694]);
    assign outputs[4967] = (layer0_outputs[3036]) ^ (layer0_outputs[47]);
    assign outputs[4968] = (layer0_outputs[1224]) ^ (layer0_outputs[203]);
    assign outputs[4969] = layer0_outputs[278];
    assign outputs[4970] = ~(layer0_outputs[4681]);
    assign outputs[4971] = ~(layer0_outputs[9248]);
    assign outputs[4972] = ~((layer0_outputs[2890]) ^ (layer0_outputs[9169]));
    assign outputs[4973] = (layer0_outputs[8601]) ^ (layer0_outputs[3522]);
    assign outputs[4974] = (layer0_outputs[276]) & ~(layer0_outputs[4806]);
    assign outputs[4975] = ~(layer0_outputs[4805]);
    assign outputs[4976] = (layer0_outputs[4169]) ^ (layer0_outputs[5440]);
    assign outputs[4977] = (layer0_outputs[8017]) & ~(layer0_outputs[7442]);
    assign outputs[4978] = layer0_outputs[7504];
    assign outputs[4979] = ~(layer0_outputs[2151]) | (layer0_outputs[5297]);
    assign outputs[4980] = ~((layer0_outputs[2133]) ^ (layer0_outputs[201]));
    assign outputs[4981] = layer0_outputs[9334];
    assign outputs[4982] = (layer0_outputs[8131]) ^ (layer0_outputs[2904]);
    assign outputs[4983] = (layer0_outputs[1640]) & ~(layer0_outputs[2030]);
    assign outputs[4984] = ~(layer0_outputs[5538]) | (layer0_outputs[4164]);
    assign outputs[4985] = ~((layer0_outputs[1881]) ^ (layer0_outputs[3553]));
    assign outputs[4986] = ~(layer0_outputs[7700]);
    assign outputs[4987] = layer0_outputs[5251];
    assign outputs[4988] = ~((layer0_outputs[9531]) ^ (layer0_outputs[4730]));
    assign outputs[4989] = layer0_outputs[9743];
    assign outputs[4990] = layer0_outputs[453];
    assign outputs[4991] = ~((layer0_outputs[4960]) ^ (layer0_outputs[7395]));
    assign outputs[4992] = ~((layer0_outputs[680]) ^ (layer0_outputs[9279]));
    assign outputs[4993] = ~((layer0_outputs[7400]) ^ (layer0_outputs[7188]));
    assign outputs[4994] = (layer0_outputs[146]) & (layer0_outputs[7712]);
    assign outputs[4995] = 1'b0;
    assign outputs[4996] = ~(layer0_outputs[234]) | (layer0_outputs[2257]);
    assign outputs[4997] = ~((layer0_outputs[2208]) ^ (layer0_outputs[7896]));
    assign outputs[4998] = (layer0_outputs[4487]) & ~(layer0_outputs[10127]);
    assign outputs[4999] = layer0_outputs[4370];
    assign outputs[5000] = layer0_outputs[8568];
    assign outputs[5001] = (layer0_outputs[2019]) & ~(layer0_outputs[5287]);
    assign outputs[5002] = ~((layer0_outputs[9536]) ^ (layer0_outputs[2679]));
    assign outputs[5003] = (layer0_outputs[4987]) & ~(layer0_outputs[4642]);
    assign outputs[5004] = ~((layer0_outputs[5530]) & (layer0_outputs[6239]));
    assign outputs[5005] = layer0_outputs[2774];
    assign outputs[5006] = ~((layer0_outputs[9443]) | (layer0_outputs[759]));
    assign outputs[5007] = ~((layer0_outputs[7367]) ^ (layer0_outputs[7385]));
    assign outputs[5008] = (layer0_outputs[146]) & ~(layer0_outputs[7768]);
    assign outputs[5009] = (layer0_outputs[9438]) ^ (layer0_outputs[1430]);
    assign outputs[5010] = layer0_outputs[7010];
    assign outputs[5011] = (layer0_outputs[1705]) ^ (layer0_outputs[381]);
    assign outputs[5012] = ~((layer0_outputs[169]) ^ (layer0_outputs[3585]));
    assign outputs[5013] = (layer0_outputs[8331]) | (layer0_outputs[5359]);
    assign outputs[5014] = layer0_outputs[1271];
    assign outputs[5015] = ~(layer0_outputs[4131]) | (layer0_outputs[3848]);
    assign outputs[5016] = ~((layer0_outputs[751]) | (layer0_outputs[2089]));
    assign outputs[5017] = ~((layer0_outputs[5827]) ^ (layer0_outputs[1789]));
    assign outputs[5018] = ~(layer0_outputs[1691]) | (layer0_outputs[5813]);
    assign outputs[5019] = ~(layer0_outputs[6302]);
    assign outputs[5020] = (layer0_outputs[2340]) ^ (layer0_outputs[738]);
    assign outputs[5021] = ~(layer0_outputs[5132]) | (layer0_outputs[1916]);
    assign outputs[5022] = ~(layer0_outputs[8505]);
    assign outputs[5023] = (layer0_outputs[5090]) & (layer0_outputs[3828]);
    assign outputs[5024] = layer0_outputs[1359];
    assign outputs[5025] = ~((layer0_outputs[6892]) ^ (layer0_outputs[4174]));
    assign outputs[5026] = (layer0_outputs[2095]) | (layer0_outputs[4558]);
    assign outputs[5027] = layer0_outputs[9308];
    assign outputs[5028] = layer0_outputs[9250];
    assign outputs[5029] = layer0_outputs[7791];
    assign outputs[5030] = layer0_outputs[2141];
    assign outputs[5031] = ~((layer0_outputs[1805]) ^ (layer0_outputs[7123]));
    assign outputs[5032] = layer0_outputs[8977];
    assign outputs[5033] = (layer0_outputs[1288]) & (layer0_outputs[6171]);
    assign outputs[5034] = (layer0_outputs[6434]) ^ (layer0_outputs[5721]);
    assign outputs[5035] = (layer0_outputs[5018]) ^ (layer0_outputs[8612]);
    assign outputs[5036] = layer0_outputs[5688];
    assign outputs[5037] = (layer0_outputs[2255]) & ~(layer0_outputs[6705]);
    assign outputs[5038] = layer0_outputs[454];
    assign outputs[5039] = ~(layer0_outputs[6908]);
    assign outputs[5040] = (layer0_outputs[4956]) | (layer0_outputs[10049]);
    assign outputs[5041] = ~(layer0_outputs[339]);
    assign outputs[5042] = ~(layer0_outputs[8221]);
    assign outputs[5043] = layer0_outputs[8885];
    assign outputs[5044] = layer0_outputs[670];
    assign outputs[5045] = ~(layer0_outputs[1920]);
    assign outputs[5046] = layer0_outputs[6101];
    assign outputs[5047] = layer0_outputs[1338];
    assign outputs[5048] = layer0_outputs[4452];
    assign outputs[5049] = (layer0_outputs[9874]) | (layer0_outputs[3680]);
    assign outputs[5050] = ~((layer0_outputs[7950]) ^ (layer0_outputs[3351]));
    assign outputs[5051] = ~(layer0_outputs[6874]);
    assign outputs[5052] = ~(layer0_outputs[7310]);
    assign outputs[5053] = (layer0_outputs[223]) ^ (layer0_outputs[5765]);
    assign outputs[5054] = layer0_outputs[3564];
    assign outputs[5055] = layer0_outputs[8480];
    assign outputs[5056] = layer0_outputs[6132];
    assign outputs[5057] = layer0_outputs[5437];
    assign outputs[5058] = (layer0_outputs[9499]) & ~(layer0_outputs[3098]);
    assign outputs[5059] = layer0_outputs[5572];
    assign outputs[5060] = ~((layer0_outputs[7038]) ^ (layer0_outputs[6535]));
    assign outputs[5061] = 1'b0;
    assign outputs[5062] = layer0_outputs[9728];
    assign outputs[5063] = ~((layer0_outputs[9196]) ^ (layer0_outputs[7195]));
    assign outputs[5064] = ~(layer0_outputs[6205]);
    assign outputs[5065] = ~(layer0_outputs[3097]) | (layer0_outputs[9433]);
    assign outputs[5066] = layer0_outputs[6545];
    assign outputs[5067] = layer0_outputs[982];
    assign outputs[5068] = (layer0_outputs[1913]) ^ (layer0_outputs[96]);
    assign outputs[5069] = ~((layer0_outputs[10013]) & (layer0_outputs[2878]));
    assign outputs[5070] = layer0_outputs[4404];
    assign outputs[5071] = (layer0_outputs[7945]) ^ (layer0_outputs[7884]);
    assign outputs[5072] = ~((layer0_outputs[97]) ^ (layer0_outputs[9164]));
    assign outputs[5073] = (layer0_outputs[6165]) & (layer0_outputs[7100]);
    assign outputs[5074] = ~(layer0_outputs[5301]);
    assign outputs[5075] = layer0_outputs[2974];
    assign outputs[5076] = ~(layer0_outputs[7858]);
    assign outputs[5077] = (layer0_outputs[9633]) ^ (layer0_outputs[10154]);
    assign outputs[5078] = layer0_outputs[4492];
    assign outputs[5079] = layer0_outputs[1234];
    assign outputs[5080] = layer0_outputs[8605];
    assign outputs[5081] = (layer0_outputs[3884]) & (layer0_outputs[742]);
    assign outputs[5082] = ~(layer0_outputs[3325]);
    assign outputs[5083] = ~(layer0_outputs[5125]) | (layer0_outputs[2317]);
    assign outputs[5084] = layer0_outputs[3265];
    assign outputs[5085] = ~((layer0_outputs[3727]) | (layer0_outputs[6988]));
    assign outputs[5086] = ~(layer0_outputs[10092]);
    assign outputs[5087] = layer0_outputs[3398];
    assign outputs[5088] = ~(layer0_outputs[7232]);
    assign outputs[5089] = (layer0_outputs[5176]) | (layer0_outputs[1939]);
    assign outputs[5090] = ~(layer0_outputs[7648]);
    assign outputs[5091] = (layer0_outputs[3993]) & ~(layer0_outputs[190]);
    assign outputs[5092] = (layer0_outputs[8353]) ^ (layer0_outputs[5044]);
    assign outputs[5093] = ~((layer0_outputs[2337]) ^ (layer0_outputs[6475]));
    assign outputs[5094] = layer0_outputs[9751];
    assign outputs[5095] = (layer0_outputs[7603]) ^ (layer0_outputs[7139]);
    assign outputs[5096] = layer0_outputs[2341];
    assign outputs[5097] = (layer0_outputs[9472]) ^ (layer0_outputs[6914]);
    assign outputs[5098] = 1'b1;
    assign outputs[5099] = (layer0_outputs[5630]) & (layer0_outputs[8792]);
    assign outputs[5100] = ~((layer0_outputs[771]) ^ (layer0_outputs[7341]));
    assign outputs[5101] = ~(layer0_outputs[1294]);
    assign outputs[5102] = (layer0_outputs[7873]) & (layer0_outputs[9014]);
    assign outputs[5103] = ~(layer0_outputs[845]);
    assign outputs[5104] = ~(layer0_outputs[9488]);
    assign outputs[5105] = ~(layer0_outputs[3894]);
    assign outputs[5106] = layer0_outputs[1004];
    assign outputs[5107] = (layer0_outputs[494]) ^ (layer0_outputs[9982]);
    assign outputs[5108] = ~(layer0_outputs[5690]);
    assign outputs[5109] = ~(layer0_outputs[2308]);
    assign outputs[5110] = layer0_outputs[1639];
    assign outputs[5111] = ~((layer0_outputs[445]) ^ (layer0_outputs[459]));
    assign outputs[5112] = (layer0_outputs[6453]) | (layer0_outputs[8065]);
    assign outputs[5113] = layer0_outputs[5911];
    assign outputs[5114] = ~(layer0_outputs[2213]);
    assign outputs[5115] = ~(layer0_outputs[9836]) | (layer0_outputs[8152]);
    assign outputs[5116] = layer0_outputs[7907];
    assign outputs[5117] = (layer0_outputs[3399]) & ~(layer0_outputs[9975]);
    assign outputs[5118] = (layer0_outputs[5686]) & ~(layer0_outputs[2996]);
    assign outputs[5119] = (layer0_outputs[5928]) & ~(layer0_outputs[4283]);
    assign outputs[5120] = layer0_outputs[5555];
    assign outputs[5121] = ~(layer0_outputs[2731]);
    assign outputs[5122] = ~((layer0_outputs[9280]) | (layer0_outputs[9890]));
    assign outputs[5123] = (layer0_outputs[8613]) ^ (layer0_outputs[2246]);
    assign outputs[5124] = ~((layer0_outputs[9919]) ^ (layer0_outputs[7863]));
    assign outputs[5125] = (layer0_outputs[2958]) & ~(layer0_outputs[7348]);
    assign outputs[5126] = ~(layer0_outputs[1436]);
    assign outputs[5127] = layer0_outputs[4505];
    assign outputs[5128] = ~(layer0_outputs[3608]);
    assign outputs[5129] = (layer0_outputs[2145]) ^ (layer0_outputs[2730]);
    assign outputs[5130] = ~((layer0_outputs[2467]) & (layer0_outputs[8800]));
    assign outputs[5131] = (layer0_outputs[1091]) & (layer0_outputs[7341]);
    assign outputs[5132] = (layer0_outputs[8046]) ^ (layer0_outputs[3563]);
    assign outputs[5133] = (layer0_outputs[9855]) ^ (layer0_outputs[3411]);
    assign outputs[5134] = ~(layer0_outputs[1106]);
    assign outputs[5135] = layer0_outputs[4599];
    assign outputs[5136] = (layer0_outputs[3280]) | (layer0_outputs[1097]);
    assign outputs[5137] = (layer0_outputs[7226]) ^ (layer0_outputs[8758]);
    assign outputs[5138] = ~(layer0_outputs[9491]);
    assign outputs[5139] = ~((layer0_outputs[9847]) ^ (layer0_outputs[8765]));
    assign outputs[5140] = ~(layer0_outputs[2202]);
    assign outputs[5141] = ~((layer0_outputs[6896]) ^ (layer0_outputs[8544]));
    assign outputs[5142] = ~(layer0_outputs[3939]);
    assign outputs[5143] = ~(layer0_outputs[834]);
    assign outputs[5144] = ~((layer0_outputs[7656]) | (layer0_outputs[2569]));
    assign outputs[5145] = ~(layer0_outputs[5208]) | (layer0_outputs[4050]);
    assign outputs[5146] = layer0_outputs[9290];
    assign outputs[5147] = ~(layer0_outputs[1751]);
    assign outputs[5148] = ~((layer0_outputs[3775]) ^ (layer0_outputs[59]));
    assign outputs[5149] = ~(layer0_outputs[4248]) | (layer0_outputs[6001]);
    assign outputs[5150] = ~(layer0_outputs[5006]);
    assign outputs[5151] = (layer0_outputs[8423]) ^ (layer0_outputs[2377]);
    assign outputs[5152] = ~((layer0_outputs[3665]) | (layer0_outputs[4062]));
    assign outputs[5153] = layer0_outputs[1849];
    assign outputs[5154] = ~(layer0_outputs[8348]);
    assign outputs[5155] = ~((layer0_outputs[1261]) ^ (layer0_outputs[7559]));
    assign outputs[5156] = layer0_outputs[682];
    assign outputs[5157] = ~((layer0_outputs[2420]) ^ (layer0_outputs[6989]));
    assign outputs[5158] = layer0_outputs[6309];
    assign outputs[5159] = ~(layer0_outputs[5472]) | (layer0_outputs[4162]);
    assign outputs[5160] = ~((layer0_outputs[5423]) ^ (layer0_outputs[5389]));
    assign outputs[5161] = ~(layer0_outputs[1466]) | (layer0_outputs[5558]);
    assign outputs[5162] = (layer0_outputs[4996]) | (layer0_outputs[3547]);
    assign outputs[5163] = ~(layer0_outputs[7445]);
    assign outputs[5164] = (layer0_outputs[9710]) ^ (layer0_outputs[3516]);
    assign outputs[5165] = ~(layer0_outputs[9197]);
    assign outputs[5166] = (layer0_outputs[1102]) ^ (layer0_outputs[2616]);
    assign outputs[5167] = layer0_outputs[5348];
    assign outputs[5168] = (layer0_outputs[4334]) & ~(layer0_outputs[5155]);
    assign outputs[5169] = layer0_outputs[4873];
    assign outputs[5170] = layer0_outputs[1160];
    assign outputs[5171] = (layer0_outputs[9229]) ^ (layer0_outputs[3362]);
    assign outputs[5172] = ~(layer0_outputs[10050]);
    assign outputs[5173] = ~((layer0_outputs[8197]) | (layer0_outputs[6954]));
    assign outputs[5174] = ~(layer0_outputs[1291]) | (layer0_outputs[4453]);
    assign outputs[5175] = ~(layer0_outputs[1412]);
    assign outputs[5176] = (layer0_outputs[7410]) ^ (layer0_outputs[9810]);
    assign outputs[5177] = ~(layer0_outputs[9730]);
    assign outputs[5178] = ~(layer0_outputs[387]);
    assign outputs[5179] = 1'b1;
    assign outputs[5180] = (layer0_outputs[642]) ^ (layer0_outputs[9766]);
    assign outputs[5181] = layer0_outputs[9837];
    assign outputs[5182] = ~((layer0_outputs[4113]) ^ (layer0_outputs[2414]));
    assign outputs[5183] = ~(layer0_outputs[9618]) | (layer0_outputs[4361]);
    assign outputs[5184] = layer0_outputs[6505];
    assign outputs[5185] = layer0_outputs[5745];
    assign outputs[5186] = layer0_outputs[7218];
    assign outputs[5187] = ~((layer0_outputs[5932]) ^ (layer0_outputs[3681]));
    assign outputs[5188] = (layer0_outputs[4871]) ^ (layer0_outputs[2948]);
    assign outputs[5189] = (layer0_outputs[5705]) ^ (layer0_outputs[406]);
    assign outputs[5190] = layer0_outputs[7516];
    assign outputs[5191] = (layer0_outputs[494]) ^ (layer0_outputs[6914]);
    assign outputs[5192] = (layer0_outputs[7698]) & (layer0_outputs[8340]);
    assign outputs[5193] = (layer0_outputs[870]) & ~(layer0_outputs[9110]);
    assign outputs[5194] = layer0_outputs[9088];
    assign outputs[5195] = ~(layer0_outputs[5674]);
    assign outputs[5196] = ~(layer0_outputs[7788]);
    assign outputs[5197] = layer0_outputs[10199];
    assign outputs[5198] = ~((layer0_outputs[8163]) & (layer0_outputs[130]));
    assign outputs[5199] = ~((layer0_outputs[5404]) ^ (layer0_outputs[3815]));
    assign outputs[5200] = layer0_outputs[6714];
    assign outputs[5201] = ~(layer0_outputs[1792]);
    assign outputs[5202] = (layer0_outputs[2939]) | (layer0_outputs[1398]);
    assign outputs[5203] = layer0_outputs[8939];
    assign outputs[5204] = ~((layer0_outputs[6058]) & (layer0_outputs[435]));
    assign outputs[5205] = (layer0_outputs[3555]) ^ (layer0_outputs[7556]);
    assign outputs[5206] = layer0_outputs[6147];
    assign outputs[5207] = ~(layer0_outputs[8604]);
    assign outputs[5208] = ~((layer0_outputs[7458]) ^ (layer0_outputs[2793]));
    assign outputs[5209] = ~((layer0_outputs[7986]) ^ (layer0_outputs[462]));
    assign outputs[5210] = ~(layer0_outputs[5910]) | (layer0_outputs[4979]);
    assign outputs[5211] = layer0_outputs[758];
    assign outputs[5212] = layer0_outputs[6147];
    assign outputs[5213] = (layer0_outputs[1715]) & (layer0_outputs[5582]);
    assign outputs[5214] = layer0_outputs[6585];
    assign outputs[5215] = ~((layer0_outputs[7148]) & (layer0_outputs[8327]));
    assign outputs[5216] = (layer0_outputs[6629]) ^ (layer0_outputs[10060]);
    assign outputs[5217] = (layer0_outputs[4522]) | (layer0_outputs[805]);
    assign outputs[5218] = ~(layer0_outputs[3586]);
    assign outputs[5219] = (layer0_outputs[1086]) | (layer0_outputs[789]);
    assign outputs[5220] = layer0_outputs[8063];
    assign outputs[5221] = ~((layer0_outputs[7901]) ^ (layer0_outputs[10170]));
    assign outputs[5222] = (layer0_outputs[5832]) ^ (layer0_outputs[3566]);
    assign outputs[5223] = (layer0_outputs[9979]) ^ (layer0_outputs[866]);
    assign outputs[5224] = (layer0_outputs[9694]) & ~(layer0_outputs[9335]);
    assign outputs[5225] = (layer0_outputs[3214]) & ~(layer0_outputs[6278]);
    assign outputs[5226] = (layer0_outputs[2619]) & ~(layer0_outputs[3511]);
    assign outputs[5227] = (layer0_outputs[7421]) ^ (layer0_outputs[5470]);
    assign outputs[5228] = ~(layer0_outputs[3343]);
    assign outputs[5229] = ~((layer0_outputs[7545]) | (layer0_outputs[3599]));
    assign outputs[5230] = layer0_outputs[930];
    assign outputs[5231] = (layer0_outputs[7752]) ^ (layer0_outputs[9116]);
    assign outputs[5232] = (layer0_outputs[9111]) ^ (layer0_outputs[652]);
    assign outputs[5233] = ~(layer0_outputs[679]);
    assign outputs[5234] = ~(layer0_outputs[4717]);
    assign outputs[5235] = ~((layer0_outputs[7729]) | (layer0_outputs[879]));
    assign outputs[5236] = ~(layer0_outputs[7306]) | (layer0_outputs[6646]);
    assign outputs[5237] = (layer0_outputs[9916]) & ~(layer0_outputs[2621]);
    assign outputs[5238] = (layer0_outputs[7402]) ^ (layer0_outputs[10062]);
    assign outputs[5239] = layer0_outputs[7314];
    assign outputs[5240] = ~((layer0_outputs[8367]) | (layer0_outputs[8752]));
    assign outputs[5241] = (layer0_outputs[9373]) ^ (layer0_outputs[1193]);
    assign outputs[5242] = (layer0_outputs[2181]) ^ (layer0_outputs[3798]);
    assign outputs[5243] = ~(layer0_outputs[1998]) | (layer0_outputs[9742]);
    assign outputs[5244] = ~((layer0_outputs[665]) ^ (layer0_outputs[9563]));
    assign outputs[5245] = (layer0_outputs[2663]) ^ (layer0_outputs[2071]);
    assign outputs[5246] = layer0_outputs[6150];
    assign outputs[5247] = ~(layer0_outputs[7434]);
    assign outputs[5248] = (layer0_outputs[3807]) ^ (layer0_outputs[7651]);
    assign outputs[5249] = layer0_outputs[7296];
    assign outputs[5250] = ~((layer0_outputs[7623]) ^ (layer0_outputs[3868]));
    assign outputs[5251] = ~(layer0_outputs[591]);
    assign outputs[5252] = ~((layer0_outputs[4527]) ^ (layer0_outputs[3877]));
    assign outputs[5253] = ~((layer0_outputs[2797]) ^ (layer0_outputs[13]));
    assign outputs[5254] = (layer0_outputs[7297]) ^ (layer0_outputs[6932]);
    assign outputs[5255] = layer0_outputs[1603];
    assign outputs[5256] = ~(layer0_outputs[7160]) | (layer0_outputs[7571]);
    assign outputs[5257] = (layer0_outputs[3950]) | (layer0_outputs[6928]);
    assign outputs[5258] = ~((layer0_outputs[420]) ^ (layer0_outputs[3267]));
    assign outputs[5259] = layer0_outputs[1595];
    assign outputs[5260] = layer0_outputs[470];
    assign outputs[5261] = layer0_outputs[6847];
    assign outputs[5262] = layer0_outputs[2715];
    assign outputs[5263] = (layer0_outputs[3843]) ^ (layer0_outputs[6021]);
    assign outputs[5264] = (layer0_outputs[3658]) & (layer0_outputs[7331]);
    assign outputs[5265] = ~(layer0_outputs[393]);
    assign outputs[5266] = layer0_outputs[8714];
    assign outputs[5267] = (layer0_outputs[3998]) ^ (layer0_outputs[9669]);
    assign outputs[5268] = layer0_outputs[5431];
    assign outputs[5269] = (layer0_outputs[430]) & ~(layer0_outputs[1012]);
    assign outputs[5270] = (layer0_outputs[8465]) ^ (layer0_outputs[2886]);
    assign outputs[5271] = ~(layer0_outputs[10130]);
    assign outputs[5272] = ~((layer0_outputs[6600]) ^ (layer0_outputs[6860]));
    assign outputs[5273] = ~(layer0_outputs[3922]);
    assign outputs[5274] = ~(layer0_outputs[3660]);
    assign outputs[5275] = (layer0_outputs[9382]) ^ (layer0_outputs[6761]);
    assign outputs[5276] = ~((layer0_outputs[3249]) ^ (layer0_outputs[14]));
    assign outputs[5277] = ~((layer0_outputs[305]) & (layer0_outputs[2847]));
    assign outputs[5278] = layer0_outputs[4153];
    assign outputs[5279] = ~((layer0_outputs[8594]) ^ (layer0_outputs[1326]));
    assign outputs[5280] = ~(layer0_outputs[2138]);
    assign outputs[5281] = 1'b1;
    assign outputs[5282] = ~(layer0_outputs[2507]);
    assign outputs[5283] = ~(layer0_outputs[4791]) | (layer0_outputs[5361]);
    assign outputs[5284] = ~((layer0_outputs[1552]) ^ (layer0_outputs[8921]));
    assign outputs[5285] = (layer0_outputs[311]) ^ (layer0_outputs[6998]);
    assign outputs[5286] = (layer0_outputs[9864]) | (layer0_outputs[1924]);
    assign outputs[5287] = ~((layer0_outputs[9749]) ^ (layer0_outputs[7951]));
    assign outputs[5288] = (layer0_outputs[6256]) & ~(layer0_outputs[9113]);
    assign outputs[5289] = layer0_outputs[1414];
    assign outputs[5290] = ~(layer0_outputs[1932]);
    assign outputs[5291] = (layer0_outputs[7324]) | (layer0_outputs[8912]);
    assign outputs[5292] = layer0_outputs[4822];
    assign outputs[5293] = layer0_outputs[2780];
    assign outputs[5294] = ~((layer0_outputs[8398]) ^ (layer0_outputs[2933]));
    assign outputs[5295] = ~(layer0_outputs[6127]) | (layer0_outputs[1438]);
    assign outputs[5296] = ~(layer0_outputs[105]);
    assign outputs[5297] = (layer0_outputs[7743]) | (layer0_outputs[9213]);
    assign outputs[5298] = layer0_outputs[9587];
    assign outputs[5299] = ~((layer0_outputs[4700]) ^ (layer0_outputs[2099]));
    assign outputs[5300] = (layer0_outputs[7737]) ^ (layer0_outputs[6587]);
    assign outputs[5301] = (layer0_outputs[4082]) & ~(layer0_outputs[977]);
    assign outputs[5302] = (layer0_outputs[1103]) & ~(layer0_outputs[349]);
    assign outputs[5303] = ~((layer0_outputs[6737]) ^ (layer0_outputs[7654]));
    assign outputs[5304] = ~((layer0_outputs[5222]) ^ (layer0_outputs[3029]));
    assign outputs[5305] = (layer0_outputs[7471]) ^ (layer0_outputs[1080]);
    assign outputs[5306] = (layer0_outputs[2755]) & ~(layer0_outputs[3346]);
    assign outputs[5307] = ~(layer0_outputs[6341]);
    assign outputs[5308] = (layer0_outputs[4758]) | (layer0_outputs[9099]);
    assign outputs[5309] = (layer0_outputs[4374]) ^ (layer0_outputs[8034]);
    assign outputs[5310] = (layer0_outputs[6458]) ^ (layer0_outputs[8629]);
    assign outputs[5311] = ~(layer0_outputs[10004]);
    assign outputs[5312] = (layer0_outputs[2711]) & ~(layer0_outputs[1478]);
    assign outputs[5313] = ~(layer0_outputs[6374]);
    assign outputs[5314] = ~(layer0_outputs[9269]);
    assign outputs[5315] = layer0_outputs[651];
    assign outputs[5316] = (layer0_outputs[9203]) ^ (layer0_outputs[8960]);
    assign outputs[5317] = ~(layer0_outputs[210]);
    assign outputs[5318] = (layer0_outputs[3182]) ^ (layer0_outputs[5572]);
    assign outputs[5319] = ~(layer0_outputs[4250]) | (layer0_outputs[2387]);
    assign outputs[5320] = layer0_outputs[1176];
    assign outputs[5321] = (layer0_outputs[3536]) ^ (layer0_outputs[3891]);
    assign outputs[5322] = ~((layer0_outputs[6697]) & (layer0_outputs[1251]));
    assign outputs[5323] = layer0_outputs[8721];
    assign outputs[5324] = (layer0_outputs[4885]) & (layer0_outputs[9265]);
    assign outputs[5325] = ~((layer0_outputs[2810]) & (layer0_outputs[7512]));
    assign outputs[5326] = (layer0_outputs[1542]) & ~(layer0_outputs[52]);
    assign outputs[5327] = ~(layer0_outputs[6363]);
    assign outputs[5328] = (layer0_outputs[4365]) | (layer0_outputs[4822]);
    assign outputs[5329] = ~(layer0_outputs[5002]);
    assign outputs[5330] = ~(layer0_outputs[4585]) | (layer0_outputs[1152]);
    assign outputs[5331] = ~(layer0_outputs[2902]);
    assign outputs[5332] = ~(layer0_outputs[2908]);
    assign outputs[5333] = ~((layer0_outputs[3470]) & (layer0_outputs[7103]));
    assign outputs[5334] = ~(layer0_outputs[4614]);
    assign outputs[5335] = (layer0_outputs[9672]) ^ (layer0_outputs[8850]);
    assign outputs[5336] = ~(layer0_outputs[748]) | (layer0_outputs[2777]);
    assign outputs[5337] = ~((layer0_outputs[5043]) ^ (layer0_outputs[1249]));
    assign outputs[5338] = ~(layer0_outputs[3010]);
    assign outputs[5339] = ~(layer0_outputs[3117]);
    assign outputs[5340] = ~((layer0_outputs[4654]) ^ (layer0_outputs[2084]));
    assign outputs[5341] = ~((layer0_outputs[1796]) ^ (layer0_outputs[6378]));
    assign outputs[5342] = ~(layer0_outputs[3085]);
    assign outputs[5343] = ~(layer0_outputs[3489]);
    assign outputs[5344] = (layer0_outputs[3012]) ^ (layer0_outputs[9490]);
    assign outputs[5345] = ~(layer0_outputs[8873]);
    assign outputs[5346] = ~((layer0_outputs[2032]) ^ (layer0_outputs[1126]));
    assign outputs[5347] = (layer0_outputs[4541]) ^ (layer0_outputs[7015]);
    assign outputs[5348] = ~((layer0_outputs[2596]) ^ (layer0_outputs[9045]));
    assign outputs[5349] = layer0_outputs[1524];
    assign outputs[5350] = layer0_outputs[1908];
    assign outputs[5351] = layer0_outputs[7584];
    assign outputs[5352] = ~(layer0_outputs[4782]);
    assign outputs[5353] = (layer0_outputs[9385]) ^ (layer0_outputs[3209]);
    assign outputs[5354] = ~(layer0_outputs[9316]);
    assign outputs[5355] = ~((layer0_outputs[5500]) ^ (layer0_outputs[8094]));
    assign outputs[5356] = ~(layer0_outputs[6146]) | (layer0_outputs[422]);
    assign outputs[5357] = ~(layer0_outputs[3367]);
    assign outputs[5358] = (layer0_outputs[1989]) & ~(layer0_outputs[4683]);
    assign outputs[5359] = ~(layer0_outputs[7681]);
    assign outputs[5360] = (layer0_outputs[1113]) | (layer0_outputs[7473]);
    assign outputs[5361] = ~((layer0_outputs[3639]) ^ (layer0_outputs[1777]));
    assign outputs[5362] = ~(layer0_outputs[9943]);
    assign outputs[5363] = ~(layer0_outputs[7634]);
    assign outputs[5364] = (layer0_outputs[1899]) & ~(layer0_outputs[8752]);
    assign outputs[5365] = ~(layer0_outputs[2782]);
    assign outputs[5366] = ~((layer0_outputs[9436]) ^ (layer0_outputs[215]));
    assign outputs[5367] = (layer0_outputs[86]) | (layer0_outputs[3737]);
    assign outputs[5368] = (layer0_outputs[8830]) ^ (layer0_outputs[1652]);
    assign outputs[5369] = ~(layer0_outputs[1432]);
    assign outputs[5370] = ~((layer0_outputs[6490]) ^ (layer0_outputs[6198]));
    assign outputs[5371] = ~(layer0_outputs[3383]);
    assign outputs[5372] = ~(layer0_outputs[5417]);
    assign outputs[5373] = ~((layer0_outputs[5973]) & (layer0_outputs[7606]));
    assign outputs[5374] = (layer0_outputs[6503]) | (layer0_outputs[9821]);
    assign outputs[5375] = ~((layer0_outputs[7197]) ^ (layer0_outputs[9243]));
    assign outputs[5376] = ~(layer0_outputs[5351]) | (layer0_outputs[2388]);
    assign outputs[5377] = ~((layer0_outputs[3374]) | (layer0_outputs[8113]));
    assign outputs[5378] = ~((layer0_outputs[8900]) ^ (layer0_outputs[6959]));
    assign outputs[5379] = ~((layer0_outputs[5480]) ^ (layer0_outputs[2593]));
    assign outputs[5380] = (layer0_outputs[896]) ^ (layer0_outputs[2568]);
    assign outputs[5381] = ~((layer0_outputs[4817]) ^ (layer0_outputs[10185]));
    assign outputs[5382] = ~((layer0_outputs[6843]) ^ (layer0_outputs[5801]));
    assign outputs[5383] = ~(layer0_outputs[9466]);
    assign outputs[5384] = layer0_outputs[9414];
    assign outputs[5385] = layer0_outputs[10156];
    assign outputs[5386] = ~((layer0_outputs[5800]) ^ (layer0_outputs[3084]));
    assign outputs[5387] = ~(layer0_outputs[9254]);
    assign outputs[5388] = ~((layer0_outputs[7910]) ^ (layer0_outputs[1639]));
    assign outputs[5389] = ~(layer0_outputs[4786]) | (layer0_outputs[1437]);
    assign outputs[5390] = ~((layer0_outputs[6921]) ^ (layer0_outputs[4766]));
    assign outputs[5391] = ~((layer0_outputs[10153]) ^ (layer0_outputs[695]));
    assign outputs[5392] = ~(layer0_outputs[9675]) | (layer0_outputs[9400]);
    assign outputs[5393] = ~((layer0_outputs[7898]) ^ (layer0_outputs[980]));
    assign outputs[5394] = ~(layer0_outputs[4297]);
    assign outputs[5395] = ~(layer0_outputs[9685]) | (layer0_outputs[6928]);
    assign outputs[5396] = ~((layer0_outputs[444]) ^ (layer0_outputs[6920]));
    assign outputs[5397] = ~(layer0_outputs[3953]) | (layer0_outputs[2836]);
    assign outputs[5398] = ~(layer0_outputs[1902]);
    assign outputs[5399] = ~(layer0_outputs[6557]);
    assign outputs[5400] = layer0_outputs[4478];
    assign outputs[5401] = ~((layer0_outputs[1759]) ^ (layer0_outputs[6273]));
    assign outputs[5402] = layer0_outputs[9224];
    assign outputs[5403] = layer0_outputs[7647];
    assign outputs[5404] = (layer0_outputs[3463]) ^ (layer0_outputs[6958]);
    assign outputs[5405] = ~(layer0_outputs[9502]);
    assign outputs[5406] = ~(layer0_outputs[9187]);
    assign outputs[5407] = ~((layer0_outputs[623]) & (layer0_outputs[5262]));
    assign outputs[5408] = layer0_outputs[6693];
    assign outputs[5409] = layer0_outputs[4569];
    assign outputs[5410] = (layer0_outputs[1819]) | (layer0_outputs[2364]);
    assign outputs[5411] = ~((layer0_outputs[9231]) ^ (layer0_outputs[5253]));
    assign outputs[5412] = ~((layer0_outputs[1896]) | (layer0_outputs[2762]));
    assign outputs[5413] = ~((layer0_outputs[4136]) & (layer0_outputs[3678]));
    assign outputs[5414] = (layer0_outputs[5407]) | (layer0_outputs[2549]);
    assign outputs[5415] = layer0_outputs[2808];
    assign outputs[5416] = ~(layer0_outputs[1698]);
    assign outputs[5417] = layer0_outputs[5026];
    assign outputs[5418] = ~(layer0_outputs[3157]);
    assign outputs[5419] = (layer0_outputs[1952]) & (layer0_outputs[2570]);
    assign outputs[5420] = ~((layer0_outputs[2857]) ^ (layer0_outputs[8570]));
    assign outputs[5421] = (layer0_outputs[6070]) | (layer0_outputs[142]);
    assign outputs[5422] = (layer0_outputs[8069]) ^ (layer0_outputs[4379]);
    assign outputs[5423] = layer0_outputs[9840];
    assign outputs[5424] = ~((layer0_outputs[6968]) ^ (layer0_outputs[8345]));
    assign outputs[5425] = ~(layer0_outputs[4824]);
    assign outputs[5426] = layer0_outputs[6674];
    assign outputs[5427] = layer0_outputs[6440];
    assign outputs[5428] = ~((layer0_outputs[8660]) ^ (layer0_outputs[323]));
    assign outputs[5429] = layer0_outputs[2947];
    assign outputs[5430] = (layer0_outputs[5546]) & (layer0_outputs[4428]);
    assign outputs[5431] = (layer0_outputs[4420]) ^ (layer0_outputs[9779]);
    assign outputs[5432] = layer0_outputs[1036];
    assign outputs[5433] = ~(layer0_outputs[5289]);
    assign outputs[5434] = layer0_outputs[983];
    assign outputs[5435] = (layer0_outputs[1279]) ^ (layer0_outputs[1270]);
    assign outputs[5436] = (layer0_outputs[8986]) ^ (layer0_outputs[6502]);
    assign outputs[5437] = (layer0_outputs[5703]) & ~(layer0_outputs[7379]);
    assign outputs[5438] = (layer0_outputs[6757]) ^ (layer0_outputs[4999]);
    assign outputs[5439] = ~((layer0_outputs[1830]) & (layer0_outputs[8026]));
    assign outputs[5440] = (layer0_outputs[8032]) ^ (layer0_outputs[1850]);
    assign outputs[5441] = ~((layer0_outputs[3173]) & (layer0_outputs[8005]));
    assign outputs[5442] = ~(layer0_outputs[4976]) | (layer0_outputs[10001]);
    assign outputs[5443] = ~(layer0_outputs[7029]) | (layer0_outputs[9506]);
    assign outputs[5444] = layer0_outputs[8193];
    assign outputs[5445] = ~(layer0_outputs[6830]);
    assign outputs[5446] = ~(layer0_outputs[3758]);
    assign outputs[5447] = (layer0_outputs[3058]) & ~(layer0_outputs[906]);
    assign outputs[5448] = (layer0_outputs[306]) & ~(layer0_outputs[3158]);
    assign outputs[5449] = ~(layer0_outputs[5217]) | (layer0_outputs[2779]);
    assign outputs[5450] = ~(layer0_outputs[2381]);
    assign outputs[5451] = ~((layer0_outputs[3294]) | (layer0_outputs[3970]));
    assign outputs[5452] = (layer0_outputs[7463]) ^ (layer0_outputs[124]);
    assign outputs[5453] = (layer0_outputs[1399]) ^ (layer0_outputs[4512]);
    assign outputs[5454] = ~((layer0_outputs[3703]) | (layer0_outputs[7407]));
    assign outputs[5455] = ~(layer0_outputs[6114]);
    assign outputs[5456] = layer0_outputs[4787];
    assign outputs[5457] = layer0_outputs[4399];
    assign outputs[5458] = ~(layer0_outputs[2105]) | (layer0_outputs[5526]);
    assign outputs[5459] = ~(layer0_outputs[4503]);
    assign outputs[5460] = 1'b1;
    assign outputs[5461] = layer0_outputs[3631];
    assign outputs[5462] = ~((layer0_outputs[2993]) ^ (layer0_outputs[9]));
    assign outputs[5463] = ~(layer0_outputs[5716]);
    assign outputs[5464] = (layer0_outputs[2835]) ^ (layer0_outputs[538]);
    assign outputs[5465] = layer0_outputs[6556];
    assign outputs[5466] = layer0_outputs[9921];
    assign outputs[5467] = ~(layer0_outputs[640]);
    assign outputs[5468] = ~((layer0_outputs[1540]) | (layer0_outputs[4685]));
    assign outputs[5469] = ~(layer0_outputs[6759]);
    assign outputs[5470] = ~((layer0_outputs[8621]) ^ (layer0_outputs[3287]));
    assign outputs[5471] = ~(layer0_outputs[6891]) | (layer0_outputs[2545]);
    assign outputs[5472] = layer0_outputs[7142];
    assign outputs[5473] = 1'b1;
    assign outputs[5474] = ~(layer0_outputs[2821]);
    assign outputs[5475] = layer0_outputs[4462];
    assign outputs[5476] = ~(layer0_outputs[5640]);
    assign outputs[5477] = layer0_outputs[5073];
    assign outputs[5478] = ~(layer0_outputs[2891]);
    assign outputs[5479] = layer0_outputs[7763];
    assign outputs[5480] = ~((layer0_outputs[2409]) ^ (layer0_outputs[671]));
    assign outputs[5481] = ~((layer0_outputs[7827]) ^ (layer0_outputs[5998]));
    assign outputs[5482] = layer0_outputs[2436];
    assign outputs[5483] = (layer0_outputs[2965]) ^ (layer0_outputs[4993]);
    assign outputs[5484] = (layer0_outputs[5363]) & ~(layer0_outputs[3954]);
    assign outputs[5485] = ~(layer0_outputs[5488]);
    assign outputs[5486] = ~((layer0_outputs[3669]) & (layer0_outputs[1772]));
    assign outputs[5487] = (layer0_outputs[9110]) & ~(layer0_outputs[6334]);
    assign outputs[5488] = layer0_outputs[9704];
    assign outputs[5489] = ~(layer0_outputs[8121]) | (layer0_outputs[9260]);
    assign outputs[5490] = ~((layer0_outputs[5159]) ^ (layer0_outputs[3571]));
    assign outputs[5491] = layer0_outputs[7959];
    assign outputs[5492] = (layer0_outputs[985]) & (layer0_outputs[2408]);
    assign outputs[5493] = ~(layer0_outputs[2165]);
    assign outputs[5494] = ~((layer0_outputs[7509]) ^ (layer0_outputs[1739]));
    assign outputs[5495] = ~(layer0_outputs[3679]) | (layer0_outputs[9639]);
    assign outputs[5496] = (layer0_outputs[3838]) ^ (layer0_outputs[2588]);
    assign outputs[5497] = ~((layer0_outputs[1838]) ^ (layer0_outputs[5362]));
    assign outputs[5498] = (layer0_outputs[8470]) | (layer0_outputs[2342]);
    assign outputs[5499] = ~(layer0_outputs[4606]);
    assign outputs[5500] = layer0_outputs[5274];
    assign outputs[5501] = (layer0_outputs[88]) & (layer0_outputs[8264]);
    assign outputs[5502] = (layer0_outputs[5296]) ^ (layer0_outputs[9693]);
    assign outputs[5503] = ~((layer0_outputs[8067]) | (layer0_outputs[483]));
    assign outputs[5504] = ~(layer0_outputs[8825]) | (layer0_outputs[2762]);
    assign outputs[5505] = ~((layer0_outputs[8761]) & (layer0_outputs[7708]));
    assign outputs[5506] = layer0_outputs[7099];
    assign outputs[5507] = ~(layer0_outputs[952]) | (layer0_outputs[5386]);
    assign outputs[5508] = ~(layer0_outputs[8206]);
    assign outputs[5509] = (layer0_outputs[4918]) & (layer0_outputs[1704]);
    assign outputs[5510] = (layer0_outputs[2627]) & ~(layer0_outputs[1622]);
    assign outputs[5511] = ~(layer0_outputs[5952]);
    assign outputs[5512] = layer0_outputs[3016];
    assign outputs[5513] = (layer0_outputs[2928]) & ~(layer0_outputs[8501]);
    assign outputs[5514] = ~((layer0_outputs[6537]) ^ (layer0_outputs[303]));
    assign outputs[5515] = (layer0_outputs[9112]) ^ (layer0_outputs[260]);
    assign outputs[5516] = layer0_outputs[5639];
    assign outputs[5517] = ~(layer0_outputs[9130]) | (layer0_outputs[833]);
    assign outputs[5518] = ~((layer0_outputs[3864]) ^ (layer0_outputs[3651]));
    assign outputs[5519] = ~(layer0_outputs[6206]);
    assign outputs[5520] = layer0_outputs[5300];
    assign outputs[5521] = ~(layer0_outputs[10056]);
    assign outputs[5522] = ~((layer0_outputs[6478]) ^ (layer0_outputs[8808]));
    assign outputs[5523] = ~(layer0_outputs[5916]);
    assign outputs[5524] = (layer0_outputs[2023]) ^ (layer0_outputs[1185]);
    assign outputs[5525] = (layer0_outputs[4216]) ^ (layer0_outputs[2530]);
    assign outputs[5526] = (layer0_outputs[6894]) ^ (layer0_outputs[6652]);
    assign outputs[5527] = (layer0_outputs[9100]) ^ (layer0_outputs[8687]);
    assign outputs[5528] = ~(layer0_outputs[6554]);
    assign outputs[5529] = (layer0_outputs[647]) | (layer0_outputs[511]);
    assign outputs[5530] = layer0_outputs[5388];
    assign outputs[5531] = ~(layer0_outputs[7208]);
    assign outputs[5532] = ~((layer0_outputs[5542]) ^ (layer0_outputs[10230]));
    assign outputs[5533] = ~(layer0_outputs[4315]);
    assign outputs[5534] = ~(layer0_outputs[9318]);
    assign outputs[5535] = (layer0_outputs[3859]) & (layer0_outputs[7885]);
    assign outputs[5536] = (layer0_outputs[6696]) ^ (layer0_outputs[5650]);
    assign outputs[5537] = (layer0_outputs[9500]) ^ (layer0_outputs[4080]);
    assign outputs[5538] = ~((layer0_outputs[9737]) | (layer0_outputs[1345]));
    assign outputs[5539] = layer0_outputs[8831];
    assign outputs[5540] = ~(layer0_outputs[705]);
    assign outputs[5541] = ~((layer0_outputs[5198]) ^ (layer0_outputs[8464]));
    assign outputs[5542] = ~((layer0_outputs[8209]) & (layer0_outputs[5785]));
    assign outputs[5543] = ~((layer0_outputs[6615]) ^ (layer0_outputs[4278]));
    assign outputs[5544] = ~(layer0_outputs[6138]);
    assign outputs[5545] = ~((layer0_outputs[9784]) ^ (layer0_outputs[8577]));
    assign outputs[5546] = ~(layer0_outputs[2039]);
    assign outputs[5547] = ~(layer0_outputs[2496]) | (layer0_outputs[1829]);
    assign outputs[5548] = ~(layer0_outputs[1834]);
    assign outputs[5549] = ~((layer0_outputs[6192]) ^ (layer0_outputs[6351]));
    assign outputs[5550] = layer0_outputs[8414];
    assign outputs[5551] = ~(layer0_outputs[9349]) | (layer0_outputs[9016]);
    assign outputs[5552] = (layer0_outputs[5765]) ^ (layer0_outputs[6566]);
    assign outputs[5553] = (layer0_outputs[1697]) ^ (layer0_outputs[8687]);
    assign outputs[5554] = (layer0_outputs[806]) | (layer0_outputs[9991]);
    assign outputs[5555] = ~(layer0_outputs[3714]) | (layer0_outputs[1900]);
    assign outputs[5556] = (layer0_outputs[5924]) | (layer0_outputs[1035]);
    assign outputs[5557] = ~(layer0_outputs[5069]);
    assign outputs[5558] = ~(layer0_outputs[9959]);
    assign outputs[5559] = ~((layer0_outputs[5005]) ^ (layer0_outputs[3896]));
    assign outputs[5560] = (layer0_outputs[8726]) | (layer0_outputs[9161]);
    assign outputs[5561] = ~((layer0_outputs[1865]) & (layer0_outputs[7591]));
    assign outputs[5562] = ~(layer0_outputs[9525]) | (layer0_outputs[8006]);
    assign outputs[5563] = (layer0_outputs[1671]) ^ (layer0_outputs[5248]);
    assign outputs[5564] = ~(layer0_outputs[9333]) | (layer0_outputs[750]);
    assign outputs[5565] = ~(layer0_outputs[6798]);
    assign outputs[5566] = (layer0_outputs[6802]) & ~(layer0_outputs[8725]);
    assign outputs[5567] = (layer0_outputs[228]) ^ (layer0_outputs[5100]);
    assign outputs[5568] = ~((layer0_outputs[9423]) ^ (layer0_outputs[6978]));
    assign outputs[5569] = ~((layer0_outputs[1946]) ^ (layer0_outputs[6883]));
    assign outputs[5570] = ~((layer0_outputs[8724]) | (layer0_outputs[1500]));
    assign outputs[5571] = ~(layer0_outputs[10094]);
    assign outputs[5572] = ~((layer0_outputs[714]) & (layer0_outputs[5317]));
    assign outputs[5573] = (layer0_outputs[5391]) ^ (layer0_outputs[7245]);
    assign outputs[5574] = ~(layer0_outputs[1490]);
    assign outputs[5575] = ~(layer0_outputs[7011]) | (layer0_outputs[9331]);
    assign outputs[5576] = ~(layer0_outputs[1770]);
    assign outputs[5577] = ~(layer0_outputs[7043]);
    assign outputs[5578] = ~((layer0_outputs[8665]) & (layer0_outputs[6771]));
    assign outputs[5579] = ~((layer0_outputs[7243]) | (layer0_outputs[3503]));
    assign outputs[5580] = ~((layer0_outputs[4639]) ^ (layer0_outputs[700]));
    assign outputs[5581] = (layer0_outputs[6432]) ^ (layer0_outputs[2584]);
    assign outputs[5582] = layer0_outputs[1816];
    assign outputs[5583] = (layer0_outputs[2292]) ^ (layer0_outputs[6495]);
    assign outputs[5584] = ~(layer0_outputs[9914]);
    assign outputs[5585] = (layer0_outputs[2287]) | (layer0_outputs[3943]);
    assign outputs[5586] = layer0_outputs[10207];
    assign outputs[5587] = ~(layer0_outputs[5724]) | (layer0_outputs[2669]);
    assign outputs[5588] = layer0_outputs[8180];
    assign outputs[5589] = ~(layer0_outputs[10078]);
    assign outputs[5590] = (layer0_outputs[8557]) ^ (layer0_outputs[10163]);
    assign outputs[5591] = layer0_outputs[6962];
    assign outputs[5592] = layer0_outputs[1842];
    assign outputs[5593] = layer0_outputs[5892];
    assign outputs[5594] = (layer0_outputs[9337]) | (layer0_outputs[8973]);
    assign outputs[5595] = ~(layer0_outputs[4367]);
    assign outputs[5596] = (layer0_outputs[6760]) & ~(layer0_outputs[9652]);
    assign outputs[5597] = ~((layer0_outputs[6448]) ^ (layer0_outputs[7276]));
    assign outputs[5598] = ~(layer0_outputs[61]);
    assign outputs[5599] = ~(layer0_outputs[10060]);
    assign outputs[5600] = ~((layer0_outputs[6800]) & (layer0_outputs[7741]));
    assign outputs[5601] = layer0_outputs[943];
    assign outputs[5602] = (layer0_outputs[1416]) ^ (layer0_outputs[8941]);
    assign outputs[5603] = (layer0_outputs[5113]) | (layer0_outputs[1543]);
    assign outputs[5604] = ~(layer0_outputs[10000]);
    assign outputs[5605] = ~(layer0_outputs[919]) | (layer0_outputs[1059]);
    assign outputs[5606] = (layer0_outputs[1532]) ^ (layer0_outputs[8648]);
    assign outputs[5607] = layer0_outputs[2843];
    assign outputs[5608] = (layer0_outputs[6815]) & (layer0_outputs[5149]);
    assign outputs[5609] = ~(layer0_outputs[6650]) | (layer0_outputs[6383]);
    assign outputs[5610] = layer0_outputs[1425];
    assign outputs[5611] = ~((layer0_outputs[280]) ^ (layer0_outputs[7645]));
    assign outputs[5612] = layer0_outputs[829];
    assign outputs[5613] = ~(layer0_outputs[10218]);
    assign outputs[5614] = ~(layer0_outputs[7103]) | (layer0_outputs[8393]);
    assign outputs[5615] = layer0_outputs[434];
    assign outputs[5616] = ~(layer0_outputs[6094]) | (layer0_outputs[4324]);
    assign outputs[5617] = layer0_outputs[7611];
    assign outputs[5618] = ~((layer0_outputs[6733]) ^ (layer0_outputs[2264]));
    assign outputs[5619] = ~((layer0_outputs[1488]) ^ (layer0_outputs[8299]));
    assign outputs[5620] = ~((layer0_outputs[4407]) ^ (layer0_outputs[5643]));
    assign outputs[5621] = ~((layer0_outputs[1232]) ^ (layer0_outputs[1954]));
    assign outputs[5622] = layer0_outputs[8776];
    assign outputs[5623] = (layer0_outputs[1811]) ^ (layer0_outputs[942]);
    assign outputs[5624] = ~((layer0_outputs[8649]) & (layer0_outputs[5376]));
    assign outputs[5625] = layer0_outputs[1360];
    assign outputs[5626] = ~(layer0_outputs[1411]) | (layer0_outputs[1469]);
    assign outputs[5627] = (layer0_outputs[3961]) ^ (layer0_outputs[7245]);
    assign outputs[5628] = (layer0_outputs[2709]) ^ (layer0_outputs[3019]);
    assign outputs[5629] = ~(layer0_outputs[5033]);
    assign outputs[5630] = ~((layer0_outputs[63]) ^ (layer0_outputs[10152]));
    assign outputs[5631] = layer0_outputs[4951];
    assign outputs[5632] = (layer0_outputs[819]) & ~(layer0_outputs[4991]);
    assign outputs[5633] = ~((layer0_outputs[4932]) | (layer0_outputs[9305]));
    assign outputs[5634] = (layer0_outputs[6116]) ^ (layer0_outputs[4627]);
    assign outputs[5635] = ~(layer0_outputs[4720]) | (layer0_outputs[4017]);
    assign outputs[5636] = ~((layer0_outputs[5989]) ^ (layer0_outputs[6392]));
    assign outputs[5637] = (layer0_outputs[6741]) ^ (layer0_outputs[914]);
    assign outputs[5638] = (layer0_outputs[6429]) & (layer0_outputs[381]);
    assign outputs[5639] = (layer0_outputs[9878]) | (layer0_outputs[8725]);
    assign outputs[5640] = layer0_outputs[6177];
    assign outputs[5641] = (layer0_outputs[7707]) ^ (layer0_outputs[2467]);
    assign outputs[5642] = (layer0_outputs[4886]) ^ (layer0_outputs[4607]);
    assign outputs[5643] = ~((layer0_outputs[6260]) & (layer0_outputs[4829]));
    assign outputs[5644] = ~((layer0_outputs[9536]) & (layer0_outputs[8807]));
    assign outputs[5645] = layer0_outputs[6685];
    assign outputs[5646] = layer0_outputs[7600];
    assign outputs[5647] = (layer0_outputs[9450]) ^ (layer0_outputs[2151]);
    assign outputs[5648] = ~((layer0_outputs[3032]) & (layer0_outputs[9017]));
    assign outputs[5649] = (layer0_outputs[2354]) ^ (layer0_outputs[1705]);
    assign outputs[5650] = ~(layer0_outputs[9045]);
    assign outputs[5651] = 1'b1;
    assign outputs[5652] = (layer0_outputs[1842]) & (layer0_outputs[3004]);
    assign outputs[5653] = ~(layer0_outputs[5882]);
    assign outputs[5654] = layer0_outputs[6746];
    assign outputs[5655] = ~(layer0_outputs[5899]) | (layer0_outputs[9544]);
    assign outputs[5656] = ~((layer0_outputs[9251]) ^ (layer0_outputs[1408]));
    assign outputs[5657] = ~(layer0_outputs[3791]) | (layer0_outputs[2827]);
    assign outputs[5658] = (layer0_outputs[3515]) & ~(layer0_outputs[6184]);
    assign outputs[5659] = ~(layer0_outputs[2170]);
    assign outputs[5660] = layer0_outputs[5047];
    assign outputs[5661] = ~(layer0_outputs[4248]);
    assign outputs[5662] = ~((layer0_outputs[9835]) | (layer0_outputs[539]));
    assign outputs[5663] = (layer0_outputs[4831]) ^ (layer0_outputs[1191]);
    assign outputs[5664] = 1'b1;
    assign outputs[5665] = layer0_outputs[3175];
    assign outputs[5666] = (layer0_outputs[3259]) ^ (layer0_outputs[3755]);
    assign outputs[5667] = (layer0_outputs[9600]) & (layer0_outputs[6315]);
    assign outputs[5668] = ~((layer0_outputs[8892]) ^ (layer0_outputs[7995]));
    assign outputs[5669] = layer0_outputs[1993];
    assign outputs[5670] = layer0_outputs[7378];
    assign outputs[5671] = (layer0_outputs[3320]) ^ (layer0_outputs[5535]);
    assign outputs[5672] = ~((layer0_outputs[246]) & (layer0_outputs[2199]));
    assign outputs[5673] = ~(layer0_outputs[361]) | (layer0_outputs[2215]);
    assign outputs[5674] = (layer0_outputs[1274]) ^ (layer0_outputs[9904]);
    assign outputs[5675] = layer0_outputs[6942];
    assign outputs[5676] = (layer0_outputs[2175]) ^ (layer0_outputs[4565]);
    assign outputs[5677] = (layer0_outputs[2514]) ^ (layer0_outputs[6319]);
    assign outputs[5678] = layer0_outputs[1159];
    assign outputs[5679] = layer0_outputs[8335];
    assign outputs[5680] = ~((layer0_outputs[6507]) ^ (layer0_outputs[9824]));
    assign outputs[5681] = ~(layer0_outputs[7843]);
    assign outputs[5682] = ~(layer0_outputs[2054]);
    assign outputs[5683] = layer0_outputs[7635];
    assign outputs[5684] = (layer0_outputs[2898]) ^ (layer0_outputs[5407]);
    assign outputs[5685] = (layer0_outputs[4009]) ^ (layer0_outputs[8558]);
    assign outputs[5686] = ~(layer0_outputs[4364]);
    assign outputs[5687] = ~(layer0_outputs[8683]) | (layer0_outputs[5274]);
    assign outputs[5688] = (layer0_outputs[9862]) & (layer0_outputs[3327]);
    assign outputs[5689] = ~(layer0_outputs[6607]);
    assign outputs[5690] = (layer0_outputs[2144]) & ~(layer0_outputs[4882]);
    assign outputs[5691] = ~((layer0_outputs[4921]) ^ (layer0_outputs[7935]));
    assign outputs[5692] = (layer0_outputs[1410]) ^ (layer0_outputs[535]);
    assign outputs[5693] = ~((layer0_outputs[9931]) | (layer0_outputs[9920]));
    assign outputs[5694] = (layer0_outputs[6464]) ^ (layer0_outputs[147]);
    assign outputs[5695] = ~((layer0_outputs[5953]) ^ (layer0_outputs[2940]));
    assign outputs[5696] = (layer0_outputs[8785]) ^ (layer0_outputs[3109]);
    assign outputs[5697] = ~(layer0_outputs[9316]);
    assign outputs[5698] = ~(layer0_outputs[698]);
    assign outputs[5699] = (layer0_outputs[8772]) ^ (layer0_outputs[7837]);
    assign outputs[5700] = ~((layer0_outputs[267]) ^ (layer0_outputs[7663]));
    assign outputs[5701] = (layer0_outputs[948]) ^ (layer0_outputs[9158]);
    assign outputs[5702] = layer0_outputs[3024];
    assign outputs[5703] = ~((layer0_outputs[460]) ^ (layer0_outputs[1864]));
    assign outputs[5704] = ~((layer0_outputs[4146]) ^ (layer0_outputs[2574]));
    assign outputs[5705] = ~(layer0_outputs[4474]) | (layer0_outputs[6849]);
    assign outputs[5706] = ~(layer0_outputs[6823]);
    assign outputs[5707] = (layer0_outputs[8652]) ^ (layer0_outputs[8922]);
    assign outputs[5708] = layer0_outputs[7844];
    assign outputs[5709] = (layer0_outputs[8627]) ^ (layer0_outputs[58]);
    assign outputs[5710] = ~(layer0_outputs[8784]);
    assign outputs[5711] = ~(layer0_outputs[7968]);
    assign outputs[5712] = layer0_outputs[5335];
    assign outputs[5713] = (layer0_outputs[405]) & ~(layer0_outputs[4958]);
    assign outputs[5714] = ~((layer0_outputs[2466]) | (layer0_outputs[7510]));
    assign outputs[5715] = layer0_outputs[9827];
    assign outputs[5716] = layer0_outputs[6484];
    assign outputs[5717] = ~((layer0_outputs[1228]) ^ (layer0_outputs[9341]));
    assign outputs[5718] = layer0_outputs[9894];
    assign outputs[5719] = (layer0_outputs[2856]) ^ (layer0_outputs[10007]);
    assign outputs[5720] = (layer0_outputs[8040]) ^ (layer0_outputs[4766]);
    assign outputs[5721] = ~(layer0_outputs[2630]);
    assign outputs[5722] = (layer0_outputs[4067]) & (layer0_outputs[4239]);
    assign outputs[5723] = layer0_outputs[5223];
    assign outputs[5724] = layer0_outputs[2879];
    assign outputs[5725] = layer0_outputs[2885];
    assign outputs[5726] = ~(layer0_outputs[6529]);
    assign outputs[5727] = ~(layer0_outputs[8645]);
    assign outputs[5728] = (layer0_outputs[9515]) ^ (layer0_outputs[615]);
    assign outputs[5729] = (layer0_outputs[4081]) & ~(layer0_outputs[3509]);
    assign outputs[5730] = ~((layer0_outputs[7533]) & (layer0_outputs[5991]));
    assign outputs[5731] = ~((layer0_outputs[393]) | (layer0_outputs[6047]));
    assign outputs[5732] = ~((layer0_outputs[2905]) ^ (layer0_outputs[9845]));
    assign outputs[5733] = ~((layer0_outputs[2571]) | (layer0_outputs[217]));
    assign outputs[5734] = layer0_outputs[7323];
    assign outputs[5735] = ~(layer0_outputs[6861]);
    assign outputs[5736] = (layer0_outputs[4848]) & (layer0_outputs[9512]);
    assign outputs[5737] = (layer0_outputs[8002]) ^ (layer0_outputs[10148]);
    assign outputs[5738] = layer0_outputs[7267];
    assign outputs[5739] = ~(layer0_outputs[8400]);
    assign outputs[5740] = layer0_outputs[347];
    assign outputs[5741] = (layer0_outputs[2723]) & ~(layer0_outputs[2562]);
    assign outputs[5742] = (layer0_outputs[2212]) ^ (layer0_outputs[6732]);
    assign outputs[5743] = ~(layer0_outputs[2687]);
    assign outputs[5744] = ~((layer0_outputs[3103]) ^ (layer0_outputs[8915]));
    assign outputs[5745] = layer0_outputs[7929];
    assign outputs[5746] = ~(layer0_outputs[4060]) | (layer0_outputs[1526]);
    assign outputs[5747] = ~(layer0_outputs[4023]);
    assign outputs[5748] = (layer0_outputs[110]) ^ (layer0_outputs[5920]);
    assign outputs[5749] = ~((layer0_outputs[2038]) & (layer0_outputs[4225]));
    assign outputs[5750] = layer0_outputs[1516];
    assign outputs[5751] = layer0_outputs[5056];
    assign outputs[5752] = ~(layer0_outputs[8852]) | (layer0_outputs[5692]);
    assign outputs[5753] = (layer0_outputs[2219]) ^ (layer0_outputs[2532]);
    assign outputs[5754] = layer0_outputs[6506];
    assign outputs[5755] = layer0_outputs[5775];
    assign outputs[5756] = ~(layer0_outputs[5592]);
    assign outputs[5757] = ~(layer0_outputs[3740]);
    assign outputs[5758] = ~(layer0_outputs[3994]);
    assign outputs[5759] = (layer0_outputs[2751]) | (layer0_outputs[1129]);
    assign outputs[5760] = (layer0_outputs[4989]) | (layer0_outputs[1107]);
    assign outputs[5761] = ~(layer0_outputs[5876]);
    assign outputs[5762] = (layer0_outputs[5833]) & (layer0_outputs[2313]);
    assign outputs[5763] = ~(layer0_outputs[6253]);
    assign outputs[5764] = ~((layer0_outputs[4926]) ^ (layer0_outputs[8608]));
    assign outputs[5765] = layer0_outputs[3112];
    assign outputs[5766] = 1'b1;
    assign outputs[5767] = ~(layer0_outputs[3508]);
    assign outputs[5768] = (layer0_outputs[9932]) | (layer0_outputs[6827]);
    assign outputs[5769] = ~((layer0_outputs[5901]) ^ (layer0_outputs[4350]));
    assign outputs[5770] = (layer0_outputs[4014]) ^ (layer0_outputs[6024]);
    assign outputs[5771] = (layer0_outputs[8195]) ^ (layer0_outputs[5589]);
    assign outputs[5772] = ~((layer0_outputs[1243]) | (layer0_outputs[6819]));
    assign outputs[5773] = ~(layer0_outputs[8257]) | (layer0_outputs[7474]);
    assign outputs[5774] = ~(layer0_outputs[1403]);
    assign outputs[5775] = (layer0_outputs[4715]) ^ (layer0_outputs[8817]);
    assign outputs[5776] = ~(layer0_outputs[6751]);
    assign outputs[5777] = layer0_outputs[9767];
    assign outputs[5778] = layer0_outputs[3908];
    assign outputs[5779] = (layer0_outputs[9611]) ^ (layer0_outputs[9477]);
    assign outputs[5780] = (layer0_outputs[5524]) ^ (layer0_outputs[6517]);
    assign outputs[5781] = ~(layer0_outputs[7514]);
    assign outputs[5782] = ~((layer0_outputs[449]) ^ (layer0_outputs[8783]));
    assign outputs[5783] = layer0_outputs[1840];
    assign outputs[5784] = ~((layer0_outputs[6028]) ^ (layer0_outputs[2184]));
    assign outputs[5785] = ~(layer0_outputs[6282]);
    assign outputs[5786] = (layer0_outputs[4202]) | (layer0_outputs[7933]);
    assign outputs[5787] = (layer0_outputs[4630]) | (layer0_outputs[3150]);
    assign outputs[5788] = ~(layer0_outputs[6879]);
    assign outputs[5789] = (layer0_outputs[4273]) ^ (layer0_outputs[3203]);
    assign outputs[5790] = layer0_outputs[7008];
    assign outputs[5791] = (layer0_outputs[506]) ^ (layer0_outputs[5946]);
    assign outputs[5792] = layer0_outputs[5167];
    assign outputs[5793] = layer0_outputs[9040];
    assign outputs[5794] = ~(layer0_outputs[2039]);
    assign outputs[5795] = ~((layer0_outputs[823]) & (layer0_outputs[9787]));
    assign outputs[5796] = layer0_outputs[10077];
    assign outputs[5797] = ~((layer0_outputs[2749]) ^ (layer0_outputs[4198]));
    assign outputs[5798] = ~(layer0_outputs[6676]) | (layer0_outputs[1288]);
    assign outputs[5799] = (layer0_outputs[2725]) ^ (layer0_outputs[4950]);
    assign outputs[5800] = ~(layer0_outputs[4597]);
    assign outputs[5801] = layer0_outputs[4470];
    assign outputs[5802] = (layer0_outputs[897]) | (layer0_outputs[5832]);
    assign outputs[5803] = (layer0_outputs[5527]) ^ (layer0_outputs[6164]);
    assign outputs[5804] = ~(layer0_outputs[401]);
    assign outputs[5805] = ~(layer0_outputs[6086]) | (layer0_outputs[9188]);
    assign outputs[5806] = ~(layer0_outputs[1247]);
    assign outputs[5807] = (layer0_outputs[2503]) ^ (layer0_outputs[3289]);
    assign outputs[5808] = ~(layer0_outputs[9614]);
    assign outputs[5809] = ~((layer0_outputs[1740]) & (layer0_outputs[3927]));
    assign outputs[5810] = layer0_outputs[2975];
    assign outputs[5811] = ~(layer0_outputs[9993]);
    assign outputs[5812] = ~((layer0_outputs[9240]) | (layer0_outputs[5330]));
    assign outputs[5813] = layer0_outputs[889];
    assign outputs[5814] = ~((layer0_outputs[10034]) ^ (layer0_outputs[3527]));
    assign outputs[5815] = ~(layer0_outputs[6945]);
    assign outputs[5816] = layer0_outputs[4331];
    assign outputs[5817] = layer0_outputs[8567];
    assign outputs[5818] = ~((layer0_outputs[5727]) & (layer0_outputs[2838]));
    assign outputs[5819] = ~((layer0_outputs[416]) ^ (layer0_outputs[2000]));
    assign outputs[5820] = ~((layer0_outputs[6646]) ^ (layer0_outputs[247]));
    assign outputs[5821] = (layer0_outputs[9188]) ^ (layer0_outputs[7847]);
    assign outputs[5822] = 1'b1;
    assign outputs[5823] = ~(layer0_outputs[7287]) | (layer0_outputs[9805]);
    assign outputs[5824] = (layer0_outputs[9015]) & ~(layer0_outputs[435]);
    assign outputs[5825] = layer0_outputs[8729];
    assign outputs[5826] = (layer0_outputs[7506]) | (layer0_outputs[10103]);
    assign outputs[5827] = ~((layer0_outputs[908]) ^ (layer0_outputs[3644]));
    assign outputs[5828] = layer0_outputs[5774];
    assign outputs[5829] = layer0_outputs[8748];
    assign outputs[5830] = ~(layer0_outputs[2685]);
    assign outputs[5831] = (layer0_outputs[6789]) & ~(layer0_outputs[2539]);
    assign outputs[5832] = (layer0_outputs[8385]) | (layer0_outputs[7815]);
    assign outputs[5833] = layer0_outputs[493];
    assign outputs[5834] = (layer0_outputs[8991]) ^ (layer0_outputs[6160]);
    assign outputs[5835] = layer0_outputs[5681];
    assign outputs[5836] = layer0_outputs[336];
    assign outputs[5837] = ~(layer0_outputs[6892]);
    assign outputs[5838] = ~((layer0_outputs[8814]) ^ (layer0_outputs[5271]));
    assign outputs[5839] = layer0_outputs[7088];
    assign outputs[5840] = ~(layer0_outputs[220]) | (layer0_outputs[565]);
    assign outputs[5841] = ~(layer0_outputs[2143]);
    assign outputs[5842] = (layer0_outputs[9594]) & (layer0_outputs[6712]);
    assign outputs[5843] = (layer0_outputs[6427]) & ~(layer0_outputs[3695]);
    assign outputs[5844] = ~(layer0_outputs[2421]) | (layer0_outputs[7028]);
    assign outputs[5845] = (layer0_outputs[5697]) & ~(layer0_outputs[317]);
    assign outputs[5846] = ~(layer0_outputs[594]);
    assign outputs[5847] = layer0_outputs[4765];
    assign outputs[5848] = ~(layer0_outputs[2281]);
    assign outputs[5849] = layer0_outputs[7549];
    assign outputs[5850] = ~((layer0_outputs[7593]) | (layer0_outputs[9571]));
    assign outputs[5851] = (layer0_outputs[7465]) | (layer0_outputs[7280]);
    assign outputs[5852] = ~(layer0_outputs[7185]);
    assign outputs[5853] = layer0_outputs[1088];
    assign outputs[5854] = ~((layer0_outputs[1738]) | (layer0_outputs[8142]));
    assign outputs[5855] = ~((layer0_outputs[2775]) ^ (layer0_outputs[6578]));
    assign outputs[5856] = ~(layer0_outputs[1555]);
    assign outputs[5857] = (layer0_outputs[5104]) ^ (layer0_outputs[9313]);
    assign outputs[5858] = ~(layer0_outputs[7481]);
    assign outputs[5859] = (layer0_outputs[4094]) & ~(layer0_outputs[9576]);
    assign outputs[5860] = ~(layer0_outputs[1845]);
    assign outputs[5861] = (layer0_outputs[5611]) ^ (layer0_outputs[1728]);
    assign outputs[5862] = ~((layer0_outputs[10135]) ^ (layer0_outputs[8038]));
    assign outputs[5863] = ~(layer0_outputs[3447]);
    assign outputs[5864] = ~((layer0_outputs[9459]) ^ (layer0_outputs[7753]));
    assign outputs[5865] = ~((layer0_outputs[2853]) ^ (layer0_outputs[3091]));
    assign outputs[5866] = (layer0_outputs[3255]) ^ (layer0_outputs[4575]);
    assign outputs[5867] = (layer0_outputs[6106]) ^ (layer0_outputs[9065]);
    assign outputs[5868] = (layer0_outputs[7983]) ^ (layer0_outputs[1836]);
    assign outputs[5869] = (layer0_outputs[5195]) & (layer0_outputs[4479]);
    assign outputs[5870] = (layer0_outputs[2777]) & (layer0_outputs[5612]);
    assign outputs[5871] = ~(layer0_outputs[5660]) | (layer0_outputs[2708]);
    assign outputs[5872] = ~((layer0_outputs[1682]) ^ (layer0_outputs[7866]));
    assign outputs[5873] = ~(layer0_outputs[2006]);
    assign outputs[5874] = (layer0_outputs[1817]) & (layer0_outputs[2628]);
    assign outputs[5875] = layer0_outputs[6756];
    assign outputs[5876] = (layer0_outputs[7224]) & (layer0_outputs[344]);
    assign outputs[5877] = layer0_outputs[5132];
    assign outputs[5878] = ~((layer0_outputs[7186]) | (layer0_outputs[6459]));
    assign outputs[5879] = layer0_outputs[1225];
    assign outputs[5880] = (layer0_outputs[1620]) | (layer0_outputs[5026]);
    assign outputs[5881] = (layer0_outputs[1358]) ^ (layer0_outputs[4648]);
    assign outputs[5882] = layer0_outputs[8823];
    assign outputs[5883] = ~(layer0_outputs[7507]) | (layer0_outputs[2353]);
    assign outputs[5884] = ~((layer0_outputs[8406]) ^ (layer0_outputs[1135]));
    assign outputs[5885] = (layer0_outputs[3822]) ^ (layer0_outputs[5539]);
    assign outputs[5886] = (layer0_outputs[4185]) ^ (layer0_outputs[7747]);
    assign outputs[5887] = (layer0_outputs[8487]) | (layer0_outputs[2595]);
    assign outputs[5888] = layer0_outputs[1819];
    assign outputs[5889] = ~(layer0_outputs[1503]) | (layer0_outputs[1805]);
    assign outputs[5890] = 1'b1;
    assign outputs[5891] = ~((layer0_outputs[7112]) ^ (layer0_outputs[4201]));
    assign outputs[5892] = layer0_outputs[1595];
    assign outputs[5893] = (layer0_outputs[894]) & (layer0_outputs[4579]);
    assign outputs[5894] = (layer0_outputs[9452]) ^ (layer0_outputs[2745]);
    assign outputs[5895] = layer0_outputs[8315];
    assign outputs[5896] = ~((layer0_outputs[2869]) & (layer0_outputs[5282]));
    assign outputs[5897] = layer0_outputs[964];
    assign outputs[5898] = ~((layer0_outputs[4424]) ^ (layer0_outputs[600]));
    assign outputs[5899] = ~(layer0_outputs[8827]) | (layer0_outputs[5709]);
    assign outputs[5900] = (layer0_outputs[171]) | (layer0_outputs[6901]);
    assign outputs[5901] = (layer0_outputs[3160]) & ~(layer0_outputs[3223]);
    assign outputs[5902] = layer0_outputs[2717];
    assign outputs[5903] = (layer0_outputs[9720]) | (layer0_outputs[9467]);
    assign outputs[5904] = ~(layer0_outputs[21]);
    assign outputs[5905] = (layer0_outputs[5221]) ^ (layer0_outputs[5050]);
    assign outputs[5906] = ~(layer0_outputs[3995]) | (layer0_outputs[990]);
    assign outputs[5907] = (layer0_outputs[118]) & (layer0_outputs[5898]);
    assign outputs[5908] = ~((layer0_outputs[143]) & (layer0_outputs[6392]));
    assign outputs[5909] = (layer0_outputs[9495]) ^ (layer0_outputs[3815]);
    assign outputs[5910] = ~(layer0_outputs[8887]);
    assign outputs[5911] = (layer0_outputs[71]) ^ (layer0_outputs[7997]);
    assign outputs[5912] = ~(layer0_outputs[3614]);
    assign outputs[5913] = ~((layer0_outputs[6211]) ^ (layer0_outputs[4323]));
    assign outputs[5914] = (layer0_outputs[1722]) & (layer0_outputs[6508]);
    assign outputs[5915] = ~((layer0_outputs[8803]) & (layer0_outputs[8373]));
    assign outputs[5916] = ~(layer0_outputs[9456]);
    assign outputs[5917] = ~((layer0_outputs[7942]) ^ (layer0_outputs[9738]));
    assign outputs[5918] = ~((layer0_outputs[6898]) ^ (layer0_outputs[4695]));
    assign outputs[5919] = ~(layer0_outputs[2585]);
    assign outputs[5920] = layer0_outputs[6066];
    assign outputs[5921] = ~(layer0_outputs[7394]);
    assign outputs[5922] = (layer0_outputs[1935]) ^ (layer0_outputs[6516]);
    assign outputs[5923] = layer0_outputs[4165];
    assign outputs[5924] = ~(layer0_outputs[6128]);
    assign outputs[5925] = ~(layer0_outputs[1953]);
    assign outputs[5926] = ~(layer0_outputs[3676]);
    assign outputs[5927] = (layer0_outputs[3992]) ^ (layer0_outputs[1140]);
    assign outputs[5928] = (layer0_outputs[3849]) ^ (layer0_outputs[2041]);
    assign outputs[5929] = layer0_outputs[4572];
    assign outputs[5930] = ~(layer0_outputs[43]);
    assign outputs[5931] = ~(layer0_outputs[1902]);
    assign outputs[5932] = ~(layer0_outputs[9945]);
    assign outputs[5933] = (layer0_outputs[270]) ^ (layer0_outputs[1750]);
    assign outputs[5934] = ~((layer0_outputs[9584]) ^ (layer0_outputs[3910]));
    assign outputs[5935] = ~((layer0_outputs[8461]) | (layer0_outputs[3114]));
    assign outputs[5936] = (layer0_outputs[5396]) ^ (layer0_outputs[40]);
    assign outputs[5937] = ~(layer0_outputs[6191]);
    assign outputs[5938] = ~((layer0_outputs[4870]) ^ (layer0_outputs[7193]));
    assign outputs[5939] = (layer0_outputs[727]) & (layer0_outputs[4205]);
    assign outputs[5940] = layer0_outputs[273];
    assign outputs[5941] = ~(layer0_outputs[718]);
    assign outputs[5942] = ~(layer0_outputs[4498]);
    assign outputs[5943] = ~((layer0_outputs[6003]) ^ (layer0_outputs[1921]));
    assign outputs[5944] = ~((layer0_outputs[9425]) | (layer0_outputs[6569]));
    assign outputs[5945] = (layer0_outputs[8988]) ^ (layer0_outputs[9649]);
    assign outputs[5946] = ~(layer0_outputs[9421]);
    assign outputs[5947] = (layer0_outputs[6983]) & ~(layer0_outputs[1564]);
    assign outputs[5948] = (layer0_outputs[5471]) ^ (layer0_outputs[6916]);
    assign outputs[5949] = ~(layer0_outputs[2635]);
    assign outputs[5950] = (layer0_outputs[3473]) ^ (layer0_outputs[9343]);
    assign outputs[5951] = ~(layer0_outputs[5230]) | (layer0_outputs[9813]);
    assign outputs[5952] = layer0_outputs[6742];
    assign outputs[5953] = layer0_outputs[1360];
    assign outputs[5954] = ~(layer0_outputs[10223]);
    assign outputs[5955] = (layer0_outputs[5156]) ^ (layer0_outputs[855]);
    assign outputs[5956] = (layer0_outputs[8317]) ^ (layer0_outputs[7496]);
    assign outputs[5957] = layer0_outputs[1544];
    assign outputs[5958] = ~((layer0_outputs[904]) ^ (layer0_outputs[1108]));
    assign outputs[5959] = ~(layer0_outputs[9883]);
    assign outputs[5960] = layer0_outputs[976];
    assign outputs[5961] = ~(layer0_outputs[9313]);
    assign outputs[5962] = ~(layer0_outputs[7642]) | (layer0_outputs[4961]);
    assign outputs[5963] = ~((layer0_outputs[8269]) & (layer0_outputs[4100]));
    assign outputs[5964] = layer0_outputs[637];
    assign outputs[5965] = (layer0_outputs[9020]) ^ (layer0_outputs[4069]);
    assign outputs[5966] = (layer0_outputs[8474]) ^ (layer0_outputs[10205]);
    assign outputs[5967] = layer0_outputs[8633];
    assign outputs[5968] = ~(layer0_outputs[4330]);
    assign outputs[5969] = ~(layer0_outputs[1886]);
    assign outputs[5970] = ~(layer0_outputs[9345]) | (layer0_outputs[341]);
    assign outputs[5971] = layer0_outputs[9028];
    assign outputs[5972] = (layer0_outputs[3705]) ^ (layer0_outputs[5193]);
    assign outputs[5973] = ~(layer0_outputs[1087]);
    assign outputs[5974] = ~(layer0_outputs[3451]);
    assign outputs[5975] = (layer0_outputs[1273]) & ~(layer0_outputs[7293]);
    assign outputs[5976] = layer0_outputs[4973];
    assign outputs[5977] = layer0_outputs[2992];
    assign outputs[5978] = ~((layer0_outputs[1926]) ^ (layer0_outputs[7833]));
    assign outputs[5979] = ~(layer0_outputs[2463]);
    assign outputs[5980] = ~(layer0_outputs[2509]);
    assign outputs[5981] = ~(layer0_outputs[8887]);
    assign outputs[5982] = ~(layer0_outputs[1624]);
    assign outputs[5983] = (layer0_outputs[8070]) ^ (layer0_outputs[9794]);
    assign outputs[5984] = (layer0_outputs[2438]) ^ (layer0_outputs[3417]);
    assign outputs[5985] = ~(layer0_outputs[3272]);
    assign outputs[5986] = ~((layer0_outputs[1685]) | (layer0_outputs[10192]));
    assign outputs[5987] = ~(layer0_outputs[8588]);
    assign outputs[5988] = ~(layer0_outputs[8416]);
    assign outputs[5989] = ~(layer0_outputs[9931]);
    assign outputs[5990] = ~(layer0_outputs[9503]);
    assign outputs[5991] = (layer0_outputs[6859]) | (layer0_outputs[3268]);
    assign outputs[5992] = ~(layer0_outputs[6120]);
    assign outputs[5993] = layer0_outputs[2050];
    assign outputs[5994] = 1'b1;
    assign outputs[5995] = ~(layer0_outputs[7219]);
    assign outputs[5996] = (layer0_outputs[7239]) & ~(layer0_outputs[723]);
    assign outputs[5997] = (layer0_outputs[10083]) | (layer0_outputs[2942]);
    assign outputs[5998] = ~((layer0_outputs[572]) ^ (layer0_outputs[8973]));
    assign outputs[5999] = (layer0_outputs[1880]) ^ (layer0_outputs[9357]);
    assign outputs[6000] = (layer0_outputs[3641]) ^ (layer0_outputs[8255]);
    assign outputs[6001] = layer0_outputs[669];
    assign outputs[6002] = ~(layer0_outputs[4387]) | (layer0_outputs[450]);
    assign outputs[6003] = ~((layer0_outputs[186]) ^ (layer0_outputs[5938]));
    assign outputs[6004] = ~((layer0_outputs[2586]) ^ (layer0_outputs[9330]));
    assign outputs[6005] = (layer0_outputs[4617]) | (layer0_outputs[5307]);
    assign outputs[6006] = ~((layer0_outputs[8635]) ^ (layer0_outputs[2370]));
    assign outputs[6007] = (layer0_outputs[778]) & ~(layer0_outputs[4621]);
    assign outputs[6008] = ~((layer0_outputs[7993]) ^ (layer0_outputs[330]));
    assign outputs[6009] = (layer0_outputs[1526]) ^ (layer0_outputs[1237]);
    assign outputs[6010] = ~((layer0_outputs[7206]) ^ (layer0_outputs[1694]));
    assign outputs[6011] = ~((layer0_outputs[2804]) ^ (layer0_outputs[1623]));
    assign outputs[6012] = layer0_outputs[6276];
    assign outputs[6013] = (layer0_outputs[4321]) | (layer0_outputs[9661]);
    assign outputs[6014] = ~((layer0_outputs[9567]) ^ (layer0_outputs[8889]));
    assign outputs[6015] = ~((layer0_outputs[5387]) ^ (layer0_outputs[1603]));
    assign outputs[6016] = layer0_outputs[6981];
    assign outputs[6017] = layer0_outputs[9156];
    assign outputs[6018] = (layer0_outputs[7400]) ^ (layer0_outputs[2740]);
    assign outputs[6019] = ~((layer0_outputs[1015]) ^ (layer0_outputs[308]));
    assign outputs[6020] = ~(layer0_outputs[5559]) | (layer0_outputs[1169]);
    assign outputs[6021] = ~((layer0_outputs[7823]) ^ (layer0_outputs[6360]));
    assign outputs[6022] = ~(layer0_outputs[8282]) | (layer0_outputs[4577]);
    assign outputs[6023] = (layer0_outputs[4646]) & ~(layer0_outputs[8761]);
    assign outputs[6024] = layer0_outputs[3987];
    assign outputs[6025] = (layer0_outputs[6112]) ^ (layer0_outputs[5922]);
    assign outputs[6026] = (layer0_outputs[3283]) ^ (layer0_outputs[1239]);
    assign outputs[6027] = layer0_outputs[1185];
    assign outputs[6028] = layer0_outputs[1236];
    assign outputs[6029] = ~(layer0_outputs[61]);
    assign outputs[6030] = ~(layer0_outputs[8004]);
    assign outputs[6031] = (layer0_outputs[1422]) | (layer0_outputs[3438]);
    assign outputs[6032] = ~((layer0_outputs[8690]) ^ (layer0_outputs[5739]));
    assign outputs[6033] = ~(layer0_outputs[10108]);
    assign outputs[6034] = ~((layer0_outputs[6211]) ^ (layer0_outputs[7902]));
    assign outputs[6035] = (layer0_outputs[5241]) | (layer0_outputs[9589]);
    assign outputs[6036] = (layer0_outputs[9910]) & (layer0_outputs[8301]);
    assign outputs[6037] = (layer0_outputs[9151]) ^ (layer0_outputs[3332]);
    assign outputs[6038] = (layer0_outputs[8836]) ^ (layer0_outputs[5091]);
    assign outputs[6039] = (layer0_outputs[2688]) ^ (layer0_outputs[4255]);
    assign outputs[6040] = ~(layer0_outputs[9448]);
    assign outputs[6041] = (layer0_outputs[6701]) & ~(layer0_outputs[4566]);
    assign outputs[6042] = (layer0_outputs[4951]) & (layer0_outputs[6985]);
    assign outputs[6043] = (layer0_outputs[2763]) ^ (layer0_outputs[4880]);
    assign outputs[6044] = layer0_outputs[1712];
    assign outputs[6045] = layer0_outputs[3055];
    assign outputs[6046] = ~(layer0_outputs[8392]) | (layer0_outputs[5732]);
    assign outputs[6047] = (layer0_outputs[4610]) & ~(layer0_outputs[1631]);
    assign outputs[6048] = ~(layer0_outputs[4811]) | (layer0_outputs[5900]);
    assign outputs[6049] = layer0_outputs[2492];
    assign outputs[6050] = layer0_outputs[8225];
    assign outputs[6051] = ~((layer0_outputs[2274]) ^ (layer0_outputs[5988]));
    assign outputs[6052] = layer0_outputs[3919];
    assign outputs[6053] = 1'b1;
    assign outputs[6054] = (layer0_outputs[8057]) | (layer0_outputs[6803]);
    assign outputs[6055] = layer0_outputs[4753];
    assign outputs[6056] = (layer0_outputs[2107]) | (layer0_outputs[395]);
    assign outputs[6057] = layer0_outputs[4404];
    assign outputs[6058] = ~((layer0_outputs[8441]) ^ (layer0_outputs[6793]));
    assign outputs[6059] = 1'b1;
    assign outputs[6060] = ~(layer0_outputs[2093]);
    assign outputs[6061] = ~(layer0_outputs[209]) | (layer0_outputs[2964]);
    assign outputs[6062] = (layer0_outputs[6882]) ^ (layer0_outputs[8482]);
    assign outputs[6063] = ~((layer0_outputs[1307]) & (layer0_outputs[3803]));
    assign outputs[6064] = ~(layer0_outputs[6749]);
    assign outputs[6065] = (layer0_outputs[8611]) ^ (layer0_outputs[5005]);
    assign outputs[6066] = ~((layer0_outputs[9722]) ^ (layer0_outputs[5039]));
    assign outputs[6067] = (layer0_outputs[4117]) & (layer0_outputs[3060]);
    assign outputs[6068] = ~(layer0_outputs[2375]);
    assign outputs[6069] = ~(layer0_outputs[1294]) | (layer0_outputs[974]);
    assign outputs[6070] = layer0_outputs[1872];
    assign outputs[6071] = ~((layer0_outputs[3975]) ^ (layer0_outputs[5445]));
    assign outputs[6072] = layer0_outputs[2058];
    assign outputs[6073] = ~(layer0_outputs[6251]);
    assign outputs[6074] = (layer0_outputs[3991]) ^ (layer0_outputs[64]);
    assign outputs[6075] = (layer0_outputs[5420]) | (layer0_outputs[6102]);
    assign outputs[6076] = (layer0_outputs[2792]) ^ (layer0_outputs[4757]);
    assign outputs[6077] = ~(layer0_outputs[610]);
    assign outputs[6078] = (layer0_outputs[3912]) ^ (layer0_outputs[2810]);
    assign outputs[6079] = layer0_outputs[9826];
    assign outputs[6080] = layer0_outputs[4682];
    assign outputs[6081] = layer0_outputs[1606];
    assign outputs[6082] = (layer0_outputs[2197]) ^ (layer0_outputs[2272]);
    assign outputs[6083] = ~((layer0_outputs[8378]) & (layer0_outputs[105]));
    assign outputs[6084] = ~(layer0_outputs[5001]);
    assign outputs[6085] = ~(layer0_outputs[3652]);
    assign outputs[6086] = (layer0_outputs[9360]) ^ (layer0_outputs[6500]);
    assign outputs[6087] = ~(layer0_outputs[6854]);
    assign outputs[6088] = ~((layer0_outputs[607]) ^ (layer0_outputs[4051]));
    assign outputs[6089] = ~(layer0_outputs[7390]);
    assign outputs[6090] = ~((layer0_outputs[221]) ^ (layer0_outputs[5718]));
    assign outputs[6091] = (layer0_outputs[3557]) & (layer0_outputs[2362]);
    assign outputs[6092] = ~(layer0_outputs[4925]);
    assign outputs[6093] = ~((layer0_outputs[2861]) ^ (layer0_outputs[3849]));
    assign outputs[6094] = ~((layer0_outputs[9966]) & (layer0_outputs[373]));
    assign outputs[6095] = layer0_outputs[9699];
    assign outputs[6096] = 1'b1;
    assign outputs[6097] = ~((layer0_outputs[1706]) & (layer0_outputs[9694]));
    assign outputs[6098] = (layer0_outputs[5315]) | (layer0_outputs[9268]);
    assign outputs[6099] = ~((layer0_outputs[6349]) | (layer0_outputs[2932]));
    assign outputs[6100] = layer0_outputs[9485];
    assign outputs[6101] = ~(layer0_outputs[5644]) | (layer0_outputs[1030]);
    assign outputs[6102] = ~(layer0_outputs[7885]) | (layer0_outputs[6986]);
    assign outputs[6103] = (layer0_outputs[7221]) ^ (layer0_outputs[773]);
    assign outputs[6104] = (layer0_outputs[2959]) ^ (layer0_outputs[2505]);
    assign outputs[6105] = ~((layer0_outputs[9232]) ^ (layer0_outputs[1586]));
    assign outputs[6106] = ~(layer0_outputs[1978]) | (layer0_outputs[3690]);
    assign outputs[6107] = layer0_outputs[9138];
    assign outputs[6108] = (layer0_outputs[2740]) ^ (layer0_outputs[8915]);
    assign outputs[6109] = ~((layer0_outputs[8424]) | (layer0_outputs[4192]));
    assign outputs[6110] = ~((layer0_outputs[660]) ^ (layer0_outputs[858]));
    assign outputs[6111] = layer0_outputs[2939];
    assign outputs[6112] = ~(layer0_outputs[8658]);
    assign outputs[6113] = (layer0_outputs[5663]) & ~(layer0_outputs[4502]);
    assign outputs[6114] = ~(layer0_outputs[960]);
    assign outputs[6115] = ~((layer0_outputs[5294]) ^ (layer0_outputs[621]));
    assign outputs[6116] = ~((layer0_outputs[3419]) ^ (layer0_outputs[8407]));
    assign outputs[6117] = ~(layer0_outputs[5664]);
    assign outputs[6118] = ~(layer0_outputs[3941]);
    assign outputs[6119] = ~(layer0_outputs[5011]);
    assign outputs[6120] = (layer0_outputs[5968]) ^ (layer0_outputs[2161]);
    assign outputs[6121] = ~(layer0_outputs[7893]);
    assign outputs[6122] = (layer0_outputs[3973]) ^ (layer0_outputs[4707]);
    assign outputs[6123] = ~((layer0_outputs[4611]) ^ (layer0_outputs[6101]));
    assign outputs[6124] = ~((layer0_outputs[7604]) ^ (layer0_outputs[8859]));
    assign outputs[6125] = ~((layer0_outputs[4190]) ^ (layer0_outputs[4322]));
    assign outputs[6126] = ~((layer0_outputs[8311]) ^ (layer0_outputs[10014]));
    assign outputs[6127] = (layer0_outputs[9532]) & ~(layer0_outputs[4188]);
    assign outputs[6128] = layer0_outputs[6142];
    assign outputs[6129] = layer0_outputs[4425];
    assign outputs[6130] = ~((layer0_outputs[9908]) | (layer0_outputs[2381]));
    assign outputs[6131] = ~(layer0_outputs[4033]) | (layer0_outputs[6546]);
    assign outputs[6132] = ~(layer0_outputs[3374]);
    assign outputs[6133] = ~(layer0_outputs[8592]);
    assign outputs[6134] = (layer0_outputs[4765]) ^ (layer0_outputs[5929]);
    assign outputs[6135] = ~(layer0_outputs[6623]);
    assign outputs[6136] = layer0_outputs[720];
    assign outputs[6137] = (layer0_outputs[8595]) | (layer0_outputs[2892]);
    assign outputs[6138] = layer0_outputs[532];
    assign outputs[6139] = (layer0_outputs[4504]) ^ (layer0_outputs[25]);
    assign outputs[6140] = ~((layer0_outputs[465]) & (layer0_outputs[537]));
    assign outputs[6141] = ~((layer0_outputs[9994]) & (layer0_outputs[1924]));
    assign outputs[6142] = layer0_outputs[6969];
    assign outputs[6143] = 1'b1;
    assign outputs[6144] = ~(layer0_outputs[5911]);
    assign outputs[6145] = (layer0_outputs[1540]) | (layer0_outputs[3221]);
    assign outputs[6146] = ~((layer0_outputs[4734]) & (layer0_outputs[1784]));
    assign outputs[6147] = (layer0_outputs[5363]) & ~(layer0_outputs[1905]);
    assign outputs[6148] = (layer0_outputs[346]) & ~(layer0_outputs[2860]);
    assign outputs[6149] = ~(layer0_outputs[1582]);
    assign outputs[6150] = ~(layer0_outputs[6151]);
    assign outputs[6151] = ~(layer0_outputs[3389]);
    assign outputs[6152] = layer0_outputs[7611];
    assign outputs[6153] = ~((layer0_outputs[1764]) | (layer0_outputs[8563]));
    assign outputs[6154] = ~(layer0_outputs[10228]);
    assign outputs[6155] = (layer0_outputs[5819]) & ~(layer0_outputs[1077]);
    assign outputs[6156] = (layer0_outputs[1745]) | (layer0_outputs[1930]);
    assign outputs[6157] = ~((layer0_outputs[10172]) ^ (layer0_outputs[6700]));
    assign outputs[6158] = ~(layer0_outputs[10166]) | (layer0_outputs[6968]);
    assign outputs[6159] = ~(layer0_outputs[2411]);
    assign outputs[6160] = ~((layer0_outputs[1100]) ^ (layer0_outputs[7209]));
    assign outputs[6161] = layer0_outputs[10155];
    assign outputs[6162] = ~(layer0_outputs[8952]) | (layer0_outputs[7595]);
    assign outputs[6163] = (layer0_outputs[3372]) ^ (layer0_outputs[925]);
    assign outputs[6164] = ~((layer0_outputs[9532]) ^ (layer0_outputs[4319]));
    assign outputs[6165] = ~((layer0_outputs[162]) ^ (layer0_outputs[6977]));
    assign outputs[6166] = ~((layer0_outputs[4793]) ^ (layer0_outputs[4966]));
    assign outputs[6167] = layer0_outputs[10061];
    assign outputs[6168] = layer0_outputs[10075];
    assign outputs[6169] = ~(layer0_outputs[817]);
    assign outputs[6170] = ~(layer0_outputs[3443]);
    assign outputs[6171] = layer0_outputs[4299];
    assign outputs[6172] = (layer0_outputs[4466]) ^ (layer0_outputs[4759]);
    assign outputs[6173] = (layer0_outputs[4479]) ^ (layer0_outputs[1992]);
    assign outputs[6174] = ~((layer0_outputs[7756]) ^ (layer0_outputs[3274]));
    assign outputs[6175] = layer0_outputs[7610];
    assign outputs[6176] = (layer0_outputs[6623]) & ~(layer0_outputs[10121]);
    assign outputs[6177] = ~((layer0_outputs[81]) & (layer0_outputs[7428]));
    assign outputs[6178] = ~(layer0_outputs[1198]);
    assign outputs[6179] = ~(layer0_outputs[484]);
    assign outputs[6180] = (layer0_outputs[4097]) ^ (layer0_outputs[7770]);
    assign outputs[6181] = ~(layer0_outputs[122]);
    assign outputs[6182] = layer0_outputs[7040];
    assign outputs[6183] = ~(layer0_outputs[4674]);
    assign outputs[6184] = (layer0_outputs[7247]) & ~(layer0_outputs[1642]);
    assign outputs[6185] = layer0_outputs[9238];
    assign outputs[6186] = layer0_outputs[1820];
    assign outputs[6187] = ~((layer0_outputs[2433]) ^ (layer0_outputs[9398]));
    assign outputs[6188] = ~((layer0_outputs[2172]) ^ (layer0_outputs[3725]));
    assign outputs[6189] = ~((layer0_outputs[4526]) ^ (layer0_outputs[2550]));
    assign outputs[6190] = ~(layer0_outputs[9064]) | (layer0_outputs[4362]);
    assign outputs[6191] = ~((layer0_outputs[3018]) | (layer0_outputs[7119]));
    assign outputs[6192] = (layer0_outputs[1539]) & ~(layer0_outputs[9692]);
    assign outputs[6193] = (layer0_outputs[8754]) & ~(layer0_outputs[1335]);
    assign outputs[6194] = layer0_outputs[8801];
    assign outputs[6195] = ~(layer0_outputs[4904]);
    assign outputs[6196] = (layer0_outputs[1611]) ^ (layer0_outputs[5943]);
    assign outputs[6197] = (layer0_outputs[3616]) & ~(layer0_outputs[3089]);
    assign outputs[6198] = ~(layer0_outputs[9751]) | (layer0_outputs[6014]);
    assign outputs[6199] = layer0_outputs[8099];
    assign outputs[6200] = ~((layer0_outputs[5328]) & (layer0_outputs[2675]));
    assign outputs[6201] = ~((layer0_outputs[5975]) | (layer0_outputs[5582]));
    assign outputs[6202] = ~(layer0_outputs[8708]);
    assign outputs[6203] = ~((layer0_outputs[7230]) & (layer0_outputs[3752]));
    assign outputs[6204] = ~(layer0_outputs[8822]);
    assign outputs[6205] = layer0_outputs[6421];
    assign outputs[6206] = (layer0_outputs[1392]) & (layer0_outputs[8094]);
    assign outputs[6207] = layer0_outputs[2198];
    assign outputs[6208] = ~(layer0_outputs[2404]) | (layer0_outputs[23]);
    assign outputs[6209] = (layer0_outputs[48]) ^ (layer0_outputs[1223]);
    assign outputs[6210] = (layer0_outputs[272]) | (layer0_outputs[9395]);
    assign outputs[6211] = ~(layer0_outputs[2159]) | (layer0_outputs[5965]);
    assign outputs[6212] = (layer0_outputs[951]) | (layer0_outputs[9603]);
    assign outputs[6213] = (layer0_outputs[8322]) ^ (layer0_outputs[4946]);
    assign outputs[6214] = ~((layer0_outputs[5992]) ^ (layer0_outputs[2132]));
    assign outputs[6215] = (layer0_outputs[4767]) & ~(layer0_outputs[2765]);
    assign outputs[6216] = ~((layer0_outputs[6254]) ^ (layer0_outputs[441]));
    assign outputs[6217] = (layer0_outputs[4489]) & ~(layer0_outputs[6591]);
    assign outputs[6218] = ~((layer0_outputs[4944]) ^ (layer0_outputs[1751]));
    assign outputs[6219] = ~(layer0_outputs[5599]);
    assign outputs[6220] = ~(layer0_outputs[6033]);
    assign outputs[6221] = ~((layer0_outputs[3541]) ^ (layer0_outputs[9487]));
    assign outputs[6222] = (layer0_outputs[7375]) ^ (layer0_outputs[5891]);
    assign outputs[6223] = layer0_outputs[2788];
    assign outputs[6224] = layer0_outputs[9208];
    assign outputs[6225] = ~(layer0_outputs[5008]);
    assign outputs[6226] = (layer0_outputs[4251]) ^ (layer0_outputs[1196]);
    assign outputs[6227] = ~((layer0_outputs[1416]) ^ (layer0_outputs[4981]));
    assign outputs[6228] = (layer0_outputs[7370]) ^ (layer0_outputs[8031]);
    assign outputs[6229] = ~(layer0_outputs[8799]) | (layer0_outputs[5174]);
    assign outputs[6230] = ~(layer0_outputs[9993]);
    assign outputs[6231] = ~((layer0_outputs[1852]) | (layer0_outputs[1906]));
    assign outputs[6232] = (layer0_outputs[5968]) & ~(layer0_outputs[900]);
    assign outputs[6233] = ~((layer0_outputs[92]) | (layer0_outputs[8760]));
    assign outputs[6234] = (layer0_outputs[1131]) | (layer0_outputs[7485]);
    assign outputs[6235] = ~((layer0_outputs[4348]) & (layer0_outputs[2873]));
    assign outputs[6236] = ~(layer0_outputs[9167]);
    assign outputs[6237] = (layer0_outputs[9580]) & (layer0_outputs[2834]);
    assign outputs[6238] = (layer0_outputs[1920]) | (layer0_outputs[9763]);
    assign outputs[6239] = (layer0_outputs[1323]) ^ (layer0_outputs[6729]);
    assign outputs[6240] = ~((layer0_outputs[1810]) | (layer0_outputs[580]));
    assign outputs[6241] = (layer0_outputs[2330]) ^ (layer0_outputs[1283]);
    assign outputs[6242] = ~(layer0_outputs[134]);
    assign outputs[6243] = (layer0_outputs[4803]) ^ (layer0_outputs[5834]);
    assign outputs[6244] = ~((layer0_outputs[1183]) ^ (layer0_outputs[10041]));
    assign outputs[6245] = layer0_outputs[6668];
    assign outputs[6246] = ~(layer0_outputs[4855]);
    assign outputs[6247] = ~(layer0_outputs[239]);
    assign outputs[6248] = ~((layer0_outputs[7242]) ^ (layer0_outputs[4655]));
    assign outputs[6249] = ~(layer0_outputs[5342]);
    assign outputs[6250] = (layer0_outputs[9986]) & (layer0_outputs[3231]);
    assign outputs[6251] = ~((layer0_outputs[6707]) & (layer0_outputs[2689]));
    assign outputs[6252] = (layer0_outputs[5050]) & ~(layer0_outputs[634]);
    assign outputs[6253] = ~(layer0_outputs[2397]);
    assign outputs[6254] = ~((layer0_outputs[9422]) ^ (layer0_outputs[10036]));
    assign outputs[6255] = ~((layer0_outputs[4440]) | (layer0_outputs[7686]));
    assign outputs[6256] = ~((layer0_outputs[9662]) & (layer0_outputs[403]));
    assign outputs[6257] = (layer0_outputs[5255]) ^ (layer0_outputs[5682]);
    assign outputs[6258] = ~(layer0_outputs[1732]);
    assign outputs[6259] = ~(layer0_outputs[10072]);
    assign outputs[6260] = ~((layer0_outputs[8437]) ^ (layer0_outputs[2266]));
    assign outputs[6261] = layer0_outputs[1718];
    assign outputs[6262] = layer0_outputs[8781];
    assign outputs[6263] = ~(layer0_outputs[6577]);
    assign outputs[6264] = (layer0_outputs[5094]) ^ (layer0_outputs[1047]);
    assign outputs[6265] = (layer0_outputs[2210]) & ~(layer0_outputs[8312]);
    assign outputs[6266] = layer0_outputs[1933];
    assign outputs[6267] = layer0_outputs[4632];
    assign outputs[6268] = ~(layer0_outputs[229]) | (layer0_outputs[5752]);
    assign outputs[6269] = ~((layer0_outputs[3049]) ^ (layer0_outputs[1960]));
    assign outputs[6270] = (layer0_outputs[7851]) & (layer0_outputs[1343]);
    assign outputs[6271] = (layer0_outputs[4183]) & ~(layer0_outputs[1022]);
    assign outputs[6272] = ~(layer0_outputs[2576]) | (layer0_outputs[2537]);
    assign outputs[6273] = ~((layer0_outputs[6761]) ^ (layer0_outputs[7710]));
    assign outputs[6274] = (layer0_outputs[5669]) ^ (layer0_outputs[8623]);
    assign outputs[6275] = layer0_outputs[2102];
    assign outputs[6276] = (layer0_outputs[6571]) ^ (layer0_outputs[358]);
    assign outputs[6277] = layer0_outputs[6397];
    assign outputs[6278] = ~(layer0_outputs[3220]);
    assign outputs[6279] = (layer0_outputs[9607]) & (layer0_outputs[3754]);
    assign outputs[6280] = ~(layer0_outputs[7726]);
    assign outputs[6281] = ~(layer0_outputs[1549]);
    assign outputs[6282] = ~((layer0_outputs[845]) ^ (layer0_outputs[5854]));
    assign outputs[6283] = ~(layer0_outputs[2252]) | (layer0_outputs[2037]);
    assign outputs[6284] = ~(layer0_outputs[2471]);
    assign outputs[6285] = layer0_outputs[568];
    assign outputs[6286] = ~(layer0_outputs[7751]);
    assign outputs[6287] = ~(layer0_outputs[4914]);
    assign outputs[6288] = (layer0_outputs[8983]) & (layer0_outputs[5571]);
    assign outputs[6289] = (layer0_outputs[1413]) ^ (layer0_outputs[4691]);
    assign outputs[6290] = (layer0_outputs[3009]) ^ (layer0_outputs[1150]);
    assign outputs[6291] = (layer0_outputs[2044]) & ~(layer0_outputs[5717]);
    assign outputs[6292] = ~(layer0_outputs[5035]) | (layer0_outputs[1197]);
    assign outputs[6293] = ~(layer0_outputs[3612]);
    assign outputs[6294] = (layer0_outputs[1207]) ^ (layer0_outputs[10032]);
    assign outputs[6295] = ~(layer0_outputs[7032]);
    assign outputs[6296] = ~((layer0_outputs[959]) | (layer0_outputs[426]));
    assign outputs[6297] = (layer0_outputs[6776]) & ~(layer0_outputs[8780]);
    assign outputs[6298] = layer0_outputs[3549];
    assign outputs[6299] = (layer0_outputs[9427]) ^ (layer0_outputs[3366]);
    assign outputs[6300] = layer0_outputs[9636];
    assign outputs[6301] = (layer0_outputs[4095]) & ~(layer0_outputs[7179]);
    assign outputs[6302] = (layer0_outputs[4760]) & ~(layer0_outputs[322]);
    assign outputs[6303] = (layer0_outputs[8940]) ^ (layer0_outputs[10238]);
    assign outputs[6304] = (layer0_outputs[6838]) ^ (layer0_outputs[882]);
    assign outputs[6305] = ~((layer0_outputs[1956]) ^ (layer0_outputs[2766]));
    assign outputs[6306] = (layer0_outputs[2108]) ^ (layer0_outputs[2]);
    assign outputs[6307] = (layer0_outputs[8294]) & ~(layer0_outputs[7425]);
    assign outputs[6308] = (layer0_outputs[5122]) ^ (layer0_outputs[10215]);
    assign outputs[6309] = (layer0_outputs[5702]) ^ (layer0_outputs[442]);
    assign outputs[6310] = (layer0_outputs[9937]) ^ (layer0_outputs[8516]);
    assign outputs[6311] = ~((layer0_outputs[5065]) ^ (layer0_outputs[5536]));
    assign outputs[6312] = layer0_outputs[23];
    assign outputs[6313] = ~((layer0_outputs[420]) & (layer0_outputs[1402]));
    assign outputs[6314] = layer0_outputs[6670];
    assign outputs[6315] = ~((layer0_outputs[3062]) ^ (layer0_outputs[2108]));
    assign outputs[6316] = 1'b1;
    assign outputs[6317] = ~(layer0_outputs[7091]);
    assign outputs[6318] = layer0_outputs[4327];
    assign outputs[6319] = (layer0_outputs[2205]) & (layer0_outputs[2193]);
    assign outputs[6320] = ~((layer0_outputs[6084]) | (layer0_outputs[3567]));
    assign outputs[6321] = (layer0_outputs[7832]) & (layer0_outputs[9296]);
    assign outputs[6322] = (layer0_outputs[3613]) ^ (layer0_outputs[723]);
    assign outputs[6323] = layer0_outputs[8681];
    assign outputs[6324] = ~(layer0_outputs[2175]);
    assign outputs[6325] = (layer0_outputs[2640]) ^ (layer0_outputs[2583]);
    assign outputs[6326] = ~((layer0_outputs[4267]) & (layer0_outputs[5600]));
    assign outputs[6327] = layer0_outputs[3490];
    assign outputs[6328] = (layer0_outputs[9266]) | (layer0_outputs[1399]);
    assign outputs[6329] = (layer0_outputs[4356]) & ~(layer0_outputs[6041]);
    assign outputs[6330] = layer0_outputs[7633];
    assign outputs[6331] = ~(layer0_outputs[6962]);
    assign outputs[6332] = layer0_outputs[1647];
    assign outputs[6333] = ~(layer0_outputs[7579]);
    assign outputs[6334] = ~(layer0_outputs[6319]);
    assign outputs[6335] = ~((layer0_outputs[8190]) ^ (layer0_outputs[28]));
    assign outputs[6336] = (layer0_outputs[7214]) ^ (layer0_outputs[5609]);
    assign outputs[6337] = ~((layer0_outputs[989]) ^ (layer0_outputs[1395]));
    assign outputs[6338] = layer0_outputs[2905];
    assign outputs[6339] = layer0_outputs[4412];
    assign outputs[6340] = (layer0_outputs[8369]) & (layer0_outputs[5257]);
    assign outputs[6341] = ~((layer0_outputs[4703]) ^ (layer0_outputs[1675]));
    assign outputs[6342] = layer0_outputs[2439];
    assign outputs[6343] = ~(layer0_outputs[7490]);
    assign outputs[6344] = (layer0_outputs[6067]) ^ (layer0_outputs[6956]);
    assign outputs[6345] = layer0_outputs[8066];
    assign outputs[6346] = ~(layer0_outputs[5278]);
    assign outputs[6347] = (layer0_outputs[1812]) ^ (layer0_outputs[8810]);
    assign outputs[6348] = ~((layer0_outputs[3708]) ^ (layer0_outputs[8023]));
    assign outputs[6349] = (layer0_outputs[7311]) & ~(layer0_outputs[9551]);
    assign outputs[6350] = ~(layer0_outputs[1972]);
    assign outputs[6351] = 1'b0;
    assign outputs[6352] = layer0_outputs[1699];
    assign outputs[6353] = ~(layer0_outputs[4790]);
    assign outputs[6354] = ~((layer0_outputs[5321]) ^ (layer0_outputs[3514]));
    assign outputs[6355] = ~(layer0_outputs[6492]) | (layer0_outputs[6813]);
    assign outputs[6356] = ~((layer0_outputs[5077]) & (layer0_outputs[1813]));
    assign outputs[6357] = layer0_outputs[9585];
    assign outputs[6358] = (layer0_outputs[1859]) & (layer0_outputs[9288]);
    assign outputs[6359] = layer0_outputs[3466];
    assign outputs[6360] = layer0_outputs[9162];
    assign outputs[6361] = (layer0_outputs[8163]) & ~(layer0_outputs[5038]);
    assign outputs[6362] = ~(layer0_outputs[9924]);
    assign outputs[6363] = (layer0_outputs[6326]) & ~(layer0_outputs[7487]);
    assign outputs[6364] = (layer0_outputs[3715]) | (layer0_outputs[4521]);
    assign outputs[6365] = (layer0_outputs[8174]) ^ (layer0_outputs[2400]);
    assign outputs[6366] = ~(layer0_outputs[442]) | (layer0_outputs[667]);
    assign outputs[6367] = (layer0_outputs[5355]) ^ (layer0_outputs[9349]);
    assign outputs[6368] = (layer0_outputs[339]) ^ (layer0_outputs[7868]);
    assign outputs[6369] = ~(layer0_outputs[2579]) | (layer0_outputs[6918]);
    assign outputs[6370] = (layer0_outputs[2925]) ^ (layer0_outputs[6701]);
    assign outputs[6371] = (layer0_outputs[1318]) & ~(layer0_outputs[1985]);
    assign outputs[6372] = layer0_outputs[5245];
    assign outputs[6373] = layer0_outputs[4363];
    assign outputs[6374] = ~(layer0_outputs[4795]);
    assign outputs[6375] = ~(layer0_outputs[8845]);
    assign outputs[6376] = ~((layer0_outputs[868]) | (layer0_outputs[743]));
    assign outputs[6377] = ~(layer0_outputs[7008]);
    assign outputs[6378] = ~(layer0_outputs[9558]);
    assign outputs[6379] = (layer0_outputs[3287]) ^ (layer0_outputs[6720]);
    assign outputs[6380] = ~((layer0_outputs[1563]) | (layer0_outputs[6414]));
    assign outputs[6381] = ~(layer0_outputs[6785]);
    assign outputs[6382] = (layer0_outputs[8793]) ^ (layer0_outputs[7042]);
    assign outputs[6383] = (layer0_outputs[9376]) & ~(layer0_outputs[1625]);
    assign outputs[6384] = ~(layer0_outputs[7597]);
    assign outputs[6385] = layer0_outputs[7368];
    assign outputs[6386] = ~((layer0_outputs[8851]) ^ (layer0_outputs[2237]));
    assign outputs[6387] = ~((layer0_outputs[107]) ^ (layer0_outputs[2432]));
    assign outputs[6388] = ~((layer0_outputs[749]) | (layer0_outputs[8330]));
    assign outputs[6389] = (layer0_outputs[6198]) & (layer0_outputs[2343]);
    assign outputs[6390] = ~(layer0_outputs[9987]);
    assign outputs[6391] = ~(layer0_outputs[7106]);
    assign outputs[6392] = ~(layer0_outputs[5585]);
    assign outputs[6393] = ~((layer0_outputs[1217]) ^ (layer0_outputs[3422]));
    assign outputs[6394] = layer0_outputs[8755];
    assign outputs[6395] = layer0_outputs[9320];
    assign outputs[6396] = (layer0_outputs[4271]) & (layer0_outputs[6891]);
    assign outputs[6397] = ~((layer0_outputs[8447]) ^ (layer0_outputs[3210]));
    assign outputs[6398] = layer0_outputs[6281];
    assign outputs[6399] = ~(layer0_outputs[4397]);
    assign outputs[6400] = ~(layer0_outputs[4409]);
    assign outputs[6401] = ~(layer0_outputs[6356]);
    assign outputs[6402] = (layer0_outputs[8261]) & ~(layer0_outputs[7749]);
    assign outputs[6403] = ~((layer0_outputs[8162]) | (layer0_outputs[4588]));
    assign outputs[6404] = ~((layer0_outputs[693]) | (layer0_outputs[4314]));
    assign outputs[6405] = layer0_outputs[244];
    assign outputs[6406] = ~((layer0_outputs[7568]) | (layer0_outputs[8714]));
    assign outputs[6407] = ~(layer0_outputs[3421]);
    assign outputs[6408] = (layer0_outputs[1366]) ^ (layer0_outputs[1452]);
    assign outputs[6409] = (layer0_outputs[1140]) & ~(layer0_outputs[10140]);
    assign outputs[6410] = ~((layer0_outputs[5369]) ^ (layer0_outputs[1738]));
    assign outputs[6411] = layer0_outputs[1783];
    assign outputs[6412] = ~(layer0_outputs[9812]);
    assign outputs[6413] = (layer0_outputs[147]) ^ (layer0_outputs[1138]);
    assign outputs[6414] = (layer0_outputs[8947]) & ~(layer0_outputs[1872]);
    assign outputs[6415] = ~(layer0_outputs[2154]) | (layer0_outputs[2910]);
    assign outputs[6416] = ~(layer0_outputs[2114]);
    assign outputs[6417] = ~(layer0_outputs[587]);
    assign outputs[6418] = layer0_outputs[1522];
    assign outputs[6419] = ~((layer0_outputs[10180]) & (layer0_outputs[6239]));
    assign outputs[6420] = ~(layer0_outputs[4669]);
    assign outputs[6421] = ~((layer0_outputs[4755]) ^ (layer0_outputs[5491]));
    assign outputs[6422] = (layer0_outputs[6204]) & ~(layer0_outputs[3497]);
    assign outputs[6423] = ~(layer0_outputs[9970]) | (layer0_outputs[5928]);
    assign outputs[6424] = ~(layer0_outputs[7190]);
    assign outputs[6425] = ~(layer0_outputs[2228]);
    assign outputs[6426] = 1'b0;
    assign outputs[6427] = (layer0_outputs[3328]) | (layer0_outputs[5591]);
    assign outputs[6428] = ~(layer0_outputs[2986]);
    assign outputs[6429] = ~(layer0_outputs[581]);
    assign outputs[6430] = (layer0_outputs[7622]) ^ (layer0_outputs[9705]);
    assign outputs[6431] = ~(layer0_outputs[2475]);
    assign outputs[6432] = layer0_outputs[9070];
    assign outputs[6433] = (layer0_outputs[707]) | (layer0_outputs[5286]);
    assign outputs[6434] = ~(layer0_outputs[9520]);
    assign outputs[6435] = (layer0_outputs[945]) | (layer0_outputs[2876]);
    assign outputs[6436] = ~(layer0_outputs[794]);
    assign outputs[6437] = (layer0_outputs[95]) & ~(layer0_outputs[4535]);
    assign outputs[6438] = ~((layer0_outputs[7565]) ^ (layer0_outputs[4369]));
    assign outputs[6439] = layer0_outputs[8833];
    assign outputs[6440] = ~(layer0_outputs[1987]);
    assign outputs[6441] = ~(layer0_outputs[6597]) | (layer0_outputs[50]);
    assign outputs[6442] = layer0_outputs[8421];
    assign outputs[6443] = ~((layer0_outputs[1152]) | (layer0_outputs[9802]));
    assign outputs[6444] = (layer0_outputs[293]) | (layer0_outputs[10168]);
    assign outputs[6445] = (layer0_outputs[3090]) & ~(layer0_outputs[7017]);
    assign outputs[6446] = (layer0_outputs[654]) & ~(layer0_outputs[3472]);
    assign outputs[6447] = (layer0_outputs[4859]) & ~(layer0_outputs[9285]);
    assign outputs[6448] = (layer0_outputs[3672]) & ~(layer0_outputs[6536]);
    assign outputs[6449] = (layer0_outputs[10089]) & ~(layer0_outputs[6236]);
    assign outputs[6450] = (layer0_outputs[6201]) & ~(layer0_outputs[776]);
    assign outputs[6451] = ~((layer0_outputs[7063]) ^ (layer0_outputs[185]));
    assign outputs[6452] = (layer0_outputs[8015]) ^ (layer0_outputs[3551]);
    assign outputs[6453] = (layer0_outputs[1251]) | (layer0_outputs[1634]);
    assign outputs[6454] = (layer0_outputs[4434]) & ~(layer0_outputs[4156]);
    assign outputs[6455] = (layer0_outputs[618]) & ~(layer0_outputs[3594]);
    assign outputs[6456] = layer0_outputs[1484];
    assign outputs[6457] = ~((layer0_outputs[7604]) ^ (layer0_outputs[5451]));
    assign outputs[6458] = ~((layer0_outputs[7459]) & (layer0_outputs[3219]));
    assign outputs[6459] = ~((layer0_outputs[7820]) | (layer0_outputs[9460]));
    assign outputs[6460] = layer0_outputs[6131];
    assign outputs[6461] = (layer0_outputs[2897]) & (layer0_outputs[4750]);
    assign outputs[6462] = ~((layer0_outputs[9719]) ^ (layer0_outputs[4667]));
    assign outputs[6463] = ~((layer0_outputs[405]) ^ (layer0_outputs[8434]));
    assign outputs[6464] = layer0_outputs[9445];
    assign outputs[6465] = ~(layer0_outputs[3348]) | (layer0_outputs[6133]);
    assign outputs[6466] = (layer0_outputs[2292]) & ~(layer0_outputs[10216]);
    assign outputs[6467] = layer0_outputs[7476];
    assign outputs[6468] = ~(layer0_outputs[4270]);
    assign outputs[6469] = (layer0_outputs[4425]) ^ (layer0_outputs[986]);
    assign outputs[6470] = ~(layer0_outputs[8777]);
    assign outputs[6471] = ~(layer0_outputs[8374]);
    assign outputs[6472] = ~(layer0_outputs[7098]);
    assign outputs[6473] = (layer0_outputs[5168]) ^ (layer0_outputs[8719]);
    assign outputs[6474] = layer0_outputs[1769];
    assign outputs[6475] = ~(layer0_outputs[5115]);
    assign outputs[6476] = layer0_outputs[7381];
    assign outputs[6477] = layer0_outputs[6259];
    assign outputs[6478] = layer0_outputs[6602];
    assign outputs[6479] = (layer0_outputs[3462]) & ~(layer0_outputs[3275]);
    assign outputs[6480] = ~((layer0_outputs[9377]) ^ (layer0_outputs[4909]));
    assign outputs[6481] = layer0_outputs[253];
    assign outputs[6482] = ~((layer0_outputs[7106]) | (layer0_outputs[4783]));
    assign outputs[6483] = ~(layer0_outputs[7058]);
    assign outputs[6484] = layer0_outputs[5170];
    assign outputs[6485] = (layer0_outputs[7783]) ^ (layer0_outputs[6382]);
    assign outputs[6486] = ~(layer0_outputs[7488]);
    assign outputs[6487] = (layer0_outputs[7446]) & (layer0_outputs[3984]);
    assign outputs[6488] = ~(layer0_outputs[6385]);
    assign outputs[6489] = ~(layer0_outputs[4149]);
    assign outputs[6490] = ~(layer0_outputs[1576]);
    assign outputs[6491] = (layer0_outputs[8525]) & ~(layer0_outputs[5865]);
    assign outputs[6492] = ~(layer0_outputs[7714]);
    assign outputs[6493] = ~((layer0_outputs[823]) ^ (layer0_outputs[5679]));
    assign outputs[6494] = ~(layer0_outputs[1593]);
    assign outputs[6495] = ~(layer0_outputs[3128]) | (layer0_outputs[3329]);
    assign outputs[6496] = (layer0_outputs[3809]) & ~(layer0_outputs[3165]);
    assign outputs[6497] = layer0_outputs[968];
    assign outputs[6498] = (layer0_outputs[2455]) ^ (layer0_outputs[9676]);
    assign outputs[6499] = (layer0_outputs[7989]) ^ (layer0_outputs[5130]);
    assign outputs[6500] = layer0_outputs[8918];
    assign outputs[6501] = (layer0_outputs[2994]) ^ (layer0_outputs[4846]);
    assign outputs[6502] = (layer0_outputs[5969]) & ~(layer0_outputs[8646]);
    assign outputs[6503] = ~(layer0_outputs[4693]);
    assign outputs[6504] = layer0_outputs[2105];
    assign outputs[6505] = layer0_outputs[5570];
    assign outputs[6506] = layer0_outputs[8189];
    assign outputs[6507] = (layer0_outputs[880]) ^ (layer0_outputs[1090]);
    assign outputs[6508] = (layer0_outputs[903]) ^ (layer0_outputs[2324]);
    assign outputs[6509] = ~(layer0_outputs[2428]);
    assign outputs[6510] = layer0_outputs[8287];
    assign outputs[6511] = 1'b0;
    assign outputs[6512] = ~(layer0_outputs[9910]) | (layer0_outputs[9509]);
    assign outputs[6513] = layer0_outputs[601];
    assign outputs[6514] = (layer0_outputs[9279]) ^ (layer0_outputs[3161]);
    assign outputs[6515] = layer0_outputs[10210];
    assign outputs[6516] = layer0_outputs[3723];
    assign outputs[6517] = ~(layer0_outputs[9350]);
    assign outputs[6518] = ~(layer0_outputs[6648]);
    assign outputs[6519] = ~((layer0_outputs[6950]) & (layer0_outputs[7284]));
    assign outputs[6520] = layer0_outputs[2982];
    assign outputs[6521] = ~(layer0_outputs[3673]);
    assign outputs[6522] = (layer0_outputs[6938]) & ~(layer0_outputs[5088]);
    assign outputs[6523] = (layer0_outputs[1689]) & (layer0_outputs[4702]);
    assign outputs[6524] = layer0_outputs[2635];
    assign outputs[6525] = ~((layer0_outputs[3675]) ^ (layer0_outputs[4789]));
    assign outputs[6526] = layer0_outputs[7760];
    assign outputs[6527] = ~((layer0_outputs[8266]) | (layer0_outputs[295]));
    assign outputs[6528] = layer0_outputs[5350];
    assign outputs[6529] = ~((layer0_outputs[10222]) ^ (layer0_outputs[5598]));
    assign outputs[6530] = ~((layer0_outputs[3601]) & (layer0_outputs[4723]));
    assign outputs[6531] = layer0_outputs[95];
    assign outputs[6532] = (layer0_outputs[4051]) & ~(layer0_outputs[8753]);
    assign outputs[6533] = layer0_outputs[9596];
    assign outputs[6534] = ~(layer0_outputs[5089]);
    assign outputs[6535] = ~(layer0_outputs[16]);
    assign outputs[6536] = (layer0_outputs[5912]) ^ (layer0_outputs[7670]);
    assign outputs[6537] = ~(layer0_outputs[5237]) | (layer0_outputs[447]);
    assign outputs[6538] = (layer0_outputs[3741]) ^ (layer0_outputs[5412]);
    assign outputs[6539] = ~(layer0_outputs[10098]) | (layer0_outputs[5525]);
    assign outputs[6540] = (layer0_outputs[8003]) & ~(layer0_outputs[1608]);
    assign outputs[6541] = layer0_outputs[8278];
    assign outputs[6542] = ~((layer0_outputs[9799]) ^ (layer0_outputs[2075]));
    assign outputs[6543] = ~(layer0_outputs[5139]);
    assign outputs[6544] = ~((layer0_outputs[8860]) ^ (layer0_outputs[889]));
    assign outputs[6545] = ~((layer0_outputs[7471]) & (layer0_outputs[8161]));
    assign outputs[6546] = ~((layer0_outputs[1915]) ^ (layer0_outputs[4550]));
    assign outputs[6547] = layer0_outputs[5602];
    assign outputs[6548] = layer0_outputs[300];
    assign outputs[6549] = layer0_outputs[6491];
    assign outputs[6550] = layer0_outputs[1050];
    assign outputs[6551] = (layer0_outputs[4781]) & (layer0_outputs[3886]);
    assign outputs[6552] = (layer0_outputs[5760]) & (layer0_outputs[8536]);
    assign outputs[6553] = (layer0_outputs[8838]) & (layer0_outputs[9318]);
    assign outputs[6554] = ~(layer0_outputs[1367]);
    assign outputs[6555] = ~(layer0_outputs[5342]);
    assign outputs[6556] = layer0_outputs[8520];
    assign outputs[6557] = ~((layer0_outputs[5883]) ^ (layer0_outputs[6122]));
    assign outputs[6558] = (layer0_outputs[2509]) & ~(layer0_outputs[8655]);
    assign outputs[6559] = (layer0_outputs[6885]) ^ (layer0_outputs[7772]);
    assign outputs[6560] = layer0_outputs[5850];
    assign outputs[6561] = layer0_outputs[166];
    assign outputs[6562] = ~((layer0_outputs[4729]) ^ (layer0_outputs[5384]));
    assign outputs[6563] = ~((layer0_outputs[9094]) & (layer0_outputs[5127]));
    assign outputs[6564] = ~(layer0_outputs[7239]) | (layer0_outputs[8175]);
    assign outputs[6565] = ~((layer0_outputs[7227]) ^ (layer0_outputs[2188]));
    assign outputs[6566] = ~(layer0_outputs[3043]);
    assign outputs[6567] = layer0_outputs[1323];
    assign outputs[6568] = (layer0_outputs[7062]) & ~(layer0_outputs[9840]);
    assign outputs[6569] = (layer0_outputs[6375]) & ~(layer0_outputs[4754]);
    assign outputs[6570] = (layer0_outputs[7814]) ^ (layer0_outputs[2774]);
    assign outputs[6571] = ~(layer0_outputs[8300]) | (layer0_outputs[9731]);
    assign outputs[6572] = layer0_outputs[3821];
    assign outputs[6573] = ~((layer0_outputs[2866]) | (layer0_outputs[2301]));
    assign outputs[6574] = ~(layer0_outputs[3702]);
    assign outputs[6575] = layer0_outputs[4329];
    assign outputs[6576] = ~(layer0_outputs[6028]);
    assign outputs[6577] = (layer0_outputs[7589]) ^ (layer0_outputs[853]);
    assign outputs[6578] = (layer0_outputs[9330]) & ~(layer0_outputs[7274]);
    assign outputs[6579] = layer0_outputs[8111];
    assign outputs[6580] = ~(layer0_outputs[623]);
    assign outputs[6581] = (layer0_outputs[1489]) & ~(layer0_outputs[7372]);
    assign outputs[6582] = ~(layer0_outputs[6865]) | (layer0_outputs[8288]);
    assign outputs[6583] = (layer0_outputs[121]) ^ (layer0_outputs[4555]);
    assign outputs[6584] = layer0_outputs[6029];
    assign outputs[6585] = ~(layer0_outputs[5994]);
    assign outputs[6586] = ~(layer0_outputs[6493]);
    assign outputs[6587] = ~((layer0_outputs[1128]) ^ (layer0_outputs[8493]));
    assign outputs[6588] = layer0_outputs[4802];
    assign outputs[6589] = ~(layer0_outputs[1468]) | (layer0_outputs[6290]);
    assign outputs[6590] = ~((layer0_outputs[2960]) ^ (layer0_outputs[7722]));
    assign outputs[6591] = (layer0_outputs[2997]) & ~(layer0_outputs[6871]);
    assign outputs[6592] = ~((layer0_outputs[1792]) | (layer0_outputs[3019]));
    assign outputs[6593] = (layer0_outputs[6919]) & (layer0_outputs[1457]);
    assign outputs[6594] = (layer0_outputs[3293]) & ~(layer0_outputs[5459]);
    assign outputs[6595] = ~(layer0_outputs[767]);
    assign outputs[6596] = ~((layer0_outputs[3892]) & (layer0_outputs[9125]));
    assign outputs[6597] = ~((layer0_outputs[3629]) | (layer0_outputs[7122]));
    assign outputs[6598] = (layer0_outputs[7555]) & ~(layer0_outputs[9799]);
    assign outputs[6599] = (layer0_outputs[784]) ^ (layer0_outputs[3159]);
    assign outputs[6600] = layer0_outputs[7781];
    assign outputs[6601] = layer0_outputs[5984];
    assign outputs[6602] = ~(layer0_outputs[6195]);
    assign outputs[6603] = ~((layer0_outputs[2262]) ^ (layer0_outputs[385]));
    assign outputs[6604] = ~((layer0_outputs[8662]) ^ (layer0_outputs[978]));
    assign outputs[6605] = (layer0_outputs[3986]) & ~(layer0_outputs[4913]);
    assign outputs[6606] = layer0_outputs[8181];
    assign outputs[6607] = ~((layer0_outputs[6865]) ^ (layer0_outputs[1173]));
    assign outputs[6608] = (layer0_outputs[948]) & ~(layer0_outputs[10182]);
    assign outputs[6609] = ~((layer0_outputs[1046]) & (layer0_outputs[6980]));
    assign outputs[6610] = (layer0_outputs[1903]) & (layer0_outputs[2238]);
    assign outputs[6611] = ~((layer0_outputs[9183]) ^ (layer0_outputs[7975]));
    assign outputs[6612] = ~((layer0_outputs[6773]) & (layer0_outputs[1011]));
    assign outputs[6613] = (layer0_outputs[1339]) & ~(layer0_outputs[2166]);
    assign outputs[6614] = (layer0_outputs[7552]) ^ (layer0_outputs[6023]);
    assign outputs[6615] = ~((layer0_outputs[5370]) ^ (layer0_outputs[8756]));
    assign outputs[6616] = layer0_outputs[9739];
    assign outputs[6617] = layer0_outputs[7282];
    assign outputs[6618] = layer0_outputs[1353];
    assign outputs[6619] = ~((layer0_outputs[3184]) ^ (layer0_outputs[5913]));
    assign outputs[6620] = ~((layer0_outputs[4828]) ^ (layer0_outputs[5057]));
    assign outputs[6621] = ~(layer0_outputs[2356]);
    assign outputs[6622] = layer0_outputs[3588];
    assign outputs[6623] = ~((layer0_outputs[3543]) | (layer0_outputs[9792]));
    assign outputs[6624] = (layer0_outputs[9594]) & ~(layer0_outputs[2075]);
    assign outputs[6625] = ~(layer0_outputs[8743]);
    assign outputs[6626] = ~(layer0_outputs[6215]);
    assign outputs[6627] = ~(layer0_outputs[6095]);
    assign outputs[6628] = layer0_outputs[2364];
    assign outputs[6629] = layer0_outputs[516];
    assign outputs[6630] = (layer0_outputs[4414]) & (layer0_outputs[7836]);
    assign outputs[6631] = ~((layer0_outputs[9559]) & (layer0_outputs[9952]));
    assign outputs[6632] = ~(layer0_outputs[6470]);
    assign outputs[6633] = ~((layer0_outputs[9076]) | (layer0_outputs[2550]));
    assign outputs[6634] = (layer0_outputs[2208]) ^ (layer0_outputs[1046]);
    assign outputs[6635] = ~((layer0_outputs[3897]) ^ (layer0_outputs[9552]));
    assign outputs[6636] = ~(layer0_outputs[8264]);
    assign outputs[6637] = (layer0_outputs[7332]) ^ (layer0_outputs[4850]);
    assign outputs[6638] = ~(layer0_outputs[852]) | (layer0_outputs[5636]);
    assign outputs[6639] = layer0_outputs[4238];
    assign outputs[6640] = ~((layer0_outputs[5691]) | (layer0_outputs[9863]));
    assign outputs[6641] = ~(layer0_outputs[3700]) | (layer0_outputs[9083]);
    assign outputs[6642] = (layer0_outputs[2989]) & ~(layer0_outputs[7795]);
    assign outputs[6643] = layer0_outputs[549];
    assign outputs[6644] = layer0_outputs[1560];
    assign outputs[6645] = (layer0_outputs[4232]) ^ (layer0_outputs[5106]);
    assign outputs[6646] = (layer0_outputs[8963]) ^ (layer0_outputs[4405]);
    assign outputs[6647] = layer0_outputs[9165];
    assign outputs[6648] = layer0_outputs[9734];
    assign outputs[6649] = layer0_outputs[2636];
    assign outputs[6650] = ~((layer0_outputs[1523]) | (layer0_outputs[8133]));
    assign outputs[6651] = layer0_outputs[6044];
    assign outputs[6652] = ~(layer0_outputs[8155]);
    assign outputs[6653] = ~(layer0_outputs[2911]);
    assign outputs[6654] = ~(layer0_outputs[1998]);
    assign outputs[6655] = (layer0_outputs[5462]) ^ (layer0_outputs[3506]);
    assign outputs[6656] = ~(layer0_outputs[8847]);
    assign outputs[6657] = (layer0_outputs[7699]) & ~(layer0_outputs[1733]);
    assign outputs[6658] = (layer0_outputs[5759]) & ~(layer0_outputs[374]);
    assign outputs[6659] = ~(layer0_outputs[6586]);
    assign outputs[6660] = ~((layer0_outputs[6724]) ^ (layer0_outputs[2452]));
    assign outputs[6661] = ~((layer0_outputs[5922]) ^ (layer0_outputs[7102]));
    assign outputs[6662] = (layer0_outputs[4265]) & ~(layer0_outputs[931]);
    assign outputs[6663] = (layer0_outputs[7192]) & (layer0_outputs[3728]);
    assign outputs[6664] = ~((layer0_outputs[2614]) | (layer0_outputs[1441]));
    assign outputs[6665] = ~((layer0_outputs[5723]) | (layer0_outputs[3812]));
    assign outputs[6666] = (layer0_outputs[9059]) & ~(layer0_outputs[4293]);
    assign outputs[6667] = ~((layer0_outputs[3650]) & (layer0_outputs[8524]));
    assign outputs[6668] = (layer0_outputs[6120]) | (layer0_outputs[5512]);
    assign outputs[6669] = (layer0_outputs[2572]) ^ (layer0_outputs[3250]);
    assign outputs[6670] = (layer0_outputs[1605]) ^ (layer0_outputs[6001]);
    assign outputs[6671] = ~((layer0_outputs[10071]) | (layer0_outputs[2085]));
    assign outputs[6672] = (layer0_outputs[9458]) ^ (layer0_outputs[6995]);
    assign outputs[6673] = layer0_outputs[8262];
    assign outputs[6674] = (layer0_outputs[1392]) ^ (layer0_outputs[2301]);
    assign outputs[6675] = layer0_outputs[4897];
    assign outputs[6676] = ~(layer0_outputs[3510]);
    assign outputs[6677] = (layer0_outputs[888]) & ~(layer0_outputs[9783]);
    assign outputs[6678] = (layer0_outputs[1026]) | (layer0_outputs[5225]);
    assign outputs[6679] = (layer0_outputs[6777]) ^ (layer0_outputs[4406]);
    assign outputs[6680] = ~(layer0_outputs[851]) | (layer0_outputs[8577]);
    assign outputs[6681] = layer0_outputs[6929];
    assign outputs[6682] = (layer0_outputs[2877]) ^ (layer0_outputs[3826]);
    assign outputs[6683] = (layer0_outputs[9201]) ^ (layer0_outputs[8523]);
    assign outputs[6684] = ~(layer0_outputs[8477]);
    assign outputs[6685] = (layer0_outputs[4369]) & (layer0_outputs[5257]);
    assign outputs[6686] = ~(layer0_outputs[1686]);
    assign outputs[6687] = ~(layer0_outputs[977]);
    assign outputs[6688] = layer0_outputs[9388];
    assign outputs[6689] = (layer0_outputs[4523]) | (layer0_outputs[9723]);
    assign outputs[6690] = layer0_outputs[3723];
    assign outputs[6691] = layer0_outputs[8522];
    assign outputs[6692] = layer0_outputs[1793];
    assign outputs[6693] = ~((layer0_outputs[3811]) ^ (layer0_outputs[9483]));
    assign outputs[6694] = ~((layer0_outputs[3486]) ^ (layer0_outputs[1032]));
    assign outputs[6695] = (layer0_outputs[8464]) & (layer0_outputs[4488]);
    assign outputs[6696] = (layer0_outputs[2124]) & (layer0_outputs[4862]);
    assign outputs[6697] = (layer0_outputs[1033]) & ~(layer0_outputs[959]);
    assign outputs[6698] = (layer0_outputs[9481]) & ~(layer0_outputs[2168]);
    assign outputs[6699] = ~((layer0_outputs[3837]) ^ (layer0_outputs[248]));
    assign outputs[6700] = ~(layer0_outputs[6545]);
    assign outputs[6701] = (layer0_outputs[6372]) & ~(layer0_outputs[4847]);
    assign outputs[6702] = (layer0_outputs[4116]) | (layer0_outputs[9112]);
    assign outputs[6703] = ~(layer0_outputs[2611]);
    assign outputs[6704] = ~((layer0_outputs[4626]) ^ (layer0_outputs[6644]));
    assign outputs[6705] = (layer0_outputs[5836]) ^ (layer0_outputs[301]);
    assign outputs[6706] = ~(layer0_outputs[5546]);
    assign outputs[6707] = (layer0_outputs[291]) & ~(layer0_outputs[2746]);
    assign outputs[6708] = ~(layer0_outputs[2608]);
    assign outputs[6709] = layer0_outputs[9744];
    assign outputs[6710] = layer0_outputs[9935];
    assign outputs[6711] = ~(layer0_outputs[4031]);
    assign outputs[6712] = layer0_outputs[514];
    assign outputs[6713] = ~(layer0_outputs[534]);
    assign outputs[6714] = ~((layer0_outputs[8307]) | (layer0_outputs[9361]));
    assign outputs[6715] = (layer0_outputs[6877]) & ~(layer0_outputs[2804]);
    assign outputs[6716] = ~((layer0_outputs[8824]) | (layer0_outputs[2178]));
    assign outputs[6717] = layer0_outputs[6911];
    assign outputs[6718] = layer0_outputs[7543];
    assign outputs[6719] = (layer0_outputs[8294]) & (layer0_outputs[5061]);
    assign outputs[6720] = (layer0_outputs[6581]) & (layer0_outputs[6931]);
    assign outputs[6721] = (layer0_outputs[7174]) & ~(layer0_outputs[8482]);
    assign outputs[6722] = ~(layer0_outputs[9374]);
    assign outputs[6723] = (layer0_outputs[8844]) & (layer0_outputs[7068]);
    assign outputs[6724] = (layer0_outputs[469]) & (layer0_outputs[9118]);
    assign outputs[6725] = ~(layer0_outputs[4063]);
    assign outputs[6726] = ~(layer0_outputs[4734]);
    assign outputs[6727] = layer0_outputs[7019];
    assign outputs[6728] = layer0_outputs[8603];
    assign outputs[6729] = ~(layer0_outputs[6209]) | (layer0_outputs[2083]);
    assign outputs[6730] = 1'b0;
    assign outputs[6731] = ~(layer0_outputs[1861]);
    assign outputs[6732] = ~(layer0_outputs[6308]);
    assign outputs[6733] = ~((layer0_outputs[1686]) | (layer0_outputs[6223]));
    assign outputs[6734] = ~(layer0_outputs[6987]);
    assign outputs[6735] = ~(layer0_outputs[1855]) | (layer0_outputs[1711]);
    assign outputs[6736] = layer0_outputs[9685];
    assign outputs[6737] = layer0_outputs[787];
    assign outputs[6738] = ~((layer0_outputs[6212]) ^ (layer0_outputs[7511]));
    assign outputs[6739] = layer0_outputs[560];
    assign outputs[6740] = (layer0_outputs[3522]) ^ (layer0_outputs[2716]);
    assign outputs[6741] = (layer0_outputs[10215]) ^ (layer0_outputs[1124]);
    assign outputs[6742] = ~(layer0_outputs[7892]);
    assign outputs[6743] = ~(layer0_outputs[3111]);
    assign outputs[6744] = (layer0_outputs[6235]) & ~(layer0_outputs[8290]);
    assign outputs[6745] = layer0_outputs[6246];
    assign outputs[6746] = (layer0_outputs[6759]) ^ (layer0_outputs[10073]);
    assign outputs[6747] = ~((layer0_outputs[1486]) & (layer0_outputs[1940]));
    assign outputs[6748] = (layer0_outputs[8192]) & ~(layer0_outputs[929]);
    assign outputs[6749] = ~(layer0_outputs[9982]);
    assign outputs[6750] = layer0_outputs[9817];
    assign outputs[6751] = ~((layer0_outputs[7151]) ^ (layer0_outputs[5959]));
    assign outputs[6752] = ~((layer0_outputs[5974]) ^ (layer0_outputs[4674]));
    assign outputs[6753] = ~((layer0_outputs[8393]) ^ (layer0_outputs[4148]));
    assign outputs[6754] = ~(layer0_outputs[5314]);
    assign outputs[6755] = ~((layer0_outputs[2260]) ^ (layer0_outputs[8100]));
    assign outputs[6756] = ~(layer0_outputs[10057]) | (layer0_outputs[8895]);
    assign outputs[6757] = layer0_outputs[8451];
    assign outputs[6758] = ~(layer0_outputs[7519]);
    assign outputs[6759] = ~((layer0_outputs[2772]) ^ (layer0_outputs[9607]));
    assign outputs[6760] = (layer0_outputs[8356]) ^ (layer0_outputs[9212]);
    assign outputs[6761] = layer0_outputs[5467];
    assign outputs[6762] = (layer0_outputs[404]) & ~(layer0_outputs[9834]);
    assign outputs[6763] = (layer0_outputs[6275]) & ~(layer0_outputs[7134]);
    assign outputs[6764] = ~((layer0_outputs[6408]) ^ (layer0_outputs[3542]));
    assign outputs[6765] = ~(layer0_outputs[262]);
    assign outputs[6766] = ~((layer0_outputs[5615]) ^ (layer0_outputs[2271]));
    assign outputs[6767] = (layer0_outputs[3515]) & ~(layer0_outputs[804]);
    assign outputs[6768] = (layer0_outputs[9415]) ^ (layer0_outputs[6733]);
    assign outputs[6769] = (layer0_outputs[2925]) & ~(layer0_outputs[4574]);
    assign outputs[6770] = layer0_outputs[3648];
    assign outputs[6771] = (layer0_outputs[8958]) ^ (layer0_outputs[1714]);
    assign outputs[6772] = (layer0_outputs[4171]) & (layer0_outputs[5646]);
    assign outputs[6773] = ~((layer0_outputs[3093]) & (layer0_outputs[214]));
    assign outputs[6774] = (layer0_outputs[8580]) & (layer0_outputs[5148]);
    assign outputs[6775] = ~(layer0_outputs[922]);
    assign outputs[6776] = ~((layer0_outputs[1385]) ^ (layer0_outputs[8007]));
    assign outputs[6777] = ~(layer0_outputs[8759]);
    assign outputs[6778] = ~((layer0_outputs[9211]) ^ (layer0_outputs[4105]));
    assign outputs[6779] = (layer0_outputs[6571]) ^ (layer0_outputs[366]);
    assign outputs[6780] = (layer0_outputs[6402]) | (layer0_outputs[8217]);
    assign outputs[6781] = layer0_outputs[6887];
    assign outputs[6782] = ~(layer0_outputs[1290]);
    assign outputs[6783] = ~(layer0_outputs[187]) | (layer0_outputs[1071]);
    assign outputs[6784] = ~(layer0_outputs[3687]);
    assign outputs[6785] = (layer0_outputs[9586]) & ~(layer0_outputs[10018]);
    assign outputs[6786] = ~((layer0_outputs[7298]) & (layer0_outputs[7128]));
    assign outputs[6787] = (layer0_outputs[8583]) & ~(layer0_outputs[5982]);
    assign outputs[6788] = (layer0_outputs[6019]) | (layer0_outputs[4640]);
    assign outputs[6789] = layer0_outputs[421];
    assign outputs[6790] = ~((layer0_outputs[5285]) ^ (layer0_outputs[1444]));
    assign outputs[6791] = ~(layer0_outputs[1674]);
    assign outputs[6792] = ~(layer0_outputs[7732]);
    assign outputs[6793] = (layer0_outputs[3232]) & (layer0_outputs[657]);
    assign outputs[6794] = 1'b0;
    assign outputs[6795] = ~(layer0_outputs[4901]);
    assign outputs[6796] = layer0_outputs[4019];
    assign outputs[6797] = (layer0_outputs[3693]) & (layer0_outputs[5411]);
    assign outputs[6798] = ~(layer0_outputs[9233]);
    assign outputs[6799] = ~((layer0_outputs[2880]) | (layer0_outputs[3877]));
    assign outputs[6800] = layer0_outputs[10196];
    assign outputs[6801] = ~(layer0_outputs[4940]);
    assign outputs[6802] = ~(layer0_outputs[9168]);
    assign outputs[6803] = ~((layer0_outputs[10147]) & (layer0_outputs[7900]));
    assign outputs[6804] = ~(layer0_outputs[8458]);
    assign outputs[6805] = (layer0_outputs[3148]) & ~(layer0_outputs[1981]);
    assign outputs[6806] = (layer0_outputs[5287]) ^ (layer0_outputs[6187]);
    assign outputs[6807] = ~((layer0_outputs[3581]) & (layer0_outputs[337]));
    assign outputs[6808] = (layer0_outputs[3655]) ^ (layer0_outputs[9683]);
    assign outputs[6809] = (layer0_outputs[7466]) ^ (layer0_outputs[9005]);
    assign outputs[6810] = layer0_outputs[2135];
    assign outputs[6811] = layer0_outputs[3090];
    assign outputs[6812] = ~(layer0_outputs[2035]);
    assign outputs[6813] = ~(layer0_outputs[608]);
    assign outputs[6814] = ~(layer0_outputs[642]);
    assign outputs[6815] = layer0_outputs[571];
    assign outputs[6816] = ~((layer0_outputs[8666]) ^ (layer0_outputs[761]));
    assign outputs[6817] = ~((layer0_outputs[7812]) | (layer0_outputs[958]));
    assign outputs[6818] = layer0_outputs[2903];
    assign outputs[6819] = ~(layer0_outputs[2832]);
    assign outputs[6820] = (layer0_outputs[4111]) & ~(layer0_outputs[5012]);
    assign outputs[6821] = (layer0_outputs[6006]) & (layer0_outputs[7414]);
    assign outputs[6822] = ~(layer0_outputs[5805]);
    assign outputs[6823] = (layer0_outputs[9768]) & (layer0_outputs[8013]);
    assign outputs[6824] = ~(layer0_outputs[1901]);
    assign outputs[6825] = layer0_outputs[3201];
    assign outputs[6826] = ~((layer0_outputs[9712]) & (layer0_outputs[6992]));
    assign outputs[6827] = (layer0_outputs[7529]) & (layer0_outputs[2818]);
    assign outputs[6828] = (layer0_outputs[7577]) & ~(layer0_outputs[9282]);
    assign outputs[6829] = ~((layer0_outputs[7735]) | (layer0_outputs[1494]));
    assign outputs[6830] = (layer0_outputs[5170]) & (layer0_outputs[3342]);
    assign outputs[6831] = ~(layer0_outputs[7911]);
    assign outputs[6832] = layer0_outputs[10155];
    assign outputs[6833] = ~(layer0_outputs[4520]);
    assign outputs[6834] = layer0_outputs[5397];
    assign outputs[6835] = ~(layer0_outputs[6366]);
    assign outputs[6836] = layer0_outputs[1330];
    assign outputs[6837] = (layer0_outputs[9996]) & (layer0_outputs[6588]);
    assign outputs[6838] = layer0_outputs[3078];
    assign outputs[6839] = ~(layer0_outputs[4229]);
    assign outputs[6840] = (layer0_outputs[9620]) & ~(layer0_outputs[7524]);
    assign outputs[6841] = ~(layer0_outputs[5346]);
    assign outputs[6842] = ~(layer0_outputs[8736]) | (layer0_outputs[8249]);
    assign outputs[6843] = ~(layer0_outputs[8211]);
    assign outputs[6844] = ~(layer0_outputs[7817]);
    assign outputs[6845] = ~(layer0_outputs[438]);
    assign outputs[6846] = ~(layer0_outputs[4486]) | (layer0_outputs[5715]);
    assign outputs[6847] = ~(layer0_outputs[5697]) | (layer0_outputs[5118]);
    assign outputs[6848] = ~(layer0_outputs[262]);
    assign outputs[6849] = (layer0_outputs[2454]) & ~(layer0_outputs[7397]);
    assign outputs[6850] = ~(layer0_outputs[7820]);
    assign outputs[6851] = layer0_outputs[4622];
    assign outputs[6852] = layer0_outputs[5659];
    assign outputs[6853] = layer0_outputs[3930];
    assign outputs[6854] = ~(layer0_outputs[971]);
    assign outputs[6855] = layer0_outputs[8144];
    assign outputs[6856] = ~(layer0_outputs[5038]);
    assign outputs[6857] = ~((layer0_outputs[8219]) ^ (layer0_outputs[7034]));
    assign outputs[6858] = ~(layer0_outputs[2014]);
    assign outputs[6859] = (layer0_outputs[8012]) | (layer0_outputs[7555]);
    assign outputs[6860] = (layer0_outputs[249]) & ~(layer0_outputs[9139]);
    assign outputs[6861] = ~((layer0_outputs[3878]) ^ (layer0_outputs[3587]));
    assign outputs[6862] = ~(layer0_outputs[6150]);
    assign outputs[6863] = (layer0_outputs[3620]) ^ (layer0_outputs[2290]);
    assign outputs[6864] = layer0_outputs[5383];
    assign outputs[6865] = (layer0_outputs[8430]) ^ (layer0_outputs[2495]);
    assign outputs[6866] = ~((layer0_outputs[2767]) ^ (layer0_outputs[5949]));
    assign outputs[6867] = ~(layer0_outputs[1161]) | (layer0_outputs[4990]);
    assign outputs[6868] = ~((layer0_outputs[3162]) | (layer0_outputs[2226]));
    assign outputs[6869] = ~(layer0_outputs[3195]) | (layer0_outputs[1495]);
    assign outputs[6870] = ~(layer0_outputs[8922]);
    assign outputs[6871] = layer0_outputs[75];
    assign outputs[6872] = ~((layer0_outputs[8267]) ^ (layer0_outputs[3256]));
    assign outputs[6873] = ~((layer0_outputs[2128]) | (layer0_outputs[1012]));
    assign outputs[6874] = ~((layer0_outputs[3763]) ^ (layer0_outputs[4834]));
    assign outputs[6875] = layer0_outputs[3011];
    assign outputs[6876] = ~(layer0_outputs[890]);
    assign outputs[6877] = (layer0_outputs[815]) ^ (layer0_outputs[9729]);
    assign outputs[6878] = layer0_outputs[8148];
    assign outputs[6879] = layer0_outputs[9414];
    assign outputs[6880] = layer0_outputs[9817];
    assign outputs[6881] = (layer0_outputs[9916]) & (layer0_outputs[6419]);
    assign outputs[6882] = ~((layer0_outputs[3180]) | (layer0_outputs[5242]));
    assign outputs[6883] = ~((layer0_outputs[9621]) ^ (layer0_outputs[7750]));
    assign outputs[6884] = layer0_outputs[3258];
    assign outputs[6885] = ~(layer0_outputs[2643]);
    assign outputs[6886] = (layer0_outputs[4738]) & ~(layer0_outputs[5508]);
    assign outputs[6887] = ~((layer0_outputs[862]) ^ (layer0_outputs[5084]));
    assign outputs[6888] = layer0_outputs[6073];
    assign outputs[6889] = (layer0_outputs[2630]) ^ (layer0_outputs[7269]);
    assign outputs[6890] = (layer0_outputs[10090]) & (layer0_outputs[233]);
    assign outputs[6891] = layer0_outputs[189];
    assign outputs[6892] = ~((layer0_outputs[8341]) | (layer0_outputs[7079]));
    assign outputs[6893] = (layer0_outputs[4295]) & (layer0_outputs[7565]);
    assign outputs[6894] = (layer0_outputs[3125]) ^ (layer0_outputs[7775]);
    assign outputs[6895] = layer0_outputs[9420];
    assign outputs[6896] = ~((layer0_outputs[8024]) ^ (layer0_outputs[9934]));
    assign outputs[6897] = (layer0_outputs[7818]) ^ (layer0_outputs[37]);
    assign outputs[6898] = ~((layer0_outputs[7605]) & (layer0_outputs[5447]));
    assign outputs[6899] = ~((layer0_outputs[3599]) ^ (layer0_outputs[83]));
    assign outputs[6900] = ~((layer0_outputs[191]) | (layer0_outputs[9956]));
    assign outputs[6901] = layer0_outputs[2451];
    assign outputs[6902] = layer0_outputs[663];
    assign outputs[6903] = (layer0_outputs[8204]) ^ (layer0_outputs[4629]);
    assign outputs[6904] = ~((layer0_outputs[322]) ^ (layer0_outputs[6195]));
    assign outputs[6905] = (layer0_outputs[9419]) ^ (layer0_outputs[2449]);
    assign outputs[6906] = ~((layer0_outputs[1997]) | (layer0_outputs[4058]));
    assign outputs[6907] = layer0_outputs[1967];
    assign outputs[6908] = ~(layer0_outputs[2430]) | (layer0_outputs[10175]);
    assign outputs[6909] = layer0_outputs[6663];
    assign outputs[6910] = layer0_outputs[6888];
    assign outputs[6911] = (layer0_outputs[9178]) & (layer0_outputs[7522]);
    assign outputs[6912] = layer0_outputs[5207];
    assign outputs[6913] = ~(layer0_outputs[8641]) | (layer0_outputs[544]);
    assign outputs[6914] = layer0_outputs[10198];
    assign outputs[6915] = ~(layer0_outputs[5807]);
    assign outputs[6916] = (layer0_outputs[4617]) ^ (layer0_outputs[9402]);
    assign outputs[6917] = ~(layer0_outputs[378]);
    assign outputs[6918] = ~(layer0_outputs[10087]);
    assign outputs[6919] = layer0_outputs[2216];
    assign outputs[6920] = ~((layer0_outputs[4643]) ^ (layer0_outputs[7299]));
    assign outputs[6921] = (layer0_outputs[90]) & ~(layer0_outputs[5059]);
    assign outputs[6922] = (layer0_outputs[8835]) & ~(layer0_outputs[3369]);
    assign outputs[6923] = (layer0_outputs[10121]) ^ (layer0_outputs[3060]);
    assign outputs[6924] = (layer0_outputs[3163]) & ~(layer0_outputs[1919]);
    assign outputs[6925] = ~((layer0_outputs[9962]) ^ (layer0_outputs[3316]));
    assign outputs[6926] = layer0_outputs[4296];
    assign outputs[6927] = (layer0_outputs[7287]) & ~(layer0_outputs[3472]);
    assign outputs[6928] = ~((layer0_outputs[2671]) | (layer0_outputs[132]));
    assign outputs[6929] = (layer0_outputs[6907]) ^ (layer0_outputs[10128]);
    assign outputs[6930] = ~(layer0_outputs[2922]) | (layer0_outputs[946]);
    assign outputs[6931] = layer0_outputs[9630];
    assign outputs[6932] = ~((layer0_outputs[3560]) | (layer0_outputs[694]));
    assign outputs[6933] = (layer0_outputs[6231]) | (layer0_outputs[5370]);
    assign outputs[6934] = (layer0_outputs[1110]) & ~(layer0_outputs[4948]);
    assign outputs[6935] = (layer0_outputs[746]) | (layer0_outputs[2156]);
    assign outputs[6936] = (layer0_outputs[8098]) ^ (layer0_outputs[6094]);
    assign outputs[6937] = ~(layer0_outputs[509]);
    assign outputs[6938] = layer0_outputs[7730];
    assign outputs[6939] = ~((layer0_outputs[7358]) | (layer0_outputs[2112]));
    assign outputs[6940] = ~(layer0_outputs[185]);
    assign outputs[6941] = layer0_outputs[5667];
    assign outputs[6942] = (layer0_outputs[7340]) | (layer0_outputs[8770]);
    assign outputs[6943] = (layer0_outputs[6458]) & (layer0_outputs[6238]);
    assign outputs[6944] = layer0_outputs[3959];
    assign outputs[6945] = ~(layer0_outputs[4591]);
    assign outputs[6946] = ~(layer0_outputs[6852]) | (layer0_outputs[5413]);
    assign outputs[6947] = (layer0_outputs[8080]) & ~(layer0_outputs[515]);
    assign outputs[6948] = ~((layer0_outputs[9037]) ^ (layer0_outputs[6994]));
    assign outputs[6949] = ~(layer0_outputs[7516]);
    assign outputs[6950] = ~(layer0_outputs[802]);
    assign outputs[6951] = ~(layer0_outputs[3966]);
    assign outputs[6952] = ~(layer0_outputs[7108]);
    assign outputs[6953] = ~((layer0_outputs[8671]) | (layer0_outputs[6699]));
    assign outputs[6954] = ~((layer0_outputs[9785]) & (layer0_outputs[7054]));
    assign outputs[6955] = (layer0_outputs[204]) & (layer0_outputs[874]);
    assign outputs[6956] = ~((layer0_outputs[8300]) | (layer0_outputs[1479]));
    assign outputs[6957] = (layer0_outputs[3857]) ^ (layer0_outputs[5285]);
    assign outputs[6958] = (layer0_outputs[4265]) & ~(layer0_outputs[6694]);
    assign outputs[6959] = ~((layer0_outputs[1656]) ^ (layer0_outputs[8275]));
    assign outputs[6960] = (layer0_outputs[7288]) ^ (layer0_outputs[9123]);
    assign outputs[6961] = layer0_outputs[8302];
    assign outputs[6962] = ~((layer0_outputs[3281]) ^ (layer0_outputs[6932]));
    assign outputs[6963] = ~(layer0_outputs[8703]);
    assign outputs[6964] = ~((layer0_outputs[6437]) ^ (layer0_outputs[8471]));
    assign outputs[6965] = (layer0_outputs[3612]) & ~(layer0_outputs[2344]);
    assign outputs[6966] = (layer0_outputs[7154]) ^ (layer0_outputs[93]);
    assign outputs[6967] = (layer0_outputs[8870]) ^ (layer0_outputs[7133]);
    assign outputs[6968] = ~(layer0_outputs[8196]);
    assign outputs[6969] = ~(layer0_outputs[3580]);
    assign outputs[6970] = layer0_outputs[9780];
    assign outputs[6971] = layer0_outputs[2003];
    assign outputs[6972] = (layer0_outputs[321]) & ~(layer0_outputs[7519]);
    assign outputs[6973] = layer0_outputs[7997];
    assign outputs[6974] = ~(layer0_outputs[6203]);
    assign outputs[6975] = ~(layer0_outputs[5420]);
    assign outputs[6976] = ~(layer0_outputs[2990]);
    assign outputs[6977] = ~((layer0_outputs[6525]) & (layer0_outputs[2373]));
    assign outputs[6978] = ~((layer0_outputs[2802]) & (layer0_outputs[5004]));
    assign outputs[6979] = layer0_outputs[4332];
    assign outputs[6980] = (layer0_outputs[4637]) ^ (layer0_outputs[93]);
    assign outputs[6981] = layer0_outputs[7247];
    assign outputs[6982] = ~(layer0_outputs[5807]) | (layer0_outputs[5185]);
    assign outputs[6983] = ~(layer0_outputs[8118]);
    assign outputs[6984] = (layer0_outputs[1191]) ^ (layer0_outputs[1123]);
    assign outputs[6985] = ~((layer0_outputs[7278]) ^ (layer0_outputs[3140]));
    assign outputs[6986] = (layer0_outputs[4145]) ^ (layer0_outputs[1896]);
    assign outputs[6987] = (layer0_outputs[2798]) & ~(layer0_outputs[6917]);
    assign outputs[6988] = ~((layer0_outputs[1378]) | (layer0_outputs[5393]));
    assign outputs[6989] = ~(layer0_outputs[1199]);
    assign outputs[6990] = layer0_outputs[4989];
    assign outputs[6991] = ~(layer0_outputs[1300]) | (layer0_outputs[5976]);
    assign outputs[6992] = layer0_outputs[1869];
    assign outputs[6993] = (layer0_outputs[6489]) ^ (layer0_outputs[8944]);
    assign outputs[6994] = ~(layer0_outputs[5455]) | (layer0_outputs[6039]);
    assign outputs[6995] = (layer0_outputs[2823]) & (layer0_outputs[6146]);
    assign outputs[6996] = ~(layer0_outputs[3513]) | (layer0_outputs[8262]);
    assign outputs[6997] = ~((layer0_outputs[2893]) & (layer0_outputs[3344]));
    assign outputs[6998] = (layer0_outputs[4008]) ^ (layer0_outputs[4891]);
    assign outputs[6999] = ~(layer0_outputs[8341]);
    assign outputs[7000] = ~(layer0_outputs[9801]);
    assign outputs[7001] = layer0_outputs[2700];
    assign outputs[7002] = layer0_outputs[2206];
    assign outputs[7003] = layer0_outputs[3852];
    assign outputs[7004] = layer0_outputs[4118];
    assign outputs[7005] = (layer0_outputs[8053]) & ~(layer0_outputs[5960]);
    assign outputs[7006] = layer0_outputs[3269];
    assign outputs[7007] = (layer0_outputs[7324]) ^ (layer0_outputs[8587]);
    assign outputs[7008] = ~(layer0_outputs[199]);
    assign outputs[7009] = layer0_outputs[5022];
    assign outputs[7010] = layer0_outputs[2093];
    assign outputs[7011] = layer0_outputs[6831];
    assign outputs[7012] = (layer0_outputs[2673]) & (layer0_outputs[9622]);
    assign outputs[7013] = layer0_outputs[9078];
    assign outputs[7014] = ~((layer0_outputs[7075]) ^ (layer0_outputs[595]));
    assign outputs[7015] = ~(layer0_outputs[6317]);
    assign outputs[7016] = ~(layer0_outputs[3967]);
    assign outputs[7017] = ~((layer0_outputs[6314]) & (layer0_outputs[4637]));
    assign outputs[7018] = ~((layer0_outputs[1080]) ^ (layer0_outputs[2866]));
    assign outputs[7019] = ~(layer0_outputs[2306]);
    assign outputs[7020] = ~(layer0_outputs[4679]) | (layer0_outputs[1931]);
    assign outputs[7021] = (layer0_outputs[1449]) ^ (layer0_outputs[10100]);
    assign outputs[7022] = layer0_outputs[6480];
    assign outputs[7023] = 1'b1;
    assign outputs[7024] = (layer0_outputs[1518]) & ~(layer0_outputs[4591]);
    assign outputs[7025] = (layer0_outputs[9052]) & ~(layer0_outputs[1727]);
    assign outputs[7026] = ~((layer0_outputs[4877]) & (layer0_outputs[9136]));
    assign outputs[7027] = ~(layer0_outputs[2367]);
    assign outputs[7028] = layer0_outputs[4978];
    assign outputs[7029] = ~(layer0_outputs[3934]);
    assign outputs[7030] = layer0_outputs[4272];
    assign outputs[7031] = layer0_outputs[10118];
    assign outputs[7032] = ~(layer0_outputs[8242]) | (layer0_outputs[904]);
    assign outputs[7033] = layer0_outputs[250];
    assign outputs[7034] = ~((layer0_outputs[4628]) ^ (layer0_outputs[8302]));
    assign outputs[7035] = ~(layer0_outputs[835]) | (layer0_outputs[3098]);
    assign outputs[7036] = ~(layer0_outputs[9144]);
    assign outputs[7037] = layer0_outputs[3520];
    assign outputs[7038] = ~((layer0_outputs[3360]) | (layer0_outputs[3401]));
    assign outputs[7039] = ~(layer0_outputs[3622]) | (layer0_outputs[6410]);
    assign outputs[7040] = ~(layer0_outputs[10071]) | (layer0_outputs[7908]);
    assign outputs[7041] = ~(layer0_outputs[2205]);
    assign outputs[7042] = layer0_outputs[4283];
    assign outputs[7043] = ~(layer0_outputs[9823]);
    assign outputs[7044] = (layer0_outputs[614]) & ~(layer0_outputs[4535]);
    assign outputs[7045] = ~(layer0_outputs[6658]) | (layer0_outputs[10080]);
    assign outputs[7046] = (layer0_outputs[8858]) ^ (layer0_outputs[8830]);
    assign outputs[7047] = layer0_outputs[577];
    assign outputs[7048] = ~((layer0_outputs[9412]) ^ (layer0_outputs[2074]));
    assign outputs[7049] = ~((layer0_outputs[4793]) | (layer0_outputs[8443]));
    assign outputs[7050] = ~(layer0_outputs[3382]);
    assign outputs[7051] = layer0_outputs[3607];
    assign outputs[7052] = ~(layer0_outputs[6854]);
    assign outputs[7053] = layer0_outputs[2506];
    assign outputs[7054] = ~((layer0_outputs[8914]) ^ (layer0_outputs[2021]));
    assign outputs[7055] = ~(layer0_outputs[10184]);
    assign outputs[7056] = layer0_outputs[6675];
    assign outputs[7057] = ~((layer0_outputs[6682]) ^ (layer0_outputs[1495]));
    assign outputs[7058] = (layer0_outputs[7891]) | (layer0_outputs[10202]);
    assign outputs[7059] = (layer0_outputs[4087]) & ~(layer0_outputs[2955]);
    assign outputs[7060] = layer0_outputs[7328];
    assign outputs[7061] = (layer0_outputs[3254]) & ~(layer0_outputs[3003]);
    assign outputs[7062] = layer0_outputs[3480];
    assign outputs[7063] = (layer0_outputs[287]) ^ (layer0_outputs[9405]);
    assign outputs[7064] = layer0_outputs[3795];
    assign outputs[7065] = (layer0_outputs[1017]) & ~(layer0_outputs[3932]);
    assign outputs[7066] = ~(layer0_outputs[1175]);
    assign outputs[7067] = (layer0_outputs[10014]) | (layer0_outputs[8826]);
    assign outputs[7068] = layer0_outputs[5853];
    assign outputs[7069] = 1'b1;
    assign outputs[7070] = (layer0_outputs[3646]) & ~(layer0_outputs[394]);
    assign outputs[7071] = layer0_outputs[7259];
    assign outputs[7072] = ~(layer0_outputs[8210]);
    assign outputs[7073] = (layer0_outputs[8450]) & ~(layer0_outputs[213]);
    assign outputs[7074] = (layer0_outputs[5023]) & ~(layer0_outputs[5277]);
    assign outputs[7075] = ~(layer0_outputs[72]);
    assign outputs[7076] = ~(layer0_outputs[1006]);
    assign outputs[7077] = layer0_outputs[7643];
    assign outputs[7078] = (layer0_outputs[8910]) | (layer0_outputs[7827]);
    assign outputs[7079] = ~((layer0_outputs[7661]) ^ (layer0_outputs[5030]));
    assign outputs[7080] = ~((layer0_outputs[8659]) ^ (layer0_outputs[4381]));
    assign outputs[7081] = layer0_outputs[8008];
    assign outputs[7082] = ~(layer0_outputs[6024]) | (layer0_outputs[8475]);
    assign outputs[7083] = ~((layer0_outputs[4206]) ^ (layer0_outputs[9557]));
    assign outputs[7084] = ~((layer0_outputs[9126]) & (layer0_outputs[6232]));
    assign outputs[7085] = (layer0_outputs[4259]) & ~(layer0_outputs[4467]);
    assign outputs[7086] = (layer0_outputs[3653]) & ~(layer0_outputs[8654]);
    assign outputs[7087] = ~(layer0_outputs[2832]);
    assign outputs[7088] = ~((layer0_outputs[5936]) ^ (layer0_outputs[3246]));
    assign outputs[7089] = layer0_outputs[5552];
    assign outputs[7090] = ~(layer0_outputs[2065]);
    assign outputs[7091] = (layer0_outputs[7403]) | (layer0_outputs[1944]);
    assign outputs[7092] = layer0_outputs[4028];
    assign outputs[7093] = ~(layer0_outputs[603]);
    assign outputs[7094] = ~(layer0_outputs[4199]);
    assign outputs[7095] = ~(layer0_outputs[6045]);
    assign outputs[7096] = (layer0_outputs[4869]) ^ (layer0_outputs[9286]);
    assign outputs[7097] = layer0_outputs[6026];
    assign outputs[7098] = (layer0_outputs[7365]) ^ (layer0_outputs[7821]);
    assign outputs[7099] = ~(layer0_outputs[8554]);
    assign outputs[7100] = (layer0_outputs[2144]) & (layer0_outputs[3185]);
    assign outputs[7101] = layer0_outputs[377];
    assign outputs[7102] = ~(layer0_outputs[378]) | (layer0_outputs[7081]);
    assign outputs[7103] = ~((layer0_outputs[2690]) | (layer0_outputs[2085]));
    assign outputs[7104] = ~((layer0_outputs[9324]) ^ (layer0_outputs[2102]));
    assign outputs[7105] = ~(layer0_outputs[3615]) | (layer0_outputs[2335]);
    assign outputs[7106] = (layer0_outputs[1503]) & ~(layer0_outputs[3354]);
    assign outputs[7107] = ~(layer0_outputs[7515]);
    assign outputs[7108] = (layer0_outputs[1061]) & ~(layer0_outputs[186]);
    assign outputs[7109] = (layer0_outputs[8543]) & (layer0_outputs[8120]);
    assign outputs[7110] = (layer0_outputs[6664]) & ~(layer0_outputs[6333]);
    assign outputs[7111] = ~(layer0_outputs[5672]);
    assign outputs[7112] = layer0_outputs[811];
    assign outputs[7113] = (layer0_outputs[8611]) ^ (layer0_outputs[2559]);
    assign outputs[7114] = layer0_outputs[7346];
    assign outputs[7115] = 1'b0;
    assign outputs[7116] = layer0_outputs[586];
    assign outputs[7117] = ~(layer0_outputs[3314]);
    assign outputs[7118] = ~((layer0_outputs[5094]) ^ (layer0_outputs[4303]));
    assign outputs[7119] = (layer0_outputs[6901]) ^ (layer0_outputs[7130]);
    assign outputs[7120] = layer0_outputs[1331];
    assign outputs[7121] = ~((layer0_outputs[8630]) ^ (layer0_outputs[10143]));
    assign outputs[7122] = ~(layer0_outputs[5856]);
    assign outputs[7123] = ~((layer0_outputs[9678]) ^ (layer0_outputs[8654]));
    assign outputs[7124] = layer0_outputs[2691];
    assign outputs[7125] = ~(layer0_outputs[4249]);
    assign outputs[7126] = ~(layer0_outputs[5356]);
    assign outputs[7127] = (layer0_outputs[5760]) & ~(layer0_outputs[3598]);
    assign outputs[7128] = (layer0_outputs[643]) & ~(layer0_outputs[10068]);
    assign outputs[7129] = (layer0_outputs[1721]) & ~(layer0_outputs[9626]);
    assign outputs[7130] = (layer0_outputs[1033]) & ~(layer0_outputs[8550]);
    assign outputs[7131] = layer0_outputs[5443];
    assign outputs[7132] = ~(layer0_outputs[5019]);
    assign outputs[7133] = ~((layer0_outputs[6791]) ^ (layer0_outputs[342]));
    assign outputs[7134] = ~(layer0_outputs[7668]);
    assign outputs[7135] = ~((layer0_outputs[2789]) & (layer0_outputs[9576]));
    assign outputs[7136] = ~((layer0_outputs[9960]) ^ (layer0_outputs[4065]));
    assign outputs[7137] = ~(layer0_outputs[2976]);
    assign outputs[7138] = layer0_outputs[7181];
    assign outputs[7139] = (layer0_outputs[5456]) & (layer0_outputs[3193]);
    assign outputs[7140] = (layer0_outputs[3268]) ^ (layer0_outputs[5446]);
    assign outputs[7141] = layer0_outputs[6243];
    assign outputs[7142] = ~((layer0_outputs[241]) ^ (layer0_outputs[7564]));
    assign outputs[7143] = layer0_outputs[7293];
    assign outputs[7144] = (layer0_outputs[3866]) ^ (layer0_outputs[3178]);
    assign outputs[7145] = ~((layer0_outputs[7357]) | (layer0_outputs[9006]));
    assign outputs[7146] = (layer0_outputs[6535]) & ~(layer0_outputs[3583]);
    assign outputs[7147] = (layer0_outputs[6071]) & ~(layer0_outputs[1186]);
    assign outputs[7148] = layer0_outputs[2005];
    assign outputs[7149] = ~(layer0_outputs[3572]);
    assign outputs[7150] = ~((layer0_outputs[1891]) ^ (layer0_outputs[1501]));
    assign outputs[7151] = ~((layer0_outputs[10128]) & (layer0_outputs[9396]));
    assign outputs[7152] = (layer0_outputs[1380]) & ~(layer0_outputs[5810]);
    assign outputs[7153] = (layer0_outputs[4374]) & ~(layer0_outputs[1151]);
    assign outputs[7154] = ~((layer0_outputs[5098]) & (layer0_outputs[954]));
    assign outputs[7155] = layer0_outputs[6662];
    assign outputs[7156] = (layer0_outputs[7283]) & ~(layer0_outputs[6586]);
    assign outputs[7157] = ~(layer0_outputs[2994]) | (layer0_outputs[1663]);
    assign outputs[7158] = ~((layer0_outputs[7614]) ^ (layer0_outputs[1994]));
    assign outputs[7159] = (layer0_outputs[7551]) & ~(layer0_outputs[975]);
    assign outputs[7160] = (layer0_outputs[9090]) & ~(layer0_outputs[6183]);
    assign outputs[7161] = layer0_outputs[8603];
    assign outputs[7162] = ~((layer0_outputs[1601]) ^ (layer0_outputs[206]));
    assign outputs[7163] = (layer0_outputs[9359]) ^ (layer0_outputs[8354]);
    assign outputs[7164] = ~(layer0_outputs[6274]);
    assign outputs[7165] = layer0_outputs[7808];
    assign outputs[7166] = ~((layer0_outputs[8232]) ^ (layer0_outputs[10227]));
    assign outputs[7167] = ~(layer0_outputs[852]);
    assign outputs[7168] = ~((layer0_outputs[4020]) | (layer0_outputs[7278]));
    assign outputs[7169] = (layer0_outputs[3177]) & ~(layer0_outputs[9138]);
    assign outputs[7170] = layer0_outputs[6779];
    assign outputs[7171] = (layer0_outputs[6709]) ^ (layer0_outputs[7785]);
    assign outputs[7172] = layer0_outputs[6199];
    assign outputs[7173] = ~(layer0_outputs[1234]);
    assign outputs[7174] = layer0_outputs[2853];
    assign outputs[7175] = layer0_outputs[4916];
    assign outputs[7176] = (layer0_outputs[9545]) & ~(layer0_outputs[2135]);
    assign outputs[7177] = (layer0_outputs[3512]) ^ (layer0_outputs[9920]);
    assign outputs[7178] = (layer0_outputs[8206]) & ~(layer0_outputs[7825]);
    assign outputs[7179] = ~(layer0_outputs[5259]);
    assign outputs[7180] = ~(layer0_outputs[466]) | (layer0_outputs[3066]);
    assign outputs[7181] = (layer0_outputs[998]) & (layer0_outputs[9921]);
    assign outputs[7182] = (layer0_outputs[1831]) ^ (layer0_outputs[633]);
    assign outputs[7183] = ~(layer0_outputs[8442]);
    assign outputs[7184] = ~(layer0_outputs[632]);
    assign outputs[7185] = ~(layer0_outputs[5429]) | (layer0_outputs[7625]);
    assign outputs[7186] = layer0_outputs[5024];
    assign outputs[7187] = ~(layer0_outputs[10087]) | (layer0_outputs[9980]);
    assign outputs[7188] = ~((layer0_outputs[3831]) ^ (layer0_outputs[2101]));
    assign outputs[7189] = ~((layer0_outputs[4967]) | (layer0_outputs[1147]));
    assign outputs[7190] = (layer0_outputs[9582]) & ~(layer0_outputs[1975]);
    assign outputs[7191] = layer0_outputs[6954];
    assign outputs[7192] = ~((layer0_outputs[8846]) ^ (layer0_outputs[6307]));
    assign outputs[7193] = ~(layer0_outputs[1261]);
    assign outputs[7194] = (layer0_outputs[2469]) & ~(layer0_outputs[410]);
    assign outputs[7195] = ~((layer0_outputs[148]) | (layer0_outputs[6025]));
    assign outputs[7196] = ~(layer0_outputs[558]);
    assign outputs[7197] = layer0_outputs[5442];
    assign outputs[7198] = ~(layer0_outputs[5552]) | (layer0_outputs[3486]);
    assign outputs[7199] = ~((layer0_outputs[9484]) | (layer0_outputs[5893]));
    assign outputs[7200] = (layer0_outputs[9886]) ^ (layer0_outputs[9971]);
    assign outputs[7201] = layer0_outputs[9182];
    assign outputs[7202] = ~((layer0_outputs[6602]) | (layer0_outputs[5174]));
    assign outputs[7203] = (layer0_outputs[5016]) & ~(layer0_outputs[2369]);
    assign outputs[7204] = layer0_outputs[4432];
    assign outputs[7205] = (layer0_outputs[434]) & ~(layer0_outputs[3869]);
    assign outputs[7206] = (layer0_outputs[7370]) & (layer0_outputs[8893]);
    assign outputs[7207] = (layer0_outputs[8696]) & ~(layer0_outputs[388]);
    assign outputs[7208] = ~(layer0_outputs[5888]) | (layer0_outputs[7564]);
    assign outputs[7209] = layer0_outputs[7708];
    assign outputs[7210] = layer0_outputs[4104];
    assign outputs[7211] = layer0_outputs[9505];
    assign outputs[7212] = ~(layer0_outputs[7566]);
    assign outputs[7213] = (layer0_outputs[3730]) & (layer0_outputs[6635]);
    assign outputs[7214] = (layer0_outputs[7542]) & ~(layer0_outputs[4500]);
    assign outputs[7215] = (layer0_outputs[8541]) & (layer0_outputs[2755]);
    assign outputs[7216] = layer0_outputs[2980];
    assign outputs[7217] = layer0_outputs[9670];
    assign outputs[7218] = layer0_outputs[731];
    assign outputs[7219] = layer0_outputs[7543];
    assign outputs[7220] = (layer0_outputs[8055]) & (layer0_outputs[8327]);
    assign outputs[7221] = ~(layer0_outputs[2127]) | (layer0_outputs[2459]);
    assign outputs[7222] = ~((layer0_outputs[8610]) & (layer0_outputs[2042]));
    assign outputs[7223] = ~(layer0_outputs[1930]);
    assign outputs[7224] = ~((layer0_outputs[342]) | (layer0_outputs[2476]));
    assign outputs[7225] = (layer0_outputs[5879]) | (layer0_outputs[4736]);
    assign outputs[7226] = ~((layer0_outputs[8295]) ^ (layer0_outputs[5013]));
    assign outputs[7227] = layer0_outputs[4600];
    assign outputs[7228] = ~(layer0_outputs[2258]) | (layer0_outputs[7076]);
    assign outputs[7229] = (layer0_outputs[8539]) ^ (layer0_outputs[3537]);
    assign outputs[7230] = ~(layer0_outputs[8653]);
    assign outputs[7231] = (layer0_outputs[5791]) & ~(layer0_outputs[2206]);
    assign outputs[7232] = (layer0_outputs[4529]) & ~(layer0_outputs[624]);
    assign outputs[7233] = ~((layer0_outputs[2353]) & (layer0_outputs[6099]));
    assign outputs[7234] = (layer0_outputs[1460]) & ~(layer0_outputs[7071]);
    assign outputs[7235] = ~(layer0_outputs[7692]);
    assign outputs[7236] = ~(layer0_outputs[4415]);
    assign outputs[7237] = ~((layer0_outputs[3729]) & (layer0_outputs[6566]));
    assign outputs[7238] = ~((layer0_outputs[9323]) ^ (layer0_outputs[10183]));
    assign outputs[7239] = ~((layer0_outputs[3638]) ^ (layer0_outputs[8712]));
    assign outputs[7240] = (layer0_outputs[8023]) ^ (layer0_outputs[10058]);
    assign outputs[7241] = ~((layer0_outputs[8981]) ^ (layer0_outputs[9711]));
    assign outputs[7242] = ~(layer0_outputs[9725]);
    assign outputs[7243] = (layer0_outputs[8083]) ^ (layer0_outputs[1372]);
    assign outputs[7244] = (layer0_outputs[7043]) & ~(layer0_outputs[4502]);
    assign outputs[7245] = (layer0_outputs[8773]) & ~(layer0_outputs[1128]);
    assign outputs[7246] = layer0_outputs[7598];
    assign outputs[7247] = ~(layer0_outputs[26]);
    assign outputs[7248] = ~((layer0_outputs[4117]) ^ (layer0_outputs[4833]));
    assign outputs[7249] = ~(layer0_outputs[8596]) | (layer0_outputs[6952]);
    assign outputs[7250] = ~(layer0_outputs[713]);
    assign outputs[7251] = layer0_outputs[349];
    assign outputs[7252] = layer0_outputs[8061];
    assign outputs[7253] = (layer0_outputs[8999]) ^ (layer0_outputs[5112]);
    assign outputs[7254] = ~((layer0_outputs[4708]) & (layer0_outputs[7621]));
    assign outputs[7255] = layer0_outputs[5144];
    assign outputs[7256] = ~((layer0_outputs[2511]) | (layer0_outputs[674]));
    assign outputs[7257] = (layer0_outputs[6985]) & (layer0_outputs[2414]);
    assign outputs[7258] = ~((layer0_outputs[3647]) | (layer0_outputs[4195]));
    assign outputs[7259] = (layer0_outputs[5209]) & (layer0_outputs[6531]);
    assign outputs[7260] = layer0_outputs[3538];
    assign outputs[7261] = (layer0_outputs[1536]) & ~(layer0_outputs[7056]);
    assign outputs[7262] = layer0_outputs[3794];
    assign outputs[7263] = ~(layer0_outputs[778]) | (layer0_outputs[1673]);
    assign outputs[7264] = ~(layer0_outputs[8647]);
    assign outputs[7265] = ~((layer0_outputs[2821]) ^ (layer0_outputs[1074]));
    assign outputs[7266] = 1'b0;
    assign outputs[7267] = layer0_outputs[1492];
    assign outputs[7268] = (layer0_outputs[6974]) & (layer0_outputs[2323]);
    assign outputs[7269] = ~(layer0_outputs[2620]);
    assign outputs[7270] = ~(layer0_outputs[6713]);
    assign outputs[7271] = ~(layer0_outputs[9016]);
    assign outputs[7272] = (layer0_outputs[77]) & (layer0_outputs[8605]);
    assign outputs[7273] = layer0_outputs[4457];
    assign outputs[7274] = ~(layer0_outputs[7330]);
    assign outputs[7275] = (layer0_outputs[2752]) ^ (layer0_outputs[370]);
    assign outputs[7276] = (layer0_outputs[4231]) | (layer0_outputs[8049]);
    assign outputs[7277] = ~((layer0_outputs[9047]) ^ (layer0_outputs[9429]));
    assign outputs[7278] = layer0_outputs[7942];
    assign outputs[7279] = ~(layer0_outputs[5300]);
    assign outputs[7280] = (layer0_outputs[3225]) ^ (layer0_outputs[4832]);
    assign outputs[7281] = layer0_outputs[2025];
    assign outputs[7282] = ~((layer0_outputs[752]) ^ (layer0_outputs[7961]));
    assign outputs[7283] = layer0_outputs[8669];
    assign outputs[7284] = ~((layer0_outputs[6441]) ^ (layer0_outputs[4972]));
    assign outputs[7285] = layer0_outputs[209];
    assign outputs[7286] = layer0_outputs[3384];
    assign outputs[7287] = ~((layer0_outputs[497]) | (layer0_outputs[282]));
    assign outputs[7288] = ~((layer0_outputs[6777]) | (layer0_outputs[2217]));
    assign outputs[7289] = (layer0_outputs[2320]) ^ (layer0_outputs[2150]);
    assign outputs[7290] = layer0_outputs[2931];
    assign outputs[7291] = (layer0_outputs[1429]) ^ (layer0_outputs[3718]);
    assign outputs[7292] = (layer0_outputs[4372]) & ~(layer0_outputs[2081]);
    assign outputs[7293] = (layer0_outputs[626]) ^ (layer0_outputs[3390]);
    assign outputs[7294] = (layer0_outputs[2917]) ^ (layer0_outputs[2969]);
    assign outputs[7295] = (layer0_outputs[4276]) & ~(layer0_outputs[4751]);
    assign outputs[7296] = layer0_outputs[2051];
    assign outputs[7297] = layer0_outputs[225];
    assign outputs[7298] = ~(layer0_outputs[1205]);
    assign outputs[7299] = ~((layer0_outputs[7799]) | (layer0_outputs[3940]));
    assign outputs[7300] = (layer0_outputs[4247]) ^ (layer0_outputs[1428]);
    assign outputs[7301] = (layer0_outputs[6102]) ^ (layer0_outputs[7526]);
    assign outputs[7302] = ~((layer0_outputs[4074]) ^ (layer0_outputs[4016]));
    assign outputs[7303] = layer0_outputs[942];
    assign outputs[7304] = ~(layer0_outputs[7594]);
    assign outputs[7305] = ~(layer0_outputs[2316]);
    assign outputs[7306] = (layer0_outputs[2929]) ^ (layer0_outputs[7290]);
    assign outputs[7307] = (layer0_outputs[6438]) & (layer0_outputs[594]);
    assign outputs[7308] = (layer0_outputs[1631]) & ~(layer0_outputs[10024]);
    assign outputs[7309] = (layer0_outputs[7936]) & (layer0_outputs[3592]);
    assign outputs[7310] = layer0_outputs[3041];
    assign outputs[7311] = 1'b1;
    assign outputs[7312] = (layer0_outputs[1938]) ^ (layer0_outputs[4476]);
    assign outputs[7313] = layer0_outputs[3787];
    assign outputs[7314] = ~(layer0_outputs[4882]) | (layer0_outputs[6949]);
    assign outputs[7315] = layer0_outputs[2634];
    assign outputs[7316] = (layer0_outputs[9329]) & ~(layer0_outputs[3105]);
    assign outputs[7317] = ~((layer0_outputs[8111]) ^ (layer0_outputs[4706]));
    assign outputs[7318] = layer0_outputs[1198];
    assign outputs[7319] = ~(layer0_outputs[2712]);
    assign outputs[7320] = (layer0_outputs[605]) & (layer0_outputs[9444]);
    assign outputs[7321] = layer0_outputs[2434];
    assign outputs[7322] = (layer0_outputs[10226]) & ~(layer0_outputs[7953]);
    assign outputs[7323] = layer0_outputs[7337];
    assign outputs[7324] = ~((layer0_outputs[2136]) ^ (layer0_outputs[1724]));
    assign outputs[7325] = ~(layer0_outputs[2186]);
    assign outputs[7326] = ~((layer0_outputs[3796]) ^ (layer0_outputs[6403]));
    assign outputs[7327] = ~(layer0_outputs[1529]);
    assign outputs[7328] = layer0_outputs[3824];
    assign outputs[7329] = ~(layer0_outputs[1764]);
    assign outputs[7330] = ~(layer0_outputs[1143]);
    assign outputs[7331] = ~((layer0_outputs[878]) ^ (layer0_outputs[9498]));
    assign outputs[7332] = ~(layer0_outputs[5470]) | (layer0_outputs[1918]);
    assign outputs[7333] = ~(layer0_outputs[2489]);
    assign outputs[7334] = (layer0_outputs[4732]) ^ (layer0_outputs[7105]);
    assign outputs[7335] = ~((layer0_outputs[3774]) ^ (layer0_outputs[2403]));
    assign outputs[7336] = ~(layer0_outputs[7172]);
    assign outputs[7337] = ~(layer0_outputs[7318]) | (layer0_outputs[4083]);
    assign outputs[7338] = ~(layer0_outputs[3462]);
    assign outputs[7339] = (layer0_outputs[8983]) & (layer0_outputs[8252]);
    assign outputs[7340] = (layer0_outputs[8191]) & ~(layer0_outputs[4574]);
    assign outputs[7341] = ~(layer0_outputs[9292]) | (layer0_outputs[6316]);
    assign outputs[7342] = ~((layer0_outputs[3869]) | (layer0_outputs[803]));
    assign outputs[7343] = ~(layer0_outputs[1649]);
    assign outputs[7344] = (layer0_outputs[7323]) & ~(layer0_outputs[2371]);
    assign outputs[7345] = ~((layer0_outputs[760]) ^ (layer0_outputs[1321]));
    assign outputs[7346] = ~(layer0_outputs[5794]) | (layer0_outputs[9183]);
    assign outputs[7347] = layer0_outputs[9159];
    assign outputs[7348] = ~((layer0_outputs[8333]) | (layer0_outputs[6208]));
    assign outputs[7349] = ~((layer0_outputs[6362]) ^ (layer0_outputs[2988]));
    assign outputs[7350] = (layer0_outputs[5824]) & ~(layer0_outputs[5523]);
    assign outputs[7351] = layer0_outputs[2297];
    assign outputs[7352] = ~((layer0_outputs[3281]) | (layer0_outputs[1438]));
    assign outputs[7353] = layer0_outputs[1342];
    assign outputs[7354] = (layer0_outputs[2854]) ^ (layer0_outputs[7964]);
    assign outputs[7355] = (layer0_outputs[5750]) & ~(layer0_outputs[9630]);
    assign outputs[7356] = layer0_outputs[8383];
    assign outputs[7357] = (layer0_outputs[8090]) & ~(layer0_outputs[5258]);
    assign outputs[7358] = (layer0_outputs[7425]) | (layer0_outputs[508]);
    assign outputs[7359] = ~((layer0_outputs[8558]) ^ (layer0_outputs[5114]));
    assign outputs[7360] = ~((layer0_outputs[8134]) ^ (layer0_outputs[1098]));
    assign outputs[7361] = (layer0_outputs[1227]) & ~(layer0_outputs[345]);
    assign outputs[7362] = (layer0_outputs[8829]) ^ (layer0_outputs[2214]);
    assign outputs[7363] = (layer0_outputs[1756]) & (layer0_outputs[3142]);
    assign outputs[7364] = layer0_outputs[6671];
    assign outputs[7365] = layer0_outputs[9348];
    assign outputs[7366] = (layer0_outputs[9991]) ^ (layer0_outputs[3467]);
    assign outputs[7367] = layer0_outputs[9992];
    assign outputs[7368] = ~(layer0_outputs[5439]);
    assign outputs[7369] = (layer0_outputs[7300]) & ~(layer0_outputs[206]);
    assign outputs[7370] = layer0_outputs[6846];
    assign outputs[7371] = ~(layer0_outputs[3597]);
    assign outputs[7372] = (layer0_outputs[1980]) & (layer0_outputs[7921]);
    assign outputs[7373] = ~(layer0_outputs[1497]) | (layer0_outputs[5901]);
    assign outputs[7374] = (layer0_outputs[5442]) & (layer0_outputs[4633]);
    assign outputs[7375] = layer0_outputs[6422];
    assign outputs[7376] = ~(layer0_outputs[419]) | (layer0_outputs[2497]);
    assign outputs[7377] = ~((layer0_outputs[5320]) | (layer0_outputs[1119]));
    assign outputs[7378] = layer0_outputs[9329];
    assign outputs[7379] = ~(layer0_outputs[8114]);
    assign outputs[7380] = ~((layer0_outputs[6062]) ^ (layer0_outputs[5822]));
    assign outputs[7381] = layer0_outputs[5520];
    assign outputs[7382] = ~(layer0_outputs[8628]) | (layer0_outputs[10180]);
    assign outputs[7383] = (layer0_outputs[1691]) & ~(layer0_outputs[8389]);
    assign outputs[7384] = ~(layer0_outputs[7785]);
    assign outputs[7385] = ~((layer0_outputs[6752]) ^ (layer0_outputs[7991]));
    assign outputs[7386] = ~(layer0_outputs[785]);
    assign outputs[7387] = (layer0_outputs[9320]) ^ (layer0_outputs[3989]);
    assign outputs[7388] = ~(layer0_outputs[3271]);
    assign outputs[7389] = (layer0_outputs[9429]) & ~(layer0_outputs[4879]);
    assign outputs[7390] = ~(layer0_outputs[1465]);
    assign outputs[7391] = layer0_outputs[9654];
    assign outputs[7392] = ~(layer0_outputs[9266]);
    assign outputs[7393] = (layer0_outputs[4624]) & ~(layer0_outputs[2523]);
    assign outputs[7394] = (layer0_outputs[2134]) ^ (layer0_outputs[7956]);
    assign outputs[7395] = (layer0_outputs[2047]) & ~(layer0_outputs[5053]);
    assign outputs[7396] = (layer0_outputs[6758]) | (layer0_outputs[1112]);
    assign outputs[7397] = (layer0_outputs[8732]) ^ (layer0_outputs[5124]);
    assign outputs[7398] = ~((layer0_outputs[539]) ^ (layer0_outputs[2757]));
    assign outputs[7399] = (layer0_outputs[8553]) & (layer0_outputs[2839]);
    assign outputs[7400] = ~((layer0_outputs[8617]) ^ (layer0_outputs[5982]));
    assign outputs[7401] = layer0_outputs[9695];
    assign outputs[7402] = ~(layer0_outputs[2773]);
    assign outputs[7403] = ~((layer0_outputs[528]) | (layer0_outputs[8953]));
    assign outputs[7404] = ~((layer0_outputs[1807]) ^ (layer0_outputs[263]));
    assign outputs[7405] = (layer0_outputs[6655]) & ~(layer0_outputs[573]);
    assign outputs[7406] = (layer0_outputs[7162]) ^ (layer0_outputs[8369]);
    assign outputs[7407] = (layer0_outputs[4871]) & ~(layer0_outputs[992]);
    assign outputs[7408] = ~((layer0_outputs[2140]) ^ (layer0_outputs[5743]));
    assign outputs[7409] = ~(layer0_outputs[7439]);
    assign outputs[7410] = (layer0_outputs[3663]) & (layer0_outputs[9772]);
    assign outputs[7411] = ~((layer0_outputs[7199]) ^ (layer0_outputs[8949]));
    assign outputs[7412] = (layer0_outputs[476]) & ~(layer0_outputs[4115]);
    assign outputs[7413] = layer0_outputs[5095];
    assign outputs[7414] = ~(layer0_outputs[46]);
    assign outputs[7415] = ~((layer0_outputs[2363]) ^ (layer0_outputs[10237]));
    assign outputs[7416] = ~((layer0_outputs[6614]) ^ (layer0_outputs[8481]));
    assign outputs[7417] = ~(layer0_outputs[7730]);
    assign outputs[7418] = ~((layer0_outputs[5806]) | (layer0_outputs[3498]));
    assign outputs[7419] = (layer0_outputs[1316]) & ~(layer0_outputs[7121]);
    assign outputs[7420] = layer0_outputs[7848];
    assign outputs[7421] = (layer0_outputs[2112]) & ~(layer0_outputs[2586]);
    assign outputs[7422] = ~((layer0_outputs[3695]) | (layer0_outputs[843]));
    assign outputs[7423] = (layer0_outputs[3145]) | (layer0_outputs[8911]);
    assign outputs[7424] = layer0_outputs[5995];
    assign outputs[7425] = (layer0_outputs[1661]) & ~(layer0_outputs[3166]);
    assign outputs[7426] = (layer0_outputs[9306]) & ~(layer0_outputs[3903]);
    assign outputs[7427] = (layer0_outputs[5123]) & (layer0_outputs[9613]);
    assign outputs[7428] = ~(layer0_outputs[4950]);
    assign outputs[7429] = (layer0_outputs[1180]) & (layer0_outputs[8491]);
    assign outputs[7430] = ~((layer0_outputs[865]) ^ (layer0_outputs[3681]));
    assign outputs[7431] = (layer0_outputs[8033]) ^ (layer0_outputs[4486]);
    assign outputs[7432] = ~(layer0_outputs[4044]);
    assign outputs[7433] = ~(layer0_outputs[3677]);
    assign outputs[7434] = layer0_outputs[1101];
    assign outputs[7435] = layer0_outputs[6161];
    assign outputs[7436] = (layer0_outputs[7167]) ^ (layer0_outputs[8740]);
    assign outputs[7437] = layer0_outputs[5597];
    assign outputs[7438] = layer0_outputs[8657];
    assign outputs[7439] = ~(layer0_outputs[6965]);
    assign outputs[7440] = ~((layer0_outputs[9923]) ^ (layer0_outputs[1151]));
    assign outputs[7441] = ~((layer0_outputs[9522]) ^ (layer0_outputs[8070]));
    assign outputs[7442] = (layer0_outputs[1121]) & ~(layer0_outputs[3042]);
    assign outputs[7443] = ~((layer0_outputs[1696]) | (layer0_outputs[7150]));
    assign outputs[7444] = ~((layer0_outputs[2750]) ^ (layer0_outputs[4893]));
    assign outputs[7445] = ~(layer0_outputs[8431]);
    assign outputs[7446] = layer0_outputs[7383];
    assign outputs[7447] = (layer0_outputs[614]) ^ (layer0_outputs[1057]);
    assign outputs[7448] = ~((layer0_outputs[9660]) & (layer0_outputs[6207]));
    assign outputs[7449] = ~(layer0_outputs[4494]);
    assign outputs[7450] = (layer0_outputs[3784]) & (layer0_outputs[9221]);
    assign outputs[7451] = ~(layer0_outputs[114]);
    assign outputs[7452] = ~((layer0_outputs[222]) | (layer0_outputs[318]));
    assign outputs[7453] = (layer0_outputs[3747]) & (layer0_outputs[8438]);
    assign outputs[7454] = layer0_outputs[4964];
    assign outputs[7455] = (layer0_outputs[1962]) ^ (layer0_outputs[3592]);
    assign outputs[7456] = ~(layer0_outputs[7970]);
    assign outputs[7457] = (layer0_outputs[6330]) ^ (layer0_outputs[3424]);
    assign outputs[7458] = (layer0_outputs[2920]) & (layer0_outputs[2591]);
    assign outputs[7459] = ~(layer0_outputs[8356]);
    assign outputs[7460] = ~((layer0_outputs[2663]) | (layer0_outputs[7460]));
    assign outputs[7461] = ~(layer0_outputs[8399]);
    assign outputs[7462] = ~((layer0_outputs[8308]) | (layer0_outputs[9393]));
    assign outputs[7463] = (layer0_outputs[9705]) & ~(layer0_outputs[9008]);
    assign outputs[7464] = ~(layer0_outputs[8838]);
    assign outputs[7465] = (layer0_outputs[732]) & (layer0_outputs[8124]);
    assign outputs[7466] = layer0_outputs[4263];
    assign outputs[7467] = (layer0_outputs[8428]) | (layer0_outputs[3014]);
    assign outputs[7468] = layer0_outputs[1130];
    assign outputs[7469] = (layer0_outputs[293]) & ~(layer0_outputs[8191]);
    assign outputs[7470] = (layer0_outputs[6213]) ^ (layer0_outputs[3851]);
    assign outputs[7471] = (layer0_outputs[5755]) & ~(layer0_outputs[9260]);
    assign outputs[7472] = layer0_outputs[6091];
    assign outputs[7473] = ~((layer0_outputs[3311]) ^ (layer0_outputs[6174]));
    assign outputs[7474] = layer0_outputs[9680];
    assign outputs[7475] = (layer0_outputs[7662]) ^ (layer0_outputs[3503]);
    assign outputs[7476] = layer0_outputs[8324];
    assign outputs[7477] = ~((layer0_outputs[8535]) | (layer0_outputs[4876]));
    assign outputs[7478] = ~((layer0_outputs[9777]) & (layer0_outputs[7999]));
    assign outputs[7479] = (layer0_outputs[3781]) & ~(layer0_outputs[3682]);
    assign outputs[7480] = (layer0_outputs[8529]) ^ (layer0_outputs[4774]);
    assign outputs[7481] = ~((layer0_outputs[1327]) ^ (layer0_outputs[5010]));
    assign outputs[7482] = layer0_outputs[7253];
    assign outputs[7483] = ~((layer0_outputs[9068]) ^ (layer0_outputs[1023]));
    assign outputs[7484] = ~(layer0_outputs[2577]);
    assign outputs[7485] = (layer0_outputs[7573]) & ~(layer0_outputs[8442]);
    assign outputs[7486] = (layer0_outputs[8404]) & (layer0_outputs[7479]);
    assign outputs[7487] = (layer0_outputs[2345]) & ~(layer0_outputs[4288]);
    assign outputs[7488] = ~((layer0_outputs[8166]) ^ (layer0_outputs[5569]));
    assign outputs[7489] = ~(layer0_outputs[9387]);
    assign outputs[7490] = layer0_outputs[938];
    assign outputs[7491] = ~(layer0_outputs[5625]) | (layer0_outputs[8384]);
    assign outputs[7492] = (layer0_outputs[944]) ^ (layer0_outputs[6497]);
    assign outputs[7493] = layer0_outputs[5019];
    assign outputs[7494] = ~(layer0_outputs[3128]);
    assign outputs[7495] = ~((layer0_outputs[8220]) ^ (layer0_outputs[2790]));
    assign outputs[7496] = ~(layer0_outputs[7553]);
    assign outputs[7497] = (layer0_outputs[2617]) | (layer0_outputs[3639]);
    assign outputs[7498] = ~((layer0_outputs[4043]) | (layer0_outputs[7152]));
    assign outputs[7499] = ~(layer0_outputs[888]);
    assign outputs[7500] = (layer0_outputs[8935]) ^ (layer0_outputs[10141]);
    assign outputs[7501] = ~((layer0_outputs[4235]) ^ (layer0_outputs[6553]));
    assign outputs[7502] = layer0_outputs[7494];
    assign outputs[7503] = (layer0_outputs[7831]) & ~(layer0_outputs[7547]);
    assign outputs[7504] = ~(layer0_outputs[8705]);
    assign outputs[7505] = (layer0_outputs[1245]) ^ (layer0_outputs[6582]);
    assign outputs[7506] = ~(layer0_outputs[7057]);
    assign outputs[7507] = layer0_outputs[7165];
    assign outputs[7508] = 1'b0;
    assign outputs[7509] = ~(layer0_outputs[7572]);
    assign outputs[7510] = layer0_outputs[8086];
    assign outputs[7511] = layer0_outputs[9220];
    assign outputs[7512] = (layer0_outputs[2881]) & ~(layer0_outputs[4311]);
    assign outputs[7513] = (layer0_outputs[426]) & ~(layer0_outputs[3685]);
    assign outputs[7514] = ~((layer0_outputs[1678]) | (layer0_outputs[7529]));
    assign outputs[7515] = layer0_outputs[7686];
    assign outputs[7516] = ~((layer0_outputs[2889]) ^ (layer0_outputs[6621]));
    assign outputs[7517] = (layer0_outputs[5012]) | (layer0_outputs[1648]);
    assign outputs[7518] = ~((layer0_outputs[6050]) ^ (layer0_outputs[5769]));
    assign outputs[7519] = ~(layer0_outputs[5732]);
    assign outputs[7520] = ~((layer0_outputs[4228]) ^ (layer0_outputs[700]));
    assign outputs[7521] = (layer0_outputs[9221]) ^ (layer0_outputs[3073]);
    assign outputs[7522] = ~((layer0_outputs[450]) ^ (layer0_outputs[712]));
    assign outputs[7523] = (layer0_outputs[111]) & ~(layer0_outputs[2474]);
    assign outputs[7524] = ~((layer0_outputs[1176]) ^ (layer0_outputs[4935]));
    assign outputs[7525] = ~(layer0_outputs[9143]);
    assign outputs[7526] = ~(layer0_outputs[7989]);
    assign outputs[7527] = ~((layer0_outputs[9560]) & (layer0_outputs[9849]));
    assign outputs[7528] = ~(layer0_outputs[2731]);
    assign outputs[7529] = ~(layer0_outputs[1107]);
    assign outputs[7530] = ~(layer0_outputs[1658]);
    assign outputs[7531] = (layer0_outputs[703]) & ~(layer0_outputs[9953]);
    assign outputs[7532] = (layer0_outputs[1521]) ^ (layer0_outputs[6412]);
    assign outputs[7533] = ~((layer0_outputs[5515]) | (layer0_outputs[3810]));
    assign outputs[7534] = (layer0_outputs[315]) & ~(layer0_outputs[7142]);
    assign outputs[7535] = ~((layer0_outputs[4378]) ^ (layer0_outputs[3475]));
    assign outputs[7536] = (layer0_outputs[4998]) & ~(layer0_outputs[7913]);
    assign outputs[7537] = ~(layer0_outputs[1039]);
    assign outputs[7538] = layer0_outputs[1868];
    assign outputs[7539] = ~(layer0_outputs[5349]);
    assign outputs[7540] = ~(layer0_outputs[4565]) | (layer0_outputs[3625]);
    assign outputs[7541] = layer0_outputs[6870];
    assign outputs[7542] = (layer0_outputs[4518]) & (layer0_outputs[2870]);
    assign outputs[7543] = layer0_outputs[6961];
    assign outputs[7544] = layer0_outputs[5879];
    assign outputs[7545] = (layer0_outputs[5543]) | (layer0_outputs[2443]);
    assign outputs[7546] = ~((layer0_outputs[1049]) ^ (layer0_outputs[4984]));
    assign outputs[7547] = layer0_outputs[2847];
    assign outputs[7548] = (layer0_outputs[2619]) & ~(layer0_outputs[3604]);
    assign outputs[7549] = ~((layer0_outputs[1589]) ^ (layer0_outputs[8820]));
    assign outputs[7550] = ~(layer0_outputs[8414]);
    assign outputs[7551] = layer0_outputs[1730];
    assign outputs[7552] = ~((layer0_outputs[2778]) ^ (layer0_outputs[3230]));
    assign outputs[7553] = ~((layer0_outputs[9882]) | (layer0_outputs[6163]));
    assign outputs[7554] = (layer0_outputs[10075]) & ~(layer0_outputs[6657]);
    assign outputs[7555] = ~(layer0_outputs[5639]);
    assign outputs[7556] = (layer0_outputs[6726]) ^ (layer0_outputs[9192]);
    assign outputs[7557] = (layer0_outputs[2048]) ^ (layer0_outputs[2429]);
    assign outputs[7558] = layer0_outputs[5895];
    assign outputs[7559] = (layer0_outputs[1788]) ^ (layer0_outputs[7371]);
    assign outputs[7560] = ~(layer0_outputs[4851]);
    assign outputs[7561] = ~((layer0_outputs[3916]) ^ (layer0_outputs[10112]));
    assign outputs[7562] = ~((layer0_outputs[2910]) & (layer0_outputs[8137]));
    assign outputs[7563] = (layer0_outputs[7659]) ^ (layer0_outputs[7830]);
    assign outputs[7564] = (layer0_outputs[4743]) ^ (layer0_outputs[6282]);
    assign outputs[7565] = ~(layer0_outputs[4151]);
    assign outputs[7566] = ~((layer0_outputs[7940]) ^ (layer0_outputs[850]));
    assign outputs[7567] = layer0_outputs[7123];
    assign outputs[7568] = ~(layer0_outputs[9053]);
    assign outputs[7569] = (layer0_outputs[5327]) & ~(layer0_outputs[4181]);
    assign outputs[7570] = ~(layer0_outputs[1311]);
    assign outputs[7571] = ~((layer0_outputs[9455]) & (layer0_outputs[8978]));
    assign outputs[7572] = ~(layer0_outputs[947]);
    assign outputs[7573] = layer0_outputs[9451];
    assign outputs[7574] = (layer0_outputs[398]) ^ (layer0_outputs[9606]);
    assign outputs[7575] = (layer0_outputs[8459]) | (layer0_outputs[608]);
    assign outputs[7576] = (layer0_outputs[5166]) & ~(layer0_outputs[7992]);
    assign outputs[7577] = layer0_outputs[7478];
    assign outputs[7578] = ~((layer0_outputs[5115]) ^ (layer0_outputs[6104]));
    assign outputs[7579] = ~(layer0_outputs[193]);
    assign outputs[7580] = (layer0_outputs[9334]) & (layer0_outputs[4398]);
    assign outputs[7581] = ~((layer0_outputs[10156]) & (layer0_outputs[8863]));
    assign outputs[7582] = ~(layer0_outputs[6269]);
    assign outputs[7583] = ~(layer0_outputs[9550]) | (layer0_outputs[9731]);
    assign outputs[7584] = layer0_outputs[718];
    assign outputs[7585] = layer0_outputs[6318];
    assign outputs[7586] = (layer0_outputs[4735]) & (layer0_outputs[3834]);
    assign outputs[7587] = (layer0_outputs[6188]) ^ (layer0_outputs[3987]);
    assign outputs[7588] = ~((layer0_outputs[211]) ^ (layer0_outputs[3029]));
    assign outputs[7589] = ~(layer0_outputs[2694]);
    assign outputs[7590] = layer0_outputs[3982];
    assign outputs[7591] = ~((layer0_outputs[6012]) ^ (layer0_outputs[8716]));
    assign outputs[7592] = (layer0_outputs[2249]) & (layer0_outputs[4447]);
    assign outputs[7593] = ~(layer0_outputs[9174]);
    assign outputs[7594] = ~((layer0_outputs[9455]) ^ (layer0_outputs[9733]));
    assign outputs[7595] = ~(layer0_outputs[7464]);
    assign outputs[7596] = ~(layer0_outputs[1897]);
    assign outputs[7597] = (layer0_outputs[6621]) & ~(layer0_outputs[1312]);
    assign outputs[7598] = ~(layer0_outputs[8555]);
    assign outputs[7599] = (layer0_outputs[1760]) & ~(layer0_outputs[3161]);
    assign outputs[7600] = (layer0_outputs[8301]) ^ (layer0_outputs[2715]);
    assign outputs[7601] = ~((layer0_outputs[4022]) ^ (layer0_outputs[2813]));
    assign outputs[7602] = ~(layer0_outputs[9781]);
    assign outputs[7603] = ~(layer0_outputs[10003]) | (layer0_outputs[8156]);
    assign outputs[7604] = ~((layer0_outputs[4853]) ^ (layer0_outputs[6053]));
    assign outputs[7605] = ~(layer0_outputs[8734]);
    assign outputs[7606] = (layer0_outputs[578]) ^ (layer0_outputs[204]);
    assign outputs[7607] = ~(layer0_outputs[7532]);
    assign outputs[7608] = (layer0_outputs[3299]) | (layer0_outputs[6253]);
    assign outputs[7609] = (layer0_outputs[3104]) & ~(layer0_outputs[4349]);
    assign outputs[7610] = ~(layer0_outputs[9523]);
    assign outputs[7611] = ~(layer0_outputs[9109]) | (layer0_outputs[5655]);
    assign outputs[7612] = (layer0_outputs[2178]) & (layer0_outputs[2505]);
    assign outputs[7613] = ~(layer0_outputs[6016]);
    assign outputs[7614] = ~(layer0_outputs[9559]) | (layer0_outputs[8]);
    assign outputs[7615] = (layer0_outputs[7531]) ^ (layer0_outputs[1627]);
    assign outputs[7616] = ~((layer0_outputs[10141]) | (layer0_outputs[8402]));
    assign outputs[7617] = ~((layer0_outputs[9666]) & (layer0_outputs[2697]));
    assign outputs[7618] = (layer0_outputs[9656]) & (layer0_outputs[8896]);
    assign outputs[7619] = layer0_outputs[3082];
    assign outputs[7620] = layer0_outputs[8764];
    assign outputs[7621] = ~((layer0_outputs[9020]) ^ (layer0_outputs[6175]));
    assign outputs[7622] = (layer0_outputs[2222]) & (layer0_outputs[4047]);
    assign outputs[7623] = layer0_outputs[2286];
    assign outputs[7624] = ~(layer0_outputs[6906]) | (layer0_outputs[5645]);
    assign outputs[7625] = ~((layer0_outputs[10195]) ^ (layer0_outputs[5209]));
    assign outputs[7626] = layer0_outputs[1227];
    assign outputs[7627] = (layer0_outputs[2343]) & ~(layer0_outputs[840]);
    assign outputs[7628] = layer0_outputs[2297];
    assign outputs[7629] = layer0_outputs[2006];
    assign outputs[7630] = (layer0_outputs[8726]) & ~(layer0_outputs[9597]);
    assign outputs[7631] = (layer0_outputs[2035]) & (layer0_outputs[5648]);
    assign outputs[7632] = (layer0_outputs[625]) & ~(layer0_outputs[8205]);
    assign outputs[7633] = (layer0_outputs[6582]) & (layer0_outputs[7993]);
    assign outputs[7634] = ~(layer0_outputs[8375]);
    assign outputs[7635] = (layer0_outputs[2689]) & ~(layer0_outputs[5495]);
    assign outputs[7636] = ~((layer0_outputs[3245]) ^ (layer0_outputs[6137]));
    assign outputs[7637] = ~(layer0_outputs[7907]);
    assign outputs[7638] = (layer0_outputs[995]) & (layer0_outputs[2291]);
    assign outputs[7639] = ~((layer0_outputs[8361]) ^ (layer0_outputs[5642]));
    assign outputs[7640] = ~(layer0_outputs[4400]);
    assign outputs[7641] = ~(layer0_outputs[2336]);
    assign outputs[7642] = (layer0_outputs[1127]) ^ (layer0_outputs[8984]);
    assign outputs[7643] = layer0_outputs[8932];
    assign outputs[7644] = ~(layer0_outputs[9446]);
    assign outputs[7645] = layer0_outputs[2808];
    assign outputs[7646] = (layer0_outputs[9154]) & ~(layer0_outputs[10052]);
    assign outputs[7647] = (layer0_outputs[7620]) & (layer0_outputs[3800]);
    assign outputs[7648] = (layer0_outputs[8203]) & ~(layer0_outputs[6522]);
    assign outputs[7649] = ~(layer0_outputs[4239]) | (layer0_outputs[6620]);
    assign outputs[7650] = ~((layer0_outputs[3248]) | (layer0_outputs[4019]));
    assign outputs[7651] = ~((layer0_outputs[7317]) & (layer0_outputs[414]));
    assign outputs[7652] = (layer0_outputs[3289]) | (layer0_outputs[4831]);
    assign outputs[7653] = ~((layer0_outputs[6866]) ^ (layer0_outputs[3464]));
    assign outputs[7654] = ~(layer0_outputs[6789]) | (layer0_outputs[6353]);
    assign outputs[7655] = layer0_outputs[3494];
    assign outputs[7656] = (layer0_outputs[7045]) & ~(layer0_outputs[6847]);
    assign outputs[7657] = layer0_outputs[2543];
    assign outputs[7658] = ~(layer0_outputs[2641]);
    assign outputs[7659] = ~(layer0_outputs[4654]);
    assign outputs[7660] = layer0_outputs[9060];
    assign outputs[7661] = (layer0_outputs[2924]) | (layer0_outputs[6632]);
    assign outputs[7662] = ~(layer0_outputs[1462]);
    assign outputs[7663] = (layer0_outputs[1599]) ^ (layer0_outputs[6339]);
    assign outputs[7664] = ~((layer0_outputs[8580]) | (layer0_outputs[497]));
    assign outputs[7665] = layer0_outputs[548];
    assign outputs[7666] = (layer0_outputs[1846]) & (layer0_outputs[8202]);
    assign outputs[7667] = layer0_outputs[9860];
    assign outputs[7668] = (layer0_outputs[1545]) & ~(layer0_outputs[9276]);
    assign outputs[7669] = ~(layer0_outputs[9193]);
    assign outputs[7670] = ~((layer0_outputs[760]) ^ (layer0_outputs[5783]));
    assign outputs[7671] = layer0_outputs[6107];
    assign outputs[7672] = ~((layer0_outputs[1604]) ^ (layer0_outputs[5135]));
    assign outputs[7673] = ~(layer0_outputs[140]);
    assign outputs[7674] = layer0_outputs[1030];
    assign outputs[7675] = (layer0_outputs[6466]) & ~(layer0_outputs[3149]);
    assign outputs[7676] = ~((layer0_outputs[7345]) | (layer0_outputs[449]));
    assign outputs[7677] = ~(layer0_outputs[7939]);
    assign outputs[7678] = (layer0_outputs[6965]) ^ (layer0_outputs[2899]);
    assign outputs[7679] = layer0_outputs[4261];
    assign outputs[7680] = ~((layer0_outputs[901]) | (layer0_outputs[8047]));
    assign outputs[7681] = ~(layer0_outputs[462]) | (layer0_outputs[9606]);
    assign outputs[7682] = ~(layer0_outputs[5929]);
    assign outputs[7683] = (layer0_outputs[3913]) | (layer0_outputs[5497]);
    assign outputs[7684] = ~(layer0_outputs[3454]);
    assign outputs[7685] = layer0_outputs[7028];
    assign outputs[7686] = (layer0_outputs[8017]) & ~(layer0_outputs[599]);
    assign outputs[7687] = ~((layer0_outputs[264]) ^ (layer0_outputs[7264]));
    assign outputs[7688] = (layer0_outputs[9869]) & ~(layer0_outputs[7671]);
    assign outputs[7689] = ~(layer0_outputs[3686]);
    assign outputs[7690] = (layer0_outputs[4629]) & ~(layer0_outputs[5932]);
    assign outputs[7691] = ~((layer0_outputs[10196]) ^ (layer0_outputs[3228]));
    assign outputs[7692] = ~((layer0_outputs[3519]) | (layer0_outputs[5871]));
    assign outputs[7693] = ~(layer0_outputs[8164]);
    assign outputs[7694] = ~((layer0_outputs[5556]) ^ (layer0_outputs[765]));
    assign outputs[7695] = layer0_outputs[1088];
    assign outputs[7696] = ~(layer0_outputs[1514]);
    assign outputs[7697] = ~(layer0_outputs[9310]);
    assign outputs[7698] = ~((layer0_outputs[3899]) ^ (layer0_outputs[2392]));
    assign outputs[7699] = ~(layer0_outputs[9584]);
    assign outputs[7700] = (layer0_outputs[8888]) & ~(layer0_outputs[5381]);
    assign outputs[7701] = layer0_outputs[5778];
    assign outputs[7702] = ~((layer0_outputs[118]) & (layer0_outputs[4939]));
    assign outputs[7703] = ~(layer0_outputs[6774]) | (layer0_outputs[6097]);
    assign outputs[7704] = layer0_outputs[74];
    assign outputs[7705] = ~((layer0_outputs[3153]) & (layer0_outputs[5069]));
    assign outputs[7706] = (layer0_outputs[4993]) | (layer0_outputs[1184]);
    assign outputs[7707] = ~(layer0_outputs[8907]);
    assign outputs[7708] = layer0_outputs[7503];
    assign outputs[7709] = ~(layer0_outputs[8051]);
    assign outputs[7710] = ~(layer0_outputs[4314]);
    assign outputs[7711] = ~((layer0_outputs[1183]) ^ (layer0_outputs[9082]));
    assign outputs[7712] = (layer0_outputs[3043]) ^ (layer0_outputs[2522]);
    assign outputs[7713] = layer0_outputs[7102];
    assign outputs[7714] = (layer0_outputs[6168]) & (layer0_outputs[7265]);
    assign outputs[7715] = ~((layer0_outputs[8021]) ^ (layer0_outputs[3217]));
    assign outputs[7716] = (layer0_outputs[5651]) & ~(layer0_outputs[9392]);
    assign outputs[7717] = ~(layer0_outputs[1031]);
    assign outputs[7718] = ~(layer0_outputs[4856]);
    assign outputs[7719] = layer0_outputs[8479];
    assign outputs[7720] = ~((layer0_outputs[2034]) & (layer0_outputs[7264]));
    assign outputs[7721] = layer0_outputs[952];
    assign outputs[7722] = (layer0_outputs[9013]) | (layer0_outputs[6249]);
    assign outputs[7723] = ~(layer0_outputs[6897]);
    assign outputs[7724] = ~(layer0_outputs[6061]);
    assign outputs[7725] = (layer0_outputs[4037]) ^ (layer0_outputs[3823]);
    assign outputs[7726] = ~((layer0_outputs[7724]) | (layer0_outputs[296]));
    assign outputs[7727] = ~(layer0_outputs[2703]) | (layer0_outputs[2380]);
    assign outputs[7728] = ~(layer0_outputs[7249]);
    assign outputs[7729] = layer0_outputs[10076];
    assign outputs[7730] = ~(layer0_outputs[321]) | (layer0_outputs[9603]);
    assign outputs[7731] = (layer0_outputs[9332]) & (layer0_outputs[621]);
    assign outputs[7732] = ~(layer0_outputs[7272]);
    assign outputs[7733] = ~(layer0_outputs[9782]) | (layer0_outputs[2922]);
    assign outputs[7734] = ~(layer0_outputs[8304]);
    assign outputs[7735] = (layer0_outputs[8976]) & ~(layer0_outputs[4524]);
    assign outputs[7736] = ~((layer0_outputs[698]) | (layer0_outputs[2549]));
    assign outputs[7737] = (layer0_outputs[5569]) ^ (layer0_outputs[8421]);
    assign outputs[7738] = (layer0_outputs[6149]) & ~(layer0_outputs[830]);
    assign outputs[7739] = ~(layer0_outputs[3920]);
    assign outputs[7740] = ~(layer0_outputs[3433]);
    assign outputs[7741] = ~((layer0_outputs[7710]) ^ (layer0_outputs[1612]));
    assign outputs[7742] = layer0_outputs[9789];
    assign outputs[7743] = (layer0_outputs[7600]) ^ (layer0_outputs[726]);
    assign outputs[7744] = ~((layer0_outputs[9819]) ^ (layer0_outputs[4371]));
    assign outputs[7745] = (layer0_outputs[1576]) & ~(layer0_outputs[5868]);
    assign outputs[7746] = ~(layer0_outputs[4662]);
    assign outputs[7747] = layer0_outputs[4439];
    assign outputs[7748] = (layer0_outputs[4511]) ^ (layer0_outputs[6378]);
    assign outputs[7749] = layer0_outputs[6155];
    assign outputs[7750] = (layer0_outputs[7362]) & (layer0_outputs[8674]);
    assign outputs[7751] = ~(layer0_outputs[7429]);
    assign outputs[7752] = (layer0_outputs[10030]) & (layer0_outputs[7213]);
    assign outputs[7753] = layer0_outputs[43];
    assign outputs[7754] = layer0_outputs[8751];
    assign outputs[7755] = layer0_outputs[7554];
    assign outputs[7756] = ~((layer0_outputs[4111]) ^ (layer0_outputs[3951]));
    assign outputs[7757] = layer0_outputs[7116];
    assign outputs[7758] = (layer0_outputs[197]) & ~(layer0_outputs[1901]);
    assign outputs[7759] = (layer0_outputs[4075]) & (layer0_outputs[784]);
    assign outputs[7760] = (layer0_outputs[4482]) ^ (layer0_outputs[2251]);
    assign outputs[7761] = (layer0_outputs[7208]) ^ (layer0_outputs[6725]);
    assign outputs[7762] = ~(layer0_outputs[6000]) | (layer0_outputs[4490]);
    assign outputs[7763] = ~((layer0_outputs[9808]) ^ (layer0_outputs[1632]));
    assign outputs[7764] = (layer0_outputs[4906]) & (layer0_outputs[5468]);
    assign outputs[7765] = ~(layer0_outputs[800]);
    assign outputs[7766] = ~(layer0_outputs[4213]) | (layer0_outputs[3366]);
    assign outputs[7767] = ~(layer0_outputs[1768]);
    assign outputs[7768] = ~(layer0_outputs[4771]) | (layer0_outputs[4281]);
    assign outputs[7769] = ~((layer0_outputs[8945]) ^ (layer0_outputs[4385]));
    assign outputs[7770] = layer0_outputs[7669];
    assign outputs[7771] = ~((layer0_outputs[2275]) ^ (layer0_outputs[7417]));
    assign outputs[7772] = ~((layer0_outputs[5824]) | (layer0_outputs[9315]));
    assign outputs[7773] = (layer0_outputs[9293]) | (layer0_outputs[3640]);
    assign outputs[7774] = layer0_outputs[5764];
    assign outputs[7775] = ~(layer0_outputs[7874]);
    assign outputs[7776] = (layer0_outputs[4811]) & ~(layer0_outputs[1299]);
    assign outputs[7777] = (layer0_outputs[765]) & ~(layer0_outputs[8103]);
    assign outputs[7778] = ~((layer0_outputs[9592]) | (layer0_outputs[8051]));
    assign outputs[7779] = 1'b1;
    assign outputs[7780] = (layer0_outputs[6358]) & (layer0_outputs[9380]);
    assign outputs[7781] = ~(layer0_outputs[1874]);
    assign outputs[7782] = (layer0_outputs[831]) & ~(layer0_outputs[5818]);
    assign outputs[7783] = (layer0_outputs[80]) ^ (layer0_outputs[109]);
    assign outputs[7784] = layer0_outputs[10198];
    assign outputs[7785] = ~((layer0_outputs[5583]) | (layer0_outputs[7681]));
    assign outputs[7786] = (layer0_outputs[5079]) & (layer0_outputs[9648]);
    assign outputs[7787] = ~(layer0_outputs[5273]);
    assign outputs[7788] = (layer0_outputs[6828]) ^ (layer0_outputs[5514]);
    assign outputs[7789] = (layer0_outputs[1729]) & ~(layer0_outputs[988]);
    assign outputs[7790] = ~((layer0_outputs[664]) | (layer0_outputs[567]));
    assign outputs[7791] = ~(layer0_outputs[4551]);
    assign outputs[7792] = (layer0_outputs[8737]) & (layer0_outputs[197]);
    assign outputs[7793] = (layer0_outputs[540]) & ~(layer0_outputs[8066]);
    assign outputs[7794] = ~((layer0_outputs[1719]) & (layer0_outputs[5985]));
    assign outputs[7795] = (layer0_outputs[9198]) ^ (layer0_outputs[8237]);
    assign outputs[7796] = (layer0_outputs[7792]) & (layer0_outputs[2873]);
    assign outputs[7797] = ~((layer0_outputs[7553]) & (layer0_outputs[3373]));
    assign outputs[7798] = (layer0_outputs[3800]) & ~(layer0_outputs[8875]);
    assign outputs[7799] = layer0_outputs[3994];
    assign outputs[7800] = (layer0_outputs[7972]) & ~(layer0_outputs[9178]);
    assign outputs[7801] = layer0_outputs[8959];
    assign outputs[7802] = ~(layer0_outputs[3854]);
    assign outputs[7803] = (layer0_outputs[3562]) | (layer0_outputs[598]);
    assign outputs[7804] = ~((layer0_outputs[1585]) ^ (layer0_outputs[5776]));
    assign outputs[7805] = (layer0_outputs[9742]) & ~(layer0_outputs[7432]);
    assign outputs[7806] = (layer0_outputs[5540]) ^ (layer0_outputs[473]);
    assign outputs[7807] = ~(layer0_outputs[7420]);
    assign outputs[7808] = (layer0_outputs[6796]) ^ (layer0_outputs[3444]);
    assign outputs[7809] = layer0_outputs[5671];
    assign outputs[7810] = layer0_outputs[34];
    assign outputs[7811] = ~(layer0_outputs[5243]);
    assign outputs[7812] = ~(layer0_outputs[9625]);
    assign outputs[7813] = (layer0_outputs[540]) & ~(layer0_outputs[9152]);
    assign outputs[7814] = ~((layer0_outputs[6184]) ^ (layer0_outputs[7143]));
    assign outputs[7815] = layer0_outputs[9507];
    assign outputs[7816] = (layer0_outputs[9243]) & (layer0_outputs[7179]);
    assign outputs[7817] = layer0_outputs[4525];
    assign outputs[7818] = ~((layer0_outputs[8174]) & (layer0_outputs[3051]));
    assign outputs[7819] = layer0_outputs[3420];
    assign outputs[7820] = ~(layer0_outputs[1023]);
    assign outputs[7821] = ~((layer0_outputs[7859]) | (layer0_outputs[8342]));
    assign outputs[7822] = layer0_outputs[1336];
    assign outputs[7823] = layer0_outputs[1135];
    assign outputs[7824] = ~((layer0_outputs[9116]) & (layer0_outputs[4151]));
    assign outputs[7825] = ~(layer0_outputs[9340]);
    assign outputs[7826] = ~(layer0_outputs[5838]) | (layer0_outputs[3298]);
    assign outputs[7827] = layer0_outputs[4234];
    assign outputs[7828] = ~(layer0_outputs[6947]);
    assign outputs[7829] = (layer0_outputs[7721]) & ~(layer0_outputs[6881]);
    assign outputs[7830] = (layer0_outputs[9957]) & ~(layer0_outputs[6411]);
    assign outputs[7831] = ~(layer0_outputs[5792]) | (layer0_outputs[881]);
    assign outputs[7832] = ~(layer0_outputs[4048]);
    assign outputs[7833] = ~((layer0_outputs[3259]) | (layer0_outputs[2031]));
    assign outputs[7834] = layer0_outputs[7876];
    assign outputs[7835] = ~(layer0_outputs[1797]);
    assign outputs[7836] = (layer0_outputs[33]) & (layer0_outputs[3621]);
    assign outputs[7837] = 1'b0;
    assign outputs[7838] = ~(layer0_outputs[4034]) | (layer0_outputs[9268]);
    assign outputs[7839] = ~(layer0_outputs[3810]);
    assign outputs[7840] = ~((layer0_outputs[584]) ^ (layer0_outputs[3393]));
    assign outputs[7841] = ~(layer0_outputs[3582]) | (layer0_outputs[213]);
    assign outputs[7842] = (layer0_outputs[10232]) & ~(layer0_outputs[2115]);
    assign outputs[7843] = ~(layer0_outputs[8337]);
    assign outputs[7844] = (layer0_outputs[757]) ^ (layer0_outputs[9009]);
    assign outputs[7845] = ~(layer0_outputs[4819]);
    assign outputs[7846] = (layer0_outputs[2319]) | (layer0_outputs[9140]);
    assign outputs[7847] = (layer0_outputs[6678]) & ~(layer0_outputs[730]);
    assign outputs[7848] = (layer0_outputs[7853]) | (layer0_outputs[966]);
    assign outputs[7849] = layer0_outputs[2280];
    assign outputs[7850] = ~((layer0_outputs[10070]) ^ (layer0_outputs[4702]));
    assign outputs[7851] = 1'b0;
    assign outputs[7852] = ~(layer0_outputs[5269]);
    assign outputs[7853] = ~((layer0_outputs[8530]) | (layer0_outputs[3665]));
    assign outputs[7854] = ~(layer0_outputs[4307]) | (layer0_outputs[2171]);
    assign outputs[7855] = ~(layer0_outputs[8769]);
    assign outputs[7856] = ~(layer0_outputs[10212]);
    assign outputs[7857] = layer0_outputs[332];
    assign outputs[7858] = (layer0_outputs[7320]) ^ (layer0_outputs[3070]);
    assign outputs[7859] = (layer0_outputs[8890]) ^ (layer0_outputs[6087]);
    assign outputs[7860] = (layer0_outputs[5201]) & ~(layer0_outputs[4683]);
    assign outputs[7861] = ~(layer0_outputs[9891]) | (layer0_outputs[2491]);
    assign outputs[7862] = ~((layer0_outputs[7180]) | (layer0_outputs[4858]));
    assign outputs[7863] = layer0_outputs[2228];
    assign outputs[7864] = (layer0_outputs[3143]) ^ (layer0_outputs[9780]);
    assign outputs[7865] = layer0_outputs[5796];
    assign outputs[7866] = (layer0_outputs[5425]) & ~(layer0_outputs[2867]);
    assign outputs[7867] = layer0_outputs[5353];
    assign outputs[7868] = ~(layer0_outputs[9819]);
    assign outputs[7869] = ~((layer0_outputs[6320]) ^ (layer0_outputs[2814]));
    assign outputs[7870] = layer0_outputs[3021];
    assign outputs[7871] = layer0_outputs[8260];
    assign outputs[7872] = layer0_outputs[4154];
    assign outputs[7873] = (layer0_outputs[3206]) ^ (layer0_outputs[3114]);
    assign outputs[7874] = (layer0_outputs[4769]) & ~(layer0_outputs[9310]);
    assign outputs[7875] = ~((layer0_outputs[135]) ^ (layer0_outputs[8259]));
    assign outputs[7876] = ~((layer0_outputs[7796]) ^ (layer0_outputs[3979]));
    assign outputs[7877] = ~((layer0_outputs[524]) | (layer0_outputs[2837]));
    assign outputs[7878] = ~(layer0_outputs[4699]);
    assign outputs[7879] = ~(layer0_outputs[5866]);
    assign outputs[7880] = ~(layer0_outputs[7628]);
    assign outputs[7881] = layer0_outputs[732];
    assign outputs[7882] = ~((layer0_outputs[1647]) | (layer0_outputs[3133]));
    assign outputs[7883] = ~(layer0_outputs[7867]);
    assign outputs[7884] = ~(layer0_outputs[1753]);
    assign outputs[7885] = layer0_outputs[1404];
    assign outputs[7886] = layer0_outputs[5476];
    assign outputs[7887] = layer0_outputs[5520];
    assign outputs[7888] = ~((layer0_outputs[5241]) ^ (layer0_outputs[1057]));
    assign outputs[7889] = ~(layer0_outputs[1715]);
    assign outputs[7890] = (layer0_outputs[3543]) & ~(layer0_outputs[6278]);
    assign outputs[7891] = (layer0_outputs[9312]) & ~(layer0_outputs[22]);
    assign outputs[7892] = layer0_outputs[1333];
    assign outputs[7893] = ~(layer0_outputs[6627]) | (layer0_outputs[7697]);
    assign outputs[7894] = ~((layer0_outputs[486]) ^ (layer0_outputs[6359]));
    assign outputs[7895] = (layer0_outputs[3509]) ^ (layer0_outputs[7537]);
    assign outputs[7896] = ~((layer0_outputs[4504]) ^ (layer0_outputs[2743]));
    assign outputs[7897] = (layer0_outputs[5750]) & (layer0_outputs[757]);
    assign outputs[7898] = ~(layer0_outputs[7095]);
    assign outputs[7899] = (layer0_outputs[9322]) & ~(layer0_outputs[2562]);
    assign outputs[7900] = ~(layer0_outputs[7580]);
    assign outputs[7901] = layer0_outputs[6479];
    assign outputs[7902] = (layer0_outputs[6857]) & ~(layer0_outputs[583]);
    assign outputs[7903] = ~((layer0_outputs[9874]) ^ (layer0_outputs[7479]));
    assign outputs[7904] = (layer0_outputs[1384]) & ~(layer0_outputs[2942]);
    assign outputs[7905] = ~((layer0_outputs[5422]) ^ (layer0_outputs[100]));
    assign outputs[7906] = ~(layer0_outputs[1487]);
    assign outputs[7907] = layer0_outputs[7906];
    assign outputs[7908] = layer0_outputs[1912];
    assign outputs[7909] = ~(layer0_outputs[867]) | (layer0_outputs[7260]);
    assign outputs[7910] = ~((layer0_outputs[4363]) | (layer0_outputs[7787]));
    assign outputs[7911] = ~(layer0_outputs[1590]);
    assign outputs[7912] = ~(layer0_outputs[4289]);
    assign outputs[7913] = ~(layer0_outputs[7085]);
    assign outputs[7914] = (layer0_outputs[2680]) & ~(layer0_outputs[4044]);
    assign outputs[7915] = ~(layer0_outputs[619]);
    assign outputs[7916] = ~(layer0_outputs[10126]);
    assign outputs[7917] = ~(layer0_outputs[5121]);
    assign outputs[7918] = layer0_outputs[2597];
    assign outputs[7919] = (layer0_outputs[4888]) ^ (layer0_outputs[5908]);
    assign outputs[7920] = ~((layer0_outputs[5985]) & (layer0_outputs[551]));
    assign outputs[7921] = ~(layer0_outputs[4778]);
    assign outputs[7922] = ~((layer0_outputs[2594]) & (layer0_outputs[4567]));
    assign outputs[7923] = layer0_outputs[892];
    assign outputs[7924] = layer0_outputs[2870];
    assign outputs[7925] = (layer0_outputs[2809]) & ~(layer0_outputs[3955]);
    assign outputs[7926] = ~(layer0_outputs[7939]);
    assign outputs[7927] = ~((layer0_outputs[1116]) | (layer0_outputs[3048]));
    assign outputs[7928] = ~(layer0_outputs[8060]);
    assign outputs[7929] = ~(layer0_outputs[9966]);
    assign outputs[7930] = layer0_outputs[4069];
    assign outputs[7931] = ~((layer0_outputs[7162]) & (layer0_outputs[604]));
    assign outputs[7932] = ~(layer0_outputs[9436]);
    assign outputs[7933] = layer0_outputs[1024];
    assign outputs[7934] = (layer0_outputs[5129]) & ~(layer0_outputs[6411]);
    assign outputs[7935] = ~(layer0_outputs[5321]);
    assign outputs[7936] = ~((layer0_outputs[6547]) | (layer0_outputs[3959]));
    assign outputs[7937] = (layer0_outputs[8313]) & (layer0_outputs[1535]);
    assign outputs[7938] = (layer0_outputs[5424]) & ~(layer0_outputs[8623]);
    assign outputs[7939] = (layer0_outputs[9829]) & ~(layer0_outputs[7562]);
    assign outputs[7940] = ~(layer0_outputs[7919]) | (layer0_outputs[2406]);
    assign outputs[7941] = layer0_outputs[4719];
    assign outputs[7942] = ~((layer0_outputs[9737]) | (layer0_outputs[5553]));
    assign outputs[7943] = (layer0_outputs[6961]) | (layer0_outputs[5134]);
    assign outputs[7944] = ~((layer0_outputs[631]) ^ (layer0_outputs[928]));
    assign outputs[7945] = layer0_outputs[6225];
    assign outputs[7946] = ~(layer0_outputs[8190]) | (layer0_outputs[648]);
    assign outputs[7947] = (layer0_outputs[7962]) & ~(layer0_outputs[3901]);
    assign outputs[7948] = ~(layer0_outputs[4690]);
    assign outputs[7949] = (layer0_outputs[3912]) & ~(layer0_outputs[7340]);
    assign outputs[7950] = layer0_outputs[5686];
    assign outputs[7951] = layer0_outputs[7107];
    assign outputs[7952] = layer0_outputs[4012];
    assign outputs[7953] = layer0_outputs[2865];
    assign outputs[7954] = ~(layer0_outputs[9995]);
    assign outputs[7955] = layer0_outputs[9190];
    assign outputs[7956] = ~((layer0_outputs[155]) ^ (layer0_outputs[5819]));
    assign outputs[7957] = layer0_outputs[5031];
    assign outputs[7958] = ~((layer0_outputs[5298]) | (layer0_outputs[4881]));
    assign outputs[7959] = ~(layer0_outputs[1285]) | (layer0_outputs[1564]);
    assign outputs[7960] = (layer0_outputs[3100]) ^ (layer0_outputs[7045]);
    assign outputs[7961] = ~((layer0_outputs[2721]) ^ (layer0_outputs[5885]));
    assign outputs[7962] = (layer0_outputs[4286]) & ~(layer0_outputs[3878]);
    assign outputs[7963] = ~(layer0_outputs[9640]);
    assign outputs[7964] = (layer0_outputs[9121]) ^ (layer0_outputs[8562]);
    assign outputs[7965] = ~(layer0_outputs[2179]);
    assign outputs[7966] = layer0_outputs[5736];
    assign outputs[7967] = ~(layer0_outputs[4936]);
    assign outputs[7968] = (layer0_outputs[1527]) & ~(layer0_outputs[8001]);
    assign outputs[7969] = layer0_outputs[4347];
    assign outputs[7970] = ~((layer0_outputs[8853]) ^ (layer0_outputs[9013]));
    assign outputs[7971] = ~((layer0_outputs[9516]) ^ (layer0_outputs[1253]));
    assign outputs[7972] = ~((layer0_outputs[9956]) ^ (layer0_outputs[3054]));
    assign outputs[7973] = layer0_outputs[9368];
    assign outputs[7974] = (layer0_outputs[6853]) ^ (layer0_outputs[9928]);
    assign outputs[7975] = (layer0_outputs[9838]) & (layer0_outputs[5921]);
    assign outputs[7976] = (layer0_outputs[5177]) ^ (layer0_outputs[3540]);
    assign outputs[7977] = (layer0_outputs[5479]) & (layer0_outputs[2127]);
    assign outputs[7978] = ~(layer0_outputs[5593]);
    assign outputs[7979] = layer0_outputs[6946];
    assign outputs[7980] = (layer0_outputs[452]) & (layer0_outputs[1302]);
    assign outputs[7981] = ~((layer0_outputs[2563]) ^ (layer0_outputs[3303]));
    assign outputs[7982] = ~(layer0_outputs[4200]);
    assign outputs[7983] = layer0_outputs[9977];
    assign outputs[7984] = ~((layer0_outputs[2772]) ^ (layer0_outputs[7240]));
    assign outputs[7985] = (layer0_outputs[6314]) ^ (layer0_outputs[7059]);
    assign outputs[7986] = (layer0_outputs[1336]) & (layer0_outputs[2554]);
    assign outputs[7987] = ~(layer0_outputs[3858]) | (layer0_outputs[8744]);
    assign outputs[7988] = ~((layer0_outputs[2425]) ^ (layer0_outputs[94]));
    assign outputs[7989] = layer0_outputs[2033];
    assign outputs[7990] = ~(layer0_outputs[8014]);
    assign outputs[7991] = layer0_outputs[4397];
    assign outputs[7992] = ~((layer0_outputs[2360]) | (layer0_outputs[3885]));
    assign outputs[7993] = ~(layer0_outputs[8487]);
    assign outputs[7994] = ~(layer0_outputs[4215]);
    assign outputs[7995] = ~(layer0_outputs[366]);
    assign outputs[7996] = ~(layer0_outputs[219]);
    assign outputs[7997] = ~(layer0_outputs[5415]);
    assign outputs[7998] = ~(layer0_outputs[1892]) | (layer0_outputs[1453]);
    assign outputs[7999] = (layer0_outputs[566]) ^ (layer0_outputs[7157]);
    assign outputs[8000] = (layer0_outputs[3443]) & ~(layer0_outputs[1409]);
    assign outputs[8001] = (layer0_outputs[1791]) & (layer0_outputs[640]);
    assign outputs[8002] = ~(layer0_outputs[5622]) | (layer0_outputs[1139]);
    assign outputs[8003] = ~((layer0_outputs[2758]) | (layer0_outputs[730]));
    assign outputs[8004] = (layer0_outputs[2176]) & ~(layer0_outputs[9158]);
    assign outputs[8005] = ~(layer0_outputs[5415]);
    assign outputs[8006] = ~(layer0_outputs[60]);
    assign outputs[8007] = layer0_outputs[6528];
    assign outputs[8008] = ~(layer0_outputs[2995]) | (layer0_outputs[42]);
    assign outputs[8009] = ~(layer0_outputs[10046]);
    assign outputs[8010] = (layer0_outputs[7996]) | (layer0_outputs[9172]);
    assign outputs[8011] = ~(layer0_outputs[5477]);
    assign outputs[8012] = layer0_outputs[2155];
    assign outputs[8013] = layer0_outputs[6223];
    assign outputs[8014] = ~((layer0_outputs[4179]) ^ (layer0_outputs[10116]));
    assign outputs[8015] = (layer0_outputs[7149]) & ~(layer0_outputs[1256]);
    assign outputs[8016] = (layer0_outputs[7584]) ^ (layer0_outputs[6661]);
    assign outputs[8017] = (layer0_outputs[6467]) ^ (layer0_outputs[4318]);
    assign outputs[8018] = ~(layer0_outputs[3357]);
    assign outputs[8019] = layer0_outputs[4609];
    assign outputs[8020] = (layer0_outputs[6794]) & (layer0_outputs[9762]);
    assign outputs[8021] = (layer0_outputs[2423]) & (layer0_outputs[1036]);
    assign outputs[8022] = ~(layer0_outputs[7867]);
    assign outputs[8023] = (layer0_outputs[9372]) ^ (layer0_outputs[9934]);
    assign outputs[8024] = (layer0_outputs[4780]) & ~(layer0_outputs[8980]);
    assign outputs[8025] = ~((layer0_outputs[7732]) ^ (layer0_outputs[4275]));
    assign outputs[8026] = layer0_outputs[7845];
    assign outputs[8027] = layer0_outputs[9843];
    assign outputs[8028] = ~(layer0_outputs[8000]);
    assign outputs[8029] = layer0_outputs[520];
    assign outputs[8030] = ~((layer0_outputs[4012]) ^ (layer0_outputs[8901]));
    assign outputs[8031] = ~((layer0_outputs[3938]) ^ (layer0_outputs[5918]));
    assign outputs[8032] = ~(layer0_outputs[8625]);
    assign outputs[8033] = (layer0_outputs[7954]) & (layer0_outputs[898]);
    assign outputs[8034] = ~((layer0_outputs[5315]) | (layer0_outputs[5141]));
    assign outputs[8035] = (layer0_outputs[8391]) & ~(layer0_outputs[440]);
    assign outputs[8036] = (layer0_outputs[5320]) ^ (layer0_outputs[10029]);
    assign outputs[8037] = layer0_outputs[8519];
    assign outputs[8038] = ~((layer0_outputs[7592]) ^ (layer0_outputs[6830]));
    assign outputs[8039] = layer0_outputs[8943];
    assign outputs[8040] = layer0_outputs[331];
    assign outputs[8041] = (layer0_outputs[7945]) | (layer0_outputs[1238]);
    assign outputs[8042] = ~(layer0_outputs[8686]);
    assign outputs[8043] = ~((layer0_outputs[6368]) & (layer0_outputs[5020]));
    assign outputs[8044] = ~(layer0_outputs[10053]);
    assign outputs[8045] = layer0_outputs[8951];
    assign outputs[8046] = layer0_outputs[9396];
    assign outputs[8047] = (layer0_outputs[2200]) & ~(layer0_outputs[1597]);
    assign outputs[8048] = layer0_outputs[8607];
    assign outputs[8049] = ~((layer0_outputs[3887]) | (layer0_outputs[521]));
    assign outputs[8050] = ~(layer0_outputs[5503]) | (layer0_outputs[9885]);
    assign outputs[8051] = (layer0_outputs[1977]) & (layer0_outputs[3809]);
    assign outputs[8052] = (layer0_outputs[5341]) & ~(layer0_outputs[5680]);
    assign outputs[8053] = ~((layer0_outputs[8836]) | (layer0_outputs[2180]));
    assign outputs[8054] = 1'b0;
    assign outputs[8055] = ~((layer0_outputs[8938]) ^ (layer0_outputs[5756]));
    assign outputs[8056] = layer0_outputs[8886];
    assign outputs[8057] = layer0_outputs[7766];
    assign outputs[8058] = ~((layer0_outputs[2667]) ^ (layer0_outputs[8828]));
    assign outputs[8059] = ~(layer0_outputs[8390]);
    assign outputs[8060] = (layer0_outputs[9207]) & ~(layer0_outputs[3701]);
    assign outputs[8061] = ~(layer0_outputs[3242]);
    assign outputs[8062] = (layer0_outputs[1153]) ^ (layer0_outputs[9854]);
    assign outputs[8063] = ~((layer0_outputs[5000]) ^ (layer0_outputs[7338]));
    assign outputs[8064] = ~((layer0_outputs[9465]) ^ (layer0_outputs[6172]));
    assign outputs[8065] = layer0_outputs[4433];
    assign outputs[8066] = ~(layer0_outputs[1164]);
    assign outputs[8067] = ~((layer0_outputs[35]) ^ (layer0_outputs[8245]));
    assign outputs[8068] = layer0_outputs[6040];
    assign outputs[8069] = (layer0_outputs[1775]) & ~(layer0_outputs[10125]);
    assign outputs[8070] = ~((layer0_outputs[3988]) ^ (layer0_outputs[127]));
    assign outputs[8071] = (layer0_outputs[367]) & ~(layer0_outputs[4576]);
    assign outputs[8072] = (layer0_outputs[9457]) & ~(layer0_outputs[5213]);
    assign outputs[8073] = layer0_outputs[3833];
    assign outputs[8074] = ~((layer0_outputs[6845]) ^ (layer0_outputs[3235]));
    assign outputs[8075] = ~((layer0_outputs[7186]) | (layer0_outputs[9947]));
    assign outputs[8076] = (layer0_outputs[5617]) & ~(layer0_outputs[4857]);
    assign outputs[8077] = (layer0_outputs[9295]) & ~(layer0_outputs[1322]);
    assign outputs[8078] = layer0_outputs[7784];
    assign outputs[8079] = layer0_outputs[245];
    assign outputs[8080] = ~((layer0_outputs[8187]) ^ (layer0_outputs[918]));
    assign outputs[8081] = 1'b1;
    assign outputs[8082] = ~((layer0_outputs[5678]) ^ (layer0_outputs[3629]));
    assign outputs[8083] = ~(layer0_outputs[2636]);
    assign outputs[8084] = ~((layer0_outputs[5822]) ^ (layer0_outputs[4903]));
    assign outputs[8085] = ~(layer0_outputs[5659]);
    assign outputs[8086] = (layer0_outputs[5130]) & ~(layer0_outputs[3751]);
    assign outputs[8087] = (layer0_outputs[9321]) | (layer0_outputs[1125]);
    assign outputs[8088] = (layer0_outputs[2902]) & ~(layer0_outputs[5566]);
    assign outputs[8089] = ~((layer0_outputs[727]) & (layer0_outputs[6446]));
    assign outputs[8090] = ~((layer0_outputs[9852]) ^ (layer0_outputs[8396]));
    assign outputs[8091] = layer0_outputs[1698];
    assign outputs[8092] = ~((layer0_outputs[8612]) | (layer0_outputs[440]));
    assign outputs[8093] = ~((layer0_outputs[9309]) ^ (layer0_outputs[4089]));
    assign outputs[8094] = ~(layer0_outputs[7465]);
    assign outputs[8095] = layer0_outputs[5781];
    assign outputs[8096] = ~((layer0_outputs[5654]) | (layer0_outputs[10026]));
    assign outputs[8097] = layer0_outputs[9403];
    assign outputs[8098] = 1'b0;
    assign outputs[8099] = (layer0_outputs[6472]) ^ (layer0_outputs[6331]);
    assign outputs[8100] = ~((layer0_outputs[3661]) ^ (layer0_outputs[1464]));
    assign outputs[8101] = (layer0_outputs[7838]) & ~(layer0_outputs[10001]);
    assign outputs[8102] = ~((layer0_outputs[5978]) ^ (layer0_outputs[4753]));
    assign outputs[8103] = layer0_outputs[3593];
    assign outputs[8104] = ~(layer0_outputs[4188]);
    assign outputs[8105] = (layer0_outputs[6613]) ^ (layer0_outputs[7691]);
    assign outputs[8106] = ~((layer0_outputs[9681]) ^ (layer0_outputs[4298]));
    assign outputs[8107] = ~(layer0_outputs[4671]);
    assign outputs[8108] = (layer0_outputs[4589]) ^ (layer0_outputs[1219]);
    assign outputs[8109] = (layer0_outputs[3119]) & ~(layer0_outputs[5846]);
    assign outputs[8110] = (layer0_outputs[7469]) & ~(layer0_outputs[4712]);
    assign outputs[8111] = ~(layer0_outputs[3788]);
    assign outputs[8112] = 1'b1;
    assign outputs[8113] = ~((layer0_outputs[10059]) | (layer0_outputs[3814]));
    assign outputs[8114] = layer0_outputs[7657];
    assign outputs[8115] = ~(layer0_outputs[4536]);
    assign outputs[8116] = ~(layer0_outputs[7998]);
    assign outputs[8117] = layer0_outputs[8551];
    assign outputs[8118] = ~(layer0_outputs[5615]);
    assign outputs[8119] = (layer0_outputs[7988]) & (layer0_outputs[3923]);
    assign outputs[8120] = layer0_outputs[4874];
    assign outputs[8121] = layer0_outputs[6082];
    assign outputs[8122] = ~(layer0_outputs[7814]);
    assign outputs[8123] = ~((layer0_outputs[5531]) & (layer0_outputs[683]));
    assign outputs[8124] = (layer0_outputs[1210]) & ~(layer0_outputs[4689]);
    assign outputs[8125] = ~(layer0_outputs[6399]) | (layer0_outputs[1300]);
    assign outputs[8126] = layer0_outputs[9081];
    assign outputs[8127] = ~((layer0_outputs[1928]) ^ (layer0_outputs[8671]));
    assign outputs[8128] = layer0_outputs[1799];
    assign outputs[8129] = ~((layer0_outputs[502]) ^ (layer0_outputs[8597]));
    assign outputs[8130] = layer0_outputs[176];
    assign outputs[8131] = ~((layer0_outputs[6869]) ^ (layer0_outputs[5152]));
    assign outputs[8132] = layer0_outputs[4624];
    assign outputs[8133] = (layer0_outputs[5628]) ^ (layer0_outputs[9054]);
    assign outputs[8134] = (layer0_outputs[8229]) ^ (layer0_outputs[4854]);
    assign outputs[8135] = (layer0_outputs[2499]) & ~(layer0_outputs[4041]);
    assign outputs[8136] = (layer0_outputs[7405]) & ~(layer0_outputs[102]);
    assign outputs[8137] = layer0_outputs[2114];
    assign outputs[8138] = layer0_outputs[5144];
    assign outputs[8139] = ~(layer0_outputs[9341]);
    assign outputs[8140] = ~((layer0_outputs[10154]) | (layer0_outputs[6117]));
    assign outputs[8141] = ~((layer0_outputs[6518]) ^ (layer0_outputs[1363]));
    assign outputs[8142] = (layer0_outputs[3640]) & ~(layer0_outputs[5334]);
    assign outputs[8143] = ~(layer0_outputs[5814]) | (layer0_outputs[1909]);
    assign outputs[8144] = (layer0_outputs[2398]) & ~(layer0_outputs[2729]);
    assign outputs[8145] = (layer0_outputs[389]) & ~(layer0_outputs[1643]);
    assign outputs[8146] = (layer0_outputs[8328]) ^ (layer0_outputs[8763]);
    assign outputs[8147] = ~((layer0_outputs[7275]) | (layer0_outputs[6237]));
    assign outputs[8148] = layer0_outputs[8084];
    assign outputs[8149] = ~((layer0_outputs[1644]) & (layer0_outputs[5078]));
    assign outputs[8150] = (layer0_outputs[3081]) ^ (layer0_outputs[2753]);
    assign outputs[8151] = (layer0_outputs[5048]) & ~(layer0_outputs[177]);
    assign outputs[8152] = layer0_outputs[7077];
    assign outputs[8153] = layer0_outputs[5845];
    assign outputs[8154] = ~(layer0_outputs[6152]) | (layer0_outputs[4261]);
    assign outputs[8155] = ~((layer0_outputs[4638]) | (layer0_outputs[2719]));
    assign outputs[8156] = ~((layer0_outputs[825]) ^ (layer0_outputs[9088]));
    assign outputs[8157] = ~(layer0_outputs[8631]);
    assign outputs[8158] = ~(layer0_outputs[956]);
    assign outputs[8159] = (layer0_outputs[2306]) & ~(layer0_outputs[1067]);
    assign outputs[8160] = ~(layer0_outputs[5844]);
    assign outputs[8161] = (layer0_outputs[3075]) & ~(layer0_outputs[8540]);
    assign outputs[8162] = ~(layer0_outputs[1907]);
    assign outputs[8163] = (layer0_outputs[319]) ^ (layer0_outputs[6973]);
    assign outputs[8164] = (layer0_outputs[1470]) & (layer0_outputs[163]);
    assign outputs[8165] = ~((layer0_outputs[7344]) | (layer0_outputs[8463]));
    assign outputs[8166] = ~(layer0_outputs[1120]) | (layer0_outputs[7912]);
    assign outputs[8167] = (layer0_outputs[7263]) ^ (layer0_outputs[2247]);
    assign outputs[8168] = ~(layer0_outputs[9894]);
    assign outputs[8169] = (layer0_outputs[8906]) & (layer0_outputs[2546]);
    assign outputs[8170] = ~((layer0_outputs[3635]) | (layer0_outputs[3507]));
    assign outputs[8171] = ~((layer0_outputs[9984]) ^ (layer0_outputs[8747]));
    assign outputs[8172] = ~((layer0_outputs[9225]) | (layer0_outputs[571]));
    assign outputs[8173] = ~((layer0_outputs[960]) ^ (layer0_outputs[2753]));
    assign outputs[8174] = ~((layer0_outputs[9815]) & (layer0_outputs[4825]));
    assign outputs[8175] = ~(layer0_outputs[7570]);
    assign outputs[8176] = (layer0_outputs[2950]) ^ (layer0_outputs[5875]);
    assign outputs[8177] = (layer0_outputs[7793]) ^ (layer0_outputs[3137]);
    assign outputs[8178] = layer0_outputs[5756];
    assign outputs[8179] = (layer0_outputs[9855]) ^ (layer0_outputs[3890]);
    assign outputs[8180] = layer0_outputs[1347];
    assign outputs[8181] = ~((layer0_outputs[171]) | (layer0_outputs[4923]));
    assign outputs[8182] = (layer0_outputs[5656]) ^ (layer0_outputs[8381]);
    assign outputs[8183] = (layer0_outputs[6116]) & ~(layer0_outputs[1206]);
    assign outputs[8184] = layer0_outputs[2520];
    assign outputs[8185] = ~(layer0_outputs[681]);
    assign outputs[8186] = (layer0_outputs[5904]) & ~(layer0_outputs[3295]);
    assign outputs[8187] = ~((layer0_outputs[1973]) | (layer0_outputs[392]));
    assign outputs[8188] = ~(layer0_outputs[7984]);
    assign outputs[8189] = layer0_outputs[374];
    assign outputs[8190] = (layer0_outputs[8923]) & (layer0_outputs[2542]);
    assign outputs[8191] = (layer0_outputs[3434]) ^ (layer0_outputs[144]);
    assign outputs[8192] = layer0_outputs[6664];
    assign outputs[8193] = ~((layer0_outputs[8309]) | (layer0_outputs[2207]));
    assign outputs[8194] = ~((layer0_outputs[4749]) | (layer0_outputs[7972]));
    assign outputs[8195] = ~(layer0_outputs[4573]);
    assign outputs[8196] = ~(layer0_outputs[5558]);
    assign outputs[8197] = layer0_outputs[2937];
    assign outputs[8198] = ~(layer0_outputs[7905]) | (layer0_outputs[4547]);
    assign outputs[8199] = layer0_outputs[634];
    assign outputs[8200] = (layer0_outputs[5239]) & ~(layer0_outputs[8560]);
    assign outputs[8201] = ~((layer0_outputs[9959]) & (layer0_outputs[2946]));
    assign outputs[8202] = ~(layer0_outputs[6468]);
    assign outputs[8203] = layer0_outputs[4787];
    assign outputs[8204] = 1'b1;
    assign outputs[8205] = layer0_outputs[320];
    assign outputs[8206] = ~(layer0_outputs[1483]);
    assign outputs[8207] = layer0_outputs[10138];
    assign outputs[8208] = ~(layer0_outputs[1101]);
    assign outputs[8209] = ~(layer0_outputs[3349]);
    assign outputs[8210] = (layer0_outputs[3896]) ^ (layer0_outputs[1774]);
    assign outputs[8211] = ~(layer0_outputs[6055]);
    assign outputs[8212] = 1'b1;
    assign outputs[8213] = ~((layer0_outputs[6237]) ^ (layer0_outputs[2513]));
    assign outputs[8214] = ~((layer0_outputs[6951]) | (layer0_outputs[9035]));
    assign outputs[8215] = layer0_outputs[8423];
    assign outputs[8216] = layer0_outputs[7911];
    assign outputs[8217] = (layer0_outputs[8045]) & ~(layer0_outputs[399]);
    assign outputs[8218] = (layer0_outputs[1641]) ^ (layer0_outputs[4618]);
    assign outputs[8219] = layer0_outputs[3194];
    assign outputs[8220] = (layer0_outputs[45]) ^ (layer0_outputs[6303]);
    assign outputs[8221] = layer0_outputs[5312];
    assign outputs[8222] = layer0_outputs[4242];
    assign outputs[8223] = (layer0_outputs[8357]) ^ (layer0_outputs[1429]);
    assign outputs[8224] = ~(layer0_outputs[8228]) | (layer0_outputs[7541]);
    assign outputs[8225] = ~((layer0_outputs[2823]) | (layer0_outputs[1929]));
    assign outputs[8226] = 1'b1;
    assign outputs[8227] = ~((layer0_outputs[5539]) | (layer0_outputs[8606]));
    assign outputs[8228] = layer0_outputs[6407];
    assign outputs[8229] = (layer0_outputs[6939]) ^ (layer0_outputs[1382]);
    assign outputs[8230] = ~((layer0_outputs[7589]) ^ (layer0_outputs[2340]));
    assign outputs[8231] = ~(layer0_outputs[5598]) | (layer0_outputs[599]);
    assign outputs[8232] = (layer0_outputs[6797]) ^ (layer0_outputs[4839]);
    assign outputs[8233] = (layer0_outputs[561]) ^ (layer0_outputs[1430]);
    assign outputs[8234] = ~(layer0_outputs[3965]);
    assign outputs[8235] = ~(layer0_outputs[116]) | (layer0_outputs[755]);
    assign outputs[8236] = layer0_outputs[8323];
    assign outputs[8237] = ~(layer0_outputs[6162]);
    assign outputs[8238] = layer0_outputs[9950];
    assign outputs[8239] = layer0_outputs[3687];
    assign outputs[8240] = ~(layer0_outputs[4932]);
    assign outputs[8241] = ~((layer0_outputs[7407]) ^ (layer0_outputs[7843]));
    assign outputs[8242] = (layer0_outputs[6996]) ^ (layer0_outputs[1041]);
    assign outputs[8243] = layer0_outputs[1397];
    assign outputs[8244] = (layer0_outputs[2693]) ^ (layer0_outputs[5136]);
    assign outputs[8245] = ~(layer0_outputs[2439]);
    assign outputs[8246] = layer0_outputs[9708];
    assign outputs[8247] = (layer0_outputs[4158]) ^ (layer0_outputs[1580]);
    assign outputs[8248] = (layer0_outputs[5841]) & ~(layer0_outputs[9416]);
    assign outputs[8249] = ~(layer0_outputs[9480]);
    assign outputs[8250] = ~(layer0_outputs[3283]) | (layer0_outputs[4432]);
    assign outputs[8251] = (layer0_outputs[747]) ^ (layer0_outputs[1417]);
    assign outputs[8252] = layer0_outputs[5816];
    assign outputs[8253] = (layer0_outputs[10134]) ^ (layer0_outputs[4593]);
    assign outputs[8254] = (layer0_outputs[920]) ^ (layer0_outputs[1934]);
    assign outputs[8255] = (layer0_outputs[7865]) & ~(layer0_outputs[9770]);
    assign outputs[8256] = (layer0_outputs[4664]) & ~(layer0_outputs[6420]);
    assign outputs[8257] = layer0_outputs[8278];
    assign outputs[8258] = layer0_outputs[6861];
    assign outputs[8259] = ~(layer0_outputs[7306]);
    assign outputs[8260] = layer0_outputs[4659];
    assign outputs[8261] = (layer0_outputs[1144]) ^ (layer0_outputs[6619]);
    assign outputs[8262] = ~(layer0_outputs[8662]);
    assign outputs[8263] = ~(layer0_outputs[5391]) | (layer0_outputs[4569]);
    assign outputs[8264] = layer0_outputs[5567];
    assign outputs[8265] = ~((layer0_outputs[499]) ^ (layer0_outputs[9357]));
    assign outputs[8266] = (layer0_outputs[3801]) ^ (layer0_outputs[5419]);
    assign outputs[8267] = ~(layer0_outputs[10091]);
    assign outputs[8268] = layer0_outputs[9317];
    assign outputs[8269] = layer0_outputs[1141];
    assign outputs[8270] = ~((layer0_outputs[6281]) | (layer0_outputs[4666]));
    assign outputs[8271] = ~((layer0_outputs[10096]) ^ (layer0_outputs[9145]));
    assign outputs[8272] = layer0_outputs[5301];
    assign outputs[8273] = ~((layer0_outputs[4235]) ^ (layer0_outputs[662]));
    assign outputs[8274] = ~((layer0_outputs[289]) | (layer0_outputs[4608]));
    assign outputs[8275] = (layer0_outputs[4738]) ^ (layer0_outputs[8965]);
    assign outputs[8276] = (layer0_outputs[4647]) ^ (layer0_outputs[8607]);
    assign outputs[8277] = ~((layer0_outputs[4182]) ^ (layer0_outputs[208]));
    assign outputs[8278] = ~((layer0_outputs[5754]) ^ (layer0_outputs[2045]));
    assign outputs[8279] = (layer0_outputs[8351]) & ~(layer0_outputs[4049]);
    assign outputs[8280] = layer0_outputs[568];
    assign outputs[8281] = ~(layer0_outputs[1405]);
    assign outputs[8282] = ~((layer0_outputs[1284]) | (layer0_outputs[1840]));
    assign outputs[8283] = ~(layer0_outputs[2270]);
    assign outputs[8284] = (layer0_outputs[3083]) ^ (layer0_outputs[5677]);
    assign outputs[8285] = ~(layer0_outputs[5785]) | (layer0_outputs[4467]);
    assign outputs[8286] = (layer0_outputs[7866]) & ~(layer0_outputs[4183]);
    assign outputs[8287] = (layer0_outputs[638]) ^ (layer0_outputs[3253]);
    assign outputs[8288] = (layer0_outputs[1474]) | (layer0_outputs[9237]);
    assign outputs[8289] = layer0_outputs[9149];
    assign outputs[8290] = (layer0_outputs[4885]) | (layer0_outputs[6427]);
    assign outputs[8291] = (layer0_outputs[6462]) ^ (layer0_outputs[3481]);
    assign outputs[8292] = ~(layer0_outputs[9981]);
    assign outputs[8293] = layer0_outputs[1084];
    assign outputs[8294] = layer0_outputs[4820];
    assign outputs[8295] = ~(layer0_outputs[6036]);
    assign outputs[8296] = ~((layer0_outputs[7742]) ^ (layer0_outputs[6911]));
    assign outputs[8297] = (layer0_outputs[299]) ^ (layer0_outputs[2027]);
    assign outputs[8298] = ~(layer0_outputs[3402]);
    assign outputs[8299] = layer0_outputs[2430];
    assign outputs[8300] = (layer0_outputs[1142]) & ~(layer0_outputs[3870]);
    assign outputs[8301] = ~(layer0_outputs[7157]) | (layer0_outputs[1086]);
    assign outputs[8302] = layer0_outputs[2148];
    assign outputs[8303] = ~((layer0_outputs[9092]) ^ (layer0_outputs[9270]));
    assign outputs[8304] = layer0_outputs[5672];
    assign outputs[8305] = (layer0_outputs[5021]) | (layer0_outputs[8582]);
    assign outputs[8306] = ~((layer0_outputs[7072]) ^ (layer0_outputs[4489]));
    assign outputs[8307] = (layer0_outputs[1761]) & (layer0_outputs[7951]);
    assign outputs[8308] = ~(layer0_outputs[5694]);
    assign outputs[8309] = layer0_outputs[2015];
    assign outputs[8310] = (layer0_outputs[5502]) & ~(layer0_outputs[9877]);
    assign outputs[8311] = layer0_outputs[9235];
    assign outputs[8312] = (layer0_outputs[7284]) ^ (layer0_outputs[5282]);
    assign outputs[8313] = ~(layer0_outputs[2454]) | (layer0_outputs[3426]);
    assign outputs[8314] = (layer0_outputs[7229]) & (layer0_outputs[6694]);
    assign outputs[8315] = ~((layer0_outputs[2690]) | (layer0_outputs[6872]));
    assign outputs[8316] = ~((layer0_outputs[4162]) ^ (layer0_outputs[7098]));
    assign outputs[8317] = ~((layer0_outputs[8270]) ^ (layer0_outputs[8695]));
    assign outputs[8318] = layer0_outputs[7765];
    assign outputs[8319] = ~(layer0_outputs[996]);
    assign outputs[8320] = (layer0_outputs[2036]) & ~(layer0_outputs[8911]);
    assign outputs[8321] = (layer0_outputs[343]) & ~(layer0_outputs[8142]);
    assign outputs[8322] = ~((layer0_outputs[1328]) ^ (layer0_outputs[3164]));
    assign outputs[8323] = (layer0_outputs[3561]) & (layer0_outputs[4147]);
    assign outputs[8324] = layer0_outputs[5564];
    assign outputs[8325] = ~((layer0_outputs[9812]) ^ (layer0_outputs[7687]));
    assign outputs[8326] = ~(layer0_outputs[7585]) | (layer0_outputs[8413]);
    assign outputs[8327] = ~(layer0_outputs[4745]);
    assign outputs[8328] = ~(layer0_outputs[3191]);
    assign outputs[8329] = ~((layer0_outputs[6145]) ^ (layer0_outputs[4308]));
    assign outputs[8330] = ~(layer0_outputs[3412]);
    assign outputs[8331] = ~((layer0_outputs[242]) & (layer0_outputs[8226]));
    assign outputs[8332] = (layer0_outputs[5441]) & (layer0_outputs[9617]);
    assign outputs[8333] = ~(layer0_outputs[7014]) | (layer0_outputs[7062]);
    assign outputs[8334] = ~(layer0_outputs[8712]);
    assign outputs[8335] = ~(layer0_outputs[604]);
    assign outputs[8336] = (layer0_outputs[4917]) ^ (layer0_outputs[327]);
    assign outputs[8337] = layer0_outputs[9286];
    assign outputs[8338] = (layer0_outputs[1007]) | (layer0_outputs[8034]);
    assign outputs[8339] = layer0_outputs[298];
    assign outputs[8340] = ~((layer0_outputs[5830]) ^ (layer0_outputs[7440]));
    assign outputs[8341] = layer0_outputs[1900];
    assign outputs[8342] = ~(layer0_outputs[3203]);
    assign outputs[8343] = layer0_outputs[10105];
    assign outputs[8344] = ~((layer0_outputs[487]) ^ (layer0_outputs[10034]));
    assign outputs[8345] = ~((layer0_outputs[4821]) ^ (layer0_outputs[6488]));
    assign outputs[8346] = layer0_outputs[10114];
    assign outputs[8347] = (layer0_outputs[9948]) ^ (layer0_outputs[8443]);
    assign outputs[8348] = ~(layer0_outputs[3334]);
    assign outputs[8349] = ~(layer0_outputs[1987]);
    assign outputs[8350] = ~(layer0_outputs[7982]) | (layer0_outputs[1102]);
    assign outputs[8351] = (layer0_outputs[1010]) ^ (layer0_outputs[1893]);
    assign outputs[8352] = layer0_outputs[3272];
    assign outputs[8353] = ~(layer0_outputs[8432]);
    assign outputs[8354] = ~((layer0_outputs[3996]) ^ (layer0_outputs[7448]));
    assign outputs[8355] = 1'b1;
    assign outputs[8356] = (layer0_outputs[8216]) & ~(layer0_outputs[9788]);
    assign outputs[8357] = ~(layer0_outputs[2165]);
    assign outputs[8358] = ~(layer0_outputs[3720]);
    assign outputs[8359] = layer0_outputs[5777];
    assign outputs[8360] = ~((layer0_outputs[3369]) ^ (layer0_outputs[7369]));
    assign outputs[8361] = (layer0_outputs[3782]) & ~(layer0_outputs[1563]);
    assign outputs[8362] = layer0_outputs[6947];
    assign outputs[8363] = (layer0_outputs[3923]) & ~(layer0_outputs[3200]);
    assign outputs[8364] = ~(layer0_outputs[4424]) | (layer0_outputs[3487]);
    assign outputs[8365] = (layer0_outputs[6842]) ^ (layer0_outputs[1320]);
    assign outputs[8366] = layer0_outputs[3381];
    assign outputs[8367] = ~(layer0_outputs[4225]);
    assign outputs[8368] = layer0_outputs[7733];
    assign outputs[8369] = (layer0_outputs[8304]) & (layer0_outputs[7484]);
    assign outputs[8370] = (layer0_outputs[5220]) ^ (layer0_outputs[6353]);
    assign outputs[8371] = ~(layer0_outputs[2436]);
    assign outputs[8372] = ~(layer0_outputs[1737]);
    assign outputs[8373] = ~(layer0_outputs[297]);
    assign outputs[8374] = ~(layer0_outputs[244]) | (layer0_outputs[2011]);
    assign outputs[8375] = layer0_outputs[724];
    assign outputs[8376] = (layer0_outputs[223]) & ~(layer0_outputs[7211]);
    assign outputs[8377] = (layer0_outputs[1109]) ^ (layer0_outputs[1404]);
    assign outputs[8378] = ~(layer0_outputs[3092]);
    assign outputs[8379] = layer0_outputs[4581];
    assign outputs[8380] = (layer0_outputs[1051]) ^ (layer0_outputs[5400]);
    assign outputs[8381] = (layer0_outputs[8996]) ^ (layer0_outputs[4798]);
    assign outputs[8382] = ~((layer0_outputs[2886]) | (layer0_outputs[9058]));
    assign outputs[8383] = ~(layer0_outputs[3668]) | (layer0_outputs[2544]);
    assign outputs[8384] = (layer0_outputs[8352]) & ~(layer0_outputs[4330]);
    assign outputs[8385] = ~(layer0_outputs[7621]);
    assign outputs[8386] = ~((layer0_outputs[6640]) ^ (layer0_outputs[729]));
    assign outputs[8387] = ~(layer0_outputs[6158]);
    assign outputs[8388] = (layer0_outputs[9692]) ^ (layer0_outputs[1419]);
    assign outputs[8389] = (layer0_outputs[9039]) | (layer0_outputs[1126]);
    assign outputs[8390] = layer0_outputs[2398];
    assign outputs[8391] = ~(layer0_outputs[8284]) | (layer0_outputs[3305]);
    assign outputs[8392] = (layer0_outputs[9326]) & ~(layer0_outputs[3731]);
    assign outputs[8393] = layer0_outputs[7794];
    assign outputs[8394] = ~((layer0_outputs[2129]) & (layer0_outputs[8825]));
    assign outputs[8395] = (layer0_outputs[6053]) ^ (layer0_outputs[1652]);
    assign outputs[8396] = layer0_outputs[6581];
    assign outputs[8397] = ~((layer0_outputs[2383]) ^ (layer0_outputs[1427]));
    assign outputs[8398] = layer0_outputs[9216];
    assign outputs[8399] = layer0_outputs[8208];
    assign outputs[8400] = ~((layer0_outputs[3378]) ^ (layer0_outputs[5604]));
    assign outputs[8401] = (layer0_outputs[6481]) | (layer0_outputs[4845]);
    assign outputs[8402] = ~(layer0_outputs[2999]) | (layer0_outputs[6809]);
    assign outputs[8403] = layer0_outputs[1412];
    assign outputs[8404] = ~(layer0_outputs[1475]);
    assign outputs[8405] = ~(layer0_outputs[6846]);
    assign outputs[8406] = 1'b1;
    assign outputs[8407] = ~((layer0_outputs[7184]) ^ (layer0_outputs[2289]));
    assign outputs[8408] = ~(layer0_outputs[8669]);
    assign outputs[8409] = (layer0_outputs[7025]) | (layer0_outputs[8349]);
    assign outputs[8410] = layer0_outputs[5566];
    assign outputs[8411] = layer0_outputs[5465];
    assign outputs[8412] = ~(layer0_outputs[2676]);
    assign outputs[8413] = ~(layer0_outputs[1310]);
    assign outputs[8414] = ~((layer0_outputs[3504]) & (layer0_outputs[8093]));
    assign outputs[8415] = (layer0_outputs[9854]) | (layer0_outputs[8496]);
    assign outputs[8416] = (layer0_outputs[375]) ^ (layer0_outputs[1133]);
    assign outputs[8417] = ~(layer0_outputs[8975]) | (layer0_outputs[4845]);
    assign outputs[8418] = ~(layer0_outputs[6867]);
    assign outputs[8419] = (layer0_outputs[8638]) & (layer0_outputs[4595]);
    assign outputs[8420] = ~(layer0_outputs[8368]);
    assign outputs[8421] = layer0_outputs[3067];
    assign outputs[8422] = (layer0_outputs[7688]) ^ (layer0_outputs[3303]);
    assign outputs[8423] = ~(layer0_outputs[5987]);
    assign outputs[8424] = ~(layer0_outputs[329]);
    assign outputs[8425] = ~(layer0_outputs[9774]);
    assign outputs[8426] = (layer0_outputs[3270]) | (layer0_outputs[5515]);
    assign outputs[8427] = ~(layer0_outputs[3630]);
    assign outputs[8428] = ~((layer0_outputs[8135]) | (layer0_outputs[7023]));
    assign outputs[8429] = layer0_outputs[6828];
    assign outputs[8430] = ~(layer0_outputs[709]);
    assign outputs[8431] = ~((layer0_outputs[1692]) ^ (layer0_outputs[9659]));
    assign outputs[8432] = ~((layer0_outputs[654]) ^ (layer0_outputs[1255]));
    assign outputs[8433] = (layer0_outputs[1271]) | (layer0_outputs[9527]);
    assign outputs[8434] = ~(layer0_outputs[3211]);
    assign outputs[8435] = layer0_outputs[3999];
    assign outputs[8436] = (layer0_outputs[4876]) & (layer0_outputs[4992]);
    assign outputs[8437] = (layer0_outputs[9663]) ^ (layer0_outputs[9945]);
    assign outputs[8438] = ~((layer0_outputs[2806]) ^ (layer0_outputs[9103]));
    assign outputs[8439] = (layer0_outputs[39]) | (layer0_outputs[8226]);
    assign outputs[8440] = ~(layer0_outputs[5967]) | (layer0_outputs[9895]);
    assign outputs[8441] = (layer0_outputs[15]) & ~(layer0_outputs[3442]);
    assign outputs[8442] = (layer0_outputs[2027]) ^ (layer0_outputs[4722]);
    assign outputs[8443] = layer0_outputs[1947];
    assign outputs[8444] = ~(layer0_outputs[492]);
    assign outputs[8445] = (layer0_outputs[6042]) & (layer0_outputs[1935]);
    assign outputs[8446] = layer0_outputs[8815];
    assign outputs[8447] = ~((layer0_outputs[3862]) & (layer0_outputs[1380]));
    assign outputs[8448] = (layer0_outputs[4018]) | (layer0_outputs[630]);
    assign outputs[8449] = layer0_outputs[10110];
    assign outputs[8450] = layer0_outputs[239];
    assign outputs[8451] = ~(layer0_outputs[2730]);
    assign outputs[8452] = ~((layer0_outputs[3821]) ^ (layer0_outputs[4336]));
    assign outputs[8453] = ~((layer0_outputs[1589]) ^ (layer0_outputs[9700]));
    assign outputs[8454] = ~(layer0_outputs[3418]) | (layer0_outputs[8037]);
    assign outputs[8455] = (layer0_outputs[2453]) & ~(layer0_outputs[2318]);
    assign outputs[8456] = (layer0_outputs[6051]) ^ (layer0_outputs[6609]);
    assign outputs[8457] = ~(layer0_outputs[10038]);
    assign outputs[8458] = layer0_outputs[6296];
    assign outputs[8459] = ~(layer0_outputs[5180]);
    assign outputs[8460] = ~(layer0_outputs[4615]);
    assign outputs[8461] = layer0_outputs[8663];
    assign outputs[8462] = ~(layer0_outputs[1498]);
    assign outputs[8463] = ~((layer0_outputs[4827]) ^ (layer0_outputs[472]));
    assign outputs[8464] = 1'b1;
    assign outputs[8465] = (layer0_outputs[5027]) ^ (layer0_outputs[9866]);
    assign outputs[8466] = ~((layer0_outputs[6270]) ^ (layer0_outputs[7770]));
    assign outputs[8467] = ~(layer0_outputs[3177]) | (layer0_outputs[875]);
    assign outputs[8468] = (layer0_outputs[8456]) & ~(layer0_outputs[9469]);
    assign outputs[8469] = ~(layer0_outputs[8285]);
    assign outputs[8470] = layer0_outputs[6099];
    assign outputs[8471] = ~(layer0_outputs[6178]);
    assign outputs[8472] = layer0_outputs[9367];
    assign outputs[8473] = (layer0_outputs[5544]) & (layer0_outputs[9535]);
    assign outputs[8474] = (layer0_outputs[1456]) ^ (layer0_outputs[7114]);
    assign outputs[8475] = layer0_outputs[8415];
    assign outputs[8476] = ~(layer0_outputs[2664]);
    assign outputs[8477] = ~(layer0_outputs[8318]);
    assign outputs[8478] = ~((layer0_outputs[5747]) ^ (layer0_outputs[6895]));
    assign outputs[8479] = ~(layer0_outputs[6304]);
    assign outputs[8480] = (layer0_outputs[7158]) ^ (layer0_outputs[9328]);
    assign outputs[8481] = ~(layer0_outputs[6043]);
    assign outputs[8482] = ~(layer0_outputs[921]);
    assign outputs[8483] = (layer0_outputs[4546]) ^ (layer0_outputs[5116]);
    assign outputs[8484] = ~((layer0_outputs[728]) ^ (layer0_outputs[877]));
    assign outputs[8485] = layer0_outputs[2230];
    assign outputs[8486] = (layer0_outputs[8684]) ^ (layer0_outputs[5277]);
    assign outputs[8487] = ~(layer0_outputs[5436]);
    assign outputs[8488] = ~(layer0_outputs[10097]) | (layer0_outputs[428]);
    assign outputs[8489] = ~(layer0_outputs[5134]);
    assign outputs[8490] = (layer0_outputs[9047]) | (layer0_outputs[2321]);
    assign outputs[8491] = ~(layer0_outputs[6633]) | (layer0_outputs[8845]);
    assign outputs[8492] = layer0_outputs[6690];
    assign outputs[8493] = ~(layer0_outputs[7900]);
    assign outputs[8494] = ~(layer0_outputs[8918]) | (layer0_outputs[10072]);
    assign outputs[8495] = ~(layer0_outputs[6149]);
    assign outputs[8496] = layer0_outputs[7608];
    assign outputs[8497] = ~(layer0_outputs[1000]) | (layer0_outputs[63]);
    assign outputs[8498] = layer0_outputs[9452];
    assign outputs[8499] = ~(layer0_outputs[893]) | (layer0_outputs[6579]);
    assign outputs[8500] = (layer0_outputs[10116]) & ~(layer0_outputs[3607]);
    assign outputs[8501] = ~(layer0_outputs[3832]);
    assign outputs[8502] = ~((layer0_outputs[8473]) ^ (layer0_outputs[1676]));
    assign outputs[8503] = layer0_outputs[3050];
    assign outputs[8504] = (layer0_outputs[1076]) & ~(layer0_outputs[10186]);
    assign outputs[8505] = (layer0_outputs[9733]) | (layer0_outputs[752]);
    assign outputs[8506] = (layer0_outputs[4834]) ^ (layer0_outputs[7288]);
    assign outputs[8507] = (layer0_outputs[2389]) ^ (layer0_outputs[8337]);
    assign outputs[8508] = ~(layer0_outputs[4861]);
    assign outputs[8509] = (layer0_outputs[8955]) ^ (layer0_outputs[7861]);
    assign outputs[8510] = ~((layer0_outputs[7444]) | (layer0_outputs[4635]));
    assign outputs[8511] = ~((layer0_outputs[5454]) ^ (layer0_outputs[3767]));
    assign outputs[8512] = ~(layer0_outputs[8682]);
    assign outputs[8513] = (layer0_outputs[9017]) ^ (layer0_outputs[8121]);
    assign outputs[8514] = (layer0_outputs[4445]) ^ (layer0_outputs[3873]);
    assign outputs[8515] = (layer0_outputs[3079]) & ~(layer0_outputs[3946]);
    assign outputs[8516] = (layer0_outputs[3333]) & ~(layer0_outputs[9146]);
    assign outputs[8517] = ~(layer0_outputs[5853]) | (layer0_outputs[8622]);
    assign outputs[8518] = ~((layer0_outputs[7819]) ^ (layer0_outputs[4296]));
    assign outputs[8519] = (layer0_outputs[1301]) ^ (layer0_outputs[7725]);
    assign outputs[8520] = ~(layer0_outputs[5541]);
    assign outputs[8521] = (layer0_outputs[9176]) & (layer0_outputs[2418]);
    assign outputs[8522] = layer0_outputs[401];
    assign outputs[8523] = ~(layer0_outputs[6305]);
    assign outputs[8524] = layer0_outputs[6679];
    assign outputs[8525] = (layer0_outputs[9538]) | (layer0_outputs[3744]);
    assign outputs[8526] = (layer0_outputs[9273]) ^ (layer0_outputs[9858]);
    assign outputs[8527] = (layer0_outputs[6751]) | (layer0_outputs[4897]);
    assign outputs[8528] = ~(layer0_outputs[9555]) | (layer0_outputs[1213]);
    assign outputs[8529] = (layer0_outputs[5532]) ^ (layer0_outputs[10144]);
    assign outputs[8530] = ~(layer0_outputs[3771]);
    assign outputs[8531] = ~((layer0_outputs[4792]) ^ (layer0_outputs[5986]));
    assign outputs[8532] = ~((layer0_outputs[3356]) ^ (layer0_outputs[1460]));
    assign outputs[8533] = (layer0_outputs[9641]) ^ (layer0_outputs[7816]);
    assign outputs[8534] = layer0_outputs[8263];
    assign outputs[8535] = ~((layer0_outputs[2469]) ^ (layer0_outputs[9619]));
    assign outputs[8536] = ~((layer0_outputs[9404]) | (layer0_outputs[8014]));
    assign outputs[8537] = ~(layer0_outputs[6174]);
    assign outputs[8538] = ~((layer0_outputs[1771]) ^ (layer0_outputs[2625]));
    assign outputs[8539] = ~(layer0_outputs[4614]);
    assign outputs[8540] = ~(layer0_outputs[5835]);
    assign outputs[8541] = ~((layer0_outputs[4029]) ^ (layer0_outputs[2116]));
    assign outputs[8542] = (layer0_outputs[121]) & ~(layer0_outputs[6750]);
    assign outputs[8543] = (layer0_outputs[9830]) ^ (layer0_outputs[7251]);
    assign outputs[8544] = (layer0_outputs[5080]) | (layer0_outputs[8929]);
    assign outputs[8545] = ~(layer0_outputs[3799]);
    assign outputs[8546] = (layer0_outputs[8039]) & ~(layer0_outputs[7086]);
    assign outputs[8547] = ~((layer0_outputs[1180]) & (layer0_outputs[1508]));
    assign outputs[8548] = ~(layer0_outputs[8168]);
    assign outputs[8549] = layer0_outputs[7459];
    assign outputs[8550] = ~(layer0_outputs[7967]);
    assign outputs[8551] = (layer0_outputs[4233]) ^ (layer0_outputs[6083]);
    assign outputs[8552] = (layer0_outputs[7454]) | (layer0_outputs[7645]);
    assign outputs[8553] = layer0_outputs[5834];
    assign outputs[8554] = ~(layer0_outputs[997]);
    assign outputs[8555] = (layer0_outputs[6702]) & ~(layer0_outputs[945]);
    assign outputs[8556] = ~((layer0_outputs[4588]) ^ (layer0_outputs[7139]));
    assign outputs[8557] = ~(layer0_outputs[7083]) | (layer0_outputs[7765]);
    assign outputs[8558] = (layer0_outputs[3764]) ^ (layer0_outputs[1182]);
    assign outputs[8559] = ~(layer0_outputs[7267]);
    assign outputs[8560] = layer0_outputs[4459];
    assign outputs[8561] = ~(layer0_outputs[7478]);
    assign outputs[8562] = layer0_outputs[70];
    assign outputs[8563] = layer0_outputs[5020];
    assign outputs[8564] = (layer0_outputs[126]) ^ (layer0_outputs[1870]);
    assign outputs[8565] = ~((layer0_outputs[3084]) & (layer0_outputs[1298]));
    assign outputs[8566] = ~(layer0_outputs[9932]) | (layer0_outputs[4089]);
    assign outputs[8567] = (layer0_outputs[2674]) ^ (layer0_outputs[3047]);
    assign outputs[8568] = layer0_outputs[8797];
    assign outputs[8569] = layer0_outputs[8979];
    assign outputs[8570] = (layer0_outputs[5884]) ^ (layer0_outputs[7430]);
    assign outputs[8571] = layer0_outputs[7933];
    assign outputs[8572] = ~(layer0_outputs[3292]) | (layer0_outputs[6763]);
    assign outputs[8573] = ~(layer0_outputs[7055]);
    assign outputs[8574] = (layer0_outputs[558]) ^ (layer0_outputs[9629]);
    assign outputs[8575] = ~(layer0_outputs[8390]) | (layer0_outputs[231]);
    assign outputs[8576] = ~((layer0_outputs[1359]) & (layer0_outputs[2223]));
    assign outputs[8577] = layer0_outputs[630];
    assign outputs[8578] = (layer0_outputs[4110]) ^ (layer0_outputs[8307]);
    assign outputs[8579] = ~(layer0_outputs[3672]);
    assign outputs[8580] = ~(layer0_outputs[8498]);
    assign outputs[8581] = ~(layer0_outputs[3260]);
    assign outputs[8582] = ~(layer0_outputs[6631]);
    assign outputs[8583] = layer0_outputs[2164];
    assign outputs[8584] = layer0_outputs[6788];
    assign outputs[8585] = ~(layer0_outputs[7085]);
    assign outputs[8586] = (layer0_outputs[6294]) ^ (layer0_outputs[9776]);
    assign outputs[8587] = ~((layer0_outputs[3301]) ^ (layer0_outputs[6431]));
    assign outputs[8588] = ~((layer0_outputs[1304]) | (layer0_outputs[6614]));
    assign outputs[8589] = layer0_outputs[456];
    assign outputs[8590] = layer0_outputs[1726];
    assign outputs[8591] = ~((layer0_outputs[10069]) & (layer0_outputs[1423]));
    assign outputs[8592] = (layer0_outputs[4649]) & (layer0_outputs[5542]);
    assign outputs[8593] = (layer0_outputs[6754]) & ~(layer0_outputs[3753]);
    assign outputs[8594] = ~((layer0_outputs[8446]) ^ (layer0_outputs[9463]));
    assign outputs[8595] = layer0_outputs[3508];
    assign outputs[8596] = ~((layer0_outputs[8817]) | (layer0_outputs[6380]));
    assign outputs[8597] = ~((layer0_outputs[3452]) & (layer0_outputs[6218]));
    assign outputs[8598] = (layer0_outputs[5153]) & (layer0_outputs[4477]);
    assign outputs[8599] = layer0_outputs[3967];
    assign outputs[8600] = (layer0_outputs[4038]) & ~(layer0_outputs[5212]);
    assign outputs[8601] = ~(layer0_outputs[4777]);
    assign outputs[8602] = (layer0_outputs[5458]) ^ (layer0_outputs[7897]);
    assign outputs[8603] = ~(layer0_outputs[557]);
    assign outputs[8604] = (layer0_outputs[1785]) & ~(layer0_outputs[4597]);
    assign outputs[8605] = (layer0_outputs[3985]) & ~(layer0_outputs[6721]);
    assign outputs[8606] = layer0_outputs[2817];
    assign outputs[8607] = layer0_outputs[7064];
    assign outputs[8608] = ~(layer0_outputs[5413]) | (layer0_outputs[7329]);
    assign outputs[8609] = ~((layer0_outputs[3714]) & (layer0_outputs[735]));
    assign outputs[8610] = ~(layer0_outputs[6109]) | (layer0_outputs[1565]);
    assign outputs[8611] = (layer0_outputs[6702]) & (layer0_outputs[6773]);
    assign outputs[8612] = layer0_outputs[9749];
    assign outputs[8613] = ~(layer0_outputs[184]);
    assign outputs[8614] = ~(layer0_outputs[1445]);
    assign outputs[8615] = ~(layer0_outputs[2484]);
    assign outputs[8616] = (layer0_outputs[8176]) ^ (layer0_outputs[7372]);
    assign outputs[8617] = layer0_outputs[2348];
    assign outputs[8618] = ~((layer0_outputs[8741]) ^ (layer0_outputs[4300]));
    assign outputs[8619] = ~(layer0_outputs[7237]);
    assign outputs[8620] = (layer0_outputs[812]) & (layer0_outputs[9717]);
    assign outputs[8621] = (layer0_outputs[7173]) & (layer0_outputs[555]);
    assign outputs[8622] = ~((layer0_outputs[11]) ^ (layer0_outputs[944]));
    assign outputs[8623] = ~(layer0_outputs[1507]);
    assign outputs[8624] = ~((layer0_outputs[5377]) ^ (layer0_outputs[3262]));
    assign outputs[8625] = (layer0_outputs[2986]) & (layer0_outputs[2279]);
    assign outputs[8626] = ~((layer0_outputs[9276]) ^ (layer0_outputs[1292]));
    assign outputs[8627] = (layer0_outputs[2087]) & ~(layer0_outputs[6904]);
    assign outputs[8628] = (layer0_outputs[1093]) ^ (layer0_outputs[6649]);
    assign outputs[8629] = ~((layer0_outputs[8292]) | (layer0_outputs[2111]));
    assign outputs[8630] = ~(layer0_outputs[9278]) | (layer0_outputs[3338]);
    assign outputs[8631] = ~((layer0_outputs[3971]) & (layer0_outputs[7508]));
    assign outputs[8632] = ~(layer0_outputs[3135]) | (layer0_outputs[3337]);
    assign outputs[8633] = ~((layer0_outputs[6048]) & (layer0_outputs[8660]));
    assign outputs[8634] = (layer0_outputs[447]) ^ (layer0_outputs[9498]);
    assign outputs[8635] = ~(layer0_outputs[8123]);
    assign outputs[8636] = ~(layer0_outputs[313]) | (layer0_outputs[1574]);
    assign outputs[8637] = layer0_outputs[4305];
    assign outputs[8638] = (layer0_outputs[7881]) | (layer0_outputs[7175]);
    assign outputs[8639] = ~(layer0_outputs[8499]);
    assign outputs[8640] = (layer0_outputs[4245]) | (layer0_outputs[3125]);
    assign outputs[8641] = ~(layer0_outputs[8542]) | (layer0_outputs[207]);
    assign outputs[8642] = layer0_outputs[371];
    assign outputs[8643] = ~(layer0_outputs[4421]) | (layer0_outputs[5696]);
    assign outputs[8644] = layer0_outputs[2738];
    assign outputs[8645] = (layer0_outputs[5917]) & ~(layer0_outputs[6222]);
    assign outputs[8646] = ~((layer0_outputs[2952]) ^ (layer0_outputs[4648]));
    assign outputs[8647] = ~(layer0_outputs[1204]);
    assign outputs[8648] = layer0_outputs[4852];
    assign outputs[8649] = layer0_outputs[569];
    assign outputs[8650] = layer0_outputs[808];
    assign outputs[8651] = layer0_outputs[9828];
    assign outputs[8652] = ~((layer0_outputs[5696]) ^ (layer0_outputs[3742]));
    assign outputs[8653] = ~((layer0_outputs[8445]) & (layer0_outputs[9765]));
    assign outputs[8654] = ~(layer0_outputs[4512]);
    assign outputs[8655] = ~((layer0_outputs[545]) ^ (layer0_outputs[2643]));
    assign outputs[8656] = ~(layer0_outputs[488]);
    assign outputs[8657] = layer0_outputs[8000];
    assign outputs[8658] = ~(layer0_outputs[1192]);
    assign outputs[8659] = ~(layer0_outputs[646]);
    assign outputs[8660] = ~(layer0_outputs[2277]);
    assign outputs[8661] = (layer0_outputs[6456]) ^ (layer0_outputs[9307]);
    assign outputs[8662] = (layer0_outputs[1542]) | (layer0_outputs[7851]);
    assign outputs[8663] = (layer0_outputs[8379]) | (layer0_outputs[5364]);
    assign outputs[8664] = (layer0_outputs[8948]) ^ (layer0_outputs[4389]);
    assign outputs[8665] = (layer0_outputs[6624]) | (layer0_outputs[3769]);
    assign outputs[8666] = (layer0_outputs[5892]) & ~(layer0_outputs[4915]);
    assign outputs[8667] = ~((layer0_outputs[7077]) & (layer0_outputs[1856]));
    assign outputs[8668] = layer0_outputs[7048];
    assign outputs[8669] = ~(layer0_outputs[6414]) | (layer0_outputs[6964]);
    assign outputs[8670] = ~(layer0_outputs[9186]);
    assign outputs[8671] = ~((layer0_outputs[8472]) ^ (layer0_outputs[2545]));
    assign outputs[8672] = ~((layer0_outputs[6235]) ^ (layer0_outputs[8902]));
    assign outputs[8673] = layer0_outputs[6658];
    assign outputs[8674] = (layer0_outputs[6447]) ^ (layer0_outputs[967]);
    assign outputs[8675] = ~(layer0_outputs[5070]);
    assign outputs[8676] = layer0_outputs[9664];
    assign outputs[8677] = layer0_outputs[2126];
    assign outputs[8678] = ~((layer0_outputs[6056]) & (layer0_outputs[6749]));
    assign outputs[8679] = layer0_outputs[3400];
    assign outputs[8680] = (layer0_outputs[4982]) & (layer0_outputs[2335]);
    assign outputs[8681] = ~(layer0_outputs[827]) | (layer0_outputs[3745]);
    assign outputs[8682] = layer0_outputs[7807];
    assign outputs[8683] = ~(layer0_outputs[1005]) | (layer0_outputs[681]);
    assign outputs[8684] = (layer0_outputs[8216]) ^ (layer0_outputs[2605]);
    assign outputs[8685] = ~(layer0_outputs[1129]) | (layer0_outputs[8969]);
    assign outputs[8686] = (layer0_outputs[3705]) | (layer0_outputs[6030]);
    assign outputs[8687] = layer0_outputs[7879];
    assign outputs[8688] = ~(layer0_outputs[4706]);
    assign outputs[8689] = ~(layer0_outputs[7411]) | (layer0_outputs[843]);
    assign outputs[8690] = ~(layer0_outputs[5995]);
    assign outputs[8691] = ~(layer0_outputs[1825]);
    assign outputs[8692] = ~(layer0_outputs[10111]) | (layer0_outputs[9073]);
    assign outputs[8693] = ~(layer0_outputs[2250]);
    assign outputs[8694] = 1'b1;
    assign outputs[8695] = ~(layer0_outputs[9161]);
    assign outputs[8696] = (layer0_outputs[8105]) & ~(layer0_outputs[9323]);
    assign outputs[8697] = (layer0_outputs[8092]) ^ (layer0_outputs[4237]);
    assign outputs[8698] = layer0_outputs[9102];
    assign outputs[8699] = ~(layer0_outputs[3837]);
    assign outputs[8700] = layer0_outputs[6794];
    assign outputs[8701] = ~((layer0_outputs[7451]) & (layer0_outputs[6153]));
    assign outputs[8702] = ~(layer0_outputs[7949]);
    assign outputs[8703] = (layer0_outputs[10039]) & (layer0_outputs[7699]);
    assign outputs[8704] = layer0_outputs[6552];
    assign outputs[8705] = 1'b1;
    assign outputs[8706] = ~((layer0_outputs[477]) | (layer0_outputs[335]));
    assign outputs[8707] = (layer0_outputs[3458]) ^ (layer0_outputs[54]);
    assign outputs[8708] = ~(layer0_outputs[2881]);
    assign outputs[8709] = ~((layer0_outputs[1034]) | (layer0_outputs[6791]));
    assign outputs[8710] = layer0_outputs[8704];
    assign outputs[8711] = ~((layer0_outputs[8667]) ^ (layer0_outputs[5100]));
    assign outputs[8712] = ~(layer0_outputs[907]);
    assign outputs[8713] = ~(layer0_outputs[3207]);
    assign outputs[8714] = 1'b0;
    assign outputs[8715] = ~(layer0_outputs[9283]) | (layer0_outputs[9823]);
    assign outputs[8716] = (layer0_outputs[5293]) ^ (layer0_outputs[7347]);
    assign outputs[8717] = layer0_outputs[9097];
    assign outputs[8718] = layer0_outputs[9634];
    assign outputs[8719] = layer0_outputs[1927];
    assign outputs[8720] = layer0_outputs[8507];
    assign outputs[8721] = (layer0_outputs[821]) & ~(layer0_outputs[2309]);
    assign outputs[8722] = ~(layer0_outputs[8112]);
    assign outputs[8723] = ~(layer0_outputs[4064]);
    assign outputs[8724] = (layer0_outputs[5684]) & ~(layer0_outputs[10099]);
    assign outputs[8725] = ~((layer0_outputs[433]) ^ (layer0_outputs[3140]));
    assign outputs[8726] = (layer0_outputs[1846]) ^ (layer0_outputs[9504]);
    assign outputs[8727] = layer0_outputs[1814];
    assign outputs[8728] = layer0_outputs[7523];
    assign outputs[8729] = layer0_outputs[2441];
    assign outputs[8730] = ~(layer0_outputs[2092]) | (layer0_outputs[657]);
    assign outputs[8731] = (layer0_outputs[324]) | (layer0_outputs[5463]);
    assign outputs[8732] = layer0_outputs[4692];
    assign outputs[8733] = ~(layer0_outputs[4409]);
    assign outputs[8734] = ~((layer0_outputs[4470]) ^ (layer0_outputs[2781]));
    assign outputs[8735] = ~(layer0_outputs[6951]) | (layer0_outputs[7316]);
    assign outputs[8736] = ~(layer0_outputs[2204]) | (layer0_outputs[1272]);
    assign outputs[8737] = layer0_outputs[78];
    assign outputs[8738] = ~(layer0_outputs[854]) | (layer0_outputs[4474]);
    assign outputs[8739] = ~((layer0_outputs[3879]) ^ (layer0_outputs[2485]));
    assign outputs[8740] = ~(layer0_outputs[9671]);
    assign outputs[8741] = (layer0_outputs[8374]) | (layer0_outputs[9734]);
    assign outputs[8742] = ~((layer0_outputs[4779]) ^ (layer0_outputs[1927]));
    assign outputs[8743] = ~((layer0_outputs[9948]) & (layer0_outputs[5636]));
    assign outputs[8744] = (layer0_outputs[1699]) ^ (layer0_outputs[9643]);
    assign outputs[8745] = ~(layer0_outputs[1970]) | (layer0_outputs[5460]);
    assign outputs[8746] = ~((layer0_outputs[7776]) ^ (layer0_outputs[4391]));
    assign outputs[8747] = layer0_outputs[4177];
    assign outputs[8748] = ~(layer0_outputs[2882]);
    assign outputs[8749] = (layer0_outputs[941]) ^ (layer0_outputs[9912]);
    assign outputs[8750] = ~(layer0_outputs[8616]);
    assign outputs[8751] = (layer0_outputs[676]) ^ (layer0_outputs[4375]);
    assign outputs[8752] = ~(layer0_outputs[7148]) | (layer0_outputs[5338]);
    assign outputs[8753] = ~((layer0_outputs[2305]) ^ (layer0_outputs[3961]));
    assign outputs[8754] = layer0_outputs[7022];
    assign outputs[8755] = ~(layer0_outputs[5559]);
    assign outputs[8756] = layer0_outputs[338];
    assign outputs[8757] = ~((layer0_outputs[5722]) ^ (layer0_outputs[8072]));
    assign outputs[8758] = (layer0_outputs[84]) ^ (layer0_outputs[4828]);
    assign outputs[8759] = (layer0_outputs[1853]) & ~(layer0_outputs[5609]);
    assign outputs[8760] = ~((layer0_outputs[4554]) ^ (layer0_outputs[6829]));
    assign outputs[8761] = ~(layer0_outputs[6670]) | (layer0_outputs[1045]);
    assign outputs[8762] = layer0_outputs[202];
    assign outputs[8763] = ~(layer0_outputs[3781]);
    assign outputs[8764] = (layer0_outputs[5175]) & ~(layer0_outputs[4377]);
    assign outputs[8765] = (layer0_outputs[4447]) & ~(layer0_outputs[6616]);
    assign outputs[8766] = ~(layer0_outputs[7060]);
    assign outputs[8767] = layer0_outputs[139];
    assign outputs[8768] = ~((layer0_outputs[8286]) ^ (layer0_outputs[9080]));
    assign outputs[8769] = (layer0_outputs[113]) | (layer0_outputs[523]);
    assign outputs[8770] = 1'b1;
    assign outputs[8771] = ~(layer0_outputs[4382]) | (layer0_outputs[20]);
    assign outputs[8772] = layer0_outputs[140];
    assign outputs[8773] = (layer0_outputs[1073]) | (layer0_outputs[4289]);
    assign outputs[8774] = layer0_outputs[1598];
    assign outputs[8775] = ~(layer0_outputs[9314]) | (layer0_outputs[6021]);
    assign outputs[8776] = ~((layer0_outputs[5344]) & (layer0_outputs[7980]));
    assign outputs[8777] = ~((layer0_outputs[1265]) ^ (layer0_outputs[6245]));
    assign outputs[8778] = layer0_outputs[6365];
    assign outputs[8779] = ~(layer0_outputs[6305]);
    assign outputs[8780] = (layer0_outputs[1511]) ^ (layer0_outputs[126]);
    assign outputs[8781] = ~(layer0_outputs[6027]) | (layer0_outputs[846]);
    assign outputs[8782] = layer0_outputs[2017];
    assign outputs[8783] = layer0_outputs[4121];
    assign outputs[8784] = (layer0_outputs[4097]) ^ (layer0_outputs[9642]);
    assign outputs[8785] = ~((layer0_outputs[5206]) ^ (layer0_outputs[873]));
    assign outputs[8786] = layer0_outputs[8036];
    assign outputs[8787] = ~((layer0_outputs[9289]) ^ (layer0_outputs[8629]));
    assign outputs[8788] = ~((layer0_outputs[491]) ^ (layer0_outputs[5773]));
    assign outputs[8789] = ~(layer0_outputs[7517]) | (layer0_outputs[3448]);
    assign outputs[8790] = layer0_outputs[1862];
    assign outputs[8791] = (layer0_outputs[7921]) & (layer0_outputs[867]);
    assign outputs[8792] = ~((layer0_outputs[5889]) ^ (layer0_outputs[5210]));
    assign outputs[8793] = ~((layer0_outputs[10123]) ^ (layer0_outputs[4201]));
    assign outputs[8794] = layer0_outputs[2700];
    assign outputs[8795] = ~((layer0_outputs[6002]) ^ (layer0_outputs[6432]));
    assign outputs[8796] = (layer0_outputs[8109]) | (layer0_outputs[9933]);
    assign outputs[8797] = layer0_outputs[1795];
    assign outputs[8798] = ~(layer0_outputs[2082]) | (layer0_outputs[2915]);
    assign outputs[8799] = (layer0_outputs[9336]) & (layer0_outputs[1461]);
    assign outputs[8800] = ~(layer0_outputs[8002]);
    assign outputs[8801] = ~((layer0_outputs[5638]) & (layer0_outputs[2502]));
    assign outputs[8802] = (layer0_outputs[6046]) | (layer0_outputs[3662]);
    assign outputs[8803] = layer0_outputs[9288];
    assign outputs[8804] = ~(layer0_outputs[5068]);
    assign outputs[8805] = (layer0_outputs[9345]) & ~(layer0_outputs[1746]);
    assign outputs[8806] = (layer0_outputs[2285]) & ~(layer0_outputs[5680]);
    assign outputs[8807] = layer0_outputs[3175];
    assign outputs[8808] = ~(layer0_outputs[2966]);
    assign outputs[8809] = ~(layer0_outputs[8701]);
    assign outputs[8810] = ~(layer0_outputs[1483]);
    assign outputs[8811] = layer0_outputs[7402];
    assign outputs[8812] = ~(layer0_outputs[9477]) | (layer0_outputs[1743]);
    assign outputs[8813] = ~((layer0_outputs[6824]) ^ (layer0_outputs[3414]));
    assign outputs[8814] = ~(layer0_outputs[6808]);
    assign outputs[8815] = ~((layer0_outputs[7183]) ^ (layer0_outputs[1832]));
    assign outputs[8816] = layer0_outputs[7321];
    assign outputs[8817] = ~((layer0_outputs[7290]) ^ (layer0_outputs[7975]));
    assign outputs[8818] = ~(layer0_outputs[7915]) | (layer0_outputs[2536]);
    assign outputs[8819] = ~((layer0_outputs[717]) ^ (layer0_outputs[6097]));
    assign outputs[8820] = ~((layer0_outputs[506]) ^ (layer0_outputs[5864]));
    assign outputs[8821] = (layer0_outputs[3904]) ^ (layer0_outputs[2486]);
    assign outputs[8822] = ~((layer0_outputs[2393]) & (layer0_outputs[5311]));
    assign outputs[8823] = layer0_outputs[6936];
    assign outputs[8824] = (layer0_outputs[8409]) ^ (layer0_outputs[7049]);
    assign outputs[8825] = (layer0_outputs[3220]) ^ (layer0_outputs[2147]);
    assign outputs[8826] = layer0_outputs[7716];
    assign outputs[8827] = ~(layer0_outputs[8297]);
    assign outputs[8828] = ~((layer0_outputs[9447]) | (layer0_outputs[4728]));
    assign outputs[8829] = (layer0_outputs[1127]) & (layer0_outputs[372]);
    assign outputs[8830] = (layer0_outputs[3432]) ^ (layer0_outputs[9763]);
    assign outputs[8831] = layer0_outputs[493];
    assign outputs[8832] = ~(layer0_outputs[3209]);
    assign outputs[8833] = ~(layer0_outputs[3646]);
    assign outputs[8834] = ~(layer0_outputs[4345]);
    assign outputs[8835] = layer0_outputs[1184];
    assign outputs[8836] = layer0_outputs[8213];
    assign outputs[8837] = ~((layer0_outputs[7636]) ^ (layer0_outputs[2117]));
    assign outputs[8838] = layer0_outputs[7747];
    assign outputs[8839] = layer0_outputs[99];
    assign outputs[8840] = ~(layer0_outputs[3563]);
    assign outputs[8841] = ~(layer0_outputs[7679]) | (layer0_outputs[3397]);
    assign outputs[8842] = ~((layer0_outputs[7018]) & (layer0_outputs[10137]));
    assign outputs[8843] = ~((layer0_outputs[10222]) | (layer0_outputs[8044]));
    assign outputs[8844] = 1'b1;
    assign outputs[8845] = (layer0_outputs[4015]) & (layer0_outputs[4507]);
    assign outputs[8846] = (layer0_outputs[2010]) | (layer0_outputs[5664]);
    assign outputs[8847] = (layer0_outputs[8059]) ^ (layer0_outputs[802]);
    assign outputs[8848] = ~((layer0_outputs[4253]) ^ (layer0_outputs[8494]));
    assign outputs[8849] = ~((layer0_outputs[3395]) | (layer0_outputs[2654]));
    assign outputs[8850] = ~((layer0_outputs[2754]) | (layer0_outputs[2298]));
    assign outputs[8851] = layer0_outputs[6121];
    assign outputs[8852] = layer0_outputs[2367];
    assign outputs[8853] = layer0_outputs[6349];
    assign outputs[8854] = ~(layer0_outputs[4238]);
    assign outputs[8855] = ~((layer0_outputs[9119]) ^ (layer0_outputs[5554]));
    assign outputs[8856] = ~(layer0_outputs[1909]) | (layer0_outputs[3570]);
    assign outputs[8857] = ~(layer0_outputs[2511]);
    assign outputs[8858] = ~(layer0_outputs[3171]) | (layer0_outputs[1618]);
    assign outputs[8859] = (layer0_outputs[8147]) & ~(layer0_outputs[7856]);
    assign outputs[8860] = ~(layer0_outputs[7202]);
    assign outputs[8861] = (layer0_outputs[1669]) & ~(layer0_outputs[5512]);
    assign outputs[8862] = ~(layer0_outputs[2848]) | (layer0_outputs[5504]);
    assign outputs[8863] = (layer0_outputs[1386]) ^ (layer0_outputs[8594]);
    assign outputs[8864] = (layer0_outputs[5082]) | (layer0_outputs[5881]);
    assign outputs[8865] = ~(layer0_outputs[7726]) | (layer0_outputs[8655]);
    assign outputs[8866] = ~((layer0_outputs[9359]) ^ (layer0_outputs[387]));
    assign outputs[8867] = ~(layer0_outputs[1374]);
    assign outputs[8868] = (layer0_outputs[7188]) & (layer0_outputs[1070]);
    assign outputs[8869] = ~(layer0_outputs[7266]);
    assign outputs[8870] = ~((layer0_outputs[3904]) ^ (layer0_outputs[5509]));
    assign outputs[8871] = layer0_outputs[4714];
    assign outputs[8872] = ~(layer0_outputs[2785]);
    assign outputs[8873] = layer0_outputs[9534];
    assign outputs[8874] = ~(layer0_outputs[8282]);
    assign outputs[8875] = (layer0_outputs[7112]) | (layer0_outputs[4664]);
    assign outputs[8876] = ~((layer0_outputs[7919]) ^ (layer0_outputs[7415]));
    assign outputs[8877] = ~(layer0_outputs[4067]) | (layer0_outputs[4083]);
    assign outputs[8878] = ~(layer0_outputs[6595]);
    assign outputs[8879] = layer0_outputs[5057];
    assign outputs[8880] = ~((layer0_outputs[5426]) & (layer0_outputs[6570]));
    assign outputs[8881] = layer0_outputs[754];
    assign outputs[8882] = layer0_outputs[8610];
    assign outputs[8883] = ~(layer0_outputs[7337]);
    assign outputs[8884] = layer0_outputs[3920];
    assign outputs[8885] = (layer0_outputs[7095]) ^ (layer0_outputs[3429]);
    assign outputs[8886] = ~(layer0_outputs[7828]);
    assign outputs[8887] = (layer0_outputs[8762]) ^ (layer0_outputs[7382]);
    assign outputs[8888] = (layer0_outputs[9338]) | (layer0_outputs[7216]);
    assign outputs[8889] = ~(layer0_outputs[8679]);
    assign outputs[8890] = (layer0_outputs[2551]) ^ (layer0_outputs[6753]);
    assign outputs[8891] = layer0_outputs[6450];
    assign outputs[8892] = 1'b1;
    assign outputs[8893] = ~(layer0_outputs[7703]);
    assign outputs[8894] = layer0_outputs[5037];
    assign outputs[8895] = layer0_outputs[4934];
    assign outputs[8896] = ~(layer0_outputs[2341]);
    assign outputs[8897] = ~((layer0_outputs[7424]) & (layer0_outputs[8867]));
    assign outputs[8898] = ~((layer0_outputs[9707]) ^ (layer0_outputs[6848]));
    assign outputs[8899] = ~((layer0_outputs[7437]) ^ (layer0_outputs[4507]));
    assign outputs[8900] = ~(layer0_outputs[377]);
    assign outputs[8901] = (layer0_outputs[4784]) & ~(layer0_outputs[1923]);
    assign outputs[8902] = (layer0_outputs[10197]) & ~(layer0_outputs[8561]);
    assign outputs[8903] = layer0_outputs[4299];
    assign outputs[8904] = ~((layer0_outputs[10005]) ^ (layer0_outputs[3468]));
    assign outputs[8905] = (layer0_outputs[9833]) | (layer0_outputs[4570]);
    assign outputs[8906] = ~(layer0_outputs[5039]) | (layer0_outputs[6774]);
    assign outputs[8907] = layer0_outputs[4187];
    assign outputs[8908] = ~(layer0_outputs[7736]);
    assign outputs[8909] = ~((layer0_outputs[4490]) | (layer0_outputs[4609]));
    assign outputs[8910] = ~(layer0_outputs[1636]) | (layer0_outputs[3667]);
    assign outputs[8911] = layer0_outputs[3683];
    assign outputs[8912] = (layer0_outputs[5298]) ^ (layer0_outputs[4143]);
    assign outputs[8913] = layer0_outputs[4506];
    assign outputs[8914] = ~((layer0_outputs[4740]) | (layer0_outputs[3529]));
    assign outputs[8915] = (layer0_outputs[9235]) | (layer0_outputs[306]);
    assign outputs[8916] = layer0_outputs[2001];
    assign outputs[8917] = (layer0_outputs[3351]) ^ (layer0_outputs[1778]);
    assign outputs[8918] = layer0_outputs[3507];
    assign outputs[8919] = layer0_outputs[175];
    assign outputs[8920] = ~(layer0_outputs[4980]);
    assign outputs[8921] = ~(layer0_outputs[368]);
    assign outputs[8922] = ~(layer0_outputs[7558]);
    assign outputs[8923] = ~(layer0_outputs[4059]);
    assign outputs[8924] = (layer0_outputs[4836]) & ~(layer0_outputs[6772]);
    assign outputs[8925] = (layer0_outputs[1567]) ^ (layer0_outputs[7156]);
    assign outputs[8926] = (layer0_outputs[1905]) ^ (layer0_outputs[3387]);
    assign outputs[8927] = layer0_outputs[7704];
    assign outputs[8928] = ~((layer0_outputs[150]) ^ (layer0_outputs[98]));
    assign outputs[8929] = layer0_outputs[6524];
    assign outputs[8930] = layer0_outputs[7472];
    assign outputs[8931] = ~(layer0_outputs[504]);
    assign outputs[8932] = ~((layer0_outputs[8127]) ^ (layer0_outputs[6326]));
    assign outputs[8933] = ~(layer0_outputs[3512]) | (layer0_outputs[3960]);
    assign outputs[8934] = (layer0_outputs[7758]) ^ (layer0_outputs[6889]);
    assign outputs[8935] = ~(layer0_outputs[6778]) | (layer0_outputs[6844]);
    assign outputs[8936] = ~((layer0_outputs[9663]) ^ (layer0_outputs[8694]));
    assign outputs[8937] = ~(layer0_outputs[157]);
    assign outputs[8938] = (layer0_outputs[7617]) ^ (layer0_outputs[1858]);
    assign outputs[8939] = layer0_outputs[6300];
    assign outputs[8940] = layer0_outputs[9069];
    assign outputs[8941] = ~((layer0_outputs[8635]) & (layer0_outputs[6246]));
    assign outputs[8942] = (layer0_outputs[9417]) ^ (layer0_outputs[9325]);
    assign outputs[8943] = ~(layer0_outputs[579]) | (layer0_outputs[3738]);
    assign outputs[8944] = (layer0_outputs[5695]) ^ (layer0_outputs[9888]);
    assign outputs[8945] = (layer0_outputs[3196]) | (layer0_outputs[5840]);
    assign outputs[8946] = (layer0_outputs[3456]) ^ (layer0_outputs[7051]);
    assign outputs[8947] = (layer0_outputs[263]) & ~(layer0_outputs[10036]);
    assign outputs[8948] = ~((layer0_outputs[5064]) & (layer0_outputs[3024]));
    assign outputs[8949] = 1'b0;
    assign outputs[8950] = ~((layer0_outputs[1894]) ^ (layer0_outputs[5856]));
    assign outputs[8951] = layer0_outputs[9086];
    assign outputs[8952] = layer0_outputs[9856];
    assign outputs[8953] = ~(layer0_outputs[7164]) | (layer0_outputs[9191]);
    assign outputs[8954] = (layer0_outputs[7349]) & ~(layer0_outputs[4116]);
    assign outputs[8955] = layer0_outputs[3891];
    assign outputs[8956] = (layer0_outputs[5874]) & ~(layer0_outputs[3892]);
    assign outputs[8957] = ~(layer0_outputs[10124]);
    assign outputs[8958] = ~((layer0_outputs[7094]) ^ (layer0_outputs[8548]));
    assign outputs[8959] = ~(layer0_outputs[5505]) | (layer0_outputs[3033]);
    assign outputs[8960] = ~((layer0_outputs[5957]) ^ (layer0_outputs[9252]));
    assign outputs[8961] = ~((layer0_outputs[3096]) ^ (layer0_outputs[5574]));
    assign outputs[8962] = layer0_outputs[9194];
    assign outputs[8963] = (layer0_outputs[3984]) | (layer0_outputs[5614]);
    assign outputs[8964] = ~((layer0_outputs[6829]) ^ (layer0_outputs[6912]));
    assign outputs[8965] = (layer0_outputs[9769]) & ~(layer0_outputs[10115]);
    assign outputs[8966] = layer0_outputs[7279];
    assign outputs[8967] = ~(layer0_outputs[3977]);
    assign outputs[8968] = ~((layer0_outputs[2749]) ^ (layer0_outputs[6684]));
    assign outputs[8969] = ~((layer0_outputs[6376]) ^ (layer0_outputs[7784]));
    assign outputs[8970] = ~(layer0_outputs[2598]) | (layer0_outputs[8621]);
    assign outputs[8971] = layer0_outputs[9248];
    assign outputs[8972] = layer0_outputs[8746];
    assign outputs[8973] = (layer0_outputs[3618]) | (layer0_outputs[6668]);
    assign outputs[8974] = layer0_outputs[7219];
    assign outputs[8975] = ~(layer0_outputs[631]) | (layer0_outputs[10166]);
    assign outputs[8976] = (layer0_outputs[2374]) | (layer0_outputs[692]);
    assign outputs[8977] = ~(layer0_outputs[9724]);
    assign outputs[8978] = (layer0_outputs[3147]) & ~(layer0_outputs[4045]);
    assign outputs[8979] = layer0_outputs[8916];
    assign outputs[8980] = layer0_outputs[7398];
    assign outputs[8981] = ~(layer0_outputs[7002]) | (layer0_outputs[4199]);
    assign outputs[8982] = layer0_outputs[5408];
    assign outputs[8983] = ~((layer0_outputs[8840]) | (layer0_outputs[3113]));
    assign outputs[8984] = ~(layer0_outputs[2287]);
    assign outputs[8985] = ~(layer0_outputs[8996]) | (layer0_outputs[7853]);
    assign outputs[8986] = ~(layer0_outputs[2697]) | (layer0_outputs[34]);
    assign outputs[8987] = ~(layer0_outputs[7524]);
    assign outputs[8988] = (layer0_outputs[2393]) & (layer0_outputs[8768]);
    assign outputs[8989] = ~((layer0_outputs[6405]) ^ (layer0_outputs[1308]));
    assign outputs[8990] = (layer0_outputs[6685]) ^ (layer0_outputs[9222]);
    assign outputs[8991] = layer0_outputs[7817];
    assign outputs[8992] = (layer0_outputs[8073]) & ~(layer0_outputs[8566]);
    assign outputs[8993] = layer0_outputs[6105];
    assign outputs[8994] = ~(layer0_outputs[6079]) | (layer0_outputs[4969]);
    assign outputs[8995] = ~(layer0_outputs[7080]) | (layer0_outputs[8427]);
    assign outputs[8996] = ~(layer0_outputs[4708]);
    assign outputs[8997] = (layer0_outputs[5605]) & ~(layer0_outputs[6764]);
    assign outputs[8998] = ~((layer0_outputs[5325]) ^ (layer0_outputs[3234]));
    assign outputs[8999] = ~(layer0_outputs[3476]);
    assign outputs[9000] = ~(layer0_outputs[1315]) | (layer0_outputs[9864]);
    assign outputs[9001] = ~(layer0_outputs[6799]);
    assign outputs[9002] = ~((layer0_outputs[7257]) ^ (layer0_outputs[4784]));
    assign outputs[9003] = ~(layer0_outputs[4087]);
    assign outputs[9004] = ~((layer0_outputs[2908]) & (layer0_outputs[4947]));
    assign outputs[9005] = ~((layer0_outputs[1134]) ^ (layer0_outputs[1904]));
    assign outputs[9006] = ~(layer0_outputs[2991]) | (layer0_outputs[9615]);
    assign outputs[9007] = ~(layer0_outputs[5961]) | (layer0_outputs[5871]);
    assign outputs[9008] = (layer0_outputs[8595]) ^ (layer0_outputs[8782]);
    assign outputs[9009] = (layer0_outputs[2733]) & ~(layer0_outputs[1928]);
    assign outputs[9010] = ~((layer0_outputs[6359]) ^ (layer0_outputs[7291]));
    assign outputs[9011] = ~(layer0_outputs[3435]);
    assign outputs[9012] = layer0_outputs[8865];
    assign outputs[9013] = ~(layer0_outputs[3557]) | (layer0_outputs[5915]);
    assign outputs[9014] = ~((layer0_outputs[3985]) ^ (layer0_outputs[5945]));
    assign outputs[9015] = (layer0_outputs[6622]) | (layer0_outputs[1607]);
    assign outputs[9016] = (layer0_outputs[2373]) ^ (layer0_outputs[7304]);
    assign outputs[9017] = ~((layer0_outputs[7534]) ^ (layer0_outputs[4107]));
    assign outputs[9018] = ~(layer0_outputs[1223]);
    assign outputs[9019] = ~((layer0_outputs[3411]) | (layer0_outputs[4106]));
    assign outputs[9020] = ~(layer0_outputs[3784]);
    assign outputs[9021] = (layer0_outputs[9078]) ^ (layer0_outputs[1216]);
    assign outputs[9022] = (layer0_outputs[6159]) | (layer0_outputs[7556]);
    assign outputs[9023] = (layer0_outputs[3818]) ^ (layer0_outputs[4465]);
    assign outputs[9024] = (layer0_outputs[3058]) | (layer0_outputs[7373]);
    assign outputs[9025] = (layer0_outputs[7787]) | (layer0_outputs[1625]);
    assign outputs[9026] = (layer0_outputs[334]) ^ (layer0_outputs[3900]);
    assign outputs[9027] = ~(layer0_outputs[5847]);
    assign outputs[9028] = layer0_outputs[8101];
    assign outputs[9029] = layer0_outputs[8068];
    assign outputs[9030] = (layer0_outputs[2849]) & ~(layer0_outputs[5608]);
    assign outputs[9031] = (layer0_outputs[3138]) ^ (layer0_outputs[3657]);
    assign outputs[9032] = (layer0_outputs[3179]) ^ (layer0_outputs[4480]);
    assign outputs[9033] = ~((layer0_outputs[3409]) & (layer0_outputs[5565]));
    assign outputs[9034] = ~(layer0_outputs[1841]);
    assign outputs[9035] = layer0_outputs[40];
    assign outputs[9036] = ~(layer0_outputs[8199]);
    assign outputs[9037] = ~((layer0_outputs[3422]) ^ (layer0_outputs[2579]));
    assign outputs[9038] = ~((layer0_outputs[10057]) | (layer0_outputs[2883]));
    assign outputs[9039] = (layer0_outputs[5309]) ^ (layer0_outputs[7401]);
    assign outputs[9040] = ~((layer0_outputs[5449]) ^ (layer0_outputs[2739]));
    assign outputs[9041] = (layer0_outputs[625]) & ~(layer0_outputs[796]);
    assign outputs[9042] = ~(layer0_outputs[2597]);
    assign outputs[9043] = ~(layer0_outputs[7047]) | (layer0_outputs[2492]);
    assign outputs[9044] = ~(layer0_outputs[2811]) | (layer0_outputs[4653]);
    assign outputs[9045] = ~((layer0_outputs[9135]) ^ (layer0_outputs[5417]));
    assign outputs[9046] = ~((layer0_outputs[4732]) ^ (layer0_outputs[1397]));
    assign outputs[9047] = ~((layer0_outputs[10035]) & (layer0_outputs[6354]));
    assign outputs[9048] = (layer0_outputs[507]) ^ (layer0_outputs[6117]);
    assign outputs[9049] = (layer0_outputs[9518]) ^ (layer0_outputs[6616]);
    assign outputs[9050] = (layer0_outputs[9353]) | (layer0_outputs[4130]);
    assign outputs[9051] = ~(layer0_outputs[9736]);
    assign outputs[9052] = (layer0_outputs[7886]) ^ (layer0_outputs[7079]);
    assign outputs[9053] = (layer0_outputs[166]) | (layer0_outputs[2811]);
    assign outputs[9054] = ~(layer0_outputs[2669]);
    assign outputs[9055] = ~((layer0_outputs[8663]) & (layer0_outputs[1221]));
    assign outputs[9056] = (layer0_outputs[2352]) | (layer0_outputs[6425]);
    assign outputs[9057] = ~(layer0_outputs[8739]) | (layer0_outputs[8113]);
    assign outputs[9058] = layer0_outputs[1200];
    assign outputs[9059] = 1'b1;
    assign outputs[9060] = ~((layer0_outputs[7739]) & (layer0_outputs[1081]));
    assign outputs[9061] = ~((layer0_outputs[1314]) ^ (layer0_outputs[2875]));
    assign outputs[9062] = (layer0_outputs[9899]) & ~(layer0_outputs[9673]);
    assign outputs[9063] = ~((layer0_outputs[249]) & (layer0_outputs[3172]));
    assign outputs[9064] = ~((layer0_outputs[6945]) & (layer0_outputs[6299]));
    assign outputs[9065] = (layer0_outputs[2042]) | (layer0_outputs[6576]);
    assign outputs[9066] = ~((layer0_outputs[7538]) | (layer0_outputs[5131]));
    assign outputs[9067] = layer0_outputs[1395];
    assign outputs[9068] = ~(layer0_outputs[6863]) | (layer0_outputs[6258]);
    assign outputs[9069] = layer0_outputs[354];
    assign outputs[9070] = ~(layer0_outputs[6033]);
    assign outputs[9071] = ~(layer0_outputs[6455]);
    assign outputs[9072] = (layer0_outputs[1544]) & ~(layer0_outputs[3569]);
    assign outputs[9073] = ~(layer0_outputs[2466]);
    assign outputs[9074] = ~((layer0_outputs[2528]) & (layer0_outputs[5478]));
    assign outputs[9075] = layer0_outputs[7871];
    assign outputs[9076] = ~(layer0_outputs[2113]);
    assign outputs[9077] = (layer0_outputs[6114]) ^ (layer0_outputs[8049]);
    assign outputs[9078] = ~(layer0_outputs[2088]) | (layer0_outputs[2830]);
    assign outputs[9079] = ~(layer0_outputs[3460]) | (layer0_outputs[10143]);
    assign outputs[9080] = (layer0_outputs[3494]) & ~(layer0_outputs[3442]);
    assign outputs[9081] = ~(layer0_outputs[8065]) | (layer0_outputs[475]);
    assign outputs[9082] = ~(layer0_outputs[748]);
    assign outputs[9083] = (layer0_outputs[1818]) & (layer0_outputs[2806]);
    assign outputs[9084] = ~((layer0_outputs[703]) & (layer0_outputs[9989]));
    assign outputs[9085] = ~((layer0_outputs[10081]) | (layer0_outputs[8162]));
    assign outputs[9086] = layer0_outputs[8347];
    assign outputs[9087] = layer0_outputs[4133];
    assign outputs[9088] = (layer0_outputs[1407]) ^ (layer0_outputs[8477]);
    assign outputs[9089] = ~((layer0_outputs[5688]) ^ (layer0_outputs[5242]));
    assign outputs[9090] = (layer0_outputs[7612]) & ~(layer0_outputs[4650]);
    assign outputs[9091] = ~(layer0_outputs[8682]);
    assign outputs[9092] = ~(layer0_outputs[3703]);
    assign outputs[9093] = ~(layer0_outputs[3107]);
    assign outputs[9094] = ~(layer0_outputs[4355]);
    assign outputs[9095] = (layer0_outputs[9526]) ^ (layer0_outputs[548]);
    assign outputs[9096] = layer0_outputs[7339];
    assign outputs[9097] = ~(layer0_outputs[3171]);
    assign outputs[9098] = ~(layer0_outputs[6489]) | (layer0_outputs[5715]);
    assign outputs[9099] = ~((layer0_outputs[1287]) ^ (layer0_outputs[856]));
    assign outputs[9100] = ~((layer0_outputs[1761]) ^ (layer0_outputs[3370]));
    assign outputs[9101] = ~(layer0_outputs[8657]);
    assign outputs[9102] = ~(layer0_outputs[9195]) | (layer0_outputs[4193]);
    assign outputs[9103] = (layer0_outputs[5162]) | (layer0_outputs[4218]);
    assign outputs[9104] = ~((layer0_outputs[4082]) | (layer0_outputs[9249]));
    assign outputs[9105] = layer0_outputs[8234];
    assign outputs[9106] = ~(layer0_outputs[1822]);
    assign outputs[9107] = ~((layer0_outputs[9189]) ^ (layer0_outputs[5432]));
    assign outputs[9108] = (layer0_outputs[5150]) ^ (layer0_outputs[256]);
    assign outputs[9109] = ~((layer0_outputs[908]) ^ (layer0_outputs[4030]));
    assign outputs[9110] = ~((layer0_outputs[4152]) | (layer0_outputs[1809]));
    assign outputs[9111] = ~(layer0_outputs[3575]) | (layer0_outputs[9358]);
    assign outputs[9112] = ~((layer0_outputs[4256]) | (layer0_outputs[4218]));
    assign outputs[9113] = ~((layer0_outputs[1034]) | (layer0_outputs[7025]));
    assign outputs[9114] = ~((layer0_outputs[6523]) | (layer0_outputs[3232]));
    assign outputs[9115] = ~((layer0_outputs[4698]) ^ (layer0_outputs[3835]));
    assign outputs[9116] = (layer0_outputs[8965]) & ~(layer0_outputs[5525]);
    assign outputs[9117] = ~((layer0_outputs[1708]) ^ (layer0_outputs[4849]));
    assign outputs[9118] = (layer0_outputs[8427]) | (layer0_outputs[191]);
    assign outputs[9119] = layer0_outputs[627];
    assign outputs[9120] = ~((layer0_outputs[489]) ^ (layer0_outputs[6821]));
    assign outputs[9121] = (layer0_outputs[5711]) ^ (layer0_outputs[2347]);
    assign outputs[9122] = (layer0_outputs[2984]) | (layer0_outputs[3152]);
    assign outputs[9123] = ~((layer0_outputs[1946]) ^ (layer0_outputs[7813]));
    assign outputs[9124] = (layer0_outputs[6196]) | (layer0_outputs[6284]);
    assign outputs[9125] = ~((layer0_outputs[5523]) & (layer0_outputs[8240]));
    assign outputs[9126] = ~(layer0_outputs[5017]) | (layer0_outputs[3944]);
    assign outputs[9127] = ~(layer0_outputs[7184]) | (layer0_outputs[8717]);
    assign outputs[9128] = layer0_outputs[8349];
    assign outputs[9129] = ~(layer0_outputs[6745]);
    assign outputs[9130] = ~((layer0_outputs[2846]) ^ (layer0_outputs[7468]));
    assign outputs[9131] = (layer0_outputs[7342]) & (layer0_outputs[5513]);
    assign outputs[9132] = (layer0_outputs[1474]) ^ (layer0_outputs[1622]);
    assign outputs[9133] = (layer0_outputs[9985]) ^ (layer0_outputs[2002]);
    assign outputs[9134] = (layer0_outputs[7118]) | (layer0_outputs[4870]);
    assign outputs[9135] = ~(layer0_outputs[7434]);
    assign outputs[9136] = (layer0_outputs[2819]) ^ (layer0_outputs[4264]);
    assign outputs[9137] = (layer0_outputs[8619]) & ~(layer0_outputs[8256]);
    assign outputs[9138] = layer0_outputs[2662];
    assign outputs[9139] = ~((layer0_outputs[9332]) ^ (layer0_outputs[8968]));
    assign outputs[9140] = ~(layer0_outputs[3144]);
    assign outputs[9141] = ~(layer0_outputs[1297]) | (layer0_outputs[5795]);
    assign outputs[9142] = ~(layer0_outputs[8454]);
    assign outputs[9143] = layer0_outputs[9153];
    assign outputs[9144] = layer0_outputs[1195];
    assign outputs[9145] = ~(layer0_outputs[3560]);
    assign outputs[9146] = layer0_outputs[10161];
    assign outputs[9147] = layer0_outputs[791];
    assign outputs[9148] = layer0_outputs[6089];
    assign outputs[9149] = (layer0_outputs[4812]) & (layer0_outputs[3453]);
    assign outputs[9150] = ~(layer0_outputs[9605]);
    assign outputs[9151] = ~((layer0_outputs[1447]) ^ (layer0_outputs[4582]));
    assign outputs[9152] = ~((layer0_outputs[2263]) ^ (layer0_outputs[3856]));
    assign outputs[9153] = (layer0_outputs[10216]) ^ (layer0_outputs[2097]);
    assign outputs[9154] = ~(layer0_outputs[9980]);
    assign outputs[9155] = layer0_outputs[4677];
    assign outputs[9156] = (layer0_outputs[7318]) & ~(layer0_outputs[4458]);
    assign outputs[9157] = ~(layer0_outputs[4606]);
    assign outputs[9158] = layer0_outputs[8820];
    assign outputs[9159] = ~(layer0_outputs[7734]);
    assign outputs[9160] = ~(layer0_outputs[6963]) | (layer0_outputs[116]);
    assign outputs[9161] = (layer0_outputs[552]) ^ (layer0_outputs[8737]);
    assign outputs[9162] = layer0_outputs[2658];
    assign outputs[9163] = ~((layer0_outputs[10203]) ^ (layer0_outputs[3410]));
    assign outputs[9164] = (layer0_outputs[1121]) & ~(layer0_outputs[2191]);
    assign outputs[9165] = ~(layer0_outputs[2155]);
    assign outputs[9166] = ~((layer0_outputs[7414]) & (layer0_outputs[6583]));
    assign outputs[9167] = ~(layer0_outputs[4957]);
    assign outputs[9168] = ~(layer0_outputs[542]);
    assign outputs[9169] = layer0_outputs[3040];
    assign outputs[9170] = (layer0_outputs[5259]) & ~(layer0_outputs[8138]);
    assign outputs[9171] = ~(layer0_outputs[1289]);
    assign outputs[9172] = 1'b1;
    assign outputs[9173] = layer0_outputs[9781];
    assign outputs[9174] = ~((layer0_outputs[1949]) | (layer0_outputs[6075]));
    assign outputs[9175] = (layer0_outputs[7579]) | (layer0_outputs[4375]);
    assign outputs[9176] = ~(layer0_outputs[2891]);
    assign outputs[9177] = layer0_outputs[8038];
    assign outputs[9178] = ~((layer0_outputs[1991]) ^ (layer0_outputs[8862]));
    assign outputs[9179] = layer0_outputs[5852];
    assign outputs[9180] = (layer0_outputs[7687]) ^ (layer0_outputs[3542]);
    assign outputs[9181] = (layer0_outputs[4056]) & ~(layer0_outputs[4975]);
    assign outputs[9182] = layer0_outputs[4411];
    assign outputs[9183] = (layer0_outputs[1295]) ^ (layer0_outputs[8615]);
    assign outputs[9184] = ~((layer0_outputs[2991]) ^ (layer0_outputs[1245]));
    assign outputs[9185] = (layer0_outputs[7238]) & ~(layer0_outputs[4558]);
    assign outputs[9186] = ~(layer0_outputs[9711]) | (layer0_outputs[5851]);
    assign outputs[9187] = (layer0_outputs[4673]) | (layer0_outputs[3769]);
    assign outputs[9188] = ~(layer0_outputs[5203]);
    assign outputs[9189] = layer0_outputs[9042];
    assign outputs[9190] = ~(layer0_outputs[3682]);
    assign outputs[9191] = (layer0_outputs[9426]) & (layer0_outputs[9796]);
    assign outputs[9192] = ~(layer0_outputs[7685]);
    assign outputs[9193] = ~(layer0_outputs[5406]);
    assign outputs[9194] = layer0_outputs[5592];
    assign outputs[9195] = ~(layer0_outputs[6131]);
    assign outputs[9196] = layer0_outputs[183];
    assign outputs[9197] = layer0_outputs[1660];
    assign outputs[9198] = layer0_outputs[3716];
    assign outputs[9199] = ~((layer0_outputs[2008]) ^ (layer0_outputs[4292]));
    assign outputs[9200] = layer0_outputs[9904];
    assign outputs[9201] = 1'b1;
    assign outputs[9202] = ~(layer0_outputs[8479]);
    assign outputs[9203] = layer0_outputs[8874];
    assign outputs[9204] = ~(layer0_outputs[2422]) | (layer0_outputs[5728]);
    assign outputs[9205] = (layer0_outputs[8214]) ^ (layer0_outputs[2570]);
    assign outputs[9206] = ~(layer0_outputs[8175]);
    assign outputs[9207] = (layer0_outputs[3048]) ^ (layer0_outputs[1062]);
    assign outputs[9208] = ~(layer0_outputs[1203]) | (layer0_outputs[4481]);
    assign outputs[9209] = (layer0_outputs[9087]) ^ (layer0_outputs[3353]);
    assign outputs[9210] = (layer0_outputs[1346]) ^ (layer0_outputs[1897]);
    assign outputs[9211] = (layer0_outputs[2338]) ^ (layer0_outputs[2004]);
    assign outputs[9212] = (layer0_outputs[7092]) ^ (layer0_outputs[5341]);
    assign outputs[9213] = (layer0_outputs[3558]) & ~(layer0_outputs[589]);
    assign outputs[9214] = ~(layer0_outputs[9354]);
    assign outputs[9215] = ~(layer0_outputs[5223]);
    assign outputs[9216] = layer0_outputs[7868];
    assign outputs[9217] = layer0_outputs[9670];
    assign outputs[9218] = ~((layer0_outputs[8092]) ^ (layer0_outputs[1684]));
    assign outputs[9219] = layer0_outputs[3637];
    assign outputs[9220] = ~(layer0_outputs[7194]);
    assign outputs[9221] = 1'b0;
    assign outputs[9222] = (layer0_outputs[4096]) & ~(layer0_outputs[8097]);
    assign outputs[9223] = layer0_outputs[9522];
    assign outputs[9224] = layer0_outputs[7461];
    assign outputs[9225] = ~((layer0_outputs[73]) & (layer0_outputs[6840]));
    assign outputs[9226] = layer0_outputs[4431];
    assign outputs[9227] = ~(layer0_outputs[3894]) | (layer0_outputs[5511]);
    assign outputs[9228] = ~((layer0_outputs[9483]) ^ (layer0_outputs[7133]));
    assign outputs[9229] = (layer0_outputs[4596]) & (layer0_outputs[1990]);
    assign outputs[9230] = ~((layer0_outputs[8681]) | (layer0_outputs[1645]));
    assign outputs[9231] = ~((layer0_outputs[7332]) & (layer0_outputs[941]));
    assign outputs[9232] = ~((layer0_outputs[6017]) | (layer0_outputs[3338]));
    assign outputs[9233] = (layer0_outputs[9093]) ^ (layer0_outputs[8132]);
    assign outputs[9234] = ~(layer0_outputs[3257]);
    assign outputs[9235] = ~(layer0_outputs[3846]);
    assign outputs[9236] = layer0_outputs[7616];
    assign outputs[9237] = ~((layer0_outputs[1260]) | (layer0_outputs[8376]));
    assign outputs[9238] = layer0_outputs[4155];
    assign outputs[9239] = ~(layer0_outputs[3044]);
    assign outputs[9240] = (layer0_outputs[3600]) ^ (layer0_outputs[10185]);
    assign outputs[9241] = (layer0_outputs[8576]) ^ (layer0_outputs[5025]);
    assign outputs[9242] = layer0_outputs[7492];
    assign outputs[9243] = (layer0_outputs[7952]) & ~(layer0_outputs[5343]);
    assign outputs[9244] = (layer0_outputs[1606]) ^ (layer0_outputs[9644]);
    assign outputs[9245] = layer0_outputs[4670];
    assign outputs[9246] = ~(layer0_outputs[485]) | (layer0_outputs[591]);
    assign outputs[9247] = ~(layer0_outputs[7183]);
    assign outputs[9248] = ~((layer0_outputs[10045]) ^ (layer0_outputs[8693]));
    assign outputs[9249] = (layer0_outputs[161]) | (layer0_outputs[7289]);
    assign outputs[9250] = layer0_outputs[8589];
    assign outputs[9251] = (layer0_outputs[1961]) & (layer0_outputs[5507]);
    assign outputs[9252] = (layer0_outputs[3072]) ^ (layer0_outputs[8582]);
    assign outputs[9253] = (layer0_outputs[7353]) ^ (layer0_outputs[6529]);
    assign outputs[9254] = (layer0_outputs[8508]) ^ (layer0_outputs[4358]);
    assign outputs[9255] = (layer0_outputs[2483]) & (layer0_outputs[5843]);
    assign outputs[9256] = layer0_outputs[363];
    assign outputs[9257] = ~(layer0_outputs[3095]);
    assign outputs[9258] = layer0_outputs[4768];
    assign outputs[9259] = ~(layer0_outputs[1950]);
    assign outputs[9260] = layer0_outputs[6088];
    assign outputs[9261] = ~((layer0_outputs[6313]) ^ (layer0_outputs[1211]));
    assign outputs[9262] = ~(layer0_outputs[9069]);
    assign outputs[9263] = layer0_outputs[2204];
    assign outputs[9264] = ~(layer0_outputs[5095]);
    assign outputs[9265] = layer0_outputs[3709];
    assign outputs[9266] = (layer0_outputs[5616]) & ~(layer0_outputs[2493]);
    assign outputs[9267] = ~((layer0_outputs[2543]) & (layer0_outputs[9557]));
    assign outputs[9268] = ~(layer0_outputs[2091]);
    assign outputs[9269] = (layer0_outputs[1635]) & (layer0_outputs[1240]);
    assign outputs[9270] = ~(layer0_outputs[3211]);
    assign outputs[9271] = (layer0_outputs[1650]) ^ (layer0_outputs[2249]);
    assign outputs[9272] = ~(layer0_outputs[2248]) | (layer0_outputs[4503]);
    assign outputs[9273] = ~(layer0_outputs[2358]);
    assign outputs[9274] = ~((layer0_outputs[5826]) | (layer0_outputs[7870]));
    assign outputs[9275] = (layer0_outputs[838]) ^ (layer0_outputs[3617]);
    assign outputs[9276] = ~((layer0_outputs[9057]) | (layer0_outputs[276]));
    assign outputs[9277] = ~(layer0_outputs[1996]) | (layer0_outputs[5855]);
    assign outputs[9278] = ~((layer0_outputs[689]) | (layer0_outputs[8816]));
    assign outputs[9279] = (layer0_outputs[7403]) & ~(layer0_outputs[4413]);
    assign outputs[9280] = (layer0_outputs[9961]) & ~(layer0_outputs[9425]);
    assign outputs[9281] = (layer0_outputs[2427]) | (layer0_outputs[4800]);
    assign outputs[9282] = (layer0_outputs[7189]) ^ (layer0_outputs[5284]);
    assign outputs[9283] = (layer0_outputs[3416]) ^ (layer0_outputs[4999]);
    assign outputs[9284] = ~(layer0_outputs[10237]);
    assign outputs[9285] = (layer0_outputs[6640]) & ~(layer0_outputs[1957]);
    assign outputs[9286] = (layer0_outputs[3116]) & (layer0_outputs[4542]);
    assign outputs[9287] = ~(layer0_outputs[5409]);
    assign outputs[9288] = ~(layer0_outputs[8293]);
    assign outputs[9289] = ~((layer0_outputs[5092]) | (layer0_outputs[6026]));
    assign outputs[9290] = ~(layer0_outputs[5939]);
    assign outputs[9291] = ~(layer0_outputs[275]);
    assign outputs[9292] = ~(layer0_outputs[2435]);
    assign outputs[9293] = ~((layer0_outputs[8640]) | (layer0_outputs[9077]));
    assign outputs[9294] = layer0_outputs[7489];
    assign outputs[9295] = layer0_outputs[9121];
    assign outputs[9296] = (layer0_outputs[2076]) ^ (layer0_outputs[8578]);
    assign outputs[9297] = (layer0_outputs[182]) & (layer0_outputs[1551]);
    assign outputs[9298] = ~(layer0_outputs[9898]);
    assign outputs[9299] = ~(layer0_outputs[637]);
    assign outputs[9300] = ~((layer0_outputs[7207]) | (layer0_outputs[1521]));
    assign outputs[9301] = ~(layer0_outputs[1656]);
    assign outputs[9302] = (layer0_outputs[2294]) & ~(layer0_outputs[4095]);
    assign outputs[9303] = ~(layer0_outputs[5548]);
    assign outputs[9304] = ~(layer0_outputs[8735]);
    assign outputs[9305] = ~(layer0_outputs[3446]);
    assign outputs[9306] = ~(layer0_outputs[7709]);
    assign outputs[9307] = (layer0_outputs[3398]) & ~(layer0_outputs[7406]);
    assign outputs[9308] = (layer0_outputs[135]) ^ (layer0_outputs[5073]);
    assign outputs[9309] = ~(layer0_outputs[2201]);
    assign outputs[9310] = ~((layer0_outputs[1597]) ^ (layer0_outputs[9082]));
    assign outputs[9311] = layer0_outputs[5980];
    assign outputs[9312] = ~((layer0_outputs[2836]) ^ (layer0_outputs[8790]));
    assign outputs[9313] = (layer0_outputs[9675]) & ~(layer0_outputs[6553]);
    assign outputs[9314] = ~((layer0_outputs[10089]) & (layer0_outputs[8303]));
    assign outputs[9315] = (layer0_outputs[2121]) ^ (layer0_outputs[7159]);
    assign outputs[9316] = (layer0_outputs[3614]) ^ (layer0_outputs[8129]);
    assign outputs[9317] = ~((layer0_outputs[5797]) ^ (layer0_outputs[4735]));
    assign outputs[9318] = (layer0_outputs[4634]) | (layer0_outputs[2026]);
    assign outputs[9319] = (layer0_outputs[2440]) ^ (layer0_outputs[1569]);
    assign outputs[9320] = ~(layer0_outputs[746]) | (layer0_outputs[3007]);
    assign outputs[9321] = ~((layer0_outputs[8136]) ^ (layer0_outputs[9995]));
    assign outputs[9322] = layer0_outputs[9773];
    assign outputs[9323] = ~(layer0_outputs[5690]);
    assign outputs[9324] = ~(layer0_outputs[6900]);
    assign outputs[9325] = ~((layer0_outputs[1759]) ^ (layer0_outputs[2508]));
    assign outputs[9326] = (layer0_outputs[7282]) & ~(layer0_outputs[6992]);
    assign outputs[9327] = ~((layer0_outputs[108]) | (layer0_outputs[1482]));
    assign outputs[9328] = ~(layer0_outputs[8904]);
    assign outputs[9329] = (layer0_outputs[4818]) & (layer0_outputs[9942]);
    assign outputs[9330] = ~(layer0_outputs[6882]);
    assign outputs[9331] = layer0_outputs[8343];
    assign outputs[9332] = ~((layer0_outputs[7482]) ^ (layer0_outputs[1964]));
    assign outputs[9333] = (layer0_outputs[9985]) & ~(layer0_outputs[9976]);
    assign outputs[9334] = layer0_outputs[2424];
    assign outputs[9335] = ~(layer0_outputs[314]) | (layer0_outputs[3307]);
    assign outputs[9336] = (layer0_outputs[7475]) & ~(layer0_outputs[8827]);
    assign outputs[9337] = ~(layer0_outputs[4229]);
    assign outputs[9338] = layer0_outputs[7599];
    assign outputs[9339] = layer0_outputs[9554];
    assign outputs[9340] = (layer0_outputs[1968]) & (layer0_outputs[6346]);
    assign outputs[9341] = ~(layer0_outputs[1890]);
    assign outputs[9342] = ~(layer0_outputs[1747]) | (layer0_outputs[4221]);
    assign outputs[9343] = ~(layer0_outputs[8533]);
    assign outputs[9344] = ~((layer0_outputs[4632]) ^ (layer0_outputs[8319]));
    assign outputs[9345] = (layer0_outputs[6999]) ^ (layer0_outputs[437]);
    assign outputs[9346] = ~((layer0_outputs[7320]) | (layer0_outputs[2856]));
    assign outputs[9347] = layer0_outputs[8528];
    assign outputs[9348] = ~((layer0_outputs[4755]) | (layer0_outputs[6704]));
    assign outputs[9349] = ~(layer0_outputs[1059]);
    assign outputs[9350] = ~(layer0_outputs[797]);
    assign outputs[9351] = ~((layer0_outputs[1646]) | (layer0_outputs[4705]));
    assign outputs[9352] = (layer0_outputs[2260]) | (layer0_outputs[5177]);
    assign outputs[9353] = (layer0_outputs[2825]) ^ (layer0_outputs[961]);
    assign outputs[9354] = ~(layer0_outputs[7137]);
    assign outputs[9355] = ~((layer0_outputs[5704]) ^ (layer0_outputs[7220]));
    assign outputs[9356] = (layer0_outputs[1917]) & (layer0_outputs[4057]);
    assign outputs[9357] = ~(layer0_outputs[5228]);
    assign outputs[9358] = ~(layer0_outputs[1984]) | (layer0_outputs[6977]);
    assign outputs[9359] = ~(layer0_outputs[9615]);
    assign outputs[9360] = (layer0_outputs[2855]) & ~(layer0_outputs[4144]);
    assign outputs[9361] = ~(layer0_outputs[7068]);
    assign outputs[9362] = ~(layer0_outputs[987]);
    assign outputs[9363] = ~((layer0_outputs[3747]) ^ (layer0_outputs[1084]));
    assign outputs[9364] = layer0_outputs[2978];
    assign outputs[9365] = layer0_outputs[1436];
    assign outputs[9366] = ~(layer0_outputs[9217]);
    assign outputs[9367] = layer0_outputs[6927];
    assign outputs[9368] = (layer0_outputs[6925]) & ~(layer0_outputs[8428]);
    assign outputs[9369] = ~(layer0_outputs[7389]);
    assign outputs[9370] = ~(layer0_outputs[601]);
    assign outputs[9371] = (layer0_outputs[8444]) & (layer0_outputs[8964]);
    assign outputs[9372] = ~(layer0_outputs[6469]) | (layer0_outputs[3731]);
    assign outputs[9373] = ~((layer0_outputs[2842]) | (layer0_outputs[987]));
    assign outputs[9374] = (layer0_outputs[5278]) & ~(layer0_outputs[6618]);
    assign outputs[9375] = (layer0_outputs[6718]) & ~(layer0_outputs[1027]);
    assign outputs[9376] = layer0_outputs[5207];
    assign outputs[9377] = layer0_outputs[2351];
    assign outputs[9378] = layer0_outputs[7468];
    assign outputs[9379] = ~(layer0_outputs[933]);
    assign outputs[9380] = ~((layer0_outputs[5992]) ^ (layer0_outputs[9134]));
    assign outputs[9381] = (layer0_outputs[6051]) ^ (layer0_outputs[7758]);
    assign outputs[9382] = layer0_outputs[9802];
    assign outputs[9383] = layer0_outputs[8587];
    assign outputs[9384] = ~(layer0_outputs[6746]) | (layer0_outputs[4203]);
    assign outputs[9385] = (layer0_outputs[1936]) ^ (layer0_outputs[5111]);
    assign outputs[9386] = layer0_outputs[3311];
    assign outputs[9387] = ~(layer0_outputs[29]);
    assign outputs[9388] = layer0_outputs[7333];
    assign outputs[9389] = ~((layer0_outputs[7355]) ^ (layer0_outputs[10174]));
    assign outputs[9390] = (layer0_outputs[1769]) & ~(layer0_outputs[5118]);
    assign outputs[9391] = ~(layer0_outputs[5236]);
    assign outputs[9392] = ~(layer0_outputs[1042]);
    assign outputs[9393] = ~(layer0_outputs[224]);
    assign outputs[9394] = layer0_outputs[10168];
    assign outputs[9395] = ~(layer0_outputs[2637]);
    assign outputs[9396] = ~((layer0_outputs[1203]) ^ (layer0_outputs[7804]));
    assign outputs[9397] = ~((layer0_outputs[9296]) ^ (layer0_outputs[5276]));
    assign outputs[9398] = layer0_outputs[814];
    assign outputs[9399] = layer0_outputs[2782];
    assign outputs[9400] = ~(layer0_outputs[1149]);
    assign outputs[9401] = (layer0_outputs[4282]) ^ (layer0_outputs[1570]);
    assign outputs[9402] = ~((layer0_outputs[409]) ^ (layer0_outputs[6808]));
    assign outputs[9403] = ~((layer0_outputs[9364]) ^ (layer0_outputs[3423]));
    assign outputs[9404] = (layer0_outputs[2932]) & ~(layer0_outputs[8658]);
    assign outputs[9405] = (layer0_outputs[6434]) & (layer0_outputs[5280]);
    assign outputs[9406] = ~((layer0_outputs[5016]) ^ (layer0_outputs[7528]));
    assign outputs[9407] = layer0_outputs[8011];
    assign outputs[9408] = ~((layer0_outputs[8342]) ^ (layer0_outputs[2363]));
    assign outputs[9409] = ~((layer0_outputs[2871]) | (layer0_outputs[6332]));
    assign outputs[9410] = layer0_outputs[3527];
    assign outputs[9411] = ~((layer0_outputs[2384]) & (layer0_outputs[10037]));
    assign outputs[9412] = ~((layer0_outputs[6636]) ^ (layer0_outputs[560]));
    assign outputs[9413] = ~((layer0_outputs[8331]) ^ (layer0_outputs[2576]));
    assign outputs[9414] = layer0_outputs[9234];
    assign outputs[9415] = (layer0_outputs[1142]) & ~(layer0_outputs[5649]);
    assign outputs[9416] = ~((layer0_outputs[1735]) | (layer0_outputs[1765]));
    assign outputs[9417] = ~((layer0_outputs[9479]) ^ (layer0_outputs[1986]));
    assign outputs[9418] = (layer0_outputs[4473]) & ~(layer0_outputs[1579]);
    assign outputs[9419] = ~((layer0_outputs[1471]) ^ (layer0_outputs[3158]));
    assign outputs[9420] = ~((layer0_outputs[7212]) & (layer0_outputs[7566]));
    assign outputs[9421] = layer0_outputs[1324];
    assign outputs[9422] = ~((layer0_outputs[1951]) | (layer0_outputs[707]));
    assign outputs[9423] = (layer0_outputs[4684]) & ~(layer0_outputs[1262]);
    assign outputs[9424] = (layer0_outputs[3051]) ^ (layer0_outputs[1892]);
    assign outputs[9425] = (layer0_outputs[1839]) ^ (layer0_outputs[229]);
    assign outputs[9426] = ~(layer0_outputs[7619]);
    assign outputs[9427] = ~(layer0_outputs[3108]);
    assign outputs[9428] = ~(layer0_outputs[8719]);
    assign outputs[9429] = (layer0_outputs[1268]) ^ (layer0_outputs[8207]);
    assign outputs[9430] = (layer0_outputs[2909]) & ~(layer0_outputs[2964]);
    assign outputs[9431] = (layer0_outputs[8151]) & ~(layer0_outputs[3104]);
    assign outputs[9432] = layer0_outputs[5066];
    assign outputs[9433] = layer0_outputs[2315];
    assign outputs[9434] = layer0_outputs[6792];
    assign outputs[9435] = layer0_outputs[4873];
    assign outputs[9436] = ~(layer0_outputs[1898]) | (layer0_outputs[8646]);
    assign outputs[9437] = (layer0_outputs[9549]) & ~(layer0_outputs[8783]);
    assign outputs[9438] = (layer0_outputs[6003]) & ~(layer0_outputs[9074]);
    assign outputs[9439] = ~(layer0_outputs[2598]);
    assign outputs[9440] = (layer0_outputs[3314]) ^ (layer0_outputs[131]);
    assign outputs[9441] = (layer0_outputs[776]) & ~(layer0_outputs[2378]);
    assign outputs[9442] = ~((layer0_outputs[8160]) ^ (layer0_outputs[1270]));
    assign outputs[9443] = ~(layer0_outputs[8404]);
    assign outputs[9444] = (layer0_outputs[9968]) & ~(layer0_outputs[5015]);
    assign outputs[9445] = (layer0_outputs[2009]) & ~(layer0_outputs[4500]);
    assign outputs[9446] = ~(layer0_outputs[7163]);
    assign outputs[9447] = layer0_outputs[6390];
    assign outputs[9448] = layer0_outputs[8087];
    assign outputs[9449] = (layer0_outputs[6826]) ^ (layer0_outputs[4491]);
    assign outputs[9450] = ~((layer0_outputs[6538]) | (layer0_outputs[279]));
    assign outputs[9451] = (layer0_outputs[1632]) ^ (layer0_outputs[3407]);
    assign outputs[9452] = ~(layer0_outputs[4777]);
    assign outputs[9453] = ~(layer0_outputs[3656]);
    assign outputs[9454] = ~((layer0_outputs[1379]) ^ (layer0_outputs[2645]));
    assign outputs[9455] = ~((layer0_outputs[9478]) ^ (layer0_outputs[9541]));
    assign outputs[9456] = ~((layer0_outputs[8538]) ^ (layer0_outputs[10022]));
    assign outputs[9457] = ~(layer0_outputs[1594]);
    assign outputs[9458] = ~((layer0_outputs[9671]) ^ (layer0_outputs[6431]));
    assign outputs[9459] = (layer0_outputs[5746]) & ~(layer0_outputs[7731]);
    assign outputs[9460] = (layer0_outputs[6477]) ^ (layer0_outputs[8553]);
    assign outputs[9461] = layer0_outputs[1303];
    assign outputs[9462] = (layer0_outputs[3077]) | (layer0_outputs[4964]);
    assign outputs[9463] = (layer0_outputs[3899]) ^ (layer0_outputs[9794]);
    assign outputs[9464] = layer0_outputs[8200];
    assign outputs[9465] = ~((layer0_outputs[6747]) | (layer0_outputs[953]));
    assign outputs[9466] = layer0_outputs[10095];
    assign outputs[9467] = ~((layer0_outputs[3931]) ^ (layer0_outputs[6087]));
    assign outputs[9468] = (layer0_outputs[5288]) ^ (layer0_outputs[8194]);
    assign outputs[9469] = (layer0_outputs[8896]) & ~(layer0_outputs[4214]);
    assign outputs[9470] = (layer0_outputs[656]) & ~(layer0_outputs[2775]);
    assign outputs[9471] = (layer0_outputs[2357]) & (layer0_outputs[3380]);
    assign outputs[9472] = ~((layer0_outputs[3851]) ^ (layer0_outputs[2057]));
    assign outputs[9473] = layer0_outputs[9907];
    assign outputs[9474] = ~(layer0_outputs[2046]) | (layer0_outputs[9967]);
    assign outputs[9475] = layer0_outputs[5101];
    assign outputs[9476] = (layer0_outputs[4142]) & (layer0_outputs[5944]);
    assign outputs[9477] = ~((layer0_outputs[3768]) ^ (layer0_outputs[5568]));
    assign outputs[9478] = ~(layer0_outputs[9786]);
    assign outputs[9479] = ~((layer0_outputs[355]) ^ (layer0_outputs[4759]));
    assign outputs[9480] = ~(layer0_outputs[7869]) | (layer0_outputs[9224]);
    assign outputs[9481] = ~((layer0_outputs[9783]) | (layer0_outputs[1396]));
    assign outputs[9482] = ~((layer0_outputs[4594]) ^ (layer0_outputs[517]));
    assign outputs[9483] = ~(layer0_outputs[4132]);
    assign outputs[9484] = layer0_outputs[4357];
    assign outputs[9485] = (layer0_outputs[2236]) & ~(layer0_outputs[4405]);
    assign outputs[9486] = ~((layer0_outputs[735]) & (layer0_outputs[10174]));
    assign outputs[9487] = ~(layer0_outputs[2262]);
    assign outputs[9488] = layer0_outputs[2720];
    assign outputs[9489] = layer0_outputs[5291];
    assign outputs[9490] = ~(layer0_outputs[3226]) | (layer0_outputs[9709]);
    assign outputs[9491] = (layer0_outputs[1885]) ^ (layer0_outputs[4198]);
    assign outputs[9492] = ~(layer0_outputs[6811]);
    assign outputs[9493] = (layer0_outputs[4264]) & ~(layer0_outputs[5340]);
    assign outputs[9494] = ~(layer0_outputs[5902]);
    assign outputs[9495] = ~(layer0_outputs[8626]);
    assign outputs[9496] = layer0_outputs[8043];
    assign outputs[9497] = layer0_outputs[3866];
    assign outputs[9498] = ~((layer0_outputs[4587]) | (layer0_outputs[1572]));
    assign outputs[9499] = ~(layer0_outputs[1522]);
    assign outputs[9500] = layer0_outputs[928];
    assign outputs[9501] = (layer0_outputs[2203]) & ~(layer0_outputs[6371]);
    assign outputs[9502] = ~((layer0_outputs[4413]) ^ (layer0_outputs[5772]));
    assign outputs[9503] = (layer0_outputs[4477]) & ~(layer0_outputs[6754]);
    assign outputs[9504] = layer0_outputs[6923];
    assign outputs[9505] = ~(layer0_outputs[9386]);
    assign outputs[9506] = ~(layer0_outputs[8493]);
    assign outputs[9507] = layer0_outputs[5980];
    assign outputs[9508] = layer0_outputs[3853];
    assign outputs[9509] = 1'b0;
    assign outputs[9510] = ~(layer0_outputs[7894]);
    assign outputs[9511] = layer0_outputs[7352];
    assign outputs[9512] = (layer0_outputs[3609]) ^ (layer0_outputs[3518]);
    assign outputs[9513] = 1'b0;
    assign outputs[9514] = ~(layer0_outputs[7030]) | (layer0_outputs[9190]);
    assign outputs[9515] = layer0_outputs[7880];
    assign outputs[9516] = ~((layer0_outputs[4208]) | (layer0_outputs[7850]));
    assign outputs[9517] = ~((layer0_outputs[3344]) | (layer0_outputs[6027]));
    assign outputs[9518] = layer0_outputs[453];
    assign outputs[9519] = ~(layer0_outputs[5726]) | (layer0_outputs[792]);
    assign outputs[9520] = ~(layer0_outputs[4899]) | (layer0_outputs[7536]);
    assign outputs[9521] = (layer0_outputs[8997]) & ~(layer0_outputs[32]);
    assign outputs[9522] = layer0_outputs[7746];
    assign outputs[9523] = layer0_outputs[5372];
    assign outputs[9524] = ~(layer0_outputs[7055]);
    assign outputs[9525] = (layer0_outputs[9654]) & ~(layer0_outputs[439]);
    assign outputs[9526] = layer0_outputs[6261];
    assign outputs[9527] = layer0_outputs[157];
    assign outputs[9528] = (layer0_outputs[6925]) & ~(layer0_outputs[4115]);
    assign outputs[9529] = layer0_outputs[9964];
    assign outputs[9530] = ~((layer0_outputs[980]) | (layer0_outputs[8277]));
    assign outputs[9531] = ~(layer0_outputs[9031]);
    assign outputs[9532] = ~((layer0_outputs[9887]) & (layer0_outputs[7018]));
    assign outputs[9533] = layer0_outputs[5742];
    assign outputs[9534] = (layer0_outputs[4444]) & ~(layer0_outputs[32]);
    assign outputs[9535] = layer0_outputs[3383];
    assign outputs[9536] = (layer0_outputs[9024]) & ~(layer0_outputs[2121]);
    assign outputs[9537] = ~((layer0_outputs[5185]) ^ (layer0_outputs[7452]));
    assign outputs[9538] = (layer0_outputs[7669]) ^ (layer0_outputs[7253]);
    assign outputs[9539] = ~((layer0_outputs[6439]) ^ (layer0_outputs[9054]));
    assign outputs[9540] = ~(layer0_outputs[10162]) | (layer0_outputs[8270]);
    assign outputs[9541] = (layer0_outputs[7822]) ^ (layer0_outputs[4561]);
    assign outputs[9542] = ~((layer0_outputs[6252]) ^ (layer0_outputs[7831]));
    assign outputs[9543] = ~((layer0_outputs[6769]) ^ (layer0_outputs[4269]));
    assign outputs[9544] = (layer0_outputs[8618]) | (layer0_outputs[7171]);
    assign outputs[9545] = ~(layer0_outputs[1498]);
    assign outputs[9546] = ~((layer0_outputs[9180]) | (layer0_outputs[2427]));
    assign outputs[9547] = ~((layer0_outputs[9209]) ^ (layer0_outputs[8879]));
    assign outputs[9548] = (layer0_outputs[1439]) & ~(layer0_outputs[2017]);
    assign outputs[9549] = ~(layer0_outputs[799]);
    assign outputs[9550] = ~(layer0_outputs[1269]) | (layer0_outputs[1478]);
    assign outputs[9551] = (layer0_outputs[1148]) & (layer0_outputs[7100]);
    assign outputs[9552] = ~(layer0_outputs[1706]);
    assign outputs[9553] = ~(layer0_outputs[7486]);
    assign outputs[9554] = (layer0_outputs[8917]) & ~(layer0_outputs[526]);
    assign outputs[9555] = (layer0_outputs[3376]) & ~(layer0_outputs[8636]);
    assign outputs[9556] = ~((layer0_outputs[6009]) | (layer0_outputs[643]));
    assign outputs[9557] = ~((layer0_outputs[5088]) | (layer0_outputs[9370]));
    assign outputs[9558] = ~((layer0_outputs[8198]) & (layer0_outputs[5102]));
    assign outputs[9559] = layer0_outputs[3982];
    assign outputs[9560] = layer0_outputs[120];
    assign outputs[9561] = (layer0_outputs[6291]) | (layer0_outputs[5633]);
    assign outputs[9562] = (layer0_outputs[1042]) ^ (layer0_outputs[6990]);
    assign outputs[9563] = layer0_outputs[3952];
    assign outputs[9564] = ~(layer0_outputs[627]);
    assign outputs[9565] = (layer0_outputs[4211]) & ~(layer0_outputs[3198]);
    assign outputs[9566] = (layer0_outputs[6316]) & ~(layer0_outputs[170]);
    assign outputs[9567] = layer0_outputs[8110];
    assign outputs[9568] = (layer0_outputs[8806]) ^ (layer0_outputs[7629]);
    assign outputs[9569] = (layer0_outputs[1965]) & ~(layer0_outputs[6274]);
    assign outputs[9570] = layer0_outputs[7937];
    assign outputs[9571] = ~(layer0_outputs[3003]);
    assign outputs[9572] = layer0_outputs[8642];
    assign outputs[9573] = ~((layer0_outputs[6666]) ^ (layer0_outputs[8597]));
    assign outputs[9574] = layer0_outputs[8168];
    assign outputs[9575] = ~(layer0_outputs[8980]);
    assign outputs[9576] = ~(layer0_outputs[1783]);
    assign outputs[9577] = ~((layer0_outputs[8767]) ^ (layer0_outputs[8195]));
    assign outputs[9578] = (layer0_outputs[3518]) & (layer0_outputs[3238]);
    assign outputs[9579] = (layer0_outputs[3805]) | (layer0_outputs[9566]);
    assign outputs[9580] = ~(layer0_outputs[9246]);
    assign outputs[9581] = ~(layer0_outputs[2718]);
    assign outputs[9582] = layer0_outputs[9195];
    assign outputs[9583] = layer0_outputs[6370];
    assign outputs[9584] = layer0_outputs[1814];
    assign outputs[9585] = layer0_outputs[4934];
    assign outputs[9586] = ~((layer0_outputs[2429]) ^ (layer0_outputs[9954]));
    assign outputs[9587] = (layer0_outputs[9648]) ^ (layer0_outputs[10119]);
    assign outputs[9588] = ~(layer0_outputs[4400]);
    assign outputs[9589] = ~((layer0_outputs[5176]) ^ (layer0_outputs[5666]));
    assign outputs[9590] = (layer0_outputs[7549]) & ~(layer0_outputs[3309]);
    assign outputs[9591] = ~((layer0_outputs[5825]) ^ (layer0_outputs[266]));
    assign outputs[9592] = layer0_outputs[2413];
    assign outputs[9593] = ~((layer0_outputs[4442]) ^ (layer0_outputs[138]));
    assign outputs[9594] = (layer0_outputs[8118]) ^ (layer0_outputs[985]);
    assign outputs[9595] = layer0_outputs[9974];
    assign outputs[9596] = (layer0_outputs[1301]) & ~(layer0_outputs[4208]);
    assign outputs[9597] = ~((layer0_outputs[4659]) ^ (layer0_outputs[4666]));
    assign outputs[9598] = (layer0_outputs[3099]) & ~(layer0_outputs[758]);
    assign outputs[9599] = layer0_outputs[3142];
    assign outputs[9600] = ~(layer0_outputs[1519]);
    assign outputs[9601] = (layer0_outputs[8015]) ^ (layer0_outputs[389]);
    assign outputs[9602] = (layer0_outputs[5029]) & (layer0_outputs[3031]);
    assign outputs[9603] = (layer0_outputs[6311]) ^ (layer0_outputs[7335]);
    assign outputs[9604] = (layer0_outputs[7416]) ^ (layer0_outputs[3188]);
    assign outputs[9605] = (layer0_outputs[9085]) & ~(layer0_outputs[7061]);
    assign outputs[9606] = ~(layer0_outputs[9417]);
    assign outputs[9607] = ~((layer0_outputs[5171]) & (layer0_outputs[9719]));
    assign outputs[9608] = ~((layer0_outputs[7373]) ^ (layer0_outputs[6159]));
    assign outputs[9609] = layer0_outputs[7015];
    assign outputs[9610] = (layer0_outputs[2442]) ^ (layer0_outputs[4036]);
    assign outputs[9611] = ~(layer0_outputs[10229]);
    assign outputs[9612] = ~(layer0_outputs[1967]);
    assign outputs[9613] = ~((layer0_outputs[10088]) ^ (layer0_outputs[8125]));
    assign outputs[9614] = ~((layer0_outputs[4568]) ^ (layer0_outputs[9706]));
    assign outputs[9615] = ~(layer0_outputs[5477]) | (layer0_outputs[3900]);
    assign outputs[9616] = layer0_outputs[6479];
    assign outputs[9617] = layer0_outputs[8960];
    assign outputs[9618] = (layer0_outputs[4955]) ^ (layer0_outputs[9492]);
    assign outputs[9619] = ~(layer0_outputs[7836]);
    assign outputs[9620] = (layer0_outputs[3352]) & (layer0_outputs[8653]);
    assign outputs[9621] = ~(layer0_outputs[8700]);
    assign outputs[9622] = ~(layer0_outputs[9680]);
    assign outputs[9623] = layer0_outputs[770];
    assign outputs[9624] = ~(layer0_outputs[7613]);
    assign outputs[9625] = (layer0_outputs[3277]) | (layer0_outputs[8173]);
    assign outputs[9626] = ~((layer0_outputs[7881]) ^ (layer0_outputs[2525]));
    assign outputs[9627] = ~((layer0_outputs[3916]) | (layer0_outputs[1298]));
    assign outputs[9628] = ~(layer0_outputs[2248]);
    assign outputs[9629] = layer0_outputs[2692];
    assign outputs[9630] = layer0_outputs[9915];
    assign outputs[9631] = layer0_outputs[24];
    assign outputs[9632] = ~(layer0_outputs[3436]);
    assign outputs[9633] = layer0_outputs[5360];
    assign outputs[9634] = (layer0_outputs[1043]) & ~(layer0_outputs[4645]);
    assign outputs[9635] = ~((layer0_outputs[6592]) ^ (layer0_outputs[2766]));
    assign outputs[9636] = ~(layer0_outputs[9366]);
    assign outputs[9637] = (layer0_outputs[8449]) & (layer0_outputs[2623]);
    assign outputs[9638] = (layer0_outputs[8536]) ^ (layer0_outputs[6400]);
    assign outputs[9639] = (layer0_outputs[5986]) & ~(layer0_outputs[864]);
    assign outputs[9640] = (layer0_outputs[1075]) ^ (layer0_outputs[1591]);
    assign outputs[9641] = (layer0_outputs[4437]) ^ (layer0_outputs[5190]);
    assign outputs[9642] = ~((layer0_outputs[8929]) ^ (layer0_outputs[7496]));
    assign outputs[9643] = (layer0_outputs[5603]) & (layer0_outputs[8933]);
    assign outputs[9644] = (layer0_outputs[3735]) ^ (layer0_outputs[618]);
    assign outputs[9645] = (layer0_outputs[8224]) & ~(layer0_outputs[9105]);
    assign outputs[9646] = ~(layer0_outputs[8967]);
    assign outputs[9647] = layer0_outputs[4018];
    assign outputs[9648] = ~((layer0_outputs[9626]) ^ (layer0_outputs[21]));
    assign outputs[9649] = (layer0_outputs[10158]) & ~(layer0_outputs[10220]);
    assign outputs[9650] = (layer0_outputs[4129]) ^ (layer0_outputs[2626]);
    assign outputs[9651] = ~((layer0_outputs[3392]) ^ (layer0_outputs[1562]));
    assign outputs[9652] = ~((layer0_outputs[2419]) & (layer0_outputs[277]));
    assign outputs[9653] = ~(layer0_outputs[1371]);
    assign outputs[9654] = layer0_outputs[763];
    assign outputs[9655] = ~(layer0_outputs[6538]);
    assign outputs[9656] = ~(layer0_outputs[9445]);
    assign outputs[9657] = layer0_outputs[6934];
    assign outputs[9658] = layer0_outputs[1];
    assign outputs[9659] = (layer0_outputs[6822]) & (layer0_outputs[530]);
    assign outputs[9660] = ~(layer0_outputs[3223]);
    assign outputs[9661] = ~(layer0_outputs[8758]);
    assign outputs[9662] = (layer0_outputs[8117]) ^ (layer0_outputs[7303]);
    assign outputs[9663] = (layer0_outputs[8261]) & (layer0_outputs[4279]);
    assign outputs[9664] = (layer0_outputs[1279]) ^ (layer0_outputs[5239]);
    assign outputs[9665] = ~((layer0_outputs[8728]) ^ (layer0_outputs[6283]));
    assign outputs[9666] = ~(layer0_outputs[2863]);
    assign outputs[9667] = (layer0_outputs[3513]) & ~(layer0_outputs[8757]);
    assign outputs[9668] = (layer0_outputs[7536]) & ~(layer0_outputs[3038]);
    assign outputs[9669] = ~(layer0_outputs[704]);
    assign outputs[9670] = (layer0_outputs[2486]) ^ (layer0_outputs[2802]);
    assign outputs[9671] = layer0_outputs[6888];
    assign outputs[9672] = ~(layer0_outputs[2813]);
    assign outputs[9673] = ~(layer0_outputs[5823]) | (layer0_outputs[9435]);
    assign outputs[9674] = (layer0_outputs[5349]) ^ (layer0_outputs[10058]);
    assign outputs[9675] = layer0_outputs[710];
    assign outputs[9676] = layer0_outputs[9957];
    assign outputs[9677] = layer0_outputs[8788];
    assign outputs[9678] = layer0_outputs[501];
    assign outputs[9679] = (layer0_outputs[7393]) & ~(layer0_outputs[6442]);
    assign outputs[9680] = (layer0_outputs[7333]) & ~(layer0_outputs[8891]);
    assign outputs[9681] = ~(layer0_outputs[8096]);
    assign outputs[9682] = ~(layer0_outputs[10068]);
    assign outputs[9683] = ~((layer0_outputs[2143]) ^ (layer0_outputs[7737]));
    assign outputs[9684] = ~((layer0_outputs[3431]) ^ (layer0_outputs[201]));
    assign outputs[9685] = ~((layer0_outputs[6637]) ^ (layer0_outputs[3396]));
    assign outputs[9686] = ~((layer0_outputs[8398]) | (layer0_outputs[7754]));
    assign outputs[9687] = ~((layer0_outputs[148]) | (layer0_outputs[8995]));
    assign outputs[9688] = ~(layer0_outputs[6618]) | (layer0_outputs[8981]);
    assign outputs[9689] = ~(layer0_outputs[1668]);
    assign outputs[9690] = (layer0_outputs[1600]) ^ (layer0_outputs[6409]);
    assign outputs[9691] = ~(layer0_outputs[2685]) | (layer0_outputs[1614]);
    assign outputs[9692] = ~(layer0_outputs[6603]);
    assign outputs[9693] = ~(layer0_outputs[1043]) | (layer0_outputs[4863]);
    assign outputs[9694] = ~(layer0_outputs[4210]);
    assign outputs[9695] = layer0_outputs[7663];
    assign outputs[9696] = ~(layer0_outputs[8992]);
    assign outputs[9697] = ~((layer0_outputs[3474]) | (layer0_outputs[6605]));
    assign outputs[9698] = layer0_outputs[54];
    assign outputs[9699] = ~(layer0_outputs[2445]);
    assign outputs[9700] = ~((layer0_outputs[8212]) ^ (layer0_outputs[2259]));
    assign outputs[9701] = (layer0_outputs[770]) & ~(layer0_outputs[8001]);
    assign outputs[9702] = layer0_outputs[6822];
    assign outputs[9703] = (layer0_outputs[8413]) | (layer0_outputs[9355]);
    assign outputs[9704] = layer0_outputs[9610];
    assign outputs[9705] = ~(layer0_outputs[7535]);
    assign outputs[9706] = ~(layer0_outputs[5978]);
    assign outputs[9707] = (layer0_outputs[4906]) ^ (layer0_outputs[1708]);
    assign outputs[9708] = (layer0_outputs[6233]) & (layer0_outputs[7408]);
    assign outputs[9709] = (layer0_outputs[1335]) & (layer0_outputs[5687]);
    assign outputs[9710] = (layer0_outputs[4194]) & (layer0_outputs[4649]);
    assign outputs[9711] = layer0_outputs[6039];
    assign outputs[9712] = ~(layer0_outputs[9698]);
    assign outputs[9713] = layer0_outputs[4266];
    assign outputs[9714] = ~(layer0_outputs[865]);
    assign outputs[9715] = (layer0_outputs[8759]) & ~(layer0_outputs[5306]);
    assign outputs[9716] = ~((layer0_outputs[1299]) & (layer0_outputs[3001]));
    assign outputs[9717] = ~(layer0_outputs[2111]);
    assign outputs[9718] = ~(layer0_outputs[7809]);
    assign outputs[9719] = ~((layer0_outputs[4168]) ^ (layer0_outputs[2602]));
    assign outputs[9720] = (layer0_outputs[7778]) & ~(layer0_outputs[5238]);
    assign outputs[9721] = (layer0_outputs[8008]) ^ (layer0_outputs[4124]);
    assign outputs[9722] = layer0_outputs[3608];
    assign outputs[9723] = ~(layer0_outputs[1209]);
    assign outputs[9724] = ~((layer0_outputs[7490]) | (layer0_outputs[4126]));
    assign outputs[9725] = layer0_outputs[10030];
    assign outputs[9726] = ~(layer0_outputs[6784]);
    assign outputs[9727] = ~(layer0_outputs[7790]);
    assign outputs[9728] = layer0_outputs[1357];
    assign outputs[9729] = layer0_outputs[4384];
    assign outputs[9730] = (layer0_outputs[8236]) & ~(layer0_outputs[5940]);
    assign outputs[9731] = (layer0_outputs[1533]) & ~(layer0_outputs[590]);
    assign outputs[9732] = layer0_outputs[733];
    assign outputs[9733] = layer0_outputs[8062];
    assign outputs[9734] = layer0_outputs[7557];
    assign outputs[9735] = ~(layer0_outputs[7976]);
    assign outputs[9736] = layer0_outputs[2945];
    assign outputs[9737] = ~((layer0_outputs[3005]) ^ (layer0_outputs[9862]));
    assign outputs[9738] = ~((layer0_outputs[6729]) & (layer0_outputs[9170]));
    assign outputs[9739] = layer0_outputs[3372];
    assign outputs[9740] = ~((layer0_outputs[1002]) ^ (layer0_outputs[1973]));
    assign outputs[9741] = (layer0_outputs[1028]) & ~(layer0_outputs[2380]);
    assign outputs[9742] = layer0_outputs[4740];
    assign outputs[9743] = (layer0_outputs[2094]) ^ (layer0_outputs[7126]);
    assign outputs[9744] = layer0_outputs[4751];
    assign outputs[9745] = (layer0_outputs[4390]) ^ (layer0_outputs[2770]);
    assign outputs[9746] = (layer0_outputs[6837]) & ~(layer0_outputs[6035]);
    assign outputs[9747] = ~(layer0_outputs[4997]);
    assign outputs[9748] = layer0_outputs[5782];
    assign outputs[9749] = ~(layer0_outputs[3196]);
    assign outputs[9750] = ~(layer0_outputs[2152]);
    assign outputs[9751] = layer0_outputs[7307];
    assign outputs[9752] = ~(layer0_outputs[3981]);
    assign outputs[9753] = layer0_outputs[8571];
    assign outputs[9754] = ~(layer0_outputs[7882]);
    assign outputs[9755] = (layer0_outputs[7537]) | (layer0_outputs[8799]);
    assign outputs[9756] = (layer0_outputs[5660]) & (layer0_outputs[2003]);
    assign outputs[9757] = (layer0_outputs[3780]) ^ (layer0_outputs[9701]);
    assign outputs[9758] = layer0_outputs[481];
    assign outputs[9759] = ~((layer0_outputs[5357]) | (layer0_outputs[913]));
    assign outputs[9760] = ~(layer0_outputs[2656]);
    assign outputs[9761] = (layer0_outputs[3895]) & ~(layer0_outputs[4098]);
    assign outputs[9762] = ~((layer0_outputs[8802]) | (layer0_outputs[779]));
    assign outputs[9763] = (layer0_outputs[3830]) ^ (layer0_outputs[6624]);
    assign outputs[9764] = ~((layer0_outputs[2572]) ^ (layer0_outputs[7128]));
    assign outputs[9765] = (layer0_outputs[2596]) ^ (layer0_outputs[1695]);
    assign outputs[9766] = (layer0_outputs[9566]) & ~(layer0_outputs[2540]);
    assign outputs[9767] = layer0_outputs[2434];
    assign outputs[9768] = layer0_outputs[1845];
    assign outputs[9769] = ~(layer0_outputs[2714]);
    assign outputs[9770] = ~(layer0_outputs[2874]);
    assign outputs[9771] = ~((layer0_outputs[739]) | (layer0_outputs[3375]));
    assign outputs[9772] = (layer0_outputs[1752]) & ~(layer0_outputs[3946]);
    assign outputs[9773] = (layer0_outputs[1361]) & ~(layer0_outputs[3361]);
    assign outputs[9774] = (layer0_outputs[2628]) ^ (layer0_outputs[3988]);
    assign outputs[9775] = ~(layer0_outputs[4705]);
    assign outputs[9776] = ~(layer0_outputs[4823]);
    assign outputs[9777] = layer0_outputs[3039];
    assign outputs[9778] = (layer0_outputs[1575]) & ~(layer0_outputs[9363]);
    assign outputs[9779] = ~((layer0_outputs[5182]) ^ (layer0_outputs[9899]));
    assign outputs[9780] = layer0_outputs[5361];
    assign outputs[9781] = layer0_outputs[5537];
    assign outputs[9782] = ~(layer0_outputs[3240]);
    assign outputs[9783] = ~(layer0_outputs[9050]);
    assign outputs[9784] = layer0_outputs[9172];
    assign outputs[9785] = ~((layer0_outputs[8650]) | (layer0_outputs[8265]));
    assign outputs[9786] = layer0_outputs[1665];
    assign outputs[9787] = (layer0_outputs[112]) & ~(layer0_outputs[2845]);
    assign outputs[9788] = (layer0_outputs[4128]) & (layer0_outputs[15]);
    assign outputs[9789] = ~((layer0_outputs[6980]) & (layer0_outputs[7764]));
    assign outputs[9790] = (layer0_outputs[9291]) | (layer0_outputs[3054]);
    assign outputs[9791] = layer0_outputs[6110];
    assign outputs[9792] = ~(layer0_outputs[1120]) | (layer0_outputs[5544]);
    assign outputs[9793] = ~((layer0_outputs[6279]) & (layer0_outputs[5744]));
    assign outputs[9794] = (layer0_outputs[3221]) ^ (layer0_outputs[4392]);
    assign outputs[9795] = (layer0_outputs[5551]) & ~(layer0_outputs[470]);
    assign outputs[9796] = ~(layer0_outputs[9827]);
    assign outputs[9797] = layer0_outputs[2815];
    assign outputs[9798] = (layer0_outputs[2444]) & ~(layer0_outputs[3536]);
    assign outputs[9799] = (layer0_outputs[207]) ^ (layer0_outputs[8698]);
    assign outputs[9800] = (layer0_outputs[7237]) & ~(layer0_outputs[7330]);
    assign outputs[9801] = layer0_outputs[8534];
    assign outputs[9802] = ~((layer0_outputs[8268]) ^ (layer0_outputs[1623]));
    assign outputs[9803] = (layer0_outputs[4855]) & (layer0_outputs[6201]);
    assign outputs[9804] = ~(layer0_outputs[7539]);
    assign outputs[9805] = ~((layer0_outputs[5007]) ^ (layer0_outputs[6324]));
    assign outputs[9806] = ~((layer0_outputs[8069]) | (layer0_outputs[1256]));
    assign outputs[9807] = ~(layer0_outputs[5933]);
    assign outputs[9808] = ~(layer0_outputs[7505]);
    assign outputs[9809] = ~(layer0_outputs[3469]);
    assign outputs[9810] = (layer0_outputs[9885]) | (layer0_outputs[3788]);
    assign outputs[9811] = (layer0_outputs[6850]) & ~(layer0_outputs[1895]);
    assign outputs[9812] = ~(layer0_outputs[7928]);
    assign outputs[9813] = ~(layer0_outputs[6221]);
    assign outputs[9814] = layer0_outputs[268];
    assign outputs[9815] = ~(layer0_outputs[7329]);
    assign outputs[9816] = (layer0_outputs[5151]) & ~(layer0_outputs[2189]);
    assign outputs[9817] = layer0_outputs[482];
    assign outputs[9818] = 1'b0;
    assign outputs[9819] = (layer0_outputs[7862]) & ~(layer0_outputs[3437]);
    assign outputs[9820] = ~(layer0_outputs[6323]);
    assign outputs[9821] = ~(layer0_outputs[3855]) | (layer0_outputs[352]);
    assign outputs[9822] = ~((layer0_outputs[2638]) ^ (layer0_outputs[3526]));
    assign outputs[9823] = ~(layer0_outputs[292]);
    assign outputs[9824] = ~(layer0_outputs[1821]);
    assign outputs[9825] = ~((layer0_outputs[3400]) | (layer0_outputs[8907]));
    assign outputs[9826] = ~(layer0_outputs[5897]);
    assign outputs[9827] = (layer0_outputs[8791]) | (layer0_outputs[8640]);
    assign outputs[9828] = ~(layer0_outputs[8899]);
    assign outputs[9829] = ~((layer0_outputs[2698]) ^ (layer0_outputs[8422]));
    assign outputs[9830] = (layer0_outputs[6698]) & (layer0_outputs[6929]);
    assign outputs[9831] = layer0_outputs[9517];
    assign outputs[9832] = ~(layer0_outputs[1725]) | (layer0_outputs[8509]);
    assign outputs[9833] = layer0_outputs[2516];
    assign outputs[9834] = layer0_outputs[203];
    assign outputs[9835] = ~(layer0_outputs[2369]) | (layer0_outputs[8210]);
    assign outputs[9836] = ~(layer0_outputs[8005]) | (layer0_outputs[3996]);
    assign outputs[9837] = layer0_outputs[5183];
    assign outputs[9838] = layer0_outputs[2072];
    assign outputs[9839] = ~(layer0_outputs[8064]);
    assign outputs[9840] = (layer0_outputs[8976]) & (layer0_outputs[1375]);
    assign outputs[9841] = ~((layer0_outputs[7932]) ^ (layer0_outputs[266]));
    assign outputs[9842] = (layer0_outputs[4668]) ^ (layer0_outputs[6983]);
    assign outputs[9843] = ~((layer0_outputs[7331]) ^ (layer0_outputs[10208]));
    assign outputs[9844] = (layer0_outputs[5102]) ^ (layer0_outputs[4029]);
    assign outputs[9845] = ~((layer0_outputs[8576]) & (layer0_outputs[9690]));
    assign outputs[9846] = (layer0_outputs[6263]) & ~(layer0_outputs[2463]);
    assign outputs[9847] = ~((layer0_outputs[6910]) ^ (layer0_outputs[2349]));
    assign outputs[9848] = ~(layer0_outputs[8710]) | (layer0_outputs[2977]);
    assign outputs[9849] = layer0_outputs[474];
    assign outputs[9850] = ~(layer0_outputs[6910]);
    assign outputs[9851] = ~((layer0_outputs[10157]) | (layer0_outputs[4385]));
    assign outputs[9852] = ~(layer0_outputs[1210]);
    assign outputs[9853] = ~(layer0_outputs[7577]);
    assign outputs[9854] = ~(layer0_outputs[4919]) | (layer0_outputs[7172]);
    assign outputs[9855] = (layer0_outputs[7502]) ^ (layer0_outputs[3875]);
    assign outputs[9856] = ~(layer0_outputs[7126]);
    assign outputs[9857] = (layer0_outputs[2981]) ^ (layer0_outputs[3623]);
    assign outputs[9858] = (layer0_outputs[4401]) & (layer0_outputs[6564]);
    assign outputs[9859] = ~((layer0_outputs[9381]) | (layer0_outputs[9211]));
    assign outputs[9860] = ~((layer0_outputs[6448]) ^ (layer0_outputs[5920]));
    assign outputs[9861] = layer0_outputs[3521];
    assign outputs[9862] = ~(layer0_outputs[5199]);
    assign outputs[9863] = ~(layer0_outputs[1473]);
    assign outputs[9864] = layer0_outputs[9171];
    assign outputs[9865] = ~((layer0_outputs[9196]) & (layer0_outputs[877]));
    assign outputs[9866] = layer0_outputs[1389];
    assign outputs[9867] = (layer0_outputs[10037]) & ~(layer0_outputs[3779]);
    assign outputs[9868] = ~((layer0_outputs[902]) ^ (layer0_outputs[9852]));
    assign outputs[9869] = (layer0_outputs[710]) & ~(layer0_outputs[5158]);
    assign outputs[9870] = ~((layer0_outputs[7887]) ^ (layer0_outputs[6244]));
    assign outputs[9871] = (layer0_outputs[9019]) ^ (layer0_outputs[114]);
    assign outputs[9872] = (layer0_outputs[4237]) ^ (layer0_outputs[5996]);
    assign outputs[9873] = ~(layer0_outputs[4126]);
    assign outputs[9874] = ~(layer0_outputs[6310]);
    assign outputs[9875] = ~((layer0_outputs[5627]) ^ (layer0_outputs[6309]));
    assign outputs[9876] = (layer0_outputs[8417]) | (layer0_outputs[3553]);
    assign outputs[9877] = layer0_outputs[6654];
    assign outputs[9878] = ~(layer0_outputs[9419]) | (layer0_outputs[5263]);
    assign outputs[9879] = (layer0_outputs[546]) ^ (layer0_outputs[5126]);
    assign outputs[9880] = (layer0_outputs[9339]) | (layer0_outputs[463]);
    assign outputs[9881] = ~(layer0_outputs[4120]);
    assign outputs[9882] = (layer0_outputs[8511]) ^ (layer0_outputs[927]);
    assign outputs[9883] = (layer0_outputs[2036]) & ~(layer0_outputs[4826]);
    assign outputs[9884] = layer0_outputs[9464];
    assign outputs[9885] = ~(layer0_outputs[7802]);
    assign outputs[9886] = ~((layer0_outputs[100]) ^ (layer0_outputs[129]));
    assign outputs[9887] = ~(layer0_outputs[5054]);
    assign outputs[9888] = (layer0_outputs[1835]) ^ (layer0_outputs[4368]);
    assign outputs[9889] = ~((layer0_outputs[3730]) ^ (layer0_outputs[7559]));
    assign outputs[9890] = layer0_outputs[5046];
    assign outputs[9891] = (layer0_outputs[1818]) & ~(layer0_outputs[5158]);
    assign outputs[9892] = (layer0_outputs[6230]) & ~(layer0_outputs[8041]);
    assign outputs[9893] = (layer0_outputs[3230]) & ~(layer0_outputs[3237]);
    assign outputs[9894] = layer0_outputs[6179];
    assign outputs[9895] = layer0_outputs[30];
    assign outputs[9896] = layer0_outputs[1108];
    assign outputs[9897] = ~((layer0_outputs[6561]) ^ (layer0_outputs[1680]));
    assign outputs[9898] = (layer0_outputs[2061]) | (layer0_outputs[4035]);
    assign outputs[9899] = (layer0_outputs[6527]) & (layer0_outputs[9897]);
    assign outputs[9900] = layer0_outputs[9415];
    assign outputs[9901] = (layer0_outputs[4253]) ^ (layer0_outputs[1172]);
    assign outputs[9902] = ~(layer0_outputs[2137]);
    assign outputs[9903] = ~(layer0_outputs[4288]);
    assign outputs[9904] = layer0_outputs[4727];
    assign outputs[9905] = ~(layer0_outputs[4598]);
    assign outputs[9906] = (layer0_outputs[3063]) ^ (layer0_outputs[5591]);
    assign outputs[9907] = (layer0_outputs[5338]) ^ (layer0_outputs[2923]);
    assign outputs[9908] = (layer0_outputs[9548]) & ~(layer0_outputs[1238]);
    assign outputs[9909] = layer0_outputs[8089];
    assign outputs[9910] = (layer0_outputs[8152]) ^ (layer0_outputs[8972]);
    assign outputs[9911] = (layer0_outputs[7231]) & ~(layer0_outputs[8510]);
    assign outputs[9912] = (layer0_outputs[1375]) & ~(layer0_outputs[9311]);
    assign outputs[9913] = (layer0_outputs[8078]) & ~(layer0_outputs[5197]);
    assign outputs[9914] = ~(layer0_outputs[990]);
    assign outputs[9915] = ~(layer0_outputs[8268]);
    assign outputs[9916] = ~(layer0_outputs[9046]);
    assign outputs[9917] = 1'b1;
    assign outputs[9918] = ~((layer0_outputs[1565]) | (layer0_outputs[2887]));
    assign outputs[9919] = (layer0_outputs[2624]) & ~(layer0_outputs[6367]);
    assign outputs[9920] = ~((layer0_outputs[8431]) | (layer0_outputs[5713]));
    assign outputs[9921] = ~((layer0_outputs[7682]) ^ (layer0_outputs[5534]));
    assign outputs[9922] = ~((layer0_outputs[3902]) ^ (layer0_outputs[575]));
    assign outputs[9923] = ~(layer0_outputs[2868]);
    assign outputs[9924] = ~(layer0_outputs[1353]);
    assign outputs[9925] = ~((layer0_outputs[6115]) | (layer0_outputs[2935]));
    assign outputs[9926] = ~(layer0_outputs[1697]);
    assign outputs[9927] = 1'b0;
    assign outputs[9928] = ~(layer0_outputs[9375]);
    assign outputs[9929] = (layer0_outputs[9511]) & (layer0_outputs[9150]);
    assign outputs[9930] = ~((layer0_outputs[3346]) | (layer0_outputs[8631]));
    assign outputs[9931] = (layer0_outputs[5534]) & ~(layer0_outputs[7594]);
    assign outputs[9932] = ~((layer0_outputs[1463]) ^ (layer0_outputs[259]));
    assign outputs[9933] = (layer0_outputs[3304]) & ~(layer0_outputs[542]);
    assign outputs[9934] = (layer0_outputs[1728]) & ~(layer0_outputs[7170]);
    assign outputs[9935] = ~(layer0_outputs[6393]);
    assign outputs[9936] = ~(layer0_outputs[2988]);
    assign outputs[9937] = ~(layer0_outputs[6639]);
    assign outputs[9938] = (layer0_outputs[2401]) & ~(layer0_outputs[2941]);
    assign outputs[9939] = layer0_outputs[1806];
    assign outputs[9940] = ~((layer0_outputs[9665]) ^ (layer0_outputs[8098]));
    assign outputs[9941] = (layer0_outputs[869]) & ~(layer0_outputs[1620]);
    assign outputs[9942] = (layer0_outputs[855]) & ~(layer0_outputs[8091]);
    assign outputs[9943] = ~(layer0_outputs[1473]);
    assign outputs[9944] = layer0_outputs[6579];
    assign outputs[9945] = ~((layer0_outputs[9294]) ^ (layer0_outputs[2037]));
    assign outputs[9946] = layer0_outputs[1599];
    assign outputs[9947] = ~((layer0_outputs[8486]) | (layer0_outputs[8807]));
    assign outputs[9948] = (layer0_outputs[1038]) | (layer0_outputs[4564]);
    assign outputs[9949] = 1'b0;
    assign outputs[9950] = (layer0_outputs[4454]) ^ (layer0_outputs[10101]);
    assign outputs[9951] = ~((layer0_outputs[9745]) ^ (layer0_outputs[5076]));
    assign outputs[9952] = (layer0_outputs[4245]) & ~(layer0_outputs[10098]);
    assign outputs[9953] = (layer0_outputs[7262]) & ~(layer0_outputs[8209]);
    assign outputs[9954] = ~(layer0_outputs[1465]);
    assign outputs[9955] = ~((layer0_outputs[7387]) | (layer0_outputs[7258]));
    assign outputs[9956] = (layer0_outputs[4317]) ^ (layer0_outputs[3761]);
    assign outputs[9957] = ~((layer0_outputs[1510]) | (layer0_outputs[1883]));
    assign outputs[9958] = (layer0_outputs[7700]) & (layer0_outputs[7230]);
    assign outputs[9959] = layer0_outputs[7561];
    assign outputs[9960] = (layer0_outputs[8281]) ^ (layer0_outputs[7410]);
    assign outputs[9961] = ~((layer0_outputs[9027]) | (layer0_outputs[669]));
    assign outputs[9962] = (layer0_outputs[6300]) & ~(layer0_outputs[4838]);
    assign outputs[9963] = (layer0_outputs[8018]) & ~(layer0_outputs[7368]);
    assign outputs[9964] = ~(layer0_outputs[3026]) | (layer0_outputs[7607]);
    assign outputs[9965] = layer0_outputs[4024];
    assign outputs[9966] = ~((layer0_outputs[8728]) ^ (layer0_outputs[8871]));
    assign outputs[9967] = layer0_outputs[343];
    assign outputs[9968] = (layer0_outputs[4461]) & ~(layer0_outputs[7117]);
    assign outputs[9969] = ~((layer0_outputs[4140]) ^ (layer0_outputs[3535]));
    assign outputs[9970] = layer0_outputs[340];
    assign outputs[9971] = layer0_outputs[2577];
    assign outputs[9972] = ~(layer0_outputs[4952]);
    assign outputs[9973] = ~((layer0_outputs[6673]) | (layer0_outputs[6085]));
    assign outputs[9974] = ~(layer0_outputs[4102]) | (layer0_outputs[408]);
    assign outputs[9975] = (layer0_outputs[362]) & ~(layer0_outputs[655]);
    assign outputs[9976] = ~(layer0_outputs[505]);
    assign outputs[9977] = layer0_outputs[1052];
    assign outputs[9978] = layer0_outputs[1866];
    assign outputs[9979] = layer0_outputs[6549];
    assign outputs[9980] = (layer0_outputs[3441]) & ~(layer0_outputs[1229]);
    assign outputs[9981] = layer0_outputs[7165];
    assign outputs[9982] = layer0_outputs[9865];
    assign outputs[9983] = layer0_outputs[8763];
    assign outputs[9984] = 1'b0;
    assign outputs[9985] = ~((layer0_outputs[5698]) | (layer0_outputs[4797]));
    assign outputs[9986] = ~((layer0_outputs[7856]) ^ (layer0_outputs[3957]));
    assign outputs[9987] = layer0_outputs[9159];
    assign outputs[9988] = ~(layer0_outputs[5233]);
    assign outputs[9989] = (layer0_outputs[307]) & ~(layer0_outputs[142]);
    assign outputs[9990] = ~(layer0_outputs[7441]) | (layer0_outputs[1239]);
    assign outputs[9991] = layer0_outputs[5791];
    assign outputs[9992] = (layer0_outputs[8808]) ^ (layer0_outputs[2169]);
    assign outputs[9993] = layer0_outputs[6062];
    assign outputs[9994] = ~((layer0_outputs[1145]) & (layer0_outputs[5430]));
    assign outputs[9995] = layer0_outputs[10082];
    assign outputs[9996] = ~(layer0_outputs[7532]);
    assign outputs[9997] = (layer0_outputs[4774]) | (layer0_outputs[589]);
    assign outputs[9998] = ~(layer0_outputs[3936]);
    assign outputs[9999] = ~((layer0_outputs[9806]) ^ (layer0_outputs[4022]));
    assign outputs[10000] = layer0_outputs[624];
    assign outputs[10001] = (layer0_outputs[6389]) & ~(layer0_outputs[7754]);
    assign outputs[10002] = layer0_outputs[9210];
    assign outputs[10003] = (layer0_outputs[7780]) & (layer0_outputs[2949]);
    assign outputs[10004] = ~((layer0_outputs[475]) ^ (layer0_outputs[10158]));
    assign outputs[10005] = ~(layer0_outputs[9581]);
    assign outputs[10006] = layer0_outputs[1832];
    assign outputs[10007] = layer0_outputs[5761];
    assign outputs[10008] = ~(layer0_outputs[5399]) | (layer0_outputs[9908]);
    assign outputs[10009] = layer0_outputs[5786];
    assign outputs[10010] = layer0_outputs[6818];
    assign outputs[10011] = layer0_outputs[3521];
    assign outputs[10012] = (layer0_outputs[5281]) | (layer0_outputs[2307]);
    assign outputs[10013] = 1'b0;
    assign outputs[10014] = ~((layer0_outputs[4675]) | (layer0_outputs[2383]));
    assign outputs[10015] = ~(layer0_outputs[2841]) | (layer0_outputs[6787]);
    assign outputs[10016] = (layer0_outputs[1959]) ^ (layer0_outputs[4455]);
    assign outputs[10017] = ~(layer0_outputs[593]);
    assign outputs[10018] = ~((layer0_outputs[1065]) ^ (layer0_outputs[2158]));
    assign outputs[10019] = layer0_outputs[10041];
    assign outputs[10020] = (layer0_outputs[563]) ^ (layer0_outputs[4968]);
    assign outputs[10021] = layer0_outputs[6671];
    assign outputs[10022] = layer0_outputs[6522];
    assign outputs[10023] = (layer0_outputs[6470]) & ~(layer0_outputs[2985]);
    assign outputs[10024] = layer0_outputs[6949];
    assign outputs[10025] = ~(layer0_outputs[4690]);
    assign outputs[10026] = ~((layer0_outputs[2656]) & (layer0_outputs[2296]));
    assign outputs[10027] = ~((layer0_outputs[1048]) ^ (layer0_outputs[6388]));
    assign outputs[10028] = layer0_outputs[3949];
    assign outputs[10029] = ~((layer0_outputs[805]) | (layer0_outputs[5860]));
    assign outputs[10030] = ~(layer0_outputs[8926]);
    assign outputs[10031] = layer0_outputs[9482];
    assign outputs[10032] = (layer0_outputs[4937]) ^ (layer0_outputs[1133]);
    assign outputs[10033] = ~((layer0_outputs[1222]) ^ (layer0_outputs[3015]));
    assign outputs[10034] = (layer0_outputs[6244]) ^ (layer0_outputs[5805]);
    assign outputs[10035] = (layer0_outputs[27]) ^ (layer0_outputs[1367]);
    assign outputs[10036] = layer0_outputs[2122];
    assign outputs[10037] = (layer0_outputs[6361]) ^ (layer0_outputs[1610]);
    assign outputs[10038] = (layer0_outputs[7598]) & ~(layer0_outputs[8150]);
    assign outputs[10039] = layer0_outputs[6176];
    assign outputs[10040] = ~(layer0_outputs[526]);
    assign outputs[10041] = layer0_outputs[6633];
    assign outputs[10042] = ~(layer0_outputs[232]);
    assign outputs[10043] = (layer0_outputs[5831]) ^ (layer0_outputs[8756]);
    assign outputs[10044] = ~((layer0_outputs[2333]) | (layer0_outputs[4527]));
    assign outputs[10045] = ~((layer0_outputs[8283]) | (layer0_outputs[8474]));
    assign outputs[10046] = (layer0_outputs[902]) & (layer0_outputs[3580]);
    assign outputs[10047] = layer0_outputs[5444];
    assign outputs[10048] = (layer0_outputs[6347]) ^ (layer0_outputs[5163]);
    assign outputs[10049] = (layer0_outputs[550]) | (layer0_outputs[9185]);
    assign outputs[10050] = ~((layer0_outputs[3660]) | (layer0_outputs[1702]));
    assign outputs[10051] = (layer0_outputs[6850]) ^ (layer0_outputs[7926]);
    assign outputs[10052] = (layer0_outputs[41]) ^ (layer0_outputs[6507]);
    assign outputs[10053] = 1'b0;
    assign outputs[10054] = layer0_outputs[2918];
    assign outputs[10055] = layer0_outputs[1295];
    assign outputs[10056] = ~((layer0_outputs[8032]) & (layer0_outputs[636]));
    assign outputs[10057] = ~(layer0_outputs[9658]);
    assign outputs[10058] = ~(layer0_outputs[9839]);
    assign outputs[10059] = (layer0_outputs[9450]) ^ (layer0_outputs[2680]);
    assign outputs[10060] = (layer0_outputs[9283]) & ~(layer0_outputs[8112]);
    assign outputs[10061] = layer0_outputs[3499];
    assign outputs[10062] = layer0_outputs[8961];
    assign outputs[10063] = layer0_outputs[6180];
    assign outputs[10064] = ~((layer0_outputs[10046]) | (layer0_outputs[1024]));
    assign outputs[10065] = ~(layer0_outputs[9591]);
    assign outputs[10066] = ~(layer0_outputs[4816]);
    assign outputs[10067] = (layer0_outputs[6088]) | (layer0_outputs[10064]);
    assign outputs[10068] = (layer0_outputs[8784]) & (layer0_outputs[456]);
    assign outputs[10069] = (layer0_outputs[8574]) & (layer0_outputs[3755]);
    assign outputs[10070] = ~(layer0_outputs[7191]);
    assign outputs[10071] = ~((layer0_outputs[3343]) ^ (layer0_outputs[7626]));
    assign outputs[10072] = ~(layer0_outputs[8400]);
    assign outputs[10073] = ~(layer0_outputs[4553]);
    assign outputs[10074] = layer0_outputs[4295];
    assign outputs[10075] = (layer0_outputs[1756]) & ~(layer0_outputs[7624]);
    assign outputs[10076] = (layer0_outputs[9482]) ^ (layer0_outputs[4707]);
    assign outputs[10077] = layer0_outputs[3414];
    assign outputs[10078] = 1'b1;
    assign outputs[10079] = (layer0_outputs[364]) & ~(layer0_outputs[2982]);
    assign outputs[10080] = ~((layer0_outputs[3591]) ^ (layer0_outputs[9242]));
    assign outputs[10081] = layer0_outputs[5208];
    assign outputs[10082] = (layer0_outputs[9075]) ^ (layer0_outputs[5577]);
    assign outputs[10083] = ~((layer0_outputs[4122]) ^ (layer0_outputs[6836]));
    assign outputs[10084] = ~((layer0_outputs[6915]) ^ (layer0_outputs[7409]));
    assign outputs[10085] = (layer0_outputs[9191]) ^ (layer0_outputs[6141]);
    assign outputs[10086] = ~((layer0_outputs[151]) & (layer0_outputs[8583]));
    assign outputs[10087] = (layer0_outputs[2698]) ^ (layer0_outputs[437]);
    assign outputs[10088] = layer0_outputs[3594];
    assign outputs[10089] = ~(layer0_outputs[326]);
    assign outputs[10090] = (layer0_outputs[4548]) ^ (layer0_outputs[6481]);
    assign outputs[10091] = ~((layer0_outputs[6222]) | (layer0_outputs[346]));
    assign outputs[10092] = (layer0_outputs[7649]) & ~(layer0_outputs[4254]);
    assign outputs[10093] = (layer0_outputs[6292]) & ~(layer0_outputs[10220]);
    assign outputs[10094] = (layer0_outputs[1885]) ^ (layer0_outputs[6373]);
    assign outputs[10095] = (layer0_outputs[2842]) & ~(layer0_outputs[1982]);
    assign outputs[10096] = layer0_outputs[3329];
    assign outputs[10097] = layer0_outputs[8202];
    assign outputs[10098] = ~((layer0_outputs[8987]) ^ (layer0_outputs[6381]));
    assign outputs[10099] = (layer0_outputs[3247]) & ~(layer0_outputs[9118]);
    assign outputs[10100] = (layer0_outputs[6648]) ^ (layer0_outputs[4580]);
    assign outputs[10101] = ~((layer0_outputs[1776]) & (layer0_outputs[1515]));
    assign outputs[10102] = (layer0_outputs[9149]) & (layer0_outputs[912]);
    assign outputs[10103] = layer0_outputs[3482];
    assign outputs[10104] = ~(layer0_outputs[2234]) | (layer0_outputs[7583]);
    assign outputs[10105] = (layer0_outputs[3911]) & (layer0_outputs[5873]);
    assign outputs[10106] = ~(layer0_outputs[3023]);
    assign outputs[10107] = (layer0_outputs[9797]) & ~(layer0_outputs[3425]);
    assign outputs[10108] = ~((layer0_outputs[424]) | (layer0_outputs[2417]));
    assign outputs[10109] = (layer0_outputs[4461]) & (layer0_outputs[9344]);
    assign outputs[10110] = (layer0_outputs[6564]) & (layer0_outputs[4339]);
    assign outputs[10111] = ~((layer0_outputs[8473]) ^ (layer0_outputs[3010]));
    assign outputs[10112] = ~(layer0_outputs[2475]);
    assign outputs[10113] = ~((layer0_outputs[9641]) | (layer0_outputs[6035]));
    assign outputs[10114] = ~(layer0_outputs[2862]) | (layer0_outputs[2665]);
    assign outputs[10115] = ~((layer0_outputs[9729]) & (layer0_outputs[1649]));
    assign outputs[10116] = layer0_outputs[2507];
    assign outputs[10117] = (layer0_outputs[6814]) & (layer0_outputs[3465]);
    assign outputs[10118] = layer0_outputs[3739];
    assign outputs[10119] = ~(layer0_outputs[7217]) | (layer0_outputs[6762]);
    assign outputs[10120] = ~(layer0_outputs[5493]);
    assign outputs[10121] = layer0_outputs[5367];
    assign outputs[10122] = layer0_outputs[8600];
    assign outputs[10123] = layer0_outputs[199];
    assign outputs[10124] = ~(layer0_outputs[709]);
    assign outputs[10125] = layer0_outputs[6343];
    assign outputs[10126] = ~(layer0_outputs[5200]);
    assign outputs[10127] = layer0_outputs[3950];
    assign outputs[10128] = layer0_outputs[6874];
    assign outputs[10129] = (layer0_outputs[3386]) ^ (layer0_outputs[1844]);
    assign outputs[10130] = ~((layer0_outputs[4611]) ^ (layer0_outputs[9623]));
    assign outputs[10131] = ~(layer0_outputs[4586]);
    assign outputs[10132] = ~(layer0_outputs[5611]);
    assign outputs[10133] = (layer0_outputs[351]) ^ (layer0_outputs[9258]);
    assign outputs[10134] = (layer0_outputs[3385]) & ~(layer0_outputs[4913]);
    assign outputs[10135] = (layer0_outputs[1415]) & (layer0_outputs[9691]);
    assign outputs[10136] = (layer0_outputs[3137]) & (layer0_outputs[8353]);
    assign outputs[10137] = ~((layer0_outputs[360]) ^ (layer0_outputs[4819]));
    assign outputs[10138] = ~(layer0_outputs[7804]);
    assign outputs[10139] = (layer0_outputs[6072]) & ~(layer0_outputs[4383]);
    assign outputs[10140] = ~(layer0_outputs[5206]);
    assign outputs[10141] = layer0_outputs[7477];
    assign outputs[10142] = (layer0_outputs[2965]) ^ (layer0_outputs[2394]);
    assign outputs[10143] = ~(layer0_outputs[1313]);
    assign outputs[10144] = ~(layer0_outputs[192]) | (layer0_outputs[8952]);
    assign outputs[10145] = (layer0_outputs[210]) & (layer0_outputs[4676]);
    assign outputs[10146] = (layer0_outputs[1825]) | (layer0_outputs[4613]);
    assign outputs[10147] = ~((layer0_outputs[8632]) ^ (layer0_outputs[6464]));
    assign outputs[10148] = ~((layer0_outputs[7049]) ^ (layer0_outputs[7971]));
    assign outputs[10149] = ~((layer0_outputs[9264]) | (layer0_outputs[6519]));
    assign outputs[10150] = ~((layer0_outputs[8688]) ^ (layer0_outputs[9406]));
    assign outputs[10151] = layer0_outputs[3342];
    assign outputs[10152] = layer0_outputs[5498];
    assign outputs[10153] = ~((layer0_outputs[3167]) & (layer0_outputs[9637]));
    assign outputs[10154] = layer0_outputs[2084];
    assign outputs[10155] = ~(layer0_outputs[7706]) | (layer0_outputs[9214]);
    assign outputs[10156] = ~(layer0_outputs[9653]);
    assign outputs[10157] = ~((layer0_outputs[8273]) ^ (layer0_outputs[2040]));
    assign outputs[10158] = ~(layer0_outputs[4419]);
    assign outputs[10159] = ~(layer0_outputs[3424]);
    assign outputs[10160] = layer0_outputs[9055];
    assign outputs[10161] = ~(layer0_outputs[4415]);
    assign outputs[10162] = ~((layer0_outputs[3404]) ^ (layer0_outputs[3965]));
    assign outputs[10163] = ~((layer0_outputs[8403]) | (layer0_outputs[1989]));
    assign outputs[10164] = ~(layer0_outputs[4102]) | (layer0_outputs[2477]);
    assign outputs[10165] = ~(layer0_outputs[4954]);
    assign outputs[10166] = ~(layer0_outputs[2132]);
    assign outputs[10167] = ~(layer0_outputs[10188]);
    assign outputs[10168] = ~(layer0_outputs[1264]);
    assign outputs[10169] = (layer0_outputs[5936]) ^ (layer0_outputs[522]);
    assign outputs[10170] = layer0_outputs[8766];
    assign outputs[10171] = layer0_outputs[5138];
    assign outputs[10172] = ~((layer0_outputs[128]) | (layer0_outputs[9405]));
    assign outputs[10173] = layer0_outputs[3189];
    assign outputs[10174] = layer0_outputs[5326];
    assign outputs[10175] = layer0_outputs[1051];
    assign outputs[10176] = ~((layer0_outputs[7762]) & (layer0_outputs[4816]));
    assign outputs[10177] = ~(layer0_outputs[3407]);
    assign outputs[10178] = (layer0_outputs[786]) & ~(layer0_outputs[10127]);
    assign outputs[10179] = 1'b1;
    assign outputs[10180] = ~((layer0_outputs[1762]) | (layer0_outputs[9760]));
    assign outputs[10181] = ~((layer0_outputs[8164]) ^ (layer0_outputs[8745]));
    assign outputs[10182] = (layer0_outputs[6967]) & (layer0_outputs[4168]);
    assign outputs[10183] = (layer0_outputs[2010]) & (layer0_outputs[4818]);
    assign outputs[10184] = ~(layer0_outputs[512]);
    assign outputs[10185] = ~(layer0_outputs[5500]);
    assign outputs[10186] = ~(layer0_outputs[1456]);
    assign outputs[10187] = ~(layer0_outputs[2761]);
    assign outputs[10188] = (layer0_outputs[6799]) & (layer0_outputs[3918]);
    assign outputs[10189] = (layer0_outputs[3805]) | (layer0_outputs[4570]);
    assign outputs[10190] = ~(layer0_outputs[6988]) | (layer0_outputs[10204]);
    assign outputs[10191] = (layer0_outputs[641]) & ~(layer0_outputs[7427]);
    assign outputs[10192] = (layer0_outputs[4020]) & (layer0_outputs[6487]);
    assign outputs[10193] = (layer0_outputs[3065]) ^ (layer0_outputs[3872]);
    assign outputs[10194] = layer0_outputs[290];
    assign outputs[10195] = (layer0_outputs[6818]) & ~(layer0_outputs[1248]);
    assign outputs[10196] = ~((layer0_outputs[1025]) | (layer0_outputs[1870]));
    assign outputs[10197] = ~(layer0_outputs[4953]);
    assign outputs[10198] = ~((layer0_outputs[1278]) ^ (layer0_outputs[8706]));
    assign outputs[10199] = layer0_outputs[856];
    assign outputs[10200] = ~(layer0_outputs[1070]);
    assign outputs[10201] = (layer0_outputs[4863]) & ~(layer0_outputs[9393]);
    assign outputs[10202] = ~(layer0_outputs[376]) | (layer0_outputs[2404]);
    assign outputs[10203] = ~(layer0_outputs[10178]);
    assign outputs[10204] = ~(layer0_outputs[503]);
    assign outputs[10205] = ~((layer0_outputs[1079]) | (layer0_outputs[106]));
    assign outputs[10206] = layer0_outputs[4070];
    assign outputs[10207] = (layer0_outputs[3654]) & (layer0_outputs[1148]);
    assign outputs[10208] = (layer0_outputs[1558]) | (layer0_outputs[3888]);
    assign outputs[10209] = ~(layer0_outputs[3439]);
    assign outputs[10210] = ~(layer0_outputs[2409]) | (layer0_outputs[1731]);
    assign outputs[10211] = (layer0_outputs[7274]) | (layer0_outputs[3417]);
    assign outputs[10212] = ~(layer0_outputs[3791]);
    assign outputs[10213] = layer0_outputs[3085];
    assign outputs[10214] = ~((layer0_outputs[4579]) ^ (layer0_outputs[2288]));
    assign outputs[10215] = ~(layer0_outputs[6758]);
    assign outputs[10216] = ~(layer0_outputs[4635]);
    assign outputs[10217] = layer0_outputs[397];
    assign outputs[10218] = layer0_outputs[6801];
    assign outputs[10219] = (layer0_outputs[6926]) & ~(layer0_outputs[2415]);
    assign outputs[10220] = layer0_outputs[578];
    assign outputs[10221] = ~((layer0_outputs[3726]) & (layer0_outputs[9926]));
    assign outputs[10222] = (layer0_outputs[4359]) ^ (layer0_outputs[9859]);
    assign outputs[10223] = ~((layer0_outputs[5314]) ^ (layer0_outputs[7439]));
    assign outputs[10224] = ~((layer0_outputs[4437]) & (layer0_outputs[1275]));
    assign outputs[10225] = ~((layer0_outputs[6424]) ^ (layer0_outputs[4562]));
    assign outputs[10226] = layer0_outputs[4081];
    assign outputs[10227] = (layer0_outputs[2894]) & ~(layer0_outputs[3737]);
    assign outputs[10228] = (layer0_outputs[9493]) & (layer0_outputs[8972]);
    assign outputs[10229] = (layer0_outputs[7819]) & ~(layer0_outputs[6393]);
    assign outputs[10230] = ~((layer0_outputs[10146]) ^ (layer0_outputs[5304]));
    assign outputs[10231] = (layer0_outputs[1344]) ^ (layer0_outputs[99]);
    assign outputs[10232] = ~((layer0_outputs[7550]) ^ (layer0_outputs[563]));
    assign outputs[10233] = ~(layer0_outputs[9875]);
    assign outputs[10234] = (layer0_outputs[9616]) ^ (layer0_outputs[7679]);
    assign outputs[10235] = (layer0_outputs[3053]) ^ (layer0_outputs[7386]);
    assign outputs[10236] = (layer0_outputs[9189]) & (layer0_outputs[5575]);
    assign outputs[10237] = ~((layer0_outputs[6657]) ^ (layer0_outputs[841]));
    assign outputs[10238] = ~((layer0_outputs[4219]) & (layer0_outputs[3364]));
    assign outputs[10239] = (layer0_outputs[6312]) & ~(layer0_outputs[4621]);
endmodule
