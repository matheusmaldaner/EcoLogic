library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(5119 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);
    signal layer1_outputs : std_logic_vector(5119 downto 0);
    signal layer2_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= not(inputs(54)) or (inputs(240));
    layer0_outputs(1) <= '1';
    layer0_outputs(2) <= not(inputs(13)) or (inputs(203));
    layer0_outputs(3) <= inputs(225);
    layer0_outputs(4) <= (inputs(152)) or (inputs(1));
    layer0_outputs(5) <= inputs(197);
    layer0_outputs(6) <= not((inputs(148)) or (inputs(239)));
    layer0_outputs(7) <= not(inputs(72));
    layer0_outputs(8) <= (inputs(56)) or (inputs(49));
    layer0_outputs(9) <= inputs(100);
    layer0_outputs(10) <= not((inputs(138)) or (inputs(102)));
    layer0_outputs(11) <= not(inputs(105));
    layer0_outputs(12) <= (inputs(189)) xor (inputs(99));
    layer0_outputs(13) <= (inputs(206)) and not (inputs(81));
    layer0_outputs(14) <= inputs(223);
    layer0_outputs(15) <= (inputs(55)) or (inputs(241));
    layer0_outputs(16) <= not((inputs(183)) or (inputs(165)));
    layer0_outputs(17) <= not(inputs(89));
    layer0_outputs(18) <= '0';
    layer0_outputs(19) <= not(inputs(47)) or (inputs(218));
    layer0_outputs(20) <= inputs(198);
    layer0_outputs(21) <= not(inputs(43));
    layer0_outputs(22) <= not(inputs(83));
    layer0_outputs(23) <= not((inputs(206)) xor (inputs(172)));
    layer0_outputs(24) <= (inputs(107)) xor (inputs(3));
    layer0_outputs(25) <= not(inputs(103));
    layer0_outputs(26) <= (inputs(36)) and not (inputs(91));
    layer0_outputs(27) <= inputs(205);
    layer0_outputs(28) <= inputs(146);
    layer0_outputs(29) <= inputs(100);
    layer0_outputs(30) <= not((inputs(217)) xor (inputs(3)));
    layer0_outputs(31) <= not(inputs(113));
    layer0_outputs(32) <= not(inputs(242));
    layer0_outputs(33) <= not(inputs(215));
    layer0_outputs(34) <= (inputs(191)) and (inputs(159));
    layer0_outputs(35) <= (inputs(244)) or (inputs(47));
    layer0_outputs(36) <= inputs(85);
    layer0_outputs(37) <= not(inputs(248));
    layer0_outputs(38) <= not(inputs(22)) or (inputs(233));
    layer0_outputs(39) <= (inputs(134)) and not (inputs(132));
    layer0_outputs(40) <= not((inputs(181)) or (inputs(217)));
    layer0_outputs(41) <= not(inputs(29));
    layer0_outputs(42) <= (inputs(155)) or (inputs(145));
    layer0_outputs(43) <= (inputs(136)) and not (inputs(245));
    layer0_outputs(44) <= (inputs(24)) and not (inputs(164));
    layer0_outputs(45) <= not((inputs(61)) or (inputs(23)));
    layer0_outputs(46) <= not(inputs(93));
    layer0_outputs(47) <= not(inputs(167));
    layer0_outputs(48) <= not((inputs(246)) or (inputs(162)));
    layer0_outputs(49) <= not((inputs(49)) or (inputs(163)));
    layer0_outputs(50) <= not((inputs(187)) or (inputs(56)));
    layer0_outputs(51) <= (inputs(16)) or (inputs(121));
    layer0_outputs(52) <= (inputs(44)) or (inputs(47));
    layer0_outputs(53) <= (inputs(173)) or (inputs(223));
    layer0_outputs(54) <= (inputs(179)) or (inputs(252));
    layer0_outputs(55) <= (inputs(106)) and not (inputs(244));
    layer0_outputs(56) <= inputs(43);
    layer0_outputs(57) <= not((inputs(7)) and (inputs(205)));
    layer0_outputs(58) <= (inputs(78)) and not (inputs(235));
    layer0_outputs(59) <= (inputs(124)) or (inputs(4));
    layer0_outputs(60) <= '0';
    layer0_outputs(61) <= (inputs(2)) or (inputs(45));
    layer0_outputs(62) <= inputs(17);
    layer0_outputs(63) <= (inputs(251)) or (inputs(149));
    layer0_outputs(64) <= not(inputs(198)) or (inputs(175));
    layer0_outputs(65) <= (inputs(15)) or (inputs(131));
    layer0_outputs(66) <= (inputs(191)) and not (inputs(11));
    layer0_outputs(67) <= (inputs(25)) or (inputs(155));
    layer0_outputs(68) <= not(inputs(221)) or (inputs(228));
    layer0_outputs(69) <= (inputs(60)) and not (inputs(70));
    layer0_outputs(70) <= (inputs(101)) and not (inputs(0));
    layer0_outputs(71) <= (inputs(128)) or (inputs(155));
    layer0_outputs(72) <= (inputs(217)) or (inputs(146));
    layer0_outputs(73) <= not(inputs(128));
    layer0_outputs(74) <= inputs(9);
    layer0_outputs(75) <= not(inputs(104));
    layer0_outputs(76) <= '1';
    layer0_outputs(77) <= (inputs(132)) and not (inputs(226));
    layer0_outputs(78) <= '1';
    layer0_outputs(79) <= (inputs(58)) and not (inputs(117));
    layer0_outputs(80) <= not(inputs(96)) or (inputs(241));
    layer0_outputs(81) <= (inputs(121)) and not (inputs(106));
    layer0_outputs(82) <= not(inputs(234));
    layer0_outputs(83) <= (inputs(151)) and not (inputs(209));
    layer0_outputs(84) <= (inputs(94)) or (inputs(24));
    layer0_outputs(85) <= (inputs(242)) or (inputs(90));
    layer0_outputs(86) <= inputs(246);
    layer0_outputs(87) <= (inputs(8)) or (inputs(179));
    layer0_outputs(88) <= not(inputs(7));
    layer0_outputs(89) <= not((inputs(108)) or (inputs(120)));
    layer0_outputs(90) <= not((inputs(192)) or (inputs(39)));
    layer0_outputs(91) <= not((inputs(198)) and (inputs(170)));
    layer0_outputs(92) <= inputs(189);
    layer0_outputs(93) <= '0';
    layer0_outputs(94) <= not(inputs(75));
    layer0_outputs(95) <= (inputs(249)) and not (inputs(29));
    layer0_outputs(96) <= (inputs(36)) xor (inputs(240));
    layer0_outputs(97) <= (inputs(61)) xor (inputs(150));
    layer0_outputs(98) <= inputs(156);
    layer0_outputs(99) <= '1';
    layer0_outputs(100) <= not(inputs(75)) or (inputs(254));
    layer0_outputs(101) <= inputs(215);
    layer0_outputs(102) <= not(inputs(247));
    layer0_outputs(103) <= not(inputs(135));
    layer0_outputs(104) <= not(inputs(133)) or (inputs(46));
    layer0_outputs(105) <= (inputs(24)) and not (inputs(194));
    layer0_outputs(106) <= not(inputs(103));
    layer0_outputs(107) <= (inputs(187)) or (inputs(243));
    layer0_outputs(108) <= inputs(180);
    layer0_outputs(109) <= '1';
    layer0_outputs(110) <= inputs(90);
    layer0_outputs(111) <= not((inputs(238)) or (inputs(188)));
    layer0_outputs(112) <= not((inputs(141)) xor (inputs(253)));
    layer0_outputs(113) <= (inputs(225)) or (inputs(210));
    layer0_outputs(114) <= inputs(104);
    layer0_outputs(115) <= inputs(90);
    layer0_outputs(116) <= (inputs(255)) or (inputs(21));
    layer0_outputs(117) <= not(inputs(92));
    layer0_outputs(118) <= (inputs(157)) or (inputs(15));
    layer0_outputs(119) <= '0';
    layer0_outputs(120) <= not((inputs(217)) xor (inputs(62)));
    layer0_outputs(121) <= not(inputs(7)) or (inputs(204));
    layer0_outputs(122) <= '0';
    layer0_outputs(123) <= (inputs(50)) and not (inputs(241));
    layer0_outputs(124) <= inputs(175);
    layer0_outputs(125) <= not((inputs(3)) or (inputs(75)));
    layer0_outputs(126) <= inputs(231);
    layer0_outputs(127) <= (inputs(59)) and not (inputs(206));
    layer0_outputs(128) <= not(inputs(132));
    layer0_outputs(129) <= inputs(193);
    layer0_outputs(130) <= not(inputs(110));
    layer0_outputs(131) <= '1';
    layer0_outputs(132) <= (inputs(29)) and not (inputs(91));
    layer0_outputs(133) <= not(inputs(94));
    layer0_outputs(134) <= '0';
    layer0_outputs(135) <= (inputs(187)) and not (inputs(92));
    layer0_outputs(136) <= not(inputs(66));
    layer0_outputs(137) <= not(inputs(22));
    layer0_outputs(138) <= (inputs(21)) or (inputs(230));
    layer0_outputs(139) <= not(inputs(180));
    layer0_outputs(140) <= '0';
    layer0_outputs(141) <= '0';
    layer0_outputs(142) <= not((inputs(43)) xor (inputs(11)));
    layer0_outputs(143) <= inputs(185);
    layer0_outputs(144) <= inputs(217);
    layer0_outputs(145) <= inputs(109);
    layer0_outputs(146) <= (inputs(149)) xor (inputs(237));
    layer0_outputs(147) <= (inputs(17)) or (inputs(208));
    layer0_outputs(148) <= '0';
    layer0_outputs(149) <= not(inputs(221));
    layer0_outputs(150) <= (inputs(217)) and not (inputs(19));
    layer0_outputs(151) <= inputs(134);
    layer0_outputs(152) <= (inputs(142)) xor (inputs(136));
    layer0_outputs(153) <= (inputs(24)) or (inputs(36));
    layer0_outputs(154) <= not((inputs(174)) or (inputs(110)));
    layer0_outputs(155) <= (inputs(100)) or (inputs(254));
    layer0_outputs(156) <= inputs(166);
    layer0_outputs(157) <= not(inputs(233)) or (inputs(200));
    layer0_outputs(158) <= not(inputs(47)) or (inputs(13));
    layer0_outputs(159) <= not(inputs(245));
    layer0_outputs(160) <= (inputs(71)) xor (inputs(50));
    layer0_outputs(161) <= not((inputs(11)) and (inputs(218)));
    layer0_outputs(162) <= not(inputs(135)) or (inputs(214));
    layer0_outputs(163) <= not(inputs(21));
    layer0_outputs(164) <= not(inputs(206));
    layer0_outputs(165) <= not(inputs(23)) or (inputs(225));
    layer0_outputs(166) <= not(inputs(102));
    layer0_outputs(167) <= (inputs(22)) and not (inputs(194));
    layer0_outputs(168) <= inputs(137);
    layer0_outputs(169) <= not(inputs(120)) or (inputs(128));
    layer0_outputs(170) <= not(inputs(164));
    layer0_outputs(171) <= not((inputs(179)) or (inputs(222)));
    layer0_outputs(172) <= inputs(237);
    layer0_outputs(173) <= not(inputs(227)) or (inputs(205));
    layer0_outputs(174) <= (inputs(125)) and not (inputs(45));
    layer0_outputs(175) <= (inputs(85)) xor (inputs(24));
    layer0_outputs(176) <= not(inputs(25));
    layer0_outputs(177) <= inputs(215);
    layer0_outputs(178) <= (inputs(166)) and not (inputs(167));
    layer0_outputs(179) <= not(inputs(182));
    layer0_outputs(180) <= (inputs(155)) or (inputs(130));
    layer0_outputs(181) <= inputs(204);
    layer0_outputs(182) <= inputs(197);
    layer0_outputs(183) <= (inputs(200)) and not (inputs(49));
    layer0_outputs(184) <= not((inputs(194)) or (inputs(160)));
    layer0_outputs(185) <= not((inputs(94)) or (inputs(124)));
    layer0_outputs(186) <= '1';
    layer0_outputs(187) <= '1';
    layer0_outputs(188) <= not((inputs(142)) or (inputs(47)));
    layer0_outputs(189) <= inputs(232);
    layer0_outputs(190) <= not((inputs(145)) xor (inputs(149)));
    layer0_outputs(191) <= (inputs(59)) or (inputs(80));
    layer0_outputs(192) <= (inputs(168)) or (inputs(66));
    layer0_outputs(193) <= inputs(166);
    layer0_outputs(194) <= (inputs(17)) and (inputs(252));
    layer0_outputs(195) <= not((inputs(91)) or (inputs(163)));
    layer0_outputs(196) <= (inputs(176)) or (inputs(194));
    layer0_outputs(197) <= (inputs(200)) and not (inputs(113));
    layer0_outputs(198) <= not((inputs(45)) xor (inputs(75)));
    layer0_outputs(199) <= not((inputs(82)) or (inputs(131)));
    layer0_outputs(200) <= not(inputs(173)) or (inputs(16));
    layer0_outputs(201) <= not(inputs(133)) or (inputs(13));
    layer0_outputs(202) <= not((inputs(64)) or (inputs(135)));
    layer0_outputs(203) <= (inputs(251)) xor (inputs(170));
    layer0_outputs(204) <= not((inputs(17)) xor (inputs(48)));
    layer0_outputs(205) <= inputs(98);
    layer0_outputs(206) <= not((inputs(129)) xor (inputs(165)));
    layer0_outputs(207) <= inputs(59);
    layer0_outputs(208) <= inputs(90);
    layer0_outputs(209) <= not((inputs(203)) or (inputs(116)));
    layer0_outputs(210) <= (inputs(92)) or (inputs(177));
    layer0_outputs(211) <= (inputs(55)) and not (inputs(133));
    layer0_outputs(212) <= inputs(80);
    layer0_outputs(213) <= not(inputs(154));
    layer0_outputs(214) <= (inputs(52)) and (inputs(151));
    layer0_outputs(215) <= '1';
    layer0_outputs(216) <= not(inputs(77));
    layer0_outputs(217) <= (inputs(49)) and not (inputs(177));
    layer0_outputs(218) <= '0';
    layer0_outputs(219) <= (inputs(37)) or (inputs(35));
    layer0_outputs(220) <= (inputs(241)) or (inputs(135));
    layer0_outputs(221) <= not((inputs(112)) or (inputs(128)));
    layer0_outputs(222) <= inputs(190);
    layer0_outputs(223) <= not(inputs(188)) or (inputs(96));
    layer0_outputs(224) <= inputs(17);
    layer0_outputs(225) <= inputs(207);
    layer0_outputs(226) <= not((inputs(185)) and (inputs(196)));
    layer0_outputs(227) <= inputs(245);
    layer0_outputs(228) <= not((inputs(45)) or (inputs(1)));
    layer0_outputs(229) <= '0';
    layer0_outputs(230) <= not(inputs(91));
    layer0_outputs(231) <= not(inputs(8)) or (inputs(162));
    layer0_outputs(232) <= not(inputs(22)) or (inputs(166));
    layer0_outputs(233) <= (inputs(165)) or (inputs(114));
    layer0_outputs(234) <= (inputs(178)) or (inputs(186));
    layer0_outputs(235) <= (inputs(244)) and not (inputs(40));
    layer0_outputs(236) <= (inputs(156)) xor (inputs(27));
    layer0_outputs(237) <= not((inputs(184)) or (inputs(80)));
    layer0_outputs(238) <= (inputs(139)) or (inputs(46));
    layer0_outputs(239) <= inputs(97);
    layer0_outputs(240) <= '1';
    layer0_outputs(241) <= not(inputs(96));
    layer0_outputs(242) <= (inputs(238)) and (inputs(62));
    layer0_outputs(243) <= not((inputs(172)) or (inputs(141)));
    layer0_outputs(244) <= (inputs(192)) and not (inputs(247));
    layer0_outputs(245) <= (inputs(255)) or (inputs(254));
    layer0_outputs(246) <= not(inputs(189)) or (inputs(162));
    layer0_outputs(247) <= inputs(163);
    layer0_outputs(248) <= '1';
    layer0_outputs(249) <= '1';
    layer0_outputs(250) <= inputs(201);
    layer0_outputs(251) <= inputs(164);
    layer0_outputs(252) <= (inputs(29)) or (inputs(31));
    layer0_outputs(253) <= (inputs(6)) xor (inputs(177));
    layer0_outputs(254) <= (inputs(116)) or (inputs(214));
    layer0_outputs(255) <= (inputs(130)) or (inputs(247));
    layer0_outputs(256) <= not(inputs(99));
    layer0_outputs(257) <= not(inputs(218));
    layer0_outputs(258) <= (inputs(193)) and not (inputs(100));
    layer0_outputs(259) <= not(inputs(114));
    layer0_outputs(260) <= (inputs(34)) xor (inputs(180));
    layer0_outputs(261) <= not(inputs(207)) or (inputs(46));
    layer0_outputs(262) <= not(inputs(227)) or (inputs(93));
    layer0_outputs(263) <= '1';
    layer0_outputs(264) <= not((inputs(77)) or (inputs(106)));
    layer0_outputs(265) <= not((inputs(92)) and (inputs(83)));
    layer0_outputs(266) <= (inputs(116)) xor (inputs(208));
    layer0_outputs(267) <= not(inputs(118)) or (inputs(49));
    layer0_outputs(268) <= inputs(119);
    layer0_outputs(269) <= (inputs(153)) and not (inputs(15));
    layer0_outputs(270) <= not(inputs(213)) or (inputs(95));
    layer0_outputs(271) <= not(inputs(230));
    layer0_outputs(272) <= not(inputs(64));
    layer0_outputs(273) <= inputs(92);
    layer0_outputs(274) <= inputs(47);
    layer0_outputs(275) <= not((inputs(90)) or (inputs(3)));
    layer0_outputs(276) <= not((inputs(168)) or (inputs(66)));
    layer0_outputs(277) <= (inputs(4)) xor (inputs(0));
    layer0_outputs(278) <= inputs(96);
    layer0_outputs(279) <= not(inputs(69)) or (inputs(48));
    layer0_outputs(280) <= not(inputs(174)) or (inputs(65));
    layer0_outputs(281) <= (inputs(176)) and not (inputs(204));
    layer0_outputs(282) <= inputs(77);
    layer0_outputs(283) <= not(inputs(117)) or (inputs(84));
    layer0_outputs(284) <= '1';
    layer0_outputs(285) <= (inputs(170)) or (inputs(247));
    layer0_outputs(286) <= (inputs(7)) and not (inputs(129));
    layer0_outputs(287) <= not((inputs(147)) and (inputs(81)));
    layer0_outputs(288) <= not((inputs(208)) or (inputs(230)));
    layer0_outputs(289) <= (inputs(171)) xor (inputs(190));
    layer0_outputs(290) <= not((inputs(245)) or (inputs(202)));
    layer0_outputs(291) <= not((inputs(19)) or (inputs(64)));
    layer0_outputs(292) <= not((inputs(203)) xor (inputs(163)));
    layer0_outputs(293) <= (inputs(57)) and not (inputs(81));
    layer0_outputs(294) <= inputs(61);
    layer0_outputs(295) <= not(inputs(222));
    layer0_outputs(296) <= '1';
    layer0_outputs(297) <= not((inputs(68)) and (inputs(25)));
    layer0_outputs(298) <= not((inputs(22)) and (inputs(90)));
    layer0_outputs(299) <= not(inputs(64));
    layer0_outputs(300) <= inputs(144);
    layer0_outputs(301) <= not(inputs(77));
    layer0_outputs(302) <= inputs(52);
    layer0_outputs(303) <= '1';
    layer0_outputs(304) <= not(inputs(253)) or (inputs(107));
    layer0_outputs(305) <= not((inputs(98)) and (inputs(14)));
    layer0_outputs(306) <= (inputs(90)) or (inputs(138));
    layer0_outputs(307) <= not(inputs(211));
    layer0_outputs(308) <= not(inputs(237));
    layer0_outputs(309) <= inputs(154);
    layer0_outputs(310) <= not(inputs(173)) or (inputs(237));
    layer0_outputs(311) <= not(inputs(178));
    layer0_outputs(312) <= (inputs(88)) and not (inputs(154));
    layer0_outputs(313) <= not(inputs(244));
    layer0_outputs(314) <= not(inputs(229));
    layer0_outputs(315) <= not((inputs(156)) or (inputs(234)));
    layer0_outputs(316) <= not(inputs(26)) or (inputs(16));
    layer0_outputs(317) <= (inputs(11)) and not (inputs(146));
    layer0_outputs(318) <= not(inputs(97)) or (inputs(149));
    layer0_outputs(319) <= not(inputs(206));
    layer0_outputs(320) <= not((inputs(52)) xor (inputs(39)));
    layer0_outputs(321) <= not(inputs(85));
    layer0_outputs(322) <= not(inputs(47));
    layer0_outputs(323) <= not(inputs(230));
    layer0_outputs(324) <= not((inputs(171)) or (inputs(124)));
    layer0_outputs(325) <= inputs(33);
    layer0_outputs(326) <= (inputs(78)) and (inputs(237));
    layer0_outputs(327) <= inputs(106);
    layer0_outputs(328) <= (inputs(69)) or (inputs(250));
    layer0_outputs(329) <= (inputs(142)) or (inputs(27));
    layer0_outputs(330) <= not(inputs(154));
    layer0_outputs(331) <= not((inputs(182)) or (inputs(162)));
    layer0_outputs(332) <= not((inputs(98)) or (inputs(47)));
    layer0_outputs(333) <= not(inputs(184)) or (inputs(161));
    layer0_outputs(334) <= not((inputs(178)) or (inputs(5)));
    layer0_outputs(335) <= '0';
    layer0_outputs(336) <= inputs(185);
    layer0_outputs(337) <= (inputs(46)) xor (inputs(91));
    layer0_outputs(338) <= not(inputs(53));
    layer0_outputs(339) <= inputs(35);
    layer0_outputs(340) <= not(inputs(167));
    layer0_outputs(341) <= not(inputs(173));
    layer0_outputs(342) <= inputs(52);
    layer0_outputs(343) <= (inputs(71)) and not (inputs(43));
    layer0_outputs(344) <= not((inputs(208)) or (inputs(38)));
    layer0_outputs(345) <= '0';
    layer0_outputs(346) <= inputs(201);
    layer0_outputs(347) <= not((inputs(159)) or (inputs(185)));
    layer0_outputs(348) <= '0';
    layer0_outputs(349) <= not(inputs(44));
    layer0_outputs(350) <= not(inputs(229));
    layer0_outputs(351) <= not(inputs(8));
    layer0_outputs(352) <= not(inputs(69)) or (inputs(54));
    layer0_outputs(353) <= '0';
    layer0_outputs(354) <= not((inputs(200)) and (inputs(70)));
    layer0_outputs(355) <= not(inputs(14)) or (inputs(150));
    layer0_outputs(356) <= (inputs(127)) or (inputs(179));
    layer0_outputs(357) <= inputs(134);
    layer0_outputs(358) <= not(inputs(129));
    layer0_outputs(359) <= (inputs(108)) xor (inputs(3));
    layer0_outputs(360) <= not(inputs(15)) or (inputs(237));
    layer0_outputs(361) <= inputs(82);
    layer0_outputs(362) <= not((inputs(198)) and (inputs(233)));
    layer0_outputs(363) <= not(inputs(36)) or (inputs(59));
    layer0_outputs(364) <= not((inputs(151)) xor (inputs(239)));
    layer0_outputs(365) <= not(inputs(27));
    layer0_outputs(366) <= not(inputs(162));
    layer0_outputs(367) <= not(inputs(201));
    layer0_outputs(368) <= (inputs(127)) and not (inputs(41));
    layer0_outputs(369) <= not(inputs(196));
    layer0_outputs(370) <= '0';
    layer0_outputs(371) <= inputs(148);
    layer0_outputs(372) <= not((inputs(162)) and (inputs(130)));
    layer0_outputs(373) <= (inputs(150)) and not (inputs(151));
    layer0_outputs(374) <= not((inputs(71)) or (inputs(40)));
    layer0_outputs(375) <= not(inputs(164));
    layer0_outputs(376) <= not((inputs(248)) and (inputs(235)));
    layer0_outputs(377) <= not(inputs(213)) or (inputs(118));
    layer0_outputs(378) <= not(inputs(113)) or (inputs(16));
    layer0_outputs(379) <= not(inputs(18));
    layer0_outputs(380) <= inputs(161);
    layer0_outputs(381) <= inputs(164);
    layer0_outputs(382) <= inputs(144);
    layer0_outputs(383) <= (inputs(235)) and (inputs(183));
    layer0_outputs(384) <= not(inputs(103));
    layer0_outputs(385) <= (inputs(202)) and (inputs(243));
    layer0_outputs(386) <= (inputs(137)) xor (inputs(86));
    layer0_outputs(387) <= not((inputs(222)) or (inputs(240)));
    layer0_outputs(388) <= '0';
    layer0_outputs(389) <= not(inputs(52)) or (inputs(114));
    layer0_outputs(390) <= not((inputs(2)) or (inputs(145)));
    layer0_outputs(391) <= not(inputs(152));
    layer0_outputs(392) <= not(inputs(154)) or (inputs(181));
    layer0_outputs(393) <= '1';
    layer0_outputs(394) <= (inputs(152)) and not (inputs(4));
    layer0_outputs(395) <= (inputs(6)) or (inputs(201));
    layer0_outputs(396) <= (inputs(137)) and (inputs(137));
    layer0_outputs(397) <= (inputs(128)) and not (inputs(181));
    layer0_outputs(398) <= (inputs(208)) and not (inputs(191));
    layer0_outputs(399) <= not(inputs(143));
    layer0_outputs(400) <= not(inputs(63));
    layer0_outputs(401) <= (inputs(110)) or (inputs(158));
    layer0_outputs(402) <= not(inputs(120));
    layer0_outputs(403) <= (inputs(20)) and not (inputs(239));
    layer0_outputs(404) <= not(inputs(40));
    layer0_outputs(405) <= not(inputs(106)) or (inputs(249));
    layer0_outputs(406) <= not(inputs(97));
    layer0_outputs(407) <= inputs(193);
    layer0_outputs(408) <= inputs(163);
    layer0_outputs(409) <= not((inputs(161)) xor (inputs(23)));
    layer0_outputs(410) <= not(inputs(98));
    layer0_outputs(411) <= not(inputs(254));
    layer0_outputs(412) <= (inputs(78)) and not (inputs(7));
    layer0_outputs(413) <= '0';
    layer0_outputs(414) <= inputs(118);
    layer0_outputs(415) <= (inputs(239)) xor (inputs(48));
    layer0_outputs(416) <= not(inputs(44));
    layer0_outputs(417) <= not(inputs(100));
    layer0_outputs(418) <= not(inputs(87));
    layer0_outputs(419) <= not(inputs(232)) or (inputs(43));
    layer0_outputs(420) <= (inputs(33)) or (inputs(237));
    layer0_outputs(421) <= (inputs(98)) or (inputs(143));
    layer0_outputs(422) <= not(inputs(169)) or (inputs(166));
    layer0_outputs(423) <= inputs(228);
    layer0_outputs(424) <= inputs(248);
    layer0_outputs(425) <= not(inputs(69));
    layer0_outputs(426) <= not((inputs(94)) or (inputs(46)));
    layer0_outputs(427) <= (inputs(93)) and not (inputs(122));
    layer0_outputs(428) <= inputs(236);
    layer0_outputs(429) <= not((inputs(49)) or (inputs(22)));
    layer0_outputs(430) <= (inputs(120)) xor (inputs(173));
    layer0_outputs(431) <= (inputs(105)) and (inputs(37));
    layer0_outputs(432) <= (inputs(206)) or (inputs(138));
    layer0_outputs(433) <= not((inputs(244)) xor (inputs(85)));
    layer0_outputs(434) <= not(inputs(109)) or (inputs(143));
    layer0_outputs(435) <= inputs(28);
    layer0_outputs(436) <= '0';
    layer0_outputs(437) <= inputs(81);
    layer0_outputs(438) <= inputs(211);
    layer0_outputs(439) <= not(inputs(84));
    layer0_outputs(440) <= (inputs(146)) and not (inputs(109));
    layer0_outputs(441) <= (inputs(103)) and not (inputs(221));
    layer0_outputs(442) <= (inputs(163)) or (inputs(1));
    layer0_outputs(443) <= (inputs(6)) and not (inputs(187));
    layer0_outputs(444) <= not((inputs(156)) or (inputs(24)));
    layer0_outputs(445) <= not(inputs(36));
    layer0_outputs(446) <= not(inputs(41));
    layer0_outputs(447) <= (inputs(69)) and not (inputs(184));
    layer0_outputs(448) <= (inputs(207)) and not (inputs(63));
    layer0_outputs(449) <= (inputs(26)) and (inputs(27));
    layer0_outputs(450) <= not((inputs(162)) or (inputs(178)));
    layer0_outputs(451) <= '0';
    layer0_outputs(452) <= (inputs(208)) xor (inputs(170));
    layer0_outputs(453) <= (inputs(31)) and not (inputs(12));
    layer0_outputs(454) <= (inputs(176)) or (inputs(180));
    layer0_outputs(455) <= not(inputs(169));
    layer0_outputs(456) <= (inputs(19)) and not (inputs(50));
    layer0_outputs(457) <= not((inputs(133)) xor (inputs(252)));
    layer0_outputs(458) <= inputs(104);
    layer0_outputs(459) <= not((inputs(84)) xor (inputs(174)));
    layer0_outputs(460) <= not(inputs(66));
    layer0_outputs(461) <= not((inputs(14)) or (inputs(149)));
    layer0_outputs(462) <= (inputs(91)) and not (inputs(127));
    layer0_outputs(463) <= not(inputs(210));
    layer0_outputs(464) <= (inputs(183)) and not (inputs(170));
    layer0_outputs(465) <= '1';
    layer0_outputs(466) <= inputs(199);
    layer0_outputs(467) <= not(inputs(230));
    layer0_outputs(468) <= inputs(139);
    layer0_outputs(469) <= '0';
    layer0_outputs(470) <= (inputs(190)) or (inputs(225));
    layer0_outputs(471) <= (inputs(48)) or (inputs(105));
    layer0_outputs(472) <= not((inputs(99)) xor (inputs(151)));
    layer0_outputs(473) <= not(inputs(96));
    layer0_outputs(474) <= (inputs(179)) xor (inputs(200));
    layer0_outputs(475) <= (inputs(253)) xor (inputs(206));
    layer0_outputs(476) <= inputs(23);
    layer0_outputs(477) <= not((inputs(19)) xor (inputs(175)));
    layer0_outputs(478) <= not(inputs(222));
    layer0_outputs(479) <= (inputs(192)) and not (inputs(254));
    layer0_outputs(480) <= not(inputs(120));
    layer0_outputs(481) <= not(inputs(36)) or (inputs(131));
    layer0_outputs(482) <= not(inputs(42));
    layer0_outputs(483) <= not((inputs(173)) or (inputs(117)));
    layer0_outputs(484) <= not(inputs(102)) or (inputs(142));
    layer0_outputs(485) <= inputs(38);
    layer0_outputs(486) <= (inputs(159)) xor (inputs(190));
    layer0_outputs(487) <= inputs(187);
    layer0_outputs(488) <= not(inputs(122)) or (inputs(82));
    layer0_outputs(489) <= (inputs(103)) xor (inputs(194));
    layer0_outputs(490) <= not((inputs(147)) or (inputs(198)));
    layer0_outputs(491) <= '1';
    layer0_outputs(492) <= not(inputs(195));
    layer0_outputs(493) <= not(inputs(84));
    layer0_outputs(494) <= not(inputs(185));
    layer0_outputs(495) <= inputs(188);
    layer0_outputs(496) <= inputs(39);
    layer0_outputs(497) <= inputs(163);
    layer0_outputs(498) <= not(inputs(178));
    layer0_outputs(499) <= inputs(204);
    layer0_outputs(500) <= inputs(114);
    layer0_outputs(501) <= not((inputs(29)) or (inputs(104)));
    layer0_outputs(502) <= not(inputs(124));
    layer0_outputs(503) <= not(inputs(174)) or (inputs(113));
    layer0_outputs(504) <= inputs(165);
    layer0_outputs(505) <= (inputs(65)) or (inputs(226));
    layer0_outputs(506) <= (inputs(168)) and not (inputs(93));
    layer0_outputs(507) <= inputs(115);
    layer0_outputs(508) <= '0';
    layer0_outputs(509) <= inputs(34);
    layer0_outputs(510) <= (inputs(190)) and (inputs(78));
    layer0_outputs(511) <= '1';
    layer0_outputs(512) <= not(inputs(221)) or (inputs(158));
    layer0_outputs(513) <= inputs(102);
    layer0_outputs(514) <= (inputs(77)) and (inputs(12));
    layer0_outputs(515) <= not(inputs(126));
    layer0_outputs(516) <= not((inputs(33)) xor (inputs(248)));
    layer0_outputs(517) <= inputs(40);
    layer0_outputs(518) <= '1';
    layer0_outputs(519) <= inputs(69);
    layer0_outputs(520) <= not(inputs(228));
    layer0_outputs(521) <= (inputs(234)) or (inputs(115));
    layer0_outputs(522) <= '1';
    layer0_outputs(523) <= (inputs(88)) and not (inputs(174));
    layer0_outputs(524) <= inputs(20);
    layer0_outputs(525) <= (inputs(233)) xor (inputs(208));
    layer0_outputs(526) <= not((inputs(75)) or (inputs(61)));
    layer0_outputs(527) <= (inputs(169)) and not (inputs(72));
    layer0_outputs(528) <= inputs(142);
    layer0_outputs(529) <= (inputs(236)) or (inputs(106));
    layer0_outputs(530) <= not((inputs(213)) or (inputs(159)));
    layer0_outputs(531) <= (inputs(163)) or (inputs(106));
    layer0_outputs(532) <= '1';
    layer0_outputs(533) <= inputs(177);
    layer0_outputs(534) <= not(inputs(87));
    layer0_outputs(535) <= not((inputs(60)) xor (inputs(106)));
    layer0_outputs(536) <= '1';
    layer0_outputs(537) <= not(inputs(26));
    layer0_outputs(538) <= not(inputs(211));
    layer0_outputs(539) <= not(inputs(131));
    layer0_outputs(540) <= inputs(64);
    layer0_outputs(541) <= not(inputs(184)) or (inputs(131));
    layer0_outputs(542) <= not(inputs(71)) or (inputs(30));
    layer0_outputs(543) <= not(inputs(73)) or (inputs(239));
    layer0_outputs(544) <= inputs(19);
    layer0_outputs(545) <= not(inputs(150)) or (inputs(203));
    layer0_outputs(546) <= not((inputs(81)) and (inputs(0)));
    layer0_outputs(547) <= (inputs(197)) and (inputs(140));
    layer0_outputs(548) <= (inputs(239)) or (inputs(87));
    layer0_outputs(549) <= (inputs(69)) or (inputs(50));
    layer0_outputs(550) <= (inputs(115)) and not (inputs(197));
    layer0_outputs(551) <= not((inputs(241)) xor (inputs(196)));
    layer0_outputs(552) <= not(inputs(109));
    layer0_outputs(553) <= (inputs(241)) or (inputs(125));
    layer0_outputs(554) <= not(inputs(247));
    layer0_outputs(555) <= not(inputs(142));
    layer0_outputs(556) <= (inputs(35)) and not (inputs(51));
    layer0_outputs(557) <= '1';
    layer0_outputs(558) <= (inputs(86)) and not (inputs(49));
    layer0_outputs(559) <= not(inputs(131));
    layer0_outputs(560) <= not(inputs(251)) or (inputs(81));
    layer0_outputs(561) <= not(inputs(228));
    layer0_outputs(562) <= (inputs(161)) xor (inputs(214));
    layer0_outputs(563) <= (inputs(159)) or (inputs(252));
    layer0_outputs(564) <= '1';
    layer0_outputs(565) <= inputs(145);
    layer0_outputs(566) <= not((inputs(233)) and (inputs(168)));
    layer0_outputs(567) <= not(inputs(224)) or (inputs(66));
    layer0_outputs(568) <= not((inputs(192)) or (inputs(255)));
    layer0_outputs(569) <= not((inputs(38)) and (inputs(220)));
    layer0_outputs(570) <= not(inputs(55)) or (inputs(34));
    layer0_outputs(571) <= not(inputs(185)) or (inputs(118));
    layer0_outputs(572) <= not(inputs(90)) or (inputs(176));
    layer0_outputs(573) <= not((inputs(219)) or (inputs(243)));
    layer0_outputs(574) <= inputs(86);
    layer0_outputs(575) <= (inputs(149)) and not (inputs(0));
    layer0_outputs(576) <= not((inputs(244)) and (inputs(76)));
    layer0_outputs(577) <= not(inputs(73)) or (inputs(201));
    layer0_outputs(578) <= not(inputs(249));
    layer0_outputs(579) <= inputs(52);
    layer0_outputs(580) <= (inputs(220)) or (inputs(185));
    layer0_outputs(581) <= inputs(117);
    layer0_outputs(582) <= not(inputs(172));
    layer0_outputs(583) <= not(inputs(83)) or (inputs(156));
    layer0_outputs(584) <= (inputs(43)) and not (inputs(205));
    layer0_outputs(585) <= (inputs(108)) xor (inputs(29));
    layer0_outputs(586) <= (inputs(180)) or (inputs(253));
    layer0_outputs(587) <= not(inputs(194));
    layer0_outputs(588) <= (inputs(48)) and (inputs(250));
    layer0_outputs(589) <= (inputs(25)) or (inputs(156));
    layer0_outputs(590) <= (inputs(91)) or (inputs(104));
    layer0_outputs(591) <= not((inputs(56)) xor (inputs(45)));
    layer0_outputs(592) <= not(inputs(218)) or (inputs(109));
    layer0_outputs(593) <= not((inputs(65)) or (inputs(31)));
    layer0_outputs(594) <= not((inputs(26)) or (inputs(3)));
    layer0_outputs(595) <= not((inputs(146)) or (inputs(149)));
    layer0_outputs(596) <= (inputs(140)) or (inputs(127));
    layer0_outputs(597) <= not(inputs(76));
    layer0_outputs(598) <= not(inputs(29));
    layer0_outputs(599) <= (inputs(34)) and not (inputs(30));
    layer0_outputs(600) <= not(inputs(131));
    layer0_outputs(601) <= not(inputs(72));
    layer0_outputs(602) <= not(inputs(141)) or (inputs(223));
    layer0_outputs(603) <= not((inputs(174)) or (inputs(112)));
    layer0_outputs(604) <= (inputs(112)) xor (inputs(84));
    layer0_outputs(605) <= not(inputs(39));
    layer0_outputs(606) <= (inputs(50)) xor (inputs(62));
    layer0_outputs(607) <= inputs(156);
    layer0_outputs(608) <= (inputs(136)) and not (inputs(31));
    layer0_outputs(609) <= (inputs(65)) and (inputs(111));
    layer0_outputs(610) <= inputs(252);
    layer0_outputs(611) <= not((inputs(22)) or (inputs(77)));
    layer0_outputs(612) <= (inputs(247)) and (inputs(166));
    layer0_outputs(613) <= (inputs(142)) and (inputs(98));
    layer0_outputs(614) <= (inputs(209)) and not (inputs(111));
    layer0_outputs(615) <= not(inputs(229)) or (inputs(166));
    layer0_outputs(616) <= not(inputs(99));
    layer0_outputs(617) <= not((inputs(154)) xor (inputs(165)));
    layer0_outputs(618) <= inputs(130);
    layer0_outputs(619) <= (inputs(40)) and not (inputs(182));
    layer0_outputs(620) <= not(inputs(246));
    layer0_outputs(621) <= (inputs(141)) or (inputs(85));
    layer0_outputs(622) <= '0';
    layer0_outputs(623) <= '0';
    layer0_outputs(624) <= not(inputs(171));
    layer0_outputs(625) <= inputs(42);
    layer0_outputs(626) <= (inputs(23)) and not (inputs(83));
    layer0_outputs(627) <= not(inputs(146));
    layer0_outputs(628) <= inputs(247);
    layer0_outputs(629) <= (inputs(213)) or (inputs(167));
    layer0_outputs(630) <= '0';
    layer0_outputs(631) <= not((inputs(145)) or (inputs(147)));
    layer0_outputs(632) <= inputs(181);
    layer0_outputs(633) <= (inputs(48)) and not (inputs(220));
    layer0_outputs(634) <= inputs(230);
    layer0_outputs(635) <= (inputs(155)) or (inputs(129));
    layer0_outputs(636) <= not(inputs(21)) or (inputs(141));
    layer0_outputs(637) <= (inputs(30)) and not (inputs(253));
    layer0_outputs(638) <= not((inputs(123)) or (inputs(44)));
    layer0_outputs(639) <= not(inputs(140));
    layer0_outputs(640) <= not((inputs(76)) or (inputs(93)));
    layer0_outputs(641) <= '0';
    layer0_outputs(642) <= (inputs(50)) and not (inputs(106));
    layer0_outputs(643) <= inputs(63);
    layer0_outputs(644) <= inputs(14);
    layer0_outputs(645) <= not(inputs(57));
    layer0_outputs(646) <= (inputs(136)) and not (inputs(0));
    layer0_outputs(647) <= not(inputs(105)) or (inputs(195));
    layer0_outputs(648) <= inputs(214);
    layer0_outputs(649) <= not(inputs(234));
    layer0_outputs(650) <= not(inputs(196)) or (inputs(158));
    layer0_outputs(651) <= (inputs(210)) and (inputs(161));
    layer0_outputs(652) <= (inputs(180)) and not (inputs(78));
    layer0_outputs(653) <= not((inputs(171)) and (inputs(184)));
    layer0_outputs(654) <= not(inputs(181)) or (inputs(58));
    layer0_outputs(655) <= inputs(18);
    layer0_outputs(656) <= (inputs(76)) and not (inputs(44));
    layer0_outputs(657) <= not((inputs(236)) and (inputs(97)));
    layer0_outputs(658) <= not(inputs(254));
    layer0_outputs(659) <= inputs(121);
    layer0_outputs(660) <= not((inputs(17)) or (inputs(179)));
    layer0_outputs(661) <= not(inputs(115));
    layer0_outputs(662) <= not(inputs(235));
    layer0_outputs(663) <= not(inputs(249));
    layer0_outputs(664) <= inputs(90);
    layer0_outputs(665) <= (inputs(158)) xor (inputs(85));
    layer0_outputs(666) <= inputs(161);
    layer0_outputs(667) <= not(inputs(180));
    layer0_outputs(668) <= inputs(2);
    layer0_outputs(669) <= (inputs(42)) and (inputs(222));
    layer0_outputs(670) <= not(inputs(117)) or (inputs(176));
    layer0_outputs(671) <= inputs(98);
    layer0_outputs(672) <= '0';
    layer0_outputs(673) <= (inputs(53)) and not (inputs(53));
    layer0_outputs(674) <= not(inputs(117));
    layer0_outputs(675) <= not((inputs(156)) and (inputs(232)));
    layer0_outputs(676) <= not(inputs(222));
    layer0_outputs(677) <= (inputs(144)) and not (inputs(12));
    layer0_outputs(678) <= (inputs(138)) and not (inputs(25));
    layer0_outputs(679) <= (inputs(59)) and (inputs(251));
    layer0_outputs(680) <= (inputs(96)) or (inputs(36));
    layer0_outputs(681) <= (inputs(86)) or (inputs(157));
    layer0_outputs(682) <= not(inputs(8)) or (inputs(200));
    layer0_outputs(683) <= not((inputs(171)) or (inputs(85)));
    layer0_outputs(684) <= '1';
    layer0_outputs(685) <= not((inputs(17)) or (inputs(222)));
    layer0_outputs(686) <= inputs(208);
    layer0_outputs(687) <= (inputs(219)) xor (inputs(162));
    layer0_outputs(688) <= not(inputs(105)) or (inputs(82));
    layer0_outputs(689) <= (inputs(95)) and not (inputs(121));
    layer0_outputs(690) <= not((inputs(83)) or (inputs(56)));
    layer0_outputs(691) <= inputs(40);
    layer0_outputs(692) <= '1';
    layer0_outputs(693) <= (inputs(228)) and (inputs(179));
    layer0_outputs(694) <= '1';
    layer0_outputs(695) <= (inputs(72)) or (inputs(198));
    layer0_outputs(696) <= not((inputs(193)) or (inputs(189)));
    layer0_outputs(697) <= '1';
    layer0_outputs(698) <= (inputs(199)) and (inputs(196));
    layer0_outputs(699) <= (inputs(36)) and not (inputs(191));
    layer0_outputs(700) <= not(inputs(28));
    layer0_outputs(701) <= (inputs(24)) and not (inputs(144));
    layer0_outputs(702) <= not(inputs(149));
    layer0_outputs(703) <= not(inputs(145));
    layer0_outputs(704) <= '1';
    layer0_outputs(705) <= not((inputs(101)) or (inputs(146)));
    layer0_outputs(706) <= '0';
    layer0_outputs(707) <= not((inputs(56)) xor (inputs(48)));
    layer0_outputs(708) <= not(inputs(43));
    layer0_outputs(709) <= '1';
    layer0_outputs(710) <= (inputs(232)) and not (inputs(50));
    layer0_outputs(711) <= (inputs(13)) xor (inputs(14));
    layer0_outputs(712) <= not(inputs(20)) or (inputs(255));
    layer0_outputs(713) <= not((inputs(3)) and (inputs(3)));
    layer0_outputs(714) <= (inputs(181)) or (inputs(127));
    layer0_outputs(715) <= not(inputs(168)) or (inputs(227));
    layer0_outputs(716) <= not(inputs(229));
    layer0_outputs(717) <= not(inputs(45)) or (inputs(101));
    layer0_outputs(718) <= not((inputs(199)) xor (inputs(225)));
    layer0_outputs(719) <= not((inputs(231)) xor (inputs(224)));
    layer0_outputs(720) <= inputs(83);
    layer0_outputs(721) <= inputs(120);
    layer0_outputs(722) <= inputs(45);
    layer0_outputs(723) <= inputs(222);
    layer0_outputs(724) <= not(inputs(150));
    layer0_outputs(725) <= (inputs(84)) and not (inputs(61));
    layer0_outputs(726) <= inputs(169);
    layer0_outputs(727) <= not(inputs(170));
    layer0_outputs(728) <= not((inputs(27)) and (inputs(247)));
    layer0_outputs(729) <= not(inputs(188)) or (inputs(254));
    layer0_outputs(730) <= not(inputs(173));
    layer0_outputs(731) <= not(inputs(75)) or (inputs(233));
    layer0_outputs(732) <= not(inputs(181));
    layer0_outputs(733) <= inputs(114);
    layer0_outputs(734) <= not(inputs(59)) or (inputs(172));
    layer0_outputs(735) <= inputs(149);
    layer0_outputs(736) <= not((inputs(240)) or (inputs(23)));
    layer0_outputs(737) <= not(inputs(219));
    layer0_outputs(738) <= (inputs(143)) or (inputs(100));
    layer0_outputs(739) <= not((inputs(8)) or (inputs(189)));
    layer0_outputs(740) <= inputs(173);
    layer0_outputs(741) <= '0';
    layer0_outputs(742) <= (inputs(245)) or (inputs(5));
    layer0_outputs(743) <= '0';
    layer0_outputs(744) <= not((inputs(88)) xor (inputs(108)));
    layer0_outputs(745) <= (inputs(130)) and not (inputs(145));
    layer0_outputs(746) <= (inputs(19)) and not (inputs(220));
    layer0_outputs(747) <= not(inputs(101));
    layer0_outputs(748) <= not(inputs(8));
    layer0_outputs(749) <= (inputs(111)) or (inputs(101));
    layer0_outputs(750) <= not((inputs(155)) or (inputs(115)));
    layer0_outputs(751) <= (inputs(247)) or (inputs(192));
    layer0_outputs(752) <= (inputs(209)) or (inputs(224));
    layer0_outputs(753) <= inputs(115);
    layer0_outputs(754) <= '1';
    layer0_outputs(755) <= not((inputs(47)) or (inputs(69)));
    layer0_outputs(756) <= (inputs(118)) and not (inputs(222));
    layer0_outputs(757) <= (inputs(220)) or (inputs(54));
    layer0_outputs(758) <= (inputs(73)) xor (inputs(170));
    layer0_outputs(759) <= not(inputs(106));
    layer0_outputs(760) <= not((inputs(92)) or (inputs(47)));
    layer0_outputs(761) <= not(inputs(76));
    layer0_outputs(762) <= (inputs(105)) and (inputs(212));
    layer0_outputs(763) <= (inputs(241)) or (inputs(103));
    layer0_outputs(764) <= (inputs(211)) and not (inputs(198));
    layer0_outputs(765) <= not((inputs(124)) or (inputs(237)));
    layer0_outputs(766) <= not((inputs(197)) or (inputs(66)));
    layer0_outputs(767) <= not(inputs(229)) or (inputs(122));
    layer0_outputs(768) <= (inputs(251)) and (inputs(211));
    layer0_outputs(769) <= not(inputs(246)) or (inputs(223));
    layer0_outputs(770) <= not(inputs(170)) or (inputs(0));
    layer0_outputs(771) <= '1';
    layer0_outputs(772) <= (inputs(147)) and (inputs(155));
    layer0_outputs(773) <= not((inputs(192)) or (inputs(173)));
    layer0_outputs(774) <= not((inputs(31)) xor (inputs(62)));
    layer0_outputs(775) <= inputs(136);
    layer0_outputs(776) <= inputs(55);
    layer0_outputs(777) <= (inputs(139)) and not (inputs(122));
    layer0_outputs(778) <= not(inputs(122)) or (inputs(15));
    layer0_outputs(779) <= not((inputs(183)) and (inputs(197)));
    layer0_outputs(780) <= not((inputs(109)) or (inputs(254)));
    layer0_outputs(781) <= (inputs(119)) and not (inputs(196));
    layer0_outputs(782) <= not(inputs(91)) or (inputs(66));
    layer0_outputs(783) <= inputs(161);
    layer0_outputs(784) <= '0';
    layer0_outputs(785) <= '0';
    layer0_outputs(786) <= not(inputs(168)) or (inputs(58));
    layer0_outputs(787) <= not(inputs(226)) or (inputs(239));
    layer0_outputs(788) <= (inputs(231)) and not (inputs(21));
    layer0_outputs(789) <= (inputs(72)) and not (inputs(208));
    layer0_outputs(790) <= not(inputs(245));
    layer0_outputs(791) <= not((inputs(33)) or (inputs(60)));
    layer0_outputs(792) <= inputs(228);
    layer0_outputs(793) <= inputs(74);
    layer0_outputs(794) <= inputs(109);
    layer0_outputs(795) <= not(inputs(40));
    layer0_outputs(796) <= not((inputs(215)) or (inputs(181)));
    layer0_outputs(797) <= not(inputs(150));
    layer0_outputs(798) <= inputs(233);
    layer0_outputs(799) <= not(inputs(209));
    layer0_outputs(800) <= not((inputs(40)) or (inputs(139)));
    layer0_outputs(801) <= '1';
    layer0_outputs(802) <= not(inputs(209));
    layer0_outputs(803) <= not((inputs(34)) or (inputs(195)));
    layer0_outputs(804) <= inputs(41);
    layer0_outputs(805) <= not(inputs(54)) or (inputs(235));
    layer0_outputs(806) <= (inputs(140)) or (inputs(35));
    layer0_outputs(807) <= '1';
    layer0_outputs(808) <= (inputs(138)) and not (inputs(102));
    layer0_outputs(809) <= (inputs(176)) and not (inputs(195));
    layer0_outputs(810) <= not((inputs(44)) and (inputs(233)));
    layer0_outputs(811) <= (inputs(178)) and not (inputs(107));
    layer0_outputs(812) <= inputs(237);
    layer0_outputs(813) <= inputs(222);
    layer0_outputs(814) <= (inputs(89)) and (inputs(158));
    layer0_outputs(815) <= (inputs(33)) or (inputs(179));
    layer0_outputs(816) <= not(inputs(102));
    layer0_outputs(817) <= (inputs(172)) xor (inputs(203));
    layer0_outputs(818) <= inputs(229);
    layer0_outputs(819) <= inputs(12);
    layer0_outputs(820) <= inputs(68);
    layer0_outputs(821) <= not(inputs(254));
    layer0_outputs(822) <= not(inputs(120)) or (inputs(181));
    layer0_outputs(823) <= (inputs(227)) or (inputs(44));
    layer0_outputs(824) <= not(inputs(43)) or (inputs(220));
    layer0_outputs(825) <= not(inputs(182));
    layer0_outputs(826) <= inputs(203);
    layer0_outputs(827) <= '0';
    layer0_outputs(828) <= (inputs(100)) and not (inputs(225));
    layer0_outputs(829) <= '0';
    layer0_outputs(830) <= '1';
    layer0_outputs(831) <= not(inputs(239));
    layer0_outputs(832) <= '0';
    layer0_outputs(833) <= not(inputs(175));
    layer0_outputs(834) <= not(inputs(138)) or (inputs(192));
    layer0_outputs(835) <= (inputs(205)) xor (inputs(189));
    layer0_outputs(836) <= inputs(214);
    layer0_outputs(837) <= not((inputs(226)) or (inputs(219)));
    layer0_outputs(838) <= (inputs(76)) and (inputs(30));
    layer0_outputs(839) <= (inputs(193)) and not (inputs(253));
    layer0_outputs(840) <= not((inputs(29)) or (inputs(160)));
    layer0_outputs(841) <= '1';
    layer0_outputs(842) <= (inputs(135)) xor (inputs(93));
    layer0_outputs(843) <= not((inputs(178)) or (inputs(162)));
    layer0_outputs(844) <= (inputs(218)) and (inputs(199));
    layer0_outputs(845) <= not(inputs(168)) or (inputs(206));
    layer0_outputs(846) <= not((inputs(138)) and (inputs(184)));
    layer0_outputs(847) <= inputs(192);
    layer0_outputs(848) <= '1';
    layer0_outputs(849) <= '1';
    layer0_outputs(850) <= '0';
    layer0_outputs(851) <= not(inputs(177));
    layer0_outputs(852) <= (inputs(168)) or (inputs(120));
    layer0_outputs(853) <= (inputs(216)) and (inputs(41));
    layer0_outputs(854) <= inputs(229);
    layer0_outputs(855) <= not(inputs(6)) or (inputs(250));
    layer0_outputs(856) <= not((inputs(17)) or (inputs(220)));
    layer0_outputs(857) <= inputs(209);
    layer0_outputs(858) <= inputs(136);
    layer0_outputs(859) <= (inputs(164)) and not (inputs(97));
    layer0_outputs(860) <= not(inputs(217));
    layer0_outputs(861) <= inputs(83);
    layer0_outputs(862) <= not(inputs(28)) or (inputs(70));
    layer0_outputs(863) <= '1';
    layer0_outputs(864) <= not((inputs(210)) or (inputs(231)));
    layer0_outputs(865) <= not(inputs(238));
    layer0_outputs(866) <= inputs(154);
    layer0_outputs(867) <= not((inputs(24)) or (inputs(179)));
    layer0_outputs(868) <= not(inputs(160));
    layer0_outputs(869) <= not(inputs(94));
    layer0_outputs(870) <= not((inputs(207)) xor (inputs(79)));
    layer0_outputs(871) <= '0';
    layer0_outputs(872) <= inputs(157);
    layer0_outputs(873) <= (inputs(30)) xor (inputs(122));
    layer0_outputs(874) <= inputs(172);
    layer0_outputs(875) <= '0';
    layer0_outputs(876) <= (inputs(67)) xor (inputs(21));
    layer0_outputs(877) <= not(inputs(4));
    layer0_outputs(878) <= (inputs(67)) and not (inputs(14));
    layer0_outputs(879) <= inputs(68);
    layer0_outputs(880) <= '0';
    layer0_outputs(881) <= (inputs(20)) xor (inputs(64));
    layer0_outputs(882) <= not((inputs(14)) or (inputs(135)));
    layer0_outputs(883) <= not(inputs(139)) or (inputs(100));
    layer0_outputs(884) <= not(inputs(109));
    layer0_outputs(885) <= not(inputs(53));
    layer0_outputs(886) <= '1';
    layer0_outputs(887) <= (inputs(149)) and not (inputs(134));
    layer0_outputs(888) <= not((inputs(182)) or (inputs(54)));
    layer0_outputs(889) <= not((inputs(0)) or (inputs(139)));
    layer0_outputs(890) <= not((inputs(11)) and (inputs(235)));
    layer0_outputs(891) <= inputs(218);
    layer0_outputs(892) <= inputs(181);
    layer0_outputs(893) <= not((inputs(124)) or (inputs(73)));
    layer0_outputs(894) <= not(inputs(89)) or (inputs(57));
    layer0_outputs(895) <= not((inputs(189)) or (inputs(226)));
    layer0_outputs(896) <= (inputs(33)) or (inputs(221));
    layer0_outputs(897) <= not((inputs(148)) or (inputs(110)));
    layer0_outputs(898) <= inputs(9);
    layer0_outputs(899) <= inputs(110);
    layer0_outputs(900) <= (inputs(23)) xor (inputs(127));
    layer0_outputs(901) <= not(inputs(197));
    layer0_outputs(902) <= not(inputs(149)) or (inputs(96));
    layer0_outputs(903) <= not(inputs(182));
    layer0_outputs(904) <= inputs(145);
    layer0_outputs(905) <= inputs(37);
    layer0_outputs(906) <= (inputs(83)) xor (inputs(177));
    layer0_outputs(907) <= not(inputs(97));
    layer0_outputs(908) <= (inputs(0)) or (inputs(48));
    layer0_outputs(909) <= not(inputs(146));
    layer0_outputs(910) <= (inputs(134)) and not (inputs(219));
    layer0_outputs(911) <= (inputs(67)) and not (inputs(192));
    layer0_outputs(912) <= not((inputs(222)) or (inputs(221)));
    layer0_outputs(913) <= inputs(57);
    layer0_outputs(914) <= inputs(149);
    layer0_outputs(915) <= inputs(84);
    layer0_outputs(916) <= inputs(219);
    layer0_outputs(917) <= (inputs(155)) and not (inputs(21));
    layer0_outputs(918) <= inputs(89);
    layer0_outputs(919) <= (inputs(60)) and not (inputs(254));
    layer0_outputs(920) <= inputs(229);
    layer0_outputs(921) <= (inputs(197)) and not (inputs(16));
    layer0_outputs(922) <= not(inputs(139));
    layer0_outputs(923) <= (inputs(83)) or (inputs(44));
    layer0_outputs(924) <= (inputs(175)) xor (inputs(145));
    layer0_outputs(925) <= '0';
    layer0_outputs(926) <= inputs(166);
    layer0_outputs(927) <= inputs(51);
    layer0_outputs(928) <= '1';
    layer0_outputs(929) <= inputs(248);
    layer0_outputs(930) <= not(inputs(17)) or (inputs(79));
    layer0_outputs(931) <= '1';
    layer0_outputs(932) <= not(inputs(170)) or (inputs(41));
    layer0_outputs(933) <= '0';
    layer0_outputs(934) <= '1';
    layer0_outputs(935) <= (inputs(221)) and not (inputs(61));
    layer0_outputs(936) <= (inputs(42)) and not (inputs(136));
    layer0_outputs(937) <= '0';
    layer0_outputs(938) <= (inputs(56)) and not (inputs(103));
    layer0_outputs(939) <= (inputs(182)) or (inputs(195));
    layer0_outputs(940) <= (inputs(20)) xor (inputs(187));
    layer0_outputs(941) <= '0';
    layer0_outputs(942) <= '1';
    layer0_outputs(943) <= (inputs(221)) and not (inputs(250));
    layer0_outputs(944) <= (inputs(204)) and not (inputs(197));
    layer0_outputs(945) <= (inputs(12)) xor (inputs(177));
    layer0_outputs(946) <= inputs(193);
    layer0_outputs(947) <= inputs(106);
    layer0_outputs(948) <= not((inputs(126)) or (inputs(34)));
    layer0_outputs(949) <= inputs(148);
    layer0_outputs(950) <= not(inputs(242));
    layer0_outputs(951) <= (inputs(183)) or (inputs(85));
    layer0_outputs(952) <= not(inputs(72));
    layer0_outputs(953) <= (inputs(22)) xor (inputs(74));
    layer0_outputs(954) <= (inputs(98)) and not (inputs(146));
    layer0_outputs(955) <= '1';
    layer0_outputs(956) <= not(inputs(119)) or (inputs(2));
    layer0_outputs(957) <= not(inputs(25));
    layer0_outputs(958) <= not(inputs(89));
    layer0_outputs(959) <= not(inputs(152));
    layer0_outputs(960) <= (inputs(3)) or (inputs(24));
    layer0_outputs(961) <= (inputs(57)) and not (inputs(102));
    layer0_outputs(962) <= not(inputs(237));
    layer0_outputs(963) <= not(inputs(253));
    layer0_outputs(964) <= not(inputs(181));
    layer0_outputs(965) <= (inputs(35)) or (inputs(59));
    layer0_outputs(966) <= not(inputs(201));
    layer0_outputs(967) <= not(inputs(212)) or (inputs(61));
    layer0_outputs(968) <= (inputs(166)) and not (inputs(192));
    layer0_outputs(969) <= not(inputs(88)) or (inputs(35));
    layer0_outputs(970) <= not((inputs(82)) xor (inputs(228)));
    layer0_outputs(971) <= (inputs(171)) or (inputs(68));
    layer0_outputs(972) <= (inputs(154)) and not (inputs(35));
    layer0_outputs(973) <= not(inputs(240)) or (inputs(216));
    layer0_outputs(974) <= not(inputs(49));
    layer0_outputs(975) <= '0';
    layer0_outputs(976) <= (inputs(170)) or (inputs(172));
    layer0_outputs(977) <= not(inputs(143));
    layer0_outputs(978) <= '1';
    layer0_outputs(979) <= (inputs(156)) and not (inputs(161));
    layer0_outputs(980) <= (inputs(119)) and not (inputs(67));
    layer0_outputs(981) <= not(inputs(38)) or (inputs(204));
    layer0_outputs(982) <= (inputs(199)) xor (inputs(14));
    layer0_outputs(983) <= inputs(162);
    layer0_outputs(984) <= inputs(220);
    layer0_outputs(985) <= inputs(211);
    layer0_outputs(986) <= not(inputs(25));
    layer0_outputs(987) <= not(inputs(100)) or (inputs(33));
    layer0_outputs(988) <= not(inputs(28)) or (inputs(161));
    layer0_outputs(989) <= not((inputs(128)) xor (inputs(205)));
    layer0_outputs(990) <= '1';
    layer0_outputs(991) <= inputs(101);
    layer0_outputs(992) <= (inputs(193)) or (inputs(220));
    layer0_outputs(993) <= not((inputs(90)) and (inputs(69)));
    layer0_outputs(994) <= not((inputs(191)) or (inputs(96)));
    layer0_outputs(995) <= not(inputs(227)) or (inputs(159));
    layer0_outputs(996) <= inputs(180);
    layer0_outputs(997) <= not((inputs(7)) or (inputs(51)));
    layer0_outputs(998) <= (inputs(46)) or (inputs(66));
    layer0_outputs(999) <= '1';
    layer0_outputs(1000) <= inputs(35);
    layer0_outputs(1001) <= '0';
    layer0_outputs(1002) <= '1';
    layer0_outputs(1003) <= not(inputs(51)) or (inputs(129));
    layer0_outputs(1004) <= not(inputs(82));
    layer0_outputs(1005) <= (inputs(60)) and not (inputs(103));
    layer0_outputs(1006) <= inputs(145);
    layer0_outputs(1007) <= not(inputs(74)) or (inputs(249));
    layer0_outputs(1008) <= (inputs(117)) and (inputs(36));
    layer0_outputs(1009) <= not(inputs(85));
    layer0_outputs(1010) <= not(inputs(201)) or (inputs(185));
    layer0_outputs(1011) <= '0';
    layer0_outputs(1012) <= inputs(48);
    layer0_outputs(1013) <= inputs(153);
    layer0_outputs(1014) <= not(inputs(74));
    layer0_outputs(1015) <= not(inputs(161));
    layer0_outputs(1016) <= inputs(62);
    layer0_outputs(1017) <= not(inputs(204)) or (inputs(64));
    layer0_outputs(1018) <= not(inputs(168));
    layer0_outputs(1019) <= inputs(193);
    layer0_outputs(1020) <= not((inputs(108)) or (inputs(84)));
    layer0_outputs(1021) <= (inputs(88)) and not (inputs(1));
    layer0_outputs(1022) <= inputs(221);
    layer0_outputs(1023) <= not(inputs(105));
    layer0_outputs(1024) <= (inputs(39)) and not (inputs(119));
    layer0_outputs(1025) <= (inputs(127)) and not (inputs(59));
    layer0_outputs(1026) <= not(inputs(139));
    layer0_outputs(1027) <= inputs(231);
    layer0_outputs(1028) <= not((inputs(60)) and (inputs(13)));
    layer0_outputs(1029) <= not(inputs(232));
    layer0_outputs(1030) <= not((inputs(69)) xor (inputs(48)));
    layer0_outputs(1031) <= (inputs(28)) and not (inputs(125));
    layer0_outputs(1032) <= (inputs(202)) xor (inputs(208));
    layer0_outputs(1033) <= not((inputs(205)) or (inputs(165)));
    layer0_outputs(1034) <= inputs(240);
    layer0_outputs(1035) <= not(inputs(150));
    layer0_outputs(1036) <= not(inputs(106)) or (inputs(96));
    layer0_outputs(1037) <= not(inputs(41));
    layer0_outputs(1038) <= inputs(91);
    layer0_outputs(1039) <= (inputs(57)) xor (inputs(58));
    layer0_outputs(1040) <= (inputs(41)) or (inputs(75));
    layer0_outputs(1041) <= not((inputs(7)) or (inputs(11)));
    layer0_outputs(1042) <= inputs(146);
    layer0_outputs(1043) <= inputs(189);
    layer0_outputs(1044) <= not(inputs(54)) or (inputs(217));
    layer0_outputs(1045) <= not((inputs(18)) xor (inputs(20)));
    layer0_outputs(1046) <= not(inputs(5)) or (inputs(178));
    layer0_outputs(1047) <= not(inputs(243));
    layer0_outputs(1048) <= (inputs(254)) or (inputs(6));
    layer0_outputs(1049) <= not(inputs(165));
    layer0_outputs(1050) <= not(inputs(212)) or (inputs(3));
    layer0_outputs(1051) <= not(inputs(142)) or (inputs(151));
    layer0_outputs(1052) <= '0';
    layer0_outputs(1053) <= not(inputs(185)) or (inputs(117));
    layer0_outputs(1054) <= '0';
    layer0_outputs(1055) <= not((inputs(163)) or (inputs(198)));
    layer0_outputs(1056) <= not(inputs(29));
    layer0_outputs(1057) <= (inputs(148)) xor (inputs(118));
    layer0_outputs(1058) <= not(inputs(240)) or (inputs(139));
    layer0_outputs(1059) <= inputs(124);
    layer0_outputs(1060) <= '0';
    layer0_outputs(1061) <= not(inputs(49));
    layer0_outputs(1062) <= '0';
    layer0_outputs(1063) <= (inputs(205)) or (inputs(4));
    layer0_outputs(1064) <= not((inputs(206)) or (inputs(188)));
    layer0_outputs(1065) <= not(inputs(143)) or (inputs(27));
    layer0_outputs(1066) <= not((inputs(178)) or (inputs(238)));
    layer0_outputs(1067) <= not((inputs(67)) or (inputs(114)));
    layer0_outputs(1068) <= not((inputs(167)) or (inputs(252)));
    layer0_outputs(1069) <= (inputs(78)) or (inputs(10));
    layer0_outputs(1070) <= (inputs(203)) and (inputs(177));
    layer0_outputs(1071) <= inputs(159);
    layer0_outputs(1072) <= not(inputs(138)) or (inputs(113));
    layer0_outputs(1073) <= (inputs(217)) and not (inputs(110));
    layer0_outputs(1074) <= '0';
    layer0_outputs(1075) <= not(inputs(236)) or (inputs(77));
    layer0_outputs(1076) <= (inputs(102)) and (inputs(69));
    layer0_outputs(1077) <= not((inputs(84)) or (inputs(110)));
    layer0_outputs(1078) <= not((inputs(224)) or (inputs(36)));
    layer0_outputs(1079) <= (inputs(68)) or (inputs(220));
    layer0_outputs(1080) <= not(inputs(62));
    layer0_outputs(1081) <= (inputs(126)) and not (inputs(207));
    layer0_outputs(1082) <= not((inputs(118)) or (inputs(133)));
    layer0_outputs(1083) <= not((inputs(138)) xor (inputs(73)));
    layer0_outputs(1084) <= not((inputs(194)) or (inputs(235)));
    layer0_outputs(1085) <= inputs(182);
    layer0_outputs(1086) <= '1';
    layer0_outputs(1087) <= '0';
    layer0_outputs(1088) <= not(inputs(2));
    layer0_outputs(1089) <= not((inputs(165)) or (inputs(18)));
    layer0_outputs(1090) <= not((inputs(5)) or (inputs(206)));
    layer0_outputs(1091) <= inputs(119);
    layer0_outputs(1092) <= '0';
    layer0_outputs(1093) <= not(inputs(162));
    layer0_outputs(1094) <= (inputs(154)) and not (inputs(169));
    layer0_outputs(1095) <= inputs(195);
    layer0_outputs(1096) <= (inputs(71)) and not (inputs(100));
    layer0_outputs(1097) <= inputs(72);
    layer0_outputs(1098) <= not(inputs(191));
    layer0_outputs(1099) <= not((inputs(72)) or (inputs(92)));
    layer0_outputs(1100) <= not((inputs(81)) or (inputs(53)));
    layer0_outputs(1101) <= (inputs(115)) and not (inputs(39));
    layer0_outputs(1102) <= not((inputs(85)) and (inputs(212)));
    layer0_outputs(1103) <= not(inputs(121));
    layer0_outputs(1104) <= (inputs(58)) and (inputs(55));
    layer0_outputs(1105) <= not(inputs(193)) or (inputs(226));
    layer0_outputs(1106) <= inputs(232);
    layer0_outputs(1107) <= (inputs(114)) or (inputs(151));
    layer0_outputs(1108) <= (inputs(232)) and not (inputs(32));
    layer0_outputs(1109) <= (inputs(4)) xor (inputs(9));
    layer0_outputs(1110) <= (inputs(160)) and (inputs(126));
    layer0_outputs(1111) <= (inputs(132)) or (inputs(38));
    layer0_outputs(1112) <= not((inputs(23)) xor (inputs(71)));
    layer0_outputs(1113) <= not((inputs(202)) or (inputs(185)));
    layer0_outputs(1114) <= not(inputs(122));
    layer0_outputs(1115) <= not(inputs(13)) or (inputs(121));
    layer0_outputs(1116) <= (inputs(118)) and not (inputs(57));
    layer0_outputs(1117) <= not(inputs(26)) or (inputs(192));
    layer0_outputs(1118) <= not((inputs(112)) or (inputs(251)));
    layer0_outputs(1119) <= not(inputs(103)) or (inputs(200));
    layer0_outputs(1120) <= inputs(196);
    layer0_outputs(1121) <= not(inputs(152));
    layer0_outputs(1122) <= not(inputs(86));
    layer0_outputs(1123) <= not(inputs(202));
    layer0_outputs(1124) <= not((inputs(26)) xor (inputs(1)));
    layer0_outputs(1125) <= inputs(115);
    layer0_outputs(1126) <= inputs(8);
    layer0_outputs(1127) <= (inputs(3)) or (inputs(5));
    layer0_outputs(1128) <= not(inputs(99));
    layer0_outputs(1129) <= not((inputs(118)) or (inputs(237)));
    layer0_outputs(1130) <= not(inputs(200));
    layer0_outputs(1131) <= not(inputs(149));
    layer0_outputs(1132) <= not((inputs(186)) and (inputs(251)));
    layer0_outputs(1133) <= inputs(109);
    layer0_outputs(1134) <= not(inputs(183));
    layer0_outputs(1135) <= (inputs(178)) or (inputs(198));
    layer0_outputs(1136) <= inputs(114);
    layer0_outputs(1137) <= not((inputs(74)) or (inputs(20)));
    layer0_outputs(1138) <= not((inputs(255)) xor (inputs(119)));
    layer0_outputs(1139) <= inputs(101);
    layer0_outputs(1140) <= (inputs(217)) or (inputs(54));
    layer0_outputs(1141) <= inputs(233);
    layer0_outputs(1142) <= not((inputs(81)) or (inputs(97)));
    layer0_outputs(1143) <= (inputs(20)) or (inputs(197));
    layer0_outputs(1144) <= inputs(24);
    layer0_outputs(1145) <= inputs(62);
    layer0_outputs(1146) <= (inputs(167)) and not (inputs(156));
    layer0_outputs(1147) <= '1';
    layer0_outputs(1148) <= '1';
    layer0_outputs(1149) <= (inputs(12)) and not (inputs(75));
    layer0_outputs(1150) <= (inputs(115)) or (inputs(116));
    layer0_outputs(1151) <= not(inputs(162));
    layer0_outputs(1152) <= (inputs(109)) or (inputs(116));
    layer0_outputs(1153) <= not(inputs(77));
    layer0_outputs(1154) <= (inputs(248)) or (inputs(195));
    layer0_outputs(1155) <= '0';
    layer0_outputs(1156) <= not(inputs(10));
    layer0_outputs(1157) <= not(inputs(201));
    layer0_outputs(1158) <= inputs(194);
    layer0_outputs(1159) <= inputs(3);
    layer0_outputs(1160) <= (inputs(183)) and not (inputs(48));
    layer0_outputs(1161) <= (inputs(152)) xor (inputs(158));
    layer0_outputs(1162) <= not((inputs(24)) or (inputs(41)));
    layer0_outputs(1163) <= (inputs(51)) and (inputs(42));
    layer0_outputs(1164) <= '1';
    layer0_outputs(1165) <= (inputs(26)) and not (inputs(162));
    layer0_outputs(1166) <= (inputs(204)) and not (inputs(67));
    layer0_outputs(1167) <= not(inputs(177)) or (inputs(113));
    layer0_outputs(1168) <= not(inputs(16));
    layer0_outputs(1169) <= inputs(60);
    layer0_outputs(1170) <= (inputs(122)) or (inputs(236));
    layer0_outputs(1171) <= (inputs(100)) and not (inputs(191));
    layer0_outputs(1172) <= inputs(136);
    layer0_outputs(1173) <= inputs(92);
    layer0_outputs(1174) <= not((inputs(23)) or (inputs(108)));
    layer0_outputs(1175) <= not(inputs(45));
    layer0_outputs(1176) <= (inputs(53)) or (inputs(61));
    layer0_outputs(1177) <= '0';
    layer0_outputs(1178) <= (inputs(188)) and not (inputs(86));
    layer0_outputs(1179) <= inputs(87);
    layer0_outputs(1180) <= inputs(45);
    layer0_outputs(1181) <= not((inputs(250)) or (inputs(206)));
    layer0_outputs(1182) <= not(inputs(101));
    layer0_outputs(1183) <= not((inputs(212)) or (inputs(211)));
    layer0_outputs(1184) <= '1';
    layer0_outputs(1185) <= not((inputs(41)) or (inputs(252)));
    layer0_outputs(1186) <= (inputs(133)) or (inputs(112));
    layer0_outputs(1187) <= (inputs(134)) and not (inputs(192));
    layer0_outputs(1188) <= inputs(196);
    layer0_outputs(1189) <= (inputs(36)) xor (inputs(21));
    layer0_outputs(1190) <= (inputs(110)) or (inputs(193));
    layer0_outputs(1191) <= '1';
    layer0_outputs(1192) <= not((inputs(163)) xor (inputs(4)));
    layer0_outputs(1193) <= (inputs(63)) or (inputs(76));
    layer0_outputs(1194) <= not(inputs(93));
    layer0_outputs(1195) <= inputs(67);
    layer0_outputs(1196) <= inputs(122);
    layer0_outputs(1197) <= '0';
    layer0_outputs(1198) <= (inputs(214)) and not (inputs(75));
    layer0_outputs(1199) <= '1';
    layer0_outputs(1200) <= inputs(119);
    layer0_outputs(1201) <= '1';
    layer0_outputs(1202) <= not(inputs(187));
    layer0_outputs(1203) <= not((inputs(149)) xor (inputs(177)));
    layer0_outputs(1204) <= not((inputs(218)) or (inputs(188)));
    layer0_outputs(1205) <= (inputs(1)) and not (inputs(224));
    layer0_outputs(1206) <= not(inputs(165)) or (inputs(170));
    layer0_outputs(1207) <= (inputs(231)) or (inputs(191));
    layer0_outputs(1208) <= '0';
    layer0_outputs(1209) <= not((inputs(91)) xor (inputs(253)));
    layer0_outputs(1210) <= not(inputs(139));
    layer0_outputs(1211) <= inputs(109);
    layer0_outputs(1212) <= not(inputs(131));
    layer0_outputs(1213) <= inputs(126);
    layer0_outputs(1214) <= not(inputs(107));
    layer0_outputs(1215) <= inputs(106);
    layer0_outputs(1216) <= not(inputs(89));
    layer0_outputs(1217) <= not(inputs(179)) or (inputs(156));
    layer0_outputs(1218) <= not((inputs(249)) or (inputs(228)));
    layer0_outputs(1219) <= (inputs(216)) and not (inputs(129));
    layer0_outputs(1220) <= not((inputs(35)) xor (inputs(93)));
    layer0_outputs(1221) <= not(inputs(38)) or (inputs(15));
    layer0_outputs(1222) <= (inputs(128)) or (inputs(164));
    layer0_outputs(1223) <= (inputs(141)) xor (inputs(107));
    layer0_outputs(1224) <= not(inputs(229)) or (inputs(150));
    layer0_outputs(1225) <= inputs(26);
    layer0_outputs(1226) <= (inputs(103)) or (inputs(122));
    layer0_outputs(1227) <= (inputs(237)) and not (inputs(187));
    layer0_outputs(1228) <= inputs(210);
    layer0_outputs(1229) <= (inputs(193)) xor (inputs(253));
    layer0_outputs(1230) <= (inputs(157)) xor (inputs(138));
    layer0_outputs(1231) <= not((inputs(36)) or (inputs(67)));
    layer0_outputs(1232) <= (inputs(243)) and not (inputs(155));
    layer0_outputs(1233) <= '0';
    layer0_outputs(1234) <= inputs(91);
    layer0_outputs(1235) <= (inputs(34)) and not (inputs(144));
    layer0_outputs(1236) <= not((inputs(28)) or (inputs(4)));
    layer0_outputs(1237) <= (inputs(175)) and (inputs(86));
    layer0_outputs(1238) <= '0';
    layer0_outputs(1239) <= not(inputs(40)) or (inputs(144));
    layer0_outputs(1240) <= inputs(16);
    layer0_outputs(1241) <= not(inputs(197)) or (inputs(130));
    layer0_outputs(1242) <= not((inputs(76)) and (inputs(172)));
    layer0_outputs(1243) <= (inputs(144)) or (inputs(211));
    layer0_outputs(1244) <= (inputs(154)) or (inputs(174));
    layer0_outputs(1245) <= inputs(62);
    layer0_outputs(1246) <= not((inputs(90)) or (inputs(61)));
    layer0_outputs(1247) <= inputs(232);
    layer0_outputs(1248) <= (inputs(102)) or (inputs(178));
    layer0_outputs(1249) <= not(inputs(246)) or (inputs(168));
    layer0_outputs(1250) <= not((inputs(174)) xor (inputs(127)));
    layer0_outputs(1251) <= '0';
    layer0_outputs(1252) <= not((inputs(124)) or (inputs(31)));
    layer0_outputs(1253) <= inputs(177);
    layer0_outputs(1254) <= inputs(253);
    layer0_outputs(1255) <= not(inputs(70));
    layer0_outputs(1256) <= inputs(97);
    layer0_outputs(1257) <= inputs(81);
    layer0_outputs(1258) <= (inputs(103)) and not (inputs(187));
    layer0_outputs(1259) <= '0';
    layer0_outputs(1260) <= not(inputs(217));
    layer0_outputs(1261) <= not((inputs(133)) and (inputs(216)));
    layer0_outputs(1262) <= '1';
    layer0_outputs(1263) <= inputs(117);
    layer0_outputs(1264) <= not((inputs(183)) xor (inputs(151)));
    layer0_outputs(1265) <= inputs(234);
    layer0_outputs(1266) <= (inputs(100)) and (inputs(41));
    layer0_outputs(1267) <= not(inputs(204)) or (inputs(47));
    layer0_outputs(1268) <= inputs(222);
    layer0_outputs(1269) <= (inputs(190)) or (inputs(173));
    layer0_outputs(1270) <= not(inputs(209));
    layer0_outputs(1271) <= (inputs(173)) or (inputs(247));
    layer0_outputs(1272) <= (inputs(197)) and not (inputs(14));
    layer0_outputs(1273) <= not((inputs(234)) and (inputs(80)));
    layer0_outputs(1274) <= (inputs(201)) xor (inputs(170));
    layer0_outputs(1275) <= inputs(135);
    layer0_outputs(1276) <= not(inputs(100));
    layer0_outputs(1277) <= not((inputs(138)) or (inputs(153)));
    layer0_outputs(1278) <= inputs(49);
    layer0_outputs(1279) <= not(inputs(54)) or (inputs(222));
    layer0_outputs(1280) <= (inputs(228)) or (inputs(127));
    layer0_outputs(1281) <= not(inputs(183)) or (inputs(48));
    layer0_outputs(1282) <= not(inputs(46)) or (inputs(248));
    layer0_outputs(1283) <= (inputs(33)) and (inputs(67));
    layer0_outputs(1284) <= not(inputs(196));
    layer0_outputs(1285) <= inputs(7);
    layer0_outputs(1286) <= inputs(107);
    layer0_outputs(1287) <= (inputs(65)) xor (inputs(10));
    layer0_outputs(1288) <= not(inputs(252));
    layer0_outputs(1289) <= (inputs(218)) and not (inputs(70));
    layer0_outputs(1290) <= not(inputs(108));
    layer0_outputs(1291) <= not(inputs(189)) or (inputs(31));
    layer0_outputs(1292) <= inputs(143);
    layer0_outputs(1293) <= (inputs(64)) or (inputs(35));
    layer0_outputs(1294) <= (inputs(91)) and not (inputs(55));
    layer0_outputs(1295) <= inputs(196);
    layer0_outputs(1296) <= (inputs(141)) or (inputs(140));
    layer0_outputs(1297) <= not((inputs(175)) or (inputs(140)));
    layer0_outputs(1298) <= not(inputs(255)) or (inputs(202));
    layer0_outputs(1299) <= not(inputs(14));
    layer0_outputs(1300) <= (inputs(88)) or (inputs(205));
    layer0_outputs(1301) <= (inputs(171)) and not (inputs(48));
    layer0_outputs(1302) <= '1';
    layer0_outputs(1303) <= (inputs(41)) and not (inputs(19));
    layer0_outputs(1304) <= inputs(198);
    layer0_outputs(1305) <= not(inputs(189));
    layer0_outputs(1306) <= not(inputs(156)) or (inputs(6));
    layer0_outputs(1307) <= inputs(136);
    layer0_outputs(1308) <= inputs(60);
    layer0_outputs(1309) <= not(inputs(127)) or (inputs(238));
    layer0_outputs(1310) <= not(inputs(187)) or (inputs(186));
    layer0_outputs(1311) <= (inputs(173)) or (inputs(21));
    layer0_outputs(1312) <= not(inputs(141));
    layer0_outputs(1313) <= inputs(60);
    layer0_outputs(1314) <= not(inputs(171));
    layer0_outputs(1315) <= not(inputs(163));
    layer0_outputs(1316) <= (inputs(244)) and (inputs(157));
    layer0_outputs(1317) <= not(inputs(233));
    layer0_outputs(1318) <= (inputs(139)) and (inputs(169));
    layer0_outputs(1319) <= inputs(122);
    layer0_outputs(1320) <= not(inputs(241)) or (inputs(172));
    layer0_outputs(1321) <= not(inputs(157));
    layer0_outputs(1322) <= '0';
    layer0_outputs(1323) <= inputs(162);
    layer0_outputs(1324) <= not(inputs(131));
    layer0_outputs(1325) <= '0';
    layer0_outputs(1326) <= inputs(162);
    layer0_outputs(1327) <= (inputs(44)) and (inputs(5));
    layer0_outputs(1328) <= not((inputs(138)) or (inputs(102)));
    layer0_outputs(1329) <= inputs(2);
    layer0_outputs(1330) <= inputs(196);
    layer0_outputs(1331) <= (inputs(12)) and (inputs(70));
    layer0_outputs(1332) <= (inputs(132)) or (inputs(134));
    layer0_outputs(1333) <= not(inputs(225));
    layer0_outputs(1334) <= not(inputs(148));
    layer0_outputs(1335) <= inputs(169);
    layer0_outputs(1336) <= (inputs(84)) and (inputs(196));
    layer0_outputs(1337) <= (inputs(135)) and not (inputs(20));
    layer0_outputs(1338) <= not(inputs(50));
    layer0_outputs(1339) <= inputs(98);
    layer0_outputs(1340) <= not(inputs(165));
    layer0_outputs(1341) <= '1';
    layer0_outputs(1342) <= '1';
    layer0_outputs(1343) <= not(inputs(133)) or (inputs(141));
    layer0_outputs(1344) <= (inputs(145)) xor (inputs(218));
    layer0_outputs(1345) <= (inputs(252)) xor (inputs(123));
    layer0_outputs(1346) <= not(inputs(186)) or (inputs(144));
    layer0_outputs(1347) <= not(inputs(94));
    layer0_outputs(1348) <= inputs(238);
    layer0_outputs(1349) <= inputs(65);
    layer0_outputs(1350) <= (inputs(24)) and not (inputs(240));
    layer0_outputs(1351) <= inputs(58);
    layer0_outputs(1352) <= (inputs(83)) and not (inputs(142));
    layer0_outputs(1353) <= not((inputs(16)) or (inputs(94)));
    layer0_outputs(1354) <= inputs(29);
    layer0_outputs(1355) <= (inputs(8)) xor (inputs(47));
    layer0_outputs(1356) <= (inputs(7)) or (inputs(225));
    layer0_outputs(1357) <= inputs(218);
    layer0_outputs(1358) <= not(inputs(32)) or (inputs(65));
    layer0_outputs(1359) <= inputs(245);
    layer0_outputs(1360) <= (inputs(49)) and not (inputs(82));
    layer0_outputs(1361) <= not((inputs(58)) and (inputs(109)));
    layer0_outputs(1362) <= not(inputs(70)) or (inputs(124));
    layer0_outputs(1363) <= '0';
    layer0_outputs(1364) <= '0';
    layer0_outputs(1365) <= inputs(237);
    layer0_outputs(1366) <= not((inputs(203)) or (inputs(154)));
    layer0_outputs(1367) <= not(inputs(228));
    layer0_outputs(1368) <= not((inputs(43)) and (inputs(40)));
    layer0_outputs(1369) <= (inputs(175)) and not (inputs(166));
    layer0_outputs(1370) <= inputs(91);
    layer0_outputs(1371) <= inputs(157);
    layer0_outputs(1372) <= not(inputs(134)) or (inputs(185));
    layer0_outputs(1373) <= inputs(75);
    layer0_outputs(1374) <= (inputs(205)) or (inputs(162));
    layer0_outputs(1375) <= (inputs(181)) xor (inputs(112));
    layer0_outputs(1376) <= not((inputs(49)) or (inputs(180)));
    layer0_outputs(1377) <= (inputs(87)) and not (inputs(159));
    layer0_outputs(1378) <= not((inputs(133)) or (inputs(130)));
    layer0_outputs(1379) <= not((inputs(85)) or (inputs(250)));
    layer0_outputs(1380) <= (inputs(37)) and not (inputs(188));
    layer0_outputs(1381) <= not(inputs(73));
    layer0_outputs(1382) <= '0';
    layer0_outputs(1383) <= not(inputs(4));
    layer0_outputs(1384) <= inputs(65);
    layer0_outputs(1385) <= not(inputs(140));
    layer0_outputs(1386) <= not(inputs(52)) or (inputs(115));
    layer0_outputs(1387) <= (inputs(164)) and not (inputs(29));
    layer0_outputs(1388) <= '1';
    layer0_outputs(1389) <= inputs(33);
    layer0_outputs(1390) <= inputs(121);
    layer0_outputs(1391) <= not(inputs(110));
    layer0_outputs(1392) <= (inputs(230)) or (inputs(193));
    layer0_outputs(1393) <= (inputs(209)) or (inputs(190));
    layer0_outputs(1394) <= not(inputs(144)) or (inputs(189));
    layer0_outputs(1395) <= not(inputs(66));
    layer0_outputs(1396) <= (inputs(59)) and not (inputs(238));
    layer0_outputs(1397) <= inputs(24);
    layer0_outputs(1398) <= not(inputs(19)) or (inputs(254));
    layer0_outputs(1399) <= not(inputs(141));
    layer0_outputs(1400) <= not(inputs(147));
    layer0_outputs(1401) <= not(inputs(111));
    layer0_outputs(1402) <= inputs(249);
    layer0_outputs(1403) <= inputs(158);
    layer0_outputs(1404) <= inputs(228);
    layer0_outputs(1405) <= not((inputs(236)) or (inputs(33)));
    layer0_outputs(1406) <= (inputs(214)) or (inputs(177));
    layer0_outputs(1407) <= not(inputs(204)) or (inputs(48));
    layer0_outputs(1408) <= (inputs(246)) or (inputs(222));
    layer0_outputs(1409) <= (inputs(208)) or (inputs(82));
    layer0_outputs(1410) <= '1';
    layer0_outputs(1411) <= not(inputs(82));
    layer0_outputs(1412) <= '1';
    layer0_outputs(1413) <= not(inputs(84));
    layer0_outputs(1414) <= inputs(235);
    layer0_outputs(1415) <= (inputs(131)) or (inputs(2));
    layer0_outputs(1416) <= (inputs(28)) or (inputs(67));
    layer0_outputs(1417) <= (inputs(131)) and not (inputs(6));
    layer0_outputs(1418) <= '1';
    layer0_outputs(1419) <= inputs(63);
    layer0_outputs(1420) <= not(inputs(34)) or (inputs(214));
    layer0_outputs(1421) <= not((inputs(15)) or (inputs(116)));
    layer0_outputs(1422) <= (inputs(161)) or (inputs(246));
    layer0_outputs(1423) <= (inputs(101)) or (inputs(133));
    layer0_outputs(1424) <= inputs(56);
    layer0_outputs(1425) <= inputs(85);
    layer0_outputs(1426) <= inputs(1);
    layer0_outputs(1427) <= inputs(52);
    layer0_outputs(1428) <= not((inputs(82)) or (inputs(68)));
    layer0_outputs(1429) <= (inputs(78)) xor (inputs(36));
    layer0_outputs(1430) <= not(inputs(128));
    layer0_outputs(1431) <= (inputs(141)) and not (inputs(203));
    layer0_outputs(1432) <= (inputs(66)) and not (inputs(99));
    layer0_outputs(1433) <= inputs(99);
    layer0_outputs(1434) <= (inputs(104)) or (inputs(130));
    layer0_outputs(1435) <= (inputs(161)) or (inputs(94));
    layer0_outputs(1436) <= '0';
    layer0_outputs(1437) <= inputs(178);
    layer0_outputs(1438) <= '1';
    layer0_outputs(1439) <= not((inputs(70)) xor (inputs(251)));
    layer0_outputs(1440) <= inputs(0);
    layer0_outputs(1441) <= (inputs(100)) and not (inputs(191));
    layer0_outputs(1442) <= not(inputs(138)) or (inputs(189));
    layer0_outputs(1443) <= not((inputs(88)) or (inputs(89)));
    layer0_outputs(1444) <= (inputs(95)) xor (inputs(123));
    layer0_outputs(1445) <= not(inputs(62)) or (inputs(182));
    layer0_outputs(1446) <= (inputs(78)) or (inputs(40));
    layer0_outputs(1447) <= (inputs(35)) xor (inputs(50));
    layer0_outputs(1448) <= (inputs(27)) or (inputs(49));
    layer0_outputs(1449) <= (inputs(247)) or (inputs(47));
    layer0_outputs(1450) <= not(inputs(103));
    layer0_outputs(1451) <= inputs(76);
    layer0_outputs(1452) <= not((inputs(226)) or (inputs(128)));
    layer0_outputs(1453) <= not(inputs(174));
    layer0_outputs(1454) <= (inputs(111)) or (inputs(59));
    layer0_outputs(1455) <= not(inputs(204));
    layer0_outputs(1456) <= inputs(78);
    layer0_outputs(1457) <= not((inputs(130)) or (inputs(129)));
    layer0_outputs(1458) <= '0';
    layer0_outputs(1459) <= not(inputs(237));
    layer0_outputs(1460) <= not(inputs(179));
    layer0_outputs(1461) <= not((inputs(186)) or (inputs(94)));
    layer0_outputs(1462) <= not((inputs(214)) or (inputs(87)));
    layer0_outputs(1463) <= not(inputs(163));
    layer0_outputs(1464) <= not(inputs(193));
    layer0_outputs(1465) <= (inputs(219)) and not (inputs(83));
    layer0_outputs(1466) <= inputs(27);
    layer0_outputs(1467) <= not(inputs(232)) or (inputs(27));
    layer0_outputs(1468) <= not((inputs(3)) or (inputs(166)));
    layer0_outputs(1469) <= not(inputs(106)) or (inputs(32));
    layer0_outputs(1470) <= (inputs(86)) and not (inputs(127));
    layer0_outputs(1471) <= inputs(211);
    layer0_outputs(1472) <= not((inputs(158)) or (inputs(3)));
    layer0_outputs(1473) <= (inputs(87)) and not (inputs(145));
    layer0_outputs(1474) <= not(inputs(89));
    layer0_outputs(1475) <= inputs(70);
    layer0_outputs(1476) <= inputs(100);
    layer0_outputs(1477) <= not((inputs(173)) or (inputs(90)));
    layer0_outputs(1478) <= not(inputs(100));
    layer0_outputs(1479) <= not(inputs(202)) or (inputs(108));
    layer0_outputs(1480) <= (inputs(215)) and not (inputs(101));
    layer0_outputs(1481) <= (inputs(98)) and (inputs(240));
    layer0_outputs(1482) <= inputs(84);
    layer0_outputs(1483) <= (inputs(57)) and not (inputs(251));
    layer0_outputs(1484) <= inputs(8);
    layer0_outputs(1485) <= inputs(136);
    layer0_outputs(1486) <= not(inputs(242)) or (inputs(77));
    layer0_outputs(1487) <= (inputs(210)) or (inputs(187));
    layer0_outputs(1488) <= (inputs(26)) or (inputs(239));
    layer0_outputs(1489) <= not(inputs(108)) or (inputs(87));
    layer0_outputs(1490) <= not((inputs(111)) xor (inputs(234)));
    layer0_outputs(1491) <= inputs(19);
    layer0_outputs(1492) <= not(inputs(25));
    layer0_outputs(1493) <= not(inputs(150));
    layer0_outputs(1494) <= '0';
    layer0_outputs(1495) <= not(inputs(234));
    layer0_outputs(1496) <= not(inputs(97)) or (inputs(251));
    layer0_outputs(1497) <= '1';
    layer0_outputs(1498) <= inputs(148);
    layer0_outputs(1499) <= (inputs(15)) and not (inputs(163));
    layer0_outputs(1500) <= inputs(167);
    layer0_outputs(1501) <= (inputs(220)) or (inputs(211));
    layer0_outputs(1502) <= (inputs(116)) or (inputs(142));
    layer0_outputs(1503) <= not((inputs(25)) or (inputs(193)));
    layer0_outputs(1504) <= (inputs(248)) and not (inputs(58));
    layer0_outputs(1505) <= inputs(219);
    layer0_outputs(1506) <= '0';
    layer0_outputs(1507) <= not(inputs(90)) or (inputs(235));
    layer0_outputs(1508) <= not(inputs(152));
    layer0_outputs(1509) <= not(inputs(166)) or (inputs(30));
    layer0_outputs(1510) <= (inputs(154)) and not (inputs(9));
    layer0_outputs(1511) <= inputs(26);
    layer0_outputs(1512) <= not(inputs(56)) or (inputs(168));
    layer0_outputs(1513) <= inputs(32);
    layer0_outputs(1514) <= not(inputs(54));
    layer0_outputs(1515) <= (inputs(176)) or (inputs(208));
    layer0_outputs(1516) <= not(inputs(2));
    layer0_outputs(1517) <= inputs(84);
    layer0_outputs(1518) <= not(inputs(98)) or (inputs(227));
    layer0_outputs(1519) <= (inputs(83)) and not (inputs(1));
    layer0_outputs(1520) <= (inputs(125)) and not (inputs(2));
    layer0_outputs(1521) <= (inputs(76)) xor (inputs(14));
    layer0_outputs(1522) <= (inputs(132)) and (inputs(183));
    layer0_outputs(1523) <= (inputs(208)) and not (inputs(253));
    layer0_outputs(1524) <= not(inputs(114));
    layer0_outputs(1525) <= not((inputs(46)) and (inputs(184)));
    layer0_outputs(1526) <= '0';
    layer0_outputs(1527) <= inputs(46);
    layer0_outputs(1528) <= not((inputs(116)) xor (inputs(101)));
    layer0_outputs(1529) <= (inputs(99)) and not (inputs(4));
    layer0_outputs(1530) <= (inputs(246)) or (inputs(171));
    layer0_outputs(1531) <= (inputs(195)) and not (inputs(172));
    layer0_outputs(1532) <= not(inputs(182)) or (inputs(133));
    layer0_outputs(1533) <= not((inputs(127)) xor (inputs(155)));
    layer0_outputs(1534) <= not((inputs(53)) xor (inputs(160)));
    layer0_outputs(1535) <= not(inputs(22));
    layer0_outputs(1536) <= not((inputs(17)) or (inputs(207)));
    layer0_outputs(1537) <= inputs(251);
    layer0_outputs(1538) <= inputs(157);
    layer0_outputs(1539) <= inputs(223);
    layer0_outputs(1540) <= inputs(76);
    layer0_outputs(1541) <= inputs(200);
    layer0_outputs(1542) <= '1';
    layer0_outputs(1543) <= inputs(122);
    layer0_outputs(1544) <= inputs(198);
    layer0_outputs(1545) <= not(inputs(246));
    layer0_outputs(1546) <= not(inputs(106)) or (inputs(112));
    layer0_outputs(1547) <= '1';
    layer0_outputs(1548) <= not(inputs(124)) or (inputs(216));
    layer0_outputs(1549) <= not((inputs(165)) or (inputs(166)));
    layer0_outputs(1550) <= inputs(26);
    layer0_outputs(1551) <= not(inputs(195)) or (inputs(63));
    layer0_outputs(1552) <= '1';
    layer0_outputs(1553) <= (inputs(86)) or (inputs(72));
    layer0_outputs(1554) <= not((inputs(42)) or (inputs(160)));
    layer0_outputs(1555) <= not(inputs(112));
    layer0_outputs(1556) <= (inputs(205)) and not (inputs(94));
    layer0_outputs(1557) <= inputs(130);
    layer0_outputs(1558) <= not(inputs(125)) or (inputs(97));
    layer0_outputs(1559) <= (inputs(30)) and not (inputs(217));
    layer0_outputs(1560) <= (inputs(5)) and not (inputs(173));
    layer0_outputs(1561) <= not((inputs(53)) or (inputs(54)));
    layer0_outputs(1562) <= not((inputs(123)) xor (inputs(141)));
    layer0_outputs(1563) <= (inputs(74)) or (inputs(107));
    layer0_outputs(1564) <= inputs(107);
    layer0_outputs(1565) <= not(inputs(101));
    layer0_outputs(1566) <= not(inputs(89)) or (inputs(34));
    layer0_outputs(1567) <= (inputs(238)) and not (inputs(249));
    layer0_outputs(1568) <= not(inputs(169));
    layer0_outputs(1569) <= not((inputs(172)) or (inputs(252)));
    layer0_outputs(1570) <= not(inputs(174));
    layer0_outputs(1571) <= (inputs(140)) and (inputs(6));
    layer0_outputs(1572) <= not(inputs(188)) or (inputs(35));
    layer0_outputs(1573) <= not(inputs(210));
    layer0_outputs(1574) <= not((inputs(254)) or (inputs(76)));
    layer0_outputs(1575) <= inputs(99);
    layer0_outputs(1576) <= not(inputs(107));
    layer0_outputs(1577) <= (inputs(207)) or (inputs(45));
    layer0_outputs(1578) <= (inputs(195)) or (inputs(72));
    layer0_outputs(1579) <= '1';
    layer0_outputs(1580) <= (inputs(0)) xor (inputs(139));
    layer0_outputs(1581) <= not(inputs(241));
    layer0_outputs(1582) <= not((inputs(61)) or (inputs(95)));
    layer0_outputs(1583) <= not((inputs(86)) or (inputs(193)));
    layer0_outputs(1584) <= (inputs(103)) and not (inputs(148));
    layer0_outputs(1585) <= not(inputs(178)) or (inputs(240));
    layer0_outputs(1586) <= not(inputs(129));
    layer0_outputs(1587) <= not((inputs(64)) or (inputs(219)));
    layer0_outputs(1588) <= (inputs(65)) or (inputs(30));
    layer0_outputs(1589) <= not(inputs(248)) or (inputs(58));
    layer0_outputs(1590) <= not(inputs(104));
    layer0_outputs(1591) <= (inputs(145)) and not (inputs(181));
    layer0_outputs(1592) <= not(inputs(99)) or (inputs(223));
    layer0_outputs(1593) <= not((inputs(94)) xor (inputs(110)));
    layer0_outputs(1594) <= not((inputs(1)) and (inputs(23)));
    layer0_outputs(1595) <= not(inputs(38));
    layer0_outputs(1596) <= not(inputs(69)) or (inputs(94));
    layer0_outputs(1597) <= '1';
    layer0_outputs(1598) <= (inputs(140)) and not (inputs(60));
    layer0_outputs(1599) <= (inputs(165)) or (inputs(218));
    layer0_outputs(1600) <= not((inputs(89)) and (inputs(240)));
    layer0_outputs(1601) <= (inputs(128)) or (inputs(125));
    layer0_outputs(1602) <= (inputs(63)) or (inputs(23));
    layer0_outputs(1603) <= not((inputs(123)) or (inputs(113)));
    layer0_outputs(1604) <= not((inputs(238)) or (inputs(166)));
    layer0_outputs(1605) <= not(inputs(90)) or (inputs(181));
    layer0_outputs(1606) <= (inputs(151)) and not (inputs(111));
    layer0_outputs(1607) <= (inputs(12)) or (inputs(134));
    layer0_outputs(1608) <= not(inputs(10));
    layer0_outputs(1609) <= not(inputs(254));
    layer0_outputs(1610) <= not(inputs(84));
    layer0_outputs(1611) <= (inputs(212)) or (inputs(195));
    layer0_outputs(1612) <= inputs(131);
    layer0_outputs(1613) <= not(inputs(163));
    layer0_outputs(1614) <= not(inputs(109));
    layer0_outputs(1615) <= not((inputs(215)) and (inputs(218)));
    layer0_outputs(1616) <= (inputs(122)) and not (inputs(243));
    layer0_outputs(1617) <= '1';
    layer0_outputs(1618) <= '0';
    layer0_outputs(1619) <= '0';
    layer0_outputs(1620) <= (inputs(125)) and (inputs(117));
    layer0_outputs(1621) <= not((inputs(113)) and (inputs(150)));
    layer0_outputs(1622) <= not(inputs(58));
    layer0_outputs(1623) <= (inputs(56)) xor (inputs(26));
    layer0_outputs(1624) <= not(inputs(5)) or (inputs(161));
    layer0_outputs(1625) <= (inputs(103)) and not (inputs(170));
    layer0_outputs(1626) <= not((inputs(11)) or (inputs(131)));
    layer0_outputs(1627) <= not(inputs(122)) or (inputs(0));
    layer0_outputs(1628) <= not(inputs(85));
    layer0_outputs(1629) <= inputs(25);
    layer0_outputs(1630) <= (inputs(58)) or (inputs(166));
    layer0_outputs(1631) <= not((inputs(56)) or (inputs(67)));
    layer0_outputs(1632) <= inputs(241);
    layer0_outputs(1633) <= (inputs(125)) xor (inputs(239));
    layer0_outputs(1634) <= not((inputs(222)) or (inputs(152)));
    layer0_outputs(1635) <= not(inputs(85));
    layer0_outputs(1636) <= (inputs(84)) or (inputs(101));
    layer0_outputs(1637) <= inputs(121);
    layer0_outputs(1638) <= '0';
    layer0_outputs(1639) <= '0';
    layer0_outputs(1640) <= not((inputs(126)) and (inputs(24)));
    layer0_outputs(1641) <= (inputs(78)) and not (inputs(188));
    layer0_outputs(1642) <= (inputs(88)) and not (inputs(224));
    layer0_outputs(1643) <= '1';
    layer0_outputs(1644) <= not((inputs(108)) or (inputs(88)));
    layer0_outputs(1645) <= inputs(62);
    layer0_outputs(1646) <= not(inputs(11)) or (inputs(15));
    layer0_outputs(1647) <= inputs(82);
    layer0_outputs(1648) <= (inputs(78)) or (inputs(148));
    layer0_outputs(1649) <= inputs(53);
    layer0_outputs(1650) <= not(inputs(37));
    layer0_outputs(1651) <= (inputs(134)) and not (inputs(130));
    layer0_outputs(1652) <= not(inputs(119));
    layer0_outputs(1653) <= (inputs(34)) xor (inputs(179));
    layer0_outputs(1654) <= (inputs(108)) or (inputs(144));
    layer0_outputs(1655) <= not((inputs(64)) xor (inputs(168)));
    layer0_outputs(1656) <= not(inputs(39));
    layer0_outputs(1657) <= (inputs(76)) or (inputs(1));
    layer0_outputs(1658) <= inputs(117);
    layer0_outputs(1659) <= not(inputs(35));
    layer0_outputs(1660) <= (inputs(223)) and not (inputs(173));
    layer0_outputs(1661) <= not((inputs(249)) or (inputs(72)));
    layer0_outputs(1662) <= inputs(25);
    layer0_outputs(1663) <= not(inputs(150));
    layer0_outputs(1664) <= (inputs(61)) and not (inputs(235));
    layer0_outputs(1665) <= not(inputs(223));
    layer0_outputs(1666) <= '1';
    layer0_outputs(1667) <= not(inputs(26)) or (inputs(128));
    layer0_outputs(1668) <= '1';
    layer0_outputs(1669) <= not((inputs(79)) or (inputs(18)));
    layer0_outputs(1670) <= (inputs(195)) and not (inputs(16));
    layer0_outputs(1671) <= not(inputs(23));
    layer0_outputs(1672) <= not(inputs(144)) or (inputs(15));
    layer0_outputs(1673) <= (inputs(193)) and not (inputs(147));
    layer0_outputs(1674) <= inputs(94);
    layer0_outputs(1675) <= inputs(34);
    layer0_outputs(1676) <= '1';
    layer0_outputs(1677) <= not(inputs(34));
    layer0_outputs(1678) <= (inputs(99)) and not (inputs(148));
    layer0_outputs(1679) <= not((inputs(140)) or (inputs(194)));
    layer0_outputs(1680) <= not(inputs(31));
    layer0_outputs(1681) <= not(inputs(242));
    layer0_outputs(1682) <= '1';
    layer0_outputs(1683) <= not((inputs(168)) or (inputs(100)));
    layer0_outputs(1684) <= not((inputs(187)) or (inputs(193)));
    layer0_outputs(1685) <= not(inputs(72));
    layer0_outputs(1686) <= not(inputs(5));
    layer0_outputs(1687) <= (inputs(176)) or (inputs(186));
    layer0_outputs(1688) <= inputs(181);
    layer0_outputs(1689) <= not(inputs(11)) or (inputs(56));
    layer0_outputs(1690) <= '0';
    layer0_outputs(1691) <= not(inputs(218)) or (inputs(54));
    layer0_outputs(1692) <= not((inputs(219)) xor (inputs(150)));
    layer0_outputs(1693) <= not(inputs(32)) or (inputs(219));
    layer0_outputs(1694) <= (inputs(238)) and not (inputs(81));
    layer0_outputs(1695) <= not(inputs(232));
    layer0_outputs(1696) <= not((inputs(111)) or (inputs(245)));
    layer0_outputs(1697) <= (inputs(238)) and not (inputs(188));
    layer0_outputs(1698) <= not(inputs(163));
    layer0_outputs(1699) <= inputs(28);
    layer0_outputs(1700) <= (inputs(36)) and not (inputs(102));
    layer0_outputs(1701) <= not(inputs(231)) or (inputs(35));
    layer0_outputs(1702) <= not((inputs(63)) xor (inputs(4)));
    layer0_outputs(1703) <= (inputs(60)) and not (inputs(175));
    layer0_outputs(1704) <= not(inputs(134)) or (inputs(155));
    layer0_outputs(1705) <= inputs(91);
    layer0_outputs(1706) <= '0';
    layer0_outputs(1707) <= not(inputs(159));
    layer0_outputs(1708) <= not((inputs(195)) or (inputs(139)));
    layer0_outputs(1709) <= '0';
    layer0_outputs(1710) <= (inputs(207)) xor (inputs(95));
    layer0_outputs(1711) <= not(inputs(80));
    layer0_outputs(1712) <= (inputs(5)) and (inputs(30));
    layer0_outputs(1713) <= inputs(22);
    layer0_outputs(1714) <= not(inputs(54)) or (inputs(236));
    layer0_outputs(1715) <= not(inputs(117));
    layer0_outputs(1716) <= (inputs(160)) or (inputs(118));
    layer0_outputs(1717) <= (inputs(248)) xor (inputs(160));
    layer0_outputs(1718) <= '1';
    layer0_outputs(1719) <= inputs(8);
    layer0_outputs(1720) <= (inputs(157)) or (inputs(207));
    layer0_outputs(1721) <= not(inputs(123));
    layer0_outputs(1722) <= not((inputs(227)) or (inputs(46)));
    layer0_outputs(1723) <= not(inputs(121));
    layer0_outputs(1724) <= not((inputs(194)) or (inputs(218)));
    layer0_outputs(1725) <= inputs(161);
    layer0_outputs(1726) <= inputs(25);
    layer0_outputs(1727) <= not(inputs(193));
    layer0_outputs(1728) <= not(inputs(73));
    layer0_outputs(1729) <= (inputs(119)) or (inputs(47));
    layer0_outputs(1730) <= inputs(228);
    layer0_outputs(1731) <= not(inputs(42));
    layer0_outputs(1732) <= not(inputs(23)) or (inputs(211));
    layer0_outputs(1733) <= '0';
    layer0_outputs(1734) <= inputs(155);
    layer0_outputs(1735) <= (inputs(161)) and not (inputs(57));
    layer0_outputs(1736) <= '1';
    layer0_outputs(1737) <= not((inputs(188)) or (inputs(133)));
    layer0_outputs(1738) <= inputs(23);
    layer0_outputs(1739) <= not((inputs(162)) or (inputs(113)));
    layer0_outputs(1740) <= inputs(52);
    layer0_outputs(1741) <= (inputs(1)) or (inputs(50));
    layer0_outputs(1742) <= not(inputs(222));
    layer0_outputs(1743) <= (inputs(152)) and not (inputs(77));
    layer0_outputs(1744) <= (inputs(90)) and not (inputs(158));
    layer0_outputs(1745) <= not(inputs(195)) or (inputs(30));
    layer0_outputs(1746) <= not((inputs(91)) or (inputs(89)));
    layer0_outputs(1747) <= inputs(110);
    layer0_outputs(1748) <= '1';
    layer0_outputs(1749) <= (inputs(223)) or (inputs(164));
    layer0_outputs(1750) <= not((inputs(76)) or (inputs(126)));
    layer0_outputs(1751) <= (inputs(155)) and not (inputs(247));
    layer0_outputs(1752) <= inputs(168);
    layer0_outputs(1753) <= not((inputs(53)) and (inputs(104)));
    layer0_outputs(1754) <= not(inputs(247)) or (inputs(19));
    layer0_outputs(1755) <= (inputs(80)) xor (inputs(156));
    layer0_outputs(1756) <= inputs(47);
    layer0_outputs(1757) <= not(inputs(187));
    layer0_outputs(1758) <= (inputs(234)) and not (inputs(54));
    layer0_outputs(1759) <= not((inputs(63)) or (inputs(37)));
    layer0_outputs(1760) <= '0';
    layer0_outputs(1761) <= not((inputs(171)) xor (inputs(140)));
    layer0_outputs(1762) <= (inputs(116)) or (inputs(129));
    layer0_outputs(1763) <= inputs(228);
    layer0_outputs(1764) <= not(inputs(52)) or (inputs(20));
    layer0_outputs(1765) <= inputs(92);
    layer0_outputs(1766) <= (inputs(45)) and (inputs(108));
    layer0_outputs(1767) <= not(inputs(211));
    layer0_outputs(1768) <= '0';
    layer0_outputs(1769) <= not(inputs(127));
    layer0_outputs(1770) <= not(inputs(233)) or (inputs(120));
    layer0_outputs(1771) <= not(inputs(167));
    layer0_outputs(1772) <= not(inputs(117)) or (inputs(17));
    layer0_outputs(1773) <= inputs(85);
    layer0_outputs(1774) <= not((inputs(243)) or (inputs(21)));
    layer0_outputs(1775) <= not(inputs(100));
    layer0_outputs(1776) <= not(inputs(69)) or (inputs(182));
    layer0_outputs(1777) <= '0';
    layer0_outputs(1778) <= '1';
    layer0_outputs(1779) <= not((inputs(152)) xor (inputs(105)));
    layer0_outputs(1780) <= not(inputs(126)) or (inputs(227));
    layer0_outputs(1781) <= inputs(93);
    layer0_outputs(1782) <= not(inputs(135));
    layer0_outputs(1783) <= not((inputs(87)) or (inputs(91)));
    layer0_outputs(1784) <= (inputs(111)) or (inputs(53));
    layer0_outputs(1785) <= not(inputs(23));
    layer0_outputs(1786) <= (inputs(99)) or (inputs(169));
    layer0_outputs(1787) <= inputs(135);
    layer0_outputs(1788) <= (inputs(199)) and not (inputs(89));
    layer0_outputs(1789) <= not(inputs(255));
    layer0_outputs(1790) <= inputs(51);
    layer0_outputs(1791) <= not(inputs(207)) or (inputs(112));
    layer0_outputs(1792) <= not(inputs(183)) or (inputs(17));
    layer0_outputs(1793) <= (inputs(136)) xor (inputs(51));
    layer0_outputs(1794) <= (inputs(101)) xor (inputs(53));
    layer0_outputs(1795) <= not(inputs(179));
    layer0_outputs(1796) <= not(inputs(26));
    layer0_outputs(1797) <= not((inputs(109)) xor (inputs(190)));
    layer0_outputs(1798) <= (inputs(11)) and not (inputs(163));
    layer0_outputs(1799) <= '0';
    layer0_outputs(1800) <= inputs(213);
    layer0_outputs(1801) <= not(inputs(132));
    layer0_outputs(1802) <= (inputs(98)) or (inputs(138));
    layer0_outputs(1803) <= '0';
    layer0_outputs(1804) <= not(inputs(145));
    layer0_outputs(1805) <= not(inputs(187)) or (inputs(238));
    layer0_outputs(1806) <= (inputs(12)) and not (inputs(60));
    layer0_outputs(1807) <= (inputs(130)) and not (inputs(220));
    layer0_outputs(1808) <= not((inputs(71)) or (inputs(224)));
    layer0_outputs(1809) <= (inputs(218)) or (inputs(239));
    layer0_outputs(1810) <= not((inputs(35)) or (inputs(33)));
    layer0_outputs(1811) <= not((inputs(211)) and (inputs(7)));
    layer0_outputs(1812) <= not(inputs(42));
    layer0_outputs(1813) <= inputs(71);
    layer0_outputs(1814) <= not((inputs(172)) or (inputs(164)));
    layer0_outputs(1815) <= (inputs(220)) and not (inputs(119));
    layer0_outputs(1816) <= not(inputs(67));
    layer0_outputs(1817) <= '0';
    layer0_outputs(1818) <= inputs(70);
    layer0_outputs(1819) <= not(inputs(9));
    layer0_outputs(1820) <= not(inputs(101));
    layer0_outputs(1821) <= not((inputs(245)) and (inputs(27)));
    layer0_outputs(1822) <= '0';
    layer0_outputs(1823) <= not((inputs(125)) xor (inputs(159)));
    layer0_outputs(1824) <= (inputs(205)) xor (inputs(34));
    layer0_outputs(1825) <= not(inputs(124));
    layer0_outputs(1826) <= not(inputs(195));
    layer0_outputs(1827) <= not(inputs(91)) or (inputs(71));
    layer0_outputs(1828) <= not((inputs(222)) xor (inputs(222)));
    layer0_outputs(1829) <= (inputs(17)) xor (inputs(12));
    layer0_outputs(1830) <= not((inputs(49)) xor (inputs(95)));
    layer0_outputs(1831) <= not((inputs(67)) and (inputs(121)));
    layer0_outputs(1832) <= not(inputs(21)) or (inputs(146));
    layer0_outputs(1833) <= (inputs(72)) and (inputs(198));
    layer0_outputs(1834) <= '1';
    layer0_outputs(1835) <= inputs(94);
    layer0_outputs(1836) <= (inputs(130)) or (inputs(215));
    layer0_outputs(1837) <= not(inputs(166)) or (inputs(252));
    layer0_outputs(1838) <= not(inputs(84));
    layer0_outputs(1839) <= inputs(102);
    layer0_outputs(1840) <= not(inputs(254)) or (inputs(96));
    layer0_outputs(1841) <= not(inputs(27));
    layer0_outputs(1842) <= (inputs(215)) and (inputs(139));
    layer0_outputs(1843) <= not(inputs(201));
    layer0_outputs(1844) <= not((inputs(208)) or (inputs(118)));
    layer0_outputs(1845) <= (inputs(25)) xor (inputs(80));
    layer0_outputs(1846) <= inputs(239);
    layer0_outputs(1847) <= not((inputs(180)) xor (inputs(181)));
    layer0_outputs(1848) <= inputs(97);
    layer0_outputs(1849) <= (inputs(50)) and not (inputs(207));
    layer0_outputs(1850) <= inputs(39);
    layer0_outputs(1851) <= not(inputs(107)) or (inputs(117));
    layer0_outputs(1852) <= not(inputs(162)) or (inputs(0));
    layer0_outputs(1853) <= not(inputs(47));
    layer0_outputs(1854) <= not(inputs(95));
    layer0_outputs(1855) <= not(inputs(19));
    layer0_outputs(1856) <= '1';
    layer0_outputs(1857) <= inputs(102);
    layer0_outputs(1858) <= not((inputs(250)) or (inputs(234)));
    layer0_outputs(1859) <= (inputs(229)) and not (inputs(123));
    layer0_outputs(1860) <= not((inputs(181)) or (inputs(61)));
    layer0_outputs(1861) <= (inputs(157)) and not (inputs(65));
    layer0_outputs(1862) <= (inputs(106)) and not (inputs(112));
    layer0_outputs(1863) <= not((inputs(238)) xor (inputs(189)));
    layer0_outputs(1864) <= not(inputs(195)) or (inputs(51));
    layer0_outputs(1865) <= inputs(115);
    layer0_outputs(1866) <= (inputs(110)) and not (inputs(154));
    layer0_outputs(1867) <= inputs(102);
    layer0_outputs(1868) <= inputs(202);
    layer0_outputs(1869) <= (inputs(234)) or (inputs(179));
    layer0_outputs(1870) <= inputs(120);
    layer0_outputs(1871) <= not(inputs(31));
    layer0_outputs(1872) <= '0';
    layer0_outputs(1873) <= not(inputs(148));
    layer0_outputs(1874) <= '0';
    layer0_outputs(1875) <= (inputs(222)) xor (inputs(94));
    layer0_outputs(1876) <= not((inputs(115)) xor (inputs(72)));
    layer0_outputs(1877) <= not(inputs(74));
    layer0_outputs(1878) <= (inputs(215)) and (inputs(13));
    layer0_outputs(1879) <= inputs(140);
    layer0_outputs(1880) <= not(inputs(177)) or (inputs(231));
    layer0_outputs(1881) <= (inputs(240)) and (inputs(5));
    layer0_outputs(1882) <= inputs(180);
    layer0_outputs(1883) <= not(inputs(165));
    layer0_outputs(1884) <= not(inputs(254));
    layer0_outputs(1885) <= '1';
    layer0_outputs(1886) <= not(inputs(168));
    layer0_outputs(1887) <= not(inputs(175)) or (inputs(234));
    layer0_outputs(1888) <= (inputs(132)) and not (inputs(34));
    layer0_outputs(1889) <= not(inputs(184)) or (inputs(115));
    layer0_outputs(1890) <= not(inputs(134));
    layer0_outputs(1891) <= not((inputs(144)) or (inputs(253)));
    layer0_outputs(1892) <= inputs(230);
    layer0_outputs(1893) <= not(inputs(137)) or (inputs(57));
    layer0_outputs(1894) <= not((inputs(32)) or (inputs(181)));
    layer0_outputs(1895) <= inputs(99);
    layer0_outputs(1896) <= (inputs(106)) and not (inputs(51));
    layer0_outputs(1897) <= (inputs(255)) and (inputs(124));
    layer0_outputs(1898) <= (inputs(107)) and not (inputs(163));
    layer0_outputs(1899) <= not((inputs(141)) or (inputs(154)));
    layer0_outputs(1900) <= not(inputs(104));
    layer0_outputs(1901) <= (inputs(66)) and not (inputs(201));
    layer0_outputs(1902) <= not(inputs(212));
    layer0_outputs(1903) <= not(inputs(190));
    layer0_outputs(1904) <= not((inputs(173)) or (inputs(98)));
    layer0_outputs(1905) <= not(inputs(227)) or (inputs(112));
    layer0_outputs(1906) <= (inputs(72)) and not (inputs(33));
    layer0_outputs(1907) <= inputs(155);
    layer0_outputs(1908) <= (inputs(123)) and (inputs(238));
    layer0_outputs(1909) <= not((inputs(137)) xor (inputs(121)));
    layer0_outputs(1910) <= inputs(130);
    layer0_outputs(1911) <= (inputs(32)) or (inputs(23));
    layer0_outputs(1912) <= not(inputs(241));
    layer0_outputs(1913) <= inputs(173);
    layer0_outputs(1914) <= not((inputs(119)) and (inputs(247)));
    layer0_outputs(1915) <= not(inputs(132)) or (inputs(10));
    layer0_outputs(1916) <= not((inputs(37)) or (inputs(34)));
    layer0_outputs(1917) <= (inputs(221)) and not (inputs(186));
    layer0_outputs(1918) <= '1';
    layer0_outputs(1919) <= inputs(73);
    layer0_outputs(1920) <= not(inputs(116));
    layer0_outputs(1921) <= '1';
    layer0_outputs(1922) <= not(inputs(178)) or (inputs(76));
    layer0_outputs(1923) <= not(inputs(130));
    layer0_outputs(1924) <= not((inputs(74)) xor (inputs(255)));
    layer0_outputs(1925) <= not((inputs(30)) or (inputs(112)));
    layer0_outputs(1926) <= (inputs(32)) or (inputs(162));
    layer0_outputs(1927) <= not((inputs(161)) or (inputs(186)));
    layer0_outputs(1928) <= (inputs(16)) or (inputs(184));
    layer0_outputs(1929) <= (inputs(9)) and not (inputs(18));
    layer0_outputs(1930) <= not(inputs(227)) or (inputs(163));
    layer0_outputs(1931) <= not((inputs(211)) xor (inputs(164)));
    layer0_outputs(1932) <= inputs(66);
    layer0_outputs(1933) <= (inputs(221)) or (inputs(106));
    layer0_outputs(1934) <= not(inputs(29));
    layer0_outputs(1935) <= (inputs(168)) or (inputs(152));
    layer0_outputs(1936) <= not(inputs(112));
    layer0_outputs(1937) <= not(inputs(153));
    layer0_outputs(1938) <= (inputs(193)) or (inputs(30));
    layer0_outputs(1939) <= (inputs(229)) and not (inputs(33));
    layer0_outputs(1940) <= not((inputs(253)) xor (inputs(1)));
    layer0_outputs(1941) <= not(inputs(165));
    layer0_outputs(1942) <= '1';
    layer0_outputs(1943) <= not((inputs(252)) xor (inputs(237)));
    layer0_outputs(1944) <= (inputs(225)) or (inputs(202));
    layer0_outputs(1945) <= not((inputs(20)) xor (inputs(64)));
    layer0_outputs(1946) <= '1';
    layer0_outputs(1947) <= not(inputs(1)) or (inputs(209));
    layer0_outputs(1948) <= (inputs(103)) and not (inputs(13));
    layer0_outputs(1949) <= not((inputs(236)) xor (inputs(151)));
    layer0_outputs(1950) <= inputs(165);
    layer0_outputs(1951) <= inputs(118);
    layer0_outputs(1952) <= not((inputs(3)) or (inputs(9)));
    layer0_outputs(1953) <= (inputs(45)) and not (inputs(137));
    layer0_outputs(1954) <= (inputs(209)) or (inputs(231));
    layer0_outputs(1955) <= not(inputs(80)) or (inputs(51));
    layer0_outputs(1956) <= not(inputs(20)) or (inputs(134));
    layer0_outputs(1957) <= not(inputs(149));
    layer0_outputs(1958) <= not((inputs(231)) and (inputs(32)));
    layer0_outputs(1959) <= not(inputs(244));
    layer0_outputs(1960) <= not(inputs(79));
    layer0_outputs(1961) <= not((inputs(209)) or (inputs(89)));
    layer0_outputs(1962) <= (inputs(181)) xor (inputs(136));
    layer0_outputs(1963) <= not(inputs(44));
    layer0_outputs(1964) <= (inputs(211)) or (inputs(63));
    layer0_outputs(1965) <= inputs(182);
    layer0_outputs(1966) <= not(inputs(138)) or (inputs(199));
    layer0_outputs(1967) <= inputs(99);
    layer0_outputs(1968) <= not((inputs(249)) and (inputs(51)));
    layer0_outputs(1969) <= not(inputs(132));
    layer0_outputs(1970) <= not(inputs(167)) or (inputs(113));
    layer0_outputs(1971) <= (inputs(230)) and not (inputs(166));
    layer0_outputs(1972) <= '1';
    layer0_outputs(1973) <= (inputs(144)) or (inputs(66));
    layer0_outputs(1974) <= not(inputs(83));
    layer0_outputs(1975) <= '0';
    layer0_outputs(1976) <= not(inputs(41));
    layer0_outputs(1977) <= inputs(244);
    layer0_outputs(1978) <= inputs(104);
    layer0_outputs(1979) <= (inputs(51)) or (inputs(45));
    layer0_outputs(1980) <= (inputs(197)) and not (inputs(31));
    layer0_outputs(1981) <= '0';
    layer0_outputs(1982) <= inputs(252);
    layer0_outputs(1983) <= not(inputs(76)) or (inputs(213));
    layer0_outputs(1984) <= not(inputs(39));
    layer0_outputs(1985) <= not(inputs(212)) or (inputs(65));
    layer0_outputs(1986) <= not(inputs(21)) or (inputs(157));
    layer0_outputs(1987) <= not(inputs(148)) or (inputs(123));
    layer0_outputs(1988) <= not(inputs(89)) or (inputs(2));
    layer0_outputs(1989) <= '1';
    layer0_outputs(1990) <= (inputs(33)) or (inputs(212));
    layer0_outputs(1991) <= (inputs(93)) or (inputs(125));
    layer0_outputs(1992) <= (inputs(11)) or (inputs(77));
    layer0_outputs(1993) <= inputs(220);
    layer0_outputs(1994) <= not(inputs(52)) or (inputs(196));
    layer0_outputs(1995) <= not((inputs(71)) and (inputs(14)));
    layer0_outputs(1996) <= inputs(113);
    layer0_outputs(1997) <= (inputs(81)) or (inputs(195));
    layer0_outputs(1998) <= (inputs(75)) and not (inputs(154));
    layer0_outputs(1999) <= (inputs(63)) and (inputs(11));
    layer0_outputs(2000) <= inputs(246);
    layer0_outputs(2001) <= not((inputs(228)) or (inputs(176)));
    layer0_outputs(2002) <= inputs(86);
    layer0_outputs(2003) <= not((inputs(121)) xor (inputs(93)));
    layer0_outputs(2004) <= inputs(114);
    layer0_outputs(2005) <= not((inputs(187)) xor (inputs(63)));
    layer0_outputs(2006) <= (inputs(221)) and not (inputs(37));
    layer0_outputs(2007) <= (inputs(54)) and (inputs(134));
    layer0_outputs(2008) <= '0';
    layer0_outputs(2009) <= '1';
    layer0_outputs(2010) <= not(inputs(172));
    layer0_outputs(2011) <= (inputs(52)) or (inputs(36));
    layer0_outputs(2012) <= (inputs(219)) and not (inputs(68));
    layer0_outputs(2013) <= inputs(146);
    layer0_outputs(2014) <= not((inputs(191)) or (inputs(166)));
    layer0_outputs(2015) <= not((inputs(238)) or (inputs(24)));
    layer0_outputs(2016) <= '0';
    layer0_outputs(2017) <= (inputs(108)) and not (inputs(86));
    layer0_outputs(2018) <= (inputs(172)) xor (inputs(220));
    layer0_outputs(2019) <= not(inputs(31));
    layer0_outputs(2020) <= '0';
    layer0_outputs(2021) <= (inputs(9)) or (inputs(9));
    layer0_outputs(2022) <= not(inputs(231));
    layer0_outputs(2023) <= not((inputs(51)) or (inputs(83)));
    layer0_outputs(2024) <= (inputs(69)) and not (inputs(216));
    layer0_outputs(2025) <= not((inputs(124)) or (inputs(64)));
    layer0_outputs(2026) <= not(inputs(212)) or (inputs(39));
    layer0_outputs(2027) <= inputs(221);
    layer0_outputs(2028) <= (inputs(196)) or (inputs(0));
    layer0_outputs(2029) <= not(inputs(213));
    layer0_outputs(2030) <= (inputs(236)) xor (inputs(21));
    layer0_outputs(2031) <= (inputs(250)) and (inputs(46));
    layer0_outputs(2032) <= not((inputs(112)) or (inputs(147)));
    layer0_outputs(2033) <= (inputs(183)) and not (inputs(213));
    layer0_outputs(2034) <= (inputs(212)) or (inputs(164));
    layer0_outputs(2035) <= not(inputs(145));
    layer0_outputs(2036) <= inputs(217);
    layer0_outputs(2037) <= inputs(195);
    layer0_outputs(2038) <= (inputs(87)) and not (inputs(155));
    layer0_outputs(2039) <= not((inputs(254)) or (inputs(127)));
    layer0_outputs(2040) <= not((inputs(161)) or (inputs(186)));
    layer0_outputs(2041) <= not(inputs(174));
    layer0_outputs(2042) <= (inputs(27)) and not (inputs(148));
    layer0_outputs(2043) <= (inputs(172)) or (inputs(242));
    layer0_outputs(2044) <= not(inputs(130));
    layer0_outputs(2045) <= not(inputs(172)) or (inputs(145));
    layer0_outputs(2046) <= inputs(233);
    layer0_outputs(2047) <= not(inputs(90));
    layer0_outputs(2048) <= not(inputs(8));
    layer0_outputs(2049) <= not(inputs(235));
    layer0_outputs(2050) <= not((inputs(238)) or (inputs(212)));
    layer0_outputs(2051) <= (inputs(81)) xor (inputs(35));
    layer0_outputs(2052) <= (inputs(28)) and not (inputs(237));
    layer0_outputs(2053) <= not(inputs(170));
    layer0_outputs(2054) <= not(inputs(7));
    layer0_outputs(2055) <= not((inputs(192)) or (inputs(209)));
    layer0_outputs(2056) <= not((inputs(167)) and (inputs(121)));
    layer0_outputs(2057) <= not((inputs(1)) and (inputs(69)));
    layer0_outputs(2058) <= (inputs(179)) or (inputs(197));
    layer0_outputs(2059) <= not(inputs(9));
    layer0_outputs(2060) <= not(inputs(33)) or (inputs(178));
    layer0_outputs(2061) <= not((inputs(224)) or (inputs(187)));
    layer0_outputs(2062) <= inputs(16);
    layer0_outputs(2063) <= not(inputs(80));
    layer0_outputs(2064) <= not(inputs(162));
    layer0_outputs(2065) <= inputs(9);
    layer0_outputs(2066) <= '1';
    layer0_outputs(2067) <= (inputs(255)) or (inputs(97));
    layer0_outputs(2068) <= inputs(71);
    layer0_outputs(2069) <= inputs(212);
    layer0_outputs(2070) <= not(inputs(14)) or (inputs(118));
    layer0_outputs(2071) <= inputs(149);
    layer0_outputs(2072) <= inputs(90);
    layer0_outputs(2073) <= not(inputs(167));
    layer0_outputs(2074) <= not((inputs(43)) or (inputs(27)));
    layer0_outputs(2075) <= (inputs(116)) and not (inputs(221));
    layer0_outputs(2076) <= not(inputs(9)) or (inputs(230));
    layer0_outputs(2077) <= (inputs(28)) and not (inputs(111));
    layer0_outputs(2078) <= (inputs(177)) and not (inputs(168));
    layer0_outputs(2079) <= not((inputs(163)) xor (inputs(95)));
    layer0_outputs(2080) <= not((inputs(75)) or (inputs(3)));
    layer0_outputs(2081) <= (inputs(36)) or (inputs(155));
    layer0_outputs(2082) <= inputs(225);
    layer0_outputs(2083) <= not(inputs(15)) or (inputs(70));
    layer0_outputs(2084) <= inputs(104);
    layer0_outputs(2085) <= (inputs(191)) and (inputs(7));
    layer0_outputs(2086) <= not(inputs(134));
    layer0_outputs(2087) <= (inputs(72)) and not (inputs(228));
    layer0_outputs(2088) <= inputs(120);
    layer0_outputs(2089) <= inputs(19);
    layer0_outputs(2090) <= (inputs(17)) or (inputs(248));
    layer0_outputs(2091) <= '1';
    layer0_outputs(2092) <= not(inputs(235));
    layer0_outputs(2093) <= inputs(109);
    layer0_outputs(2094) <= not((inputs(114)) or (inputs(46)));
    layer0_outputs(2095) <= inputs(28);
    layer0_outputs(2096) <= (inputs(122)) xor (inputs(31));
    layer0_outputs(2097) <= (inputs(206)) or (inputs(189));
    layer0_outputs(2098) <= not(inputs(146)) or (inputs(58));
    layer0_outputs(2099) <= not(inputs(89)) or (inputs(210));
    layer0_outputs(2100) <= '0';
    layer0_outputs(2101) <= not((inputs(174)) or (inputs(147)));
    layer0_outputs(2102) <= inputs(55);
    layer0_outputs(2103) <= not(inputs(105));
    layer0_outputs(2104) <= (inputs(60)) and not (inputs(198));
    layer0_outputs(2105) <= (inputs(87)) and (inputs(75));
    layer0_outputs(2106) <= not(inputs(195));
    layer0_outputs(2107) <= not(inputs(75)) or (inputs(220));
    layer0_outputs(2108) <= '0';
    layer0_outputs(2109) <= not((inputs(28)) xor (inputs(45)));
    layer0_outputs(2110) <= (inputs(15)) and not (inputs(251));
    layer0_outputs(2111) <= inputs(137);
    layer0_outputs(2112) <= not(inputs(30));
    layer0_outputs(2113) <= inputs(125);
    layer0_outputs(2114) <= inputs(119);
    layer0_outputs(2115) <= not((inputs(123)) or (inputs(28)));
    layer0_outputs(2116) <= '1';
    layer0_outputs(2117) <= not((inputs(143)) or (inputs(211)));
    layer0_outputs(2118) <= (inputs(79)) or (inputs(158));
    layer0_outputs(2119) <= (inputs(6)) and not (inputs(26));
    layer0_outputs(2120) <= not(inputs(240));
    layer0_outputs(2121) <= (inputs(219)) and not (inputs(216));
    layer0_outputs(2122) <= not((inputs(68)) xor (inputs(128)));
    layer0_outputs(2123) <= not(inputs(169));
    layer0_outputs(2124) <= not(inputs(84)) or (inputs(159));
    layer0_outputs(2125) <= inputs(23);
    layer0_outputs(2126) <= inputs(101);
    layer0_outputs(2127) <= (inputs(46)) or (inputs(146));
    layer0_outputs(2128) <= (inputs(180)) or (inputs(234));
    layer0_outputs(2129) <= inputs(40);
    layer0_outputs(2130) <= not((inputs(95)) xor (inputs(175)));
    layer0_outputs(2131) <= (inputs(190)) and not (inputs(20));
    layer0_outputs(2132) <= (inputs(183)) and not (inputs(82));
    layer0_outputs(2133) <= '0';
    layer0_outputs(2134) <= inputs(23);
    layer0_outputs(2135) <= (inputs(147)) and not (inputs(115));
    layer0_outputs(2136) <= inputs(170);
    layer0_outputs(2137) <= inputs(58);
    layer0_outputs(2138) <= not(inputs(115));
    layer0_outputs(2139) <= (inputs(65)) or (inputs(131));
    layer0_outputs(2140) <= not(inputs(9));
    layer0_outputs(2141) <= not(inputs(89));
    layer0_outputs(2142) <= '0';
    layer0_outputs(2143) <= not(inputs(224));
    layer0_outputs(2144) <= not(inputs(142));
    layer0_outputs(2145) <= inputs(167);
    layer0_outputs(2146) <= not(inputs(164)) or (inputs(20));
    layer0_outputs(2147) <= (inputs(19)) and not (inputs(145));
    layer0_outputs(2148) <= not(inputs(42));
    layer0_outputs(2149) <= not(inputs(219)) or (inputs(67));
    layer0_outputs(2150) <= inputs(205);
    layer0_outputs(2151) <= not(inputs(84)) or (inputs(94));
    layer0_outputs(2152) <= inputs(21);
    layer0_outputs(2153) <= inputs(179);
    layer0_outputs(2154) <= not((inputs(238)) or (inputs(74)));
    layer0_outputs(2155) <= not(inputs(154)) or (inputs(50));
    layer0_outputs(2156) <= not(inputs(141));
    layer0_outputs(2157) <= not(inputs(133));
    layer0_outputs(2158) <= (inputs(240)) or (inputs(203));
    layer0_outputs(2159) <= (inputs(62)) and (inputs(205));
    layer0_outputs(2160) <= not(inputs(62));
    layer0_outputs(2161) <= (inputs(77)) and (inputs(114));
    layer0_outputs(2162) <= not(inputs(119)) or (inputs(238));
    layer0_outputs(2163) <= not(inputs(41));
    layer0_outputs(2164) <= not((inputs(43)) and (inputs(29)));
    layer0_outputs(2165) <= not((inputs(1)) xor (inputs(124)));
    layer0_outputs(2166) <= not(inputs(81));
    layer0_outputs(2167) <= (inputs(57)) or (inputs(235));
    layer0_outputs(2168) <= not(inputs(49)) or (inputs(212));
    layer0_outputs(2169) <= (inputs(18)) and (inputs(77));
    layer0_outputs(2170) <= inputs(56);
    layer0_outputs(2171) <= inputs(43);
    layer0_outputs(2172) <= not(inputs(213)) or (inputs(95));
    layer0_outputs(2173) <= '1';
    layer0_outputs(2174) <= (inputs(57)) or (inputs(43));
    layer0_outputs(2175) <= '1';
    layer0_outputs(2176) <= not(inputs(107)) or (inputs(151));
    layer0_outputs(2177) <= not(inputs(175));
    layer0_outputs(2178) <= not(inputs(164));
    layer0_outputs(2179) <= not((inputs(239)) or (inputs(194)));
    layer0_outputs(2180) <= (inputs(106)) and not (inputs(1));
    layer0_outputs(2181) <= (inputs(74)) and not (inputs(205));
    layer0_outputs(2182) <= (inputs(56)) and not (inputs(155));
    layer0_outputs(2183) <= not((inputs(172)) or (inputs(155)));
    layer0_outputs(2184) <= not((inputs(127)) and (inputs(154)));
    layer0_outputs(2185) <= inputs(249);
    layer0_outputs(2186) <= not(inputs(212));
    layer0_outputs(2187) <= (inputs(201)) or (inputs(244));
    layer0_outputs(2188) <= (inputs(188)) or (inputs(80));
    layer0_outputs(2189) <= not((inputs(78)) xor (inputs(206)));
    layer0_outputs(2190) <= inputs(115);
    layer0_outputs(2191) <= not(inputs(85));
    layer0_outputs(2192) <= inputs(115);
    layer0_outputs(2193) <= inputs(41);
    layer0_outputs(2194) <= '0';
    layer0_outputs(2195) <= not(inputs(232));
    layer0_outputs(2196) <= (inputs(135)) and not (inputs(58));
    layer0_outputs(2197) <= not(inputs(18));
    layer0_outputs(2198) <= (inputs(101)) and not (inputs(89));
    layer0_outputs(2199) <= inputs(40);
    layer0_outputs(2200) <= (inputs(135)) and not (inputs(220));
    layer0_outputs(2201) <= (inputs(236)) or (inputs(118));
    layer0_outputs(2202) <= inputs(71);
    layer0_outputs(2203) <= (inputs(122)) and not (inputs(5));
    layer0_outputs(2204) <= not((inputs(203)) and (inputs(61)));
    layer0_outputs(2205) <= not((inputs(105)) or (inputs(105)));
    layer0_outputs(2206) <= (inputs(212)) or (inputs(96));
    layer0_outputs(2207) <= not(inputs(120));
    layer0_outputs(2208) <= '0';
    layer0_outputs(2209) <= inputs(20);
    layer0_outputs(2210) <= not((inputs(110)) xor (inputs(66)));
    layer0_outputs(2211) <= not((inputs(197)) or (inputs(229)));
    layer0_outputs(2212) <= inputs(152);
    layer0_outputs(2213) <= inputs(28);
    layer0_outputs(2214) <= (inputs(137)) and not (inputs(96));
    layer0_outputs(2215) <= not(inputs(26)) or (inputs(112));
    layer0_outputs(2216) <= (inputs(57)) and not (inputs(200));
    layer0_outputs(2217) <= not(inputs(184));
    layer0_outputs(2218) <= (inputs(104)) or (inputs(152));
    layer0_outputs(2219) <= '1';
    layer0_outputs(2220) <= not((inputs(32)) or (inputs(2)));
    layer0_outputs(2221) <= not(inputs(141));
    layer0_outputs(2222) <= (inputs(203)) or (inputs(231));
    layer0_outputs(2223) <= not(inputs(164));
    layer0_outputs(2224) <= not(inputs(18));
    layer0_outputs(2225) <= (inputs(155)) and not (inputs(163));
    layer0_outputs(2226) <= not((inputs(244)) or (inputs(186)));
    layer0_outputs(2227) <= inputs(69);
    layer0_outputs(2228) <= not((inputs(69)) or (inputs(226)));
    layer0_outputs(2229) <= (inputs(107)) xor (inputs(1));
    layer0_outputs(2230) <= (inputs(111)) and not (inputs(40));
    layer0_outputs(2231) <= inputs(28);
    layer0_outputs(2232) <= not(inputs(232));
    layer0_outputs(2233) <= not(inputs(238)) or (inputs(253));
    layer0_outputs(2234) <= not(inputs(124)) or (inputs(228));
    layer0_outputs(2235) <= inputs(121);
    layer0_outputs(2236) <= inputs(40);
    layer0_outputs(2237) <= (inputs(203)) or (inputs(234));
    layer0_outputs(2238) <= (inputs(158)) and not (inputs(224));
    layer0_outputs(2239) <= (inputs(216)) and (inputs(211));
    layer0_outputs(2240) <= not(inputs(199)) or (inputs(63));
    layer0_outputs(2241) <= inputs(115);
    layer0_outputs(2242) <= (inputs(200)) xor (inputs(12));
    layer0_outputs(2243) <= inputs(21);
    layer0_outputs(2244) <= (inputs(49)) or (inputs(0));
    layer0_outputs(2245) <= not((inputs(106)) or (inputs(191)));
    layer0_outputs(2246) <= (inputs(13)) or (inputs(18));
    layer0_outputs(2247) <= inputs(84);
    layer0_outputs(2248) <= not(inputs(126)) or (inputs(17));
    layer0_outputs(2249) <= (inputs(83)) or (inputs(118));
    layer0_outputs(2250) <= not(inputs(152)) or (inputs(213));
    layer0_outputs(2251) <= '0';
    layer0_outputs(2252) <= not(inputs(179));
    layer0_outputs(2253) <= not((inputs(249)) xor (inputs(6)));
    layer0_outputs(2254) <= (inputs(220)) xor (inputs(177));
    layer0_outputs(2255) <= (inputs(186)) or (inputs(118));
    layer0_outputs(2256) <= not((inputs(1)) or (inputs(76)));
    layer0_outputs(2257) <= not((inputs(150)) or (inputs(105)));
    layer0_outputs(2258) <= not((inputs(209)) xor (inputs(5)));
    layer0_outputs(2259) <= (inputs(171)) or (inputs(20));
    layer0_outputs(2260) <= not(inputs(72)) or (inputs(31));
    layer0_outputs(2261) <= inputs(190);
    layer0_outputs(2262) <= not(inputs(96));
    layer0_outputs(2263) <= inputs(88);
    layer0_outputs(2264) <= (inputs(136)) and (inputs(241));
    layer0_outputs(2265) <= not(inputs(82));
    layer0_outputs(2266) <= inputs(153);
    layer0_outputs(2267) <= inputs(53);
    layer0_outputs(2268) <= '0';
    layer0_outputs(2269) <= not(inputs(194));
    layer0_outputs(2270) <= (inputs(204)) and not (inputs(31));
    layer0_outputs(2271) <= not(inputs(199));
    layer0_outputs(2272) <= (inputs(206)) and (inputs(14));
    layer0_outputs(2273) <= not(inputs(142)) or (inputs(12));
    layer0_outputs(2274) <= not(inputs(230));
    layer0_outputs(2275) <= inputs(131);
    layer0_outputs(2276) <= (inputs(170)) and not (inputs(250));
    layer0_outputs(2277) <= not(inputs(210));
    layer0_outputs(2278) <= (inputs(91)) and not (inputs(223));
    layer0_outputs(2279) <= not((inputs(82)) xor (inputs(102)));
    layer0_outputs(2280) <= not(inputs(89)) or (inputs(128));
    layer0_outputs(2281) <= not(inputs(37)) or (inputs(192));
    layer0_outputs(2282) <= not(inputs(160));
    layer0_outputs(2283) <= inputs(132);
    layer0_outputs(2284) <= not((inputs(172)) and (inputs(209)));
    layer0_outputs(2285) <= not(inputs(150)) or (inputs(127));
    layer0_outputs(2286) <= '0';
    layer0_outputs(2287) <= (inputs(132)) xor (inputs(190));
    layer0_outputs(2288) <= not(inputs(245)) or (inputs(72));
    layer0_outputs(2289) <= not((inputs(35)) or (inputs(64)));
    layer0_outputs(2290) <= not(inputs(222));
    layer0_outputs(2291) <= not((inputs(126)) or (inputs(21)));
    layer0_outputs(2292) <= not((inputs(254)) or (inputs(65)));
    layer0_outputs(2293) <= not((inputs(245)) and (inputs(132)));
    layer0_outputs(2294) <= not((inputs(157)) or (inputs(130)));
    layer0_outputs(2295) <= not(inputs(137));
    layer0_outputs(2296) <= inputs(104);
    layer0_outputs(2297) <= (inputs(103)) and not (inputs(65));
    layer0_outputs(2298) <= not(inputs(195));
    layer0_outputs(2299) <= (inputs(195)) xor (inputs(195));
    layer0_outputs(2300) <= (inputs(161)) and not (inputs(205));
    layer0_outputs(2301) <= not((inputs(18)) xor (inputs(56)));
    layer0_outputs(2302) <= '1';
    layer0_outputs(2303) <= not(inputs(26)) or (inputs(16));
    layer0_outputs(2304) <= (inputs(128)) or (inputs(197));
    layer0_outputs(2305) <= not(inputs(149));
    layer0_outputs(2306) <= inputs(104);
    layer0_outputs(2307) <= '0';
    layer0_outputs(2308) <= not((inputs(115)) or (inputs(171)));
    layer0_outputs(2309) <= not(inputs(54));
    layer0_outputs(2310) <= (inputs(106)) and (inputs(124));
    layer0_outputs(2311) <= not((inputs(170)) or (inputs(243)));
    layer0_outputs(2312) <= '0';
    layer0_outputs(2313) <= '1';
    layer0_outputs(2314) <= (inputs(174)) or (inputs(11));
    layer0_outputs(2315) <= not((inputs(232)) xor (inputs(204)));
    layer0_outputs(2316) <= inputs(247);
    layer0_outputs(2317) <= (inputs(153)) or (inputs(105));
    layer0_outputs(2318) <= inputs(62);
    layer0_outputs(2319) <= not(inputs(156)) or (inputs(167));
    layer0_outputs(2320) <= inputs(85);
    layer0_outputs(2321) <= inputs(95);
    layer0_outputs(2322) <= '0';
    layer0_outputs(2323) <= (inputs(26)) or (inputs(238));
    layer0_outputs(2324) <= not((inputs(140)) or (inputs(114)));
    layer0_outputs(2325) <= (inputs(249)) or (inputs(247));
    layer0_outputs(2326) <= (inputs(220)) xor (inputs(253));
    layer0_outputs(2327) <= (inputs(200)) or (inputs(35));
    layer0_outputs(2328) <= not(inputs(134));
    layer0_outputs(2329) <= not(inputs(130));
    layer0_outputs(2330) <= not(inputs(236)) or (inputs(95));
    layer0_outputs(2331) <= not(inputs(212));
    layer0_outputs(2332) <= not(inputs(107));
    layer0_outputs(2333) <= inputs(253);
    layer0_outputs(2334) <= not(inputs(123));
    layer0_outputs(2335) <= not((inputs(62)) or (inputs(79)));
    layer0_outputs(2336) <= (inputs(104)) and not (inputs(53));
    layer0_outputs(2337) <= not(inputs(46)) or (inputs(70));
    layer0_outputs(2338) <= not(inputs(210)) or (inputs(249));
    layer0_outputs(2339) <= inputs(49);
    layer0_outputs(2340) <= inputs(76);
    layer0_outputs(2341) <= not(inputs(2)) or (inputs(112));
    layer0_outputs(2342) <= not(inputs(116));
    layer0_outputs(2343) <= (inputs(12)) and (inputs(173));
    layer0_outputs(2344) <= not((inputs(64)) or (inputs(135)));
    layer0_outputs(2345) <= not(inputs(219));
    layer0_outputs(2346) <= not(inputs(21));
    layer0_outputs(2347) <= inputs(48);
    layer0_outputs(2348) <= inputs(156);
    layer0_outputs(2349) <= inputs(177);
    layer0_outputs(2350) <= (inputs(69)) or (inputs(64));
    layer0_outputs(2351) <= not(inputs(8));
    layer0_outputs(2352) <= '1';
    layer0_outputs(2353) <= not((inputs(54)) and (inputs(92)));
    layer0_outputs(2354) <= not(inputs(83)) or (inputs(6));
    layer0_outputs(2355) <= (inputs(219)) and not (inputs(223));
    layer0_outputs(2356) <= inputs(174);
    layer0_outputs(2357) <= not(inputs(58)) or (inputs(196));
    layer0_outputs(2358) <= not((inputs(163)) and (inputs(87)));
    layer0_outputs(2359) <= not(inputs(117)) or (inputs(2));
    layer0_outputs(2360) <= (inputs(127)) or (inputs(147));
    layer0_outputs(2361) <= (inputs(249)) or (inputs(130));
    layer0_outputs(2362) <= not((inputs(133)) xor (inputs(194)));
    layer0_outputs(2363) <= not(inputs(42));
    layer0_outputs(2364) <= not(inputs(81)) or (inputs(53));
    layer0_outputs(2365) <= not(inputs(106));
    layer0_outputs(2366) <= not(inputs(182));
    layer0_outputs(2367) <= not(inputs(119)) or (inputs(144));
    layer0_outputs(2368) <= not(inputs(24)) or (inputs(97));
    layer0_outputs(2369) <= not(inputs(247));
    layer0_outputs(2370) <= (inputs(23)) xor (inputs(26));
    layer0_outputs(2371) <= not(inputs(79));
    layer0_outputs(2372) <= not(inputs(98)) or (inputs(110));
    layer0_outputs(2373) <= not((inputs(123)) or (inputs(93)));
    layer0_outputs(2374) <= not(inputs(68));
    layer0_outputs(2375) <= not(inputs(221));
    layer0_outputs(2376) <= inputs(232);
    layer0_outputs(2377) <= not(inputs(14));
    layer0_outputs(2378) <= not(inputs(170));
    layer0_outputs(2379) <= not((inputs(240)) and (inputs(229)));
    layer0_outputs(2380) <= not((inputs(93)) or (inputs(2)));
    layer0_outputs(2381) <= not(inputs(11));
    layer0_outputs(2382) <= (inputs(84)) and not (inputs(142));
    layer0_outputs(2383) <= not((inputs(6)) and (inputs(235)));
    layer0_outputs(2384) <= not(inputs(130));
    layer0_outputs(2385) <= not(inputs(51)) or (inputs(47));
    layer0_outputs(2386) <= inputs(170);
    layer0_outputs(2387) <= not(inputs(50));
    layer0_outputs(2388) <= not((inputs(240)) and (inputs(46)));
    layer0_outputs(2389) <= (inputs(39)) xor (inputs(30));
    layer0_outputs(2390) <= not((inputs(10)) and (inputs(114)));
    layer0_outputs(2391) <= not((inputs(139)) or (inputs(201)));
    layer0_outputs(2392) <= '0';
    layer0_outputs(2393) <= inputs(181);
    layer0_outputs(2394) <= inputs(120);
    layer0_outputs(2395) <= '1';
    layer0_outputs(2396) <= (inputs(156)) xor (inputs(206));
    layer0_outputs(2397) <= inputs(136);
    layer0_outputs(2398) <= not((inputs(42)) and (inputs(29)));
    layer0_outputs(2399) <= not((inputs(213)) or (inputs(38)));
    layer0_outputs(2400) <= inputs(139);
    layer0_outputs(2401) <= not(inputs(177));
    layer0_outputs(2402) <= not(inputs(235)) or (inputs(58));
    layer0_outputs(2403) <= not(inputs(104));
    layer0_outputs(2404) <= (inputs(67)) and not (inputs(30));
    layer0_outputs(2405) <= not(inputs(55)) or (inputs(14));
    layer0_outputs(2406) <= '1';
    layer0_outputs(2407) <= not((inputs(143)) or (inputs(214)));
    layer0_outputs(2408) <= not(inputs(68));
    layer0_outputs(2409) <= not(inputs(234));
    layer0_outputs(2410) <= '0';
    layer0_outputs(2411) <= (inputs(234)) or (inputs(97));
    layer0_outputs(2412) <= (inputs(157)) and (inputs(120));
    layer0_outputs(2413) <= not((inputs(50)) or (inputs(149)));
    layer0_outputs(2414) <= not(inputs(11)) or (inputs(83));
    layer0_outputs(2415) <= inputs(199);
    layer0_outputs(2416) <= not(inputs(228));
    layer0_outputs(2417) <= not((inputs(204)) or (inputs(10)));
    layer0_outputs(2418) <= not(inputs(128));
    layer0_outputs(2419) <= inputs(203);
    layer0_outputs(2420) <= (inputs(116)) or (inputs(113));
    layer0_outputs(2421) <= (inputs(77)) or (inputs(76));
    layer0_outputs(2422) <= inputs(146);
    layer0_outputs(2423) <= not(inputs(108)) or (inputs(207));
    layer0_outputs(2424) <= not(inputs(7));
    layer0_outputs(2425) <= not((inputs(173)) or (inputs(7)));
    layer0_outputs(2426) <= not(inputs(158));
    layer0_outputs(2427) <= not(inputs(235));
    layer0_outputs(2428) <= inputs(87);
    layer0_outputs(2429) <= not((inputs(89)) and (inputs(255)));
    layer0_outputs(2430) <= inputs(40);
    layer0_outputs(2431) <= inputs(176);
    layer0_outputs(2432) <= (inputs(202)) xor (inputs(178));
    layer0_outputs(2433) <= not((inputs(40)) or (inputs(193)));
    layer0_outputs(2434) <= inputs(104);
    layer0_outputs(2435) <= '1';
    layer0_outputs(2436) <= (inputs(68)) and not (inputs(140));
    layer0_outputs(2437) <= (inputs(199)) or (inputs(197));
    layer0_outputs(2438) <= inputs(115);
    layer0_outputs(2439) <= (inputs(192)) or (inputs(227));
    layer0_outputs(2440) <= (inputs(237)) xor (inputs(173));
    layer0_outputs(2441) <= not(inputs(156));
    layer0_outputs(2442) <= inputs(72);
    layer0_outputs(2443) <= not(inputs(5)) or (inputs(78));
    layer0_outputs(2444) <= not(inputs(178)) or (inputs(30));
    layer0_outputs(2445) <= not(inputs(53)) or (inputs(73));
    layer0_outputs(2446) <= not(inputs(189)) or (inputs(52));
    layer0_outputs(2447) <= (inputs(243)) or (inputs(231));
    layer0_outputs(2448) <= not(inputs(130));
    layer0_outputs(2449) <= not(inputs(230));
    layer0_outputs(2450) <= not((inputs(237)) or (inputs(234)));
    layer0_outputs(2451) <= (inputs(194)) or (inputs(191));
    layer0_outputs(2452) <= inputs(9);
    layer0_outputs(2453) <= not(inputs(84));
    layer0_outputs(2454) <= (inputs(231)) and (inputs(226));
    layer0_outputs(2455) <= not(inputs(80)) or (inputs(169));
    layer0_outputs(2456) <= '1';
    layer0_outputs(2457) <= not(inputs(138)) or (inputs(189));
    layer0_outputs(2458) <= (inputs(244)) and not (inputs(51));
    layer0_outputs(2459) <= (inputs(19)) or (inputs(148));
    layer0_outputs(2460) <= not(inputs(202));
    layer0_outputs(2461) <= (inputs(232)) and not (inputs(19));
    layer0_outputs(2462) <= (inputs(56)) and not (inputs(74));
    layer0_outputs(2463) <= not(inputs(128));
    layer0_outputs(2464) <= inputs(53);
    layer0_outputs(2465) <= not(inputs(9));
    layer0_outputs(2466) <= inputs(90);
    layer0_outputs(2467) <= inputs(132);
    layer0_outputs(2468) <= (inputs(43)) and not (inputs(254));
    layer0_outputs(2469) <= not(inputs(118)) or (inputs(174));
    layer0_outputs(2470) <= '0';
    layer0_outputs(2471) <= not((inputs(67)) or (inputs(47)));
    layer0_outputs(2472) <= not((inputs(145)) or (inputs(167)));
    layer0_outputs(2473) <= '1';
    layer0_outputs(2474) <= inputs(39);
    layer0_outputs(2475) <= not(inputs(119));
    layer0_outputs(2476) <= not((inputs(180)) or (inputs(163)));
    layer0_outputs(2477) <= (inputs(80)) and not (inputs(93));
    layer0_outputs(2478) <= '0';
    layer0_outputs(2479) <= '1';
    layer0_outputs(2480) <= not(inputs(194)) or (inputs(34));
    layer0_outputs(2481) <= (inputs(141)) and (inputs(37));
    layer0_outputs(2482) <= not(inputs(150)) or (inputs(137));
    layer0_outputs(2483) <= inputs(74);
    layer0_outputs(2484) <= (inputs(124)) and not (inputs(23));
    layer0_outputs(2485) <= inputs(203);
    layer0_outputs(2486) <= not(inputs(49)) or (inputs(210));
    layer0_outputs(2487) <= not(inputs(29));
    layer0_outputs(2488) <= not((inputs(223)) or (inputs(95)));
    layer0_outputs(2489) <= (inputs(123)) and not (inputs(161));
    layer0_outputs(2490) <= inputs(216);
    layer0_outputs(2491) <= inputs(73);
    layer0_outputs(2492) <= not(inputs(67));
    layer0_outputs(2493) <= not(inputs(242)) or (inputs(129));
    layer0_outputs(2494) <= (inputs(6)) or (inputs(32));
    layer0_outputs(2495) <= not(inputs(200));
    layer0_outputs(2496) <= inputs(70);
    layer0_outputs(2497) <= not((inputs(179)) or (inputs(5)));
    layer0_outputs(2498) <= '1';
    layer0_outputs(2499) <= not(inputs(101));
    layer0_outputs(2500) <= (inputs(53)) xor (inputs(184));
    layer0_outputs(2501) <= (inputs(186)) and not (inputs(78));
    layer0_outputs(2502) <= (inputs(229)) or (inputs(159));
    layer0_outputs(2503) <= not(inputs(87)) or (inputs(127));
    layer0_outputs(2504) <= (inputs(79)) and not (inputs(33));
    layer0_outputs(2505) <= inputs(10);
    layer0_outputs(2506) <= not((inputs(25)) or (inputs(36)));
    layer0_outputs(2507) <= not(inputs(228));
    layer0_outputs(2508) <= '1';
    layer0_outputs(2509) <= not(inputs(116)) or (inputs(237));
    layer0_outputs(2510) <= not(inputs(242));
    layer0_outputs(2511) <= (inputs(190)) and not (inputs(232));
    layer0_outputs(2512) <= not(inputs(162));
    layer0_outputs(2513) <= not(inputs(115)) or (inputs(255));
    layer0_outputs(2514) <= not(inputs(51));
    layer0_outputs(2515) <= (inputs(154)) and not (inputs(210));
    layer0_outputs(2516) <= not(inputs(134)) or (inputs(242));
    layer0_outputs(2517) <= not((inputs(166)) xor (inputs(212)));
    layer0_outputs(2518) <= not((inputs(61)) or (inputs(94)));
    layer0_outputs(2519) <= not(inputs(83));
    layer0_outputs(2520) <= (inputs(176)) xor (inputs(12));
    layer0_outputs(2521) <= inputs(144);
    layer0_outputs(2522) <= '0';
    layer0_outputs(2523) <= not(inputs(133));
    layer0_outputs(2524) <= (inputs(74)) and not (inputs(112));
    layer0_outputs(2525) <= inputs(206);
    layer0_outputs(2526) <= inputs(178);
    layer0_outputs(2527) <= not((inputs(141)) and (inputs(188)));
    layer0_outputs(2528) <= (inputs(103)) or (inputs(174));
    layer0_outputs(2529) <= '1';
    layer0_outputs(2530) <= not(inputs(232));
    layer0_outputs(2531) <= inputs(236);
    layer0_outputs(2532) <= (inputs(140)) and not (inputs(201));
    layer0_outputs(2533) <= not(inputs(87));
    layer0_outputs(2534) <= not(inputs(57));
    layer0_outputs(2535) <= (inputs(10)) and not (inputs(125));
    layer0_outputs(2536) <= inputs(67);
    layer0_outputs(2537) <= not(inputs(35));
    layer0_outputs(2538) <= not(inputs(249));
    layer0_outputs(2539) <= inputs(209);
    layer0_outputs(2540) <= not(inputs(188));
    layer0_outputs(2541) <= not(inputs(110));
    layer0_outputs(2542) <= (inputs(72)) and not (inputs(142));
    layer0_outputs(2543) <= inputs(50);
    layer0_outputs(2544) <= not((inputs(180)) or (inputs(232)));
    layer0_outputs(2545) <= inputs(218);
    layer0_outputs(2546) <= (inputs(42)) and (inputs(247));
    layer0_outputs(2547) <= not(inputs(177));
    layer0_outputs(2548) <= inputs(10);
    layer0_outputs(2549) <= (inputs(222)) or (inputs(169));
    layer0_outputs(2550) <= not(inputs(181)) or (inputs(32));
    layer0_outputs(2551) <= (inputs(196)) or (inputs(129));
    layer0_outputs(2552) <= not(inputs(103));
    layer0_outputs(2553) <= (inputs(142)) or (inputs(113));
    layer0_outputs(2554) <= inputs(41);
    layer0_outputs(2555) <= inputs(131);
    layer0_outputs(2556) <= (inputs(172)) and not (inputs(240));
    layer0_outputs(2557) <= '1';
    layer0_outputs(2558) <= inputs(68);
    layer0_outputs(2559) <= (inputs(215)) or (inputs(1));
    layer0_outputs(2560) <= not(inputs(166));
    layer0_outputs(2561) <= not(inputs(179)) or (inputs(63));
    layer0_outputs(2562) <= inputs(137);
    layer0_outputs(2563) <= not(inputs(99));
    layer0_outputs(2564) <= not(inputs(226));
    layer0_outputs(2565) <= inputs(117);
    layer0_outputs(2566) <= '0';
    layer0_outputs(2567) <= not((inputs(241)) or (inputs(14)));
    layer0_outputs(2568) <= not(inputs(25));
    layer0_outputs(2569) <= not(inputs(240));
    layer0_outputs(2570) <= inputs(41);
    layer0_outputs(2571) <= not((inputs(14)) and (inputs(66)));
    layer0_outputs(2572) <= not(inputs(179));
    layer0_outputs(2573) <= (inputs(188)) or (inputs(32));
    layer0_outputs(2574) <= not(inputs(75)) or (inputs(242));
    layer0_outputs(2575) <= not(inputs(113));
    layer0_outputs(2576) <= not(inputs(39));
    layer0_outputs(2577) <= '0';
    layer0_outputs(2578) <= not(inputs(155)) or (inputs(61));
    layer0_outputs(2579) <= not(inputs(156)) or (inputs(222));
    layer0_outputs(2580) <= (inputs(136)) xor (inputs(106));
    layer0_outputs(2581) <= '1';
    layer0_outputs(2582) <= not(inputs(62));
    layer0_outputs(2583) <= (inputs(253)) or (inputs(90));
    layer0_outputs(2584) <= (inputs(58)) and not (inputs(13));
    layer0_outputs(2585) <= not(inputs(210));
    layer0_outputs(2586) <= not(inputs(117)) or (inputs(105));
    layer0_outputs(2587) <= not((inputs(207)) xor (inputs(178)));
    layer0_outputs(2588) <= not(inputs(71));
    layer0_outputs(2589) <= not(inputs(132));
    layer0_outputs(2590) <= not(inputs(69));
    layer0_outputs(2591) <= (inputs(37)) and (inputs(32));
    layer0_outputs(2592) <= (inputs(169)) and not (inputs(80));
    layer0_outputs(2593) <= inputs(209);
    layer0_outputs(2594) <= (inputs(146)) and not (inputs(242));
    layer0_outputs(2595) <= inputs(106);
    layer0_outputs(2596) <= (inputs(90)) and (inputs(157));
    layer0_outputs(2597) <= inputs(142);
    layer0_outputs(2598) <= (inputs(194)) or (inputs(50));
    layer0_outputs(2599) <= not(inputs(59));
    layer0_outputs(2600) <= not(inputs(249)) or (inputs(214));
    layer0_outputs(2601) <= '0';
    layer0_outputs(2602) <= (inputs(111)) and not (inputs(33));
    layer0_outputs(2603) <= not(inputs(45));
    layer0_outputs(2604) <= '1';
    layer0_outputs(2605) <= '0';
    layer0_outputs(2606) <= not((inputs(213)) and (inputs(164)));
    layer0_outputs(2607) <= (inputs(248)) or (inputs(193));
    layer0_outputs(2608) <= '1';
    layer0_outputs(2609) <= (inputs(56)) and not (inputs(81));
    layer0_outputs(2610) <= not((inputs(66)) xor (inputs(84)));
    layer0_outputs(2611) <= not((inputs(39)) or (inputs(214)));
    layer0_outputs(2612) <= (inputs(195)) and not (inputs(32));
    layer0_outputs(2613) <= not(inputs(219));
    layer0_outputs(2614) <= not(inputs(148));
    layer0_outputs(2615) <= inputs(167);
    layer0_outputs(2616) <= inputs(249);
    layer0_outputs(2617) <= '1';
    layer0_outputs(2618) <= not(inputs(90)) or (inputs(81));
    layer0_outputs(2619) <= inputs(111);
    layer0_outputs(2620) <= not((inputs(4)) or (inputs(41)));
    layer0_outputs(2621) <= (inputs(214)) and not (inputs(105));
    layer0_outputs(2622) <= not(inputs(79));
    layer0_outputs(2623) <= not((inputs(207)) or (inputs(215)));
    layer0_outputs(2624) <= not(inputs(46)) or (inputs(192));
    layer0_outputs(2625) <= (inputs(191)) or (inputs(209));
    layer0_outputs(2626) <= not(inputs(249));
    layer0_outputs(2627) <= not(inputs(185));
    layer0_outputs(2628) <= not((inputs(159)) xor (inputs(92)));
    layer0_outputs(2629) <= (inputs(7)) or (inputs(228));
    layer0_outputs(2630) <= not(inputs(109));
    layer0_outputs(2631) <= not((inputs(58)) or (inputs(136)));
    layer0_outputs(2632) <= (inputs(201)) xor (inputs(52));
    layer0_outputs(2633) <= not(inputs(157));
    layer0_outputs(2634) <= '0';
    layer0_outputs(2635) <= '1';
    layer0_outputs(2636) <= not((inputs(40)) or (inputs(191)));
    layer0_outputs(2637) <= inputs(220);
    layer0_outputs(2638) <= (inputs(78)) or (inputs(107));
    layer0_outputs(2639) <= (inputs(232)) and (inputs(76));
    layer0_outputs(2640) <= (inputs(104)) or (inputs(151));
    layer0_outputs(2641) <= inputs(9);
    layer0_outputs(2642) <= not((inputs(238)) or (inputs(9)));
    layer0_outputs(2643) <= (inputs(115)) xor (inputs(209));
    layer0_outputs(2644) <= not(inputs(195)) or (inputs(65));
    layer0_outputs(2645) <= not((inputs(110)) or (inputs(125)));
    layer0_outputs(2646) <= inputs(34);
    layer0_outputs(2647) <= (inputs(248)) xor (inputs(54));
    layer0_outputs(2648) <= inputs(106);
    layer0_outputs(2649) <= not(inputs(81));
    layer0_outputs(2650) <= not(inputs(165));
    layer0_outputs(2651) <= inputs(229);
    layer0_outputs(2652) <= not(inputs(87));
    layer0_outputs(2653) <= inputs(232);
    layer0_outputs(2654) <= not(inputs(6));
    layer0_outputs(2655) <= (inputs(224)) and (inputs(154));
    layer0_outputs(2656) <= not(inputs(242));
    layer0_outputs(2657) <= not(inputs(197)) or (inputs(74));
    layer0_outputs(2658) <= not(inputs(215));
    layer0_outputs(2659) <= (inputs(197)) and not (inputs(11));
    layer0_outputs(2660) <= inputs(104);
    layer0_outputs(2661) <= not((inputs(245)) and (inputs(53)));
    layer0_outputs(2662) <= not(inputs(178));
    layer0_outputs(2663) <= (inputs(7)) and not (inputs(112));
    layer0_outputs(2664) <= (inputs(206)) and not (inputs(171));
    layer0_outputs(2665) <= not(inputs(219)) or (inputs(146));
    layer0_outputs(2666) <= not(inputs(168)) or (inputs(118));
    layer0_outputs(2667) <= (inputs(173)) and (inputs(199));
    layer0_outputs(2668) <= not((inputs(74)) and (inputs(35)));
    layer0_outputs(2669) <= (inputs(9)) and not (inputs(172));
    layer0_outputs(2670) <= inputs(103);
    layer0_outputs(2671) <= (inputs(53)) xor (inputs(20));
    layer0_outputs(2672) <= '1';
    layer0_outputs(2673) <= inputs(142);
    layer0_outputs(2674) <= (inputs(176)) or (inputs(86));
    layer0_outputs(2675) <= not((inputs(29)) xor (inputs(19)));
    layer0_outputs(2676) <= (inputs(65)) or (inputs(243));
    layer0_outputs(2677) <= inputs(219);
    layer0_outputs(2678) <= (inputs(186)) or (inputs(221));
    layer0_outputs(2679) <= not(inputs(140)) or (inputs(93));
    layer0_outputs(2680) <= (inputs(198)) and not (inputs(250));
    layer0_outputs(2681) <= not(inputs(225)) or (inputs(0));
    layer0_outputs(2682) <= inputs(71);
    layer0_outputs(2683) <= inputs(20);
    layer0_outputs(2684) <= inputs(66);
    layer0_outputs(2685) <= inputs(24);
    layer0_outputs(2686) <= not((inputs(0)) xor (inputs(155)));
    layer0_outputs(2687) <= inputs(27);
    layer0_outputs(2688) <= (inputs(97)) or (inputs(166));
    layer0_outputs(2689) <= (inputs(18)) and (inputs(111));
    layer0_outputs(2690) <= not(inputs(230));
    layer0_outputs(2691) <= not(inputs(64));
    layer0_outputs(2692) <= not((inputs(104)) and (inputs(73)));
    layer0_outputs(2693) <= not((inputs(59)) or (inputs(61)));
    layer0_outputs(2694) <= not(inputs(171));
    layer0_outputs(2695) <= inputs(110);
    layer0_outputs(2696) <= not(inputs(150)) or (inputs(141));
    layer0_outputs(2697) <= not(inputs(11));
    layer0_outputs(2698) <= not(inputs(194));
    layer0_outputs(2699) <= (inputs(25)) and not (inputs(174));
    layer0_outputs(2700) <= inputs(210);
    layer0_outputs(2701) <= '1';
    layer0_outputs(2702) <= not(inputs(154)) or (inputs(193));
    layer0_outputs(2703) <= (inputs(61)) or (inputs(107));
    layer0_outputs(2704) <= (inputs(62)) or (inputs(104));
    layer0_outputs(2705) <= (inputs(46)) or (inputs(114));
    layer0_outputs(2706) <= inputs(20);
    layer0_outputs(2707) <= not(inputs(230));
    layer0_outputs(2708) <= (inputs(119)) or (inputs(89));
    layer0_outputs(2709) <= not((inputs(8)) or (inputs(143)));
    layer0_outputs(2710) <= not(inputs(194)) or (inputs(239));
    layer0_outputs(2711) <= not((inputs(18)) or (inputs(120)));
    layer0_outputs(2712) <= not((inputs(26)) or (inputs(143)));
    layer0_outputs(2713) <= (inputs(233)) or (inputs(142));
    layer0_outputs(2714) <= inputs(161);
    layer0_outputs(2715) <= not(inputs(196));
    layer0_outputs(2716) <= (inputs(182)) or (inputs(125));
    layer0_outputs(2717) <= '1';
    layer0_outputs(2718) <= (inputs(38)) and not (inputs(202));
    layer0_outputs(2719) <= not((inputs(3)) xor (inputs(65)));
    layer0_outputs(2720) <= not(inputs(71)) or (inputs(5));
    layer0_outputs(2721) <= not(inputs(36)) or (inputs(4));
    layer0_outputs(2722) <= inputs(219);
    layer0_outputs(2723) <= not(inputs(225));
    layer0_outputs(2724) <= not((inputs(160)) xor (inputs(22)));
    layer0_outputs(2725) <= inputs(124);
    layer0_outputs(2726) <= not((inputs(136)) or (inputs(198)));
    layer0_outputs(2727) <= not((inputs(143)) or (inputs(72)));
    layer0_outputs(2728) <= inputs(97);
    layer0_outputs(2729) <= inputs(49);
    layer0_outputs(2730) <= (inputs(150)) and not (inputs(115));
    layer0_outputs(2731) <= not(inputs(23)) or (inputs(190));
    layer0_outputs(2732) <= not(inputs(73));
    layer0_outputs(2733) <= inputs(198);
    layer0_outputs(2734) <= not((inputs(103)) or (inputs(118)));
    layer0_outputs(2735) <= (inputs(255)) or (inputs(235));
    layer0_outputs(2736) <= '1';
    layer0_outputs(2737) <= inputs(37);
    layer0_outputs(2738) <= not((inputs(118)) or (inputs(93)));
    layer0_outputs(2739) <= not((inputs(221)) or (inputs(65)));
    layer0_outputs(2740) <= not((inputs(200)) or (inputs(2)));
    layer0_outputs(2741) <= inputs(222);
    layer0_outputs(2742) <= not(inputs(169)) or (inputs(172));
    layer0_outputs(2743) <= inputs(98);
    layer0_outputs(2744) <= not((inputs(162)) or (inputs(218)));
    layer0_outputs(2745) <= not(inputs(154)) or (inputs(22));
    layer0_outputs(2746) <= (inputs(131)) and (inputs(171));
    layer0_outputs(2747) <= (inputs(83)) xor (inputs(81));
    layer0_outputs(2748) <= '0';
    layer0_outputs(2749) <= (inputs(150)) or (inputs(89));
    layer0_outputs(2750) <= not((inputs(217)) or (inputs(100)));
    layer0_outputs(2751) <= (inputs(234)) and not (inputs(185));
    layer0_outputs(2752) <= (inputs(129)) and not (inputs(173));
    layer0_outputs(2753) <= not(inputs(95));
    layer0_outputs(2754) <= (inputs(108)) and not (inputs(14));
    layer0_outputs(2755) <= not(inputs(27));
    layer0_outputs(2756) <= not((inputs(68)) or (inputs(97)));
    layer0_outputs(2757) <= not(inputs(230)) or (inputs(104));
    layer0_outputs(2758) <= not((inputs(73)) and (inputs(80)));
    layer0_outputs(2759) <= not(inputs(68)) or (inputs(242));
    layer0_outputs(2760) <= not(inputs(11));
    layer0_outputs(2761) <= inputs(135);
    layer0_outputs(2762) <= (inputs(218)) or (inputs(140));
    layer0_outputs(2763) <= not(inputs(120)) or (inputs(18));
    layer0_outputs(2764) <= (inputs(136)) and not (inputs(172));
    layer0_outputs(2765) <= inputs(149);
    layer0_outputs(2766) <= not(inputs(52)) or (inputs(78));
    layer0_outputs(2767) <= (inputs(253)) or (inputs(199));
    layer0_outputs(2768) <= '0';
    layer0_outputs(2769) <= (inputs(7)) or (inputs(78));
    layer0_outputs(2770) <= not((inputs(35)) and (inputs(241)));
    layer0_outputs(2771) <= not(inputs(244));
    layer0_outputs(2772) <= '1';
    layer0_outputs(2773) <= (inputs(138)) and not (inputs(131));
    layer0_outputs(2774) <= not((inputs(225)) or (inputs(104)));
    layer0_outputs(2775) <= not(inputs(190));
    layer0_outputs(2776) <= not(inputs(220)) or (inputs(130));
    layer0_outputs(2777) <= not(inputs(123)) or (inputs(131));
    layer0_outputs(2778) <= '0';
    layer0_outputs(2779) <= inputs(120);
    layer0_outputs(2780) <= inputs(21);
    layer0_outputs(2781) <= not((inputs(88)) xor (inputs(88)));
    layer0_outputs(2782) <= not((inputs(134)) and (inputs(160)));
    layer0_outputs(2783) <= not(inputs(203));
    layer0_outputs(2784) <= not(inputs(221));
    layer0_outputs(2785) <= not((inputs(99)) or (inputs(208)));
    layer0_outputs(2786) <= not((inputs(31)) or (inputs(139)));
    layer0_outputs(2787) <= not(inputs(152)) or (inputs(202));
    layer0_outputs(2788) <= (inputs(73)) and not (inputs(81));
    layer0_outputs(2789) <= not(inputs(223)) or (inputs(142));
    layer0_outputs(2790) <= (inputs(18)) and not (inputs(200));
    layer0_outputs(2791) <= not(inputs(119)) or (inputs(186));
    layer0_outputs(2792) <= (inputs(37)) and not (inputs(71));
    layer0_outputs(2793) <= (inputs(154)) and not (inputs(107));
    layer0_outputs(2794) <= not(inputs(67));
    layer0_outputs(2795) <= not(inputs(73));
    layer0_outputs(2796) <= not(inputs(77));
    layer0_outputs(2797) <= (inputs(50)) and not (inputs(191));
    layer0_outputs(2798) <= not((inputs(229)) or (inputs(174)));
    layer0_outputs(2799) <= inputs(211);
    layer0_outputs(2800) <= inputs(33);
    layer0_outputs(2801) <= (inputs(108)) or (inputs(83));
    layer0_outputs(2802) <= (inputs(61)) and not (inputs(124));
    layer0_outputs(2803) <= not(inputs(24)) or (inputs(155));
    layer0_outputs(2804) <= not((inputs(215)) or (inputs(76)));
    layer0_outputs(2805) <= not(inputs(9)) or (inputs(65));
    layer0_outputs(2806) <= not((inputs(31)) or (inputs(19)));
    layer0_outputs(2807) <= not(inputs(120));
    layer0_outputs(2808) <= inputs(99);
    layer0_outputs(2809) <= not(inputs(137));
    layer0_outputs(2810) <= not(inputs(58));
    layer0_outputs(2811) <= not((inputs(7)) or (inputs(212)));
    layer0_outputs(2812) <= inputs(156);
    layer0_outputs(2813) <= not(inputs(64));
    layer0_outputs(2814) <= (inputs(234)) and not (inputs(72));
    layer0_outputs(2815) <= (inputs(252)) and not (inputs(80));
    layer0_outputs(2816) <= not((inputs(116)) or (inputs(246)));
    layer0_outputs(2817) <= not(inputs(109)) or (inputs(78));
    layer0_outputs(2818) <= not(inputs(142));
    layer0_outputs(2819) <= not(inputs(104)) or (inputs(48));
    layer0_outputs(2820) <= (inputs(42)) and not (inputs(111));
    layer0_outputs(2821) <= (inputs(112)) xor (inputs(133));
    layer0_outputs(2822) <= not(inputs(130));
    layer0_outputs(2823) <= not((inputs(161)) or (inputs(195)));
    layer0_outputs(2824) <= '0';
    layer0_outputs(2825) <= inputs(242);
    layer0_outputs(2826) <= (inputs(156)) or (inputs(186));
    layer0_outputs(2827) <= not(inputs(136));
    layer0_outputs(2828) <= (inputs(71)) and (inputs(254));
    layer0_outputs(2829) <= inputs(232);
    layer0_outputs(2830) <= inputs(167);
    layer0_outputs(2831) <= '0';
    layer0_outputs(2832) <= not(inputs(62)) or (inputs(187));
    layer0_outputs(2833) <= not((inputs(10)) or (inputs(78)));
    layer0_outputs(2834) <= not(inputs(231));
    layer0_outputs(2835) <= not(inputs(83));
    layer0_outputs(2836) <= not(inputs(204)) or (inputs(14));
    layer0_outputs(2837) <= (inputs(78)) or (inputs(246));
    layer0_outputs(2838) <= (inputs(157)) or (inputs(143));
    layer0_outputs(2839) <= inputs(110);
    layer0_outputs(2840) <= not((inputs(71)) xor (inputs(70)));
    layer0_outputs(2841) <= (inputs(145)) xor (inputs(157));
    layer0_outputs(2842) <= inputs(34);
    layer0_outputs(2843) <= not(inputs(244)) or (inputs(9));
    layer0_outputs(2844) <= '1';
    layer0_outputs(2845) <= (inputs(223)) or (inputs(178));
    layer0_outputs(2846) <= '1';
    layer0_outputs(2847) <= not((inputs(164)) or (inputs(19)));
    layer0_outputs(2848) <= inputs(210);
    layer0_outputs(2849) <= not(inputs(120));
    layer0_outputs(2850) <= not(inputs(0)) or (inputs(96));
    layer0_outputs(2851) <= (inputs(190)) or (inputs(189));
    layer0_outputs(2852) <= (inputs(137)) and not (inputs(214));
    layer0_outputs(2853) <= not(inputs(22));
    layer0_outputs(2854) <= not((inputs(45)) or (inputs(22)));
    layer0_outputs(2855) <= (inputs(198)) and not (inputs(115));
    layer0_outputs(2856) <= (inputs(82)) and not (inputs(111));
    layer0_outputs(2857) <= '0';
    layer0_outputs(2858) <= not(inputs(211)) or (inputs(9));
    layer0_outputs(2859) <= not((inputs(216)) and (inputs(28)));
    layer0_outputs(2860) <= not((inputs(24)) or (inputs(34)));
    layer0_outputs(2861) <= not(inputs(221)) or (inputs(127));
    layer0_outputs(2862) <= not(inputs(88)) or (inputs(159));
    layer0_outputs(2863) <= not(inputs(77));
    layer0_outputs(2864) <= not((inputs(4)) or (inputs(79)));
    layer0_outputs(2865) <= not(inputs(64)) or (inputs(38));
    layer0_outputs(2866) <= inputs(104);
    layer0_outputs(2867) <= not(inputs(139)) or (inputs(246));
    layer0_outputs(2868) <= '1';
    layer0_outputs(2869) <= not(inputs(70)) or (inputs(189));
    layer0_outputs(2870) <= (inputs(42)) and not (inputs(57));
    layer0_outputs(2871) <= inputs(27);
    layer0_outputs(2872) <= inputs(83);
    layer0_outputs(2873) <= inputs(201);
    layer0_outputs(2874) <= (inputs(103)) and not (inputs(198));
    layer0_outputs(2875) <= (inputs(153)) or (inputs(136));
    layer0_outputs(2876) <= not((inputs(204)) or (inputs(127)));
    layer0_outputs(2877) <= inputs(74);
    layer0_outputs(2878) <= '1';
    layer0_outputs(2879) <= not(inputs(138)) or (inputs(243));
    layer0_outputs(2880) <= inputs(249);
    layer0_outputs(2881) <= not(inputs(37)) or (inputs(144));
    layer0_outputs(2882) <= (inputs(162)) xor (inputs(234));
    layer0_outputs(2883) <= not(inputs(163));
    layer0_outputs(2884) <= not(inputs(167)) or (inputs(67));
    layer0_outputs(2885) <= not(inputs(196)) or (inputs(63));
    layer0_outputs(2886) <= '1';
    layer0_outputs(2887) <= (inputs(91)) and not (inputs(236));
    layer0_outputs(2888) <= inputs(182);
    layer0_outputs(2889) <= (inputs(12)) and not (inputs(93));
    layer0_outputs(2890) <= not((inputs(39)) or (inputs(86)));
    layer0_outputs(2891) <= inputs(29);
    layer0_outputs(2892) <= not(inputs(222));
    layer0_outputs(2893) <= not(inputs(109));
    layer0_outputs(2894) <= not(inputs(23));
    layer0_outputs(2895) <= not(inputs(77));
    layer0_outputs(2896) <= not((inputs(210)) and (inputs(18)));
    layer0_outputs(2897) <= not((inputs(214)) or (inputs(84)));
    layer0_outputs(2898) <= inputs(215);
    layer0_outputs(2899) <= inputs(50);
    layer0_outputs(2900) <= not(inputs(169)) or (inputs(103));
    layer0_outputs(2901) <= not((inputs(207)) xor (inputs(218)));
    layer0_outputs(2902) <= (inputs(236)) and (inputs(36));
    layer0_outputs(2903) <= not(inputs(161)) or (inputs(9));
    layer0_outputs(2904) <= not(inputs(23));
    layer0_outputs(2905) <= (inputs(203)) or (inputs(140));
    layer0_outputs(2906) <= (inputs(228)) or (inputs(170));
    layer0_outputs(2907) <= not(inputs(88)) or (inputs(125));
    layer0_outputs(2908) <= (inputs(161)) or (inputs(209));
    layer0_outputs(2909) <= '0';
    layer0_outputs(2910) <= (inputs(17)) or (inputs(125));
    layer0_outputs(2911) <= (inputs(83)) and not (inputs(227));
    layer0_outputs(2912) <= (inputs(192)) or (inputs(126));
    layer0_outputs(2913) <= not(inputs(66));
    layer0_outputs(2914) <= not(inputs(98));
    layer0_outputs(2915) <= not((inputs(123)) or (inputs(252)));
    layer0_outputs(2916) <= not(inputs(31)) or (inputs(93));
    layer0_outputs(2917) <= (inputs(125)) or (inputs(190));
    layer0_outputs(2918) <= not(inputs(139)) or (inputs(55));
    layer0_outputs(2919) <= not(inputs(85)) or (inputs(180));
    layer0_outputs(2920) <= (inputs(165)) or (inputs(148));
    layer0_outputs(2921) <= not(inputs(169));
    layer0_outputs(2922) <= (inputs(211)) or (inputs(139));
    layer0_outputs(2923) <= '1';
    layer0_outputs(2924) <= (inputs(44)) xor (inputs(0));
    layer0_outputs(2925) <= not((inputs(193)) or (inputs(179)));
    layer0_outputs(2926) <= not(inputs(120));
    layer0_outputs(2927) <= (inputs(227)) or (inputs(239));
    layer0_outputs(2928) <= not((inputs(192)) or (inputs(173)));
    layer0_outputs(2929) <= (inputs(82)) or (inputs(75));
    layer0_outputs(2930) <= not(inputs(177)) or (inputs(167));
    layer0_outputs(2931) <= inputs(68);
    layer0_outputs(2932) <= (inputs(246)) and not (inputs(43));
    layer0_outputs(2933) <= (inputs(16)) xor (inputs(12));
    layer0_outputs(2934) <= (inputs(183)) and not (inputs(157));
    layer0_outputs(2935) <= (inputs(128)) or (inputs(232));
    layer0_outputs(2936) <= (inputs(235)) or (inputs(208));
    layer0_outputs(2937) <= inputs(140);
    layer0_outputs(2938) <= '0';
    layer0_outputs(2939) <= inputs(121);
    layer0_outputs(2940) <= (inputs(251)) or (inputs(140));
    layer0_outputs(2941) <= (inputs(52)) or (inputs(94));
    layer0_outputs(2942) <= not(inputs(69));
    layer0_outputs(2943) <= not((inputs(65)) xor (inputs(20)));
    layer0_outputs(2944) <= not((inputs(80)) xor (inputs(74)));
    layer0_outputs(2945) <= not((inputs(76)) and (inputs(119)));
    layer0_outputs(2946) <= not((inputs(8)) and (inputs(10)));
    layer0_outputs(2947) <= not((inputs(161)) xor (inputs(190)));
    layer0_outputs(2948) <= (inputs(151)) or (inputs(111));
    layer0_outputs(2949) <= not(inputs(13)) or (inputs(80));
    layer0_outputs(2950) <= not((inputs(96)) or (inputs(154)));
    layer0_outputs(2951) <= not((inputs(112)) xor (inputs(162)));
    layer0_outputs(2952) <= (inputs(68)) and not (inputs(22));
    layer0_outputs(2953) <= not(inputs(113));
    layer0_outputs(2954) <= not(inputs(44));
    layer0_outputs(2955) <= (inputs(226)) or (inputs(148));
    layer0_outputs(2956) <= '0';
    layer0_outputs(2957) <= inputs(87);
    layer0_outputs(2958) <= not((inputs(75)) and (inputs(10)));
    layer0_outputs(2959) <= not((inputs(149)) or (inputs(251)));
    layer0_outputs(2960) <= not(inputs(49)) or (inputs(82));
    layer0_outputs(2961) <= not((inputs(245)) and (inputs(217)));
    layer0_outputs(2962) <= '1';
    layer0_outputs(2963) <= not(inputs(90)) or (inputs(86));
    layer0_outputs(2964) <= not(inputs(79));
    layer0_outputs(2965) <= inputs(143);
    layer0_outputs(2966) <= '0';
    layer0_outputs(2967) <= '1';
    layer0_outputs(2968) <= '0';
    layer0_outputs(2969) <= (inputs(19)) and not (inputs(83));
    layer0_outputs(2970) <= (inputs(182)) and not (inputs(200));
    layer0_outputs(2971) <= not((inputs(211)) or (inputs(189)));
    layer0_outputs(2972) <= not((inputs(108)) or (inputs(3)));
    layer0_outputs(2973) <= not(inputs(53));
    layer0_outputs(2974) <= (inputs(63)) or (inputs(95));
    layer0_outputs(2975) <= (inputs(229)) and (inputs(243));
    layer0_outputs(2976) <= not(inputs(79)) or (inputs(192));
    layer0_outputs(2977) <= inputs(52);
    layer0_outputs(2978) <= not(inputs(17));
    layer0_outputs(2979) <= not(inputs(170));
    layer0_outputs(2980) <= (inputs(38)) or (inputs(117));
    layer0_outputs(2981) <= not(inputs(183)) or (inputs(75));
    layer0_outputs(2982) <= (inputs(212)) or (inputs(67));
    layer0_outputs(2983) <= not((inputs(170)) xor (inputs(219)));
    layer0_outputs(2984) <= not(inputs(42)) or (inputs(88));
    layer0_outputs(2985) <= not(inputs(55));
    layer0_outputs(2986) <= '0';
    layer0_outputs(2987) <= not(inputs(170));
    layer0_outputs(2988) <= (inputs(174)) xor (inputs(243));
    layer0_outputs(2989) <= not((inputs(145)) or (inputs(231)));
    layer0_outputs(2990) <= (inputs(147)) and not (inputs(0));
    layer0_outputs(2991) <= not((inputs(243)) or (inputs(108)));
    layer0_outputs(2992) <= inputs(105);
    layer0_outputs(2993) <= not(inputs(124));
    layer0_outputs(2994) <= (inputs(67)) or (inputs(83));
    layer0_outputs(2995) <= inputs(246);
    layer0_outputs(2996) <= not(inputs(163));
    layer0_outputs(2997) <= not(inputs(90));
    layer0_outputs(2998) <= (inputs(139)) or (inputs(187));
    layer0_outputs(2999) <= not(inputs(18)) or (inputs(174));
    layer0_outputs(3000) <= not((inputs(160)) or (inputs(216)));
    layer0_outputs(3001) <= not((inputs(189)) or (inputs(211)));
    layer0_outputs(3002) <= '1';
    layer0_outputs(3003) <= inputs(205);
    layer0_outputs(3004) <= not(inputs(161));
    layer0_outputs(3005) <= (inputs(232)) xor (inputs(78));
    layer0_outputs(3006) <= (inputs(19)) xor (inputs(47));
    layer0_outputs(3007) <= inputs(65);
    layer0_outputs(3008) <= (inputs(147)) and not (inputs(49));
    layer0_outputs(3009) <= inputs(233);
    layer0_outputs(3010) <= inputs(113);
    layer0_outputs(3011) <= (inputs(38)) and not (inputs(159));
    layer0_outputs(3012) <= not(inputs(151));
    layer0_outputs(3013) <= not(inputs(143)) or (inputs(10));
    layer0_outputs(3014) <= not((inputs(200)) xor (inputs(248)));
    layer0_outputs(3015) <= not(inputs(138));
    layer0_outputs(3016) <= inputs(248);
    layer0_outputs(3017) <= not(inputs(227));
    layer0_outputs(3018) <= (inputs(205)) or (inputs(216));
    layer0_outputs(3019) <= '1';
    layer0_outputs(3020) <= not(inputs(116));
    layer0_outputs(3021) <= inputs(143);
    layer0_outputs(3022) <= not(inputs(8)) or (inputs(176));
    layer0_outputs(3023) <= (inputs(172)) xor (inputs(217));
    layer0_outputs(3024) <= not(inputs(178));
    layer0_outputs(3025) <= not(inputs(78));
    layer0_outputs(3026) <= inputs(146);
    layer0_outputs(3027) <= not(inputs(24)) or (inputs(183));
    layer0_outputs(3028) <= (inputs(222)) or (inputs(171));
    layer0_outputs(3029) <= not(inputs(83));
    layer0_outputs(3030) <= not(inputs(245)) or (inputs(45));
    layer0_outputs(3031) <= not(inputs(100)) or (inputs(95));
    layer0_outputs(3032) <= not((inputs(196)) or (inputs(1)));
    layer0_outputs(3033) <= not(inputs(64)) or (inputs(251));
    layer0_outputs(3034) <= not(inputs(171));
    layer0_outputs(3035) <= '1';
    layer0_outputs(3036) <= not(inputs(124)) or (inputs(213));
    layer0_outputs(3037) <= not(inputs(22)) or (inputs(249));
    layer0_outputs(3038) <= not(inputs(225));
    layer0_outputs(3039) <= '1';
    layer0_outputs(3040) <= not(inputs(239));
    layer0_outputs(3041) <= (inputs(66)) and (inputs(234));
    layer0_outputs(3042) <= not(inputs(71)) or (inputs(110));
    layer0_outputs(3043) <= inputs(212);
    layer0_outputs(3044) <= inputs(55);
    layer0_outputs(3045) <= (inputs(186)) and not (inputs(147));
    layer0_outputs(3046) <= inputs(232);
    layer0_outputs(3047) <= (inputs(9)) and not (inputs(129));
    layer0_outputs(3048) <= (inputs(230)) and not (inputs(90));
    layer0_outputs(3049) <= not((inputs(238)) xor (inputs(202)));
    layer0_outputs(3050) <= not(inputs(176)) or (inputs(139));
    layer0_outputs(3051) <= (inputs(246)) or (inputs(0));
    layer0_outputs(3052) <= (inputs(197)) and not (inputs(98));
    layer0_outputs(3053) <= inputs(177);
    layer0_outputs(3054) <= not(inputs(32)) or (inputs(134));
    layer0_outputs(3055) <= not(inputs(44)) or (inputs(226));
    layer0_outputs(3056) <= not(inputs(100)) or (inputs(16));
    layer0_outputs(3057) <= not(inputs(213));
    layer0_outputs(3058) <= not(inputs(23));
    layer0_outputs(3059) <= (inputs(243)) and not (inputs(71));
    layer0_outputs(3060) <= not(inputs(44));
    layer0_outputs(3061) <= inputs(205);
    layer0_outputs(3062) <= inputs(30);
    layer0_outputs(3063) <= not(inputs(64));
    layer0_outputs(3064) <= inputs(62);
    layer0_outputs(3065) <= (inputs(116)) and not (inputs(221));
    layer0_outputs(3066) <= (inputs(226)) or (inputs(129));
    layer0_outputs(3067) <= (inputs(169)) or (inputs(31));
    layer0_outputs(3068) <= not(inputs(179));
    layer0_outputs(3069) <= not(inputs(24)) or (inputs(248));
    layer0_outputs(3070) <= inputs(125);
    layer0_outputs(3071) <= '1';
    layer0_outputs(3072) <= inputs(144);
    layer0_outputs(3073) <= not(inputs(160));
    layer0_outputs(3074) <= not(inputs(233)) or (inputs(27));
    layer0_outputs(3075) <= not((inputs(74)) or (inputs(5)));
    layer0_outputs(3076) <= not((inputs(60)) or (inputs(225)));
    layer0_outputs(3077) <= '1';
    layer0_outputs(3078) <= (inputs(202)) and (inputs(214));
    layer0_outputs(3079) <= not(inputs(59)) or (inputs(222));
    layer0_outputs(3080) <= (inputs(123)) and not (inputs(63));
    layer0_outputs(3081) <= '1';
    layer0_outputs(3082) <= (inputs(198)) or (inputs(207));
    layer0_outputs(3083) <= inputs(163);
    layer0_outputs(3084) <= inputs(110);
    layer0_outputs(3085) <= not(inputs(69)) or (inputs(149));
    layer0_outputs(3086) <= (inputs(249)) or (inputs(213));
    layer0_outputs(3087) <= not(inputs(51)) or (inputs(26));
    layer0_outputs(3088) <= '0';
    layer0_outputs(3089) <= inputs(148);
    layer0_outputs(3090) <= not(inputs(22));
    layer0_outputs(3091) <= not((inputs(97)) or (inputs(42)));
    layer0_outputs(3092) <= (inputs(125)) or (inputs(113));
    layer0_outputs(3093) <= not((inputs(63)) xor (inputs(129)));
    layer0_outputs(3094) <= not((inputs(118)) or (inputs(223)));
    layer0_outputs(3095) <= inputs(64);
    layer0_outputs(3096) <= not(inputs(134));
    layer0_outputs(3097) <= (inputs(84)) and not (inputs(33));
    layer0_outputs(3098) <= (inputs(93)) or (inputs(23));
    layer0_outputs(3099) <= inputs(20);
    layer0_outputs(3100) <= not(inputs(228));
    layer0_outputs(3101) <= not(inputs(207));
    layer0_outputs(3102) <= not(inputs(122));
    layer0_outputs(3103) <= inputs(238);
    layer0_outputs(3104) <= not((inputs(44)) or (inputs(61)));
    layer0_outputs(3105) <= (inputs(44)) and (inputs(108));
    layer0_outputs(3106) <= not(inputs(61));
    layer0_outputs(3107) <= (inputs(127)) or (inputs(231));
    layer0_outputs(3108) <= not(inputs(58)) or (inputs(166));
    layer0_outputs(3109) <= (inputs(58)) or (inputs(87));
    layer0_outputs(3110) <= not((inputs(20)) or (inputs(125)));
    layer0_outputs(3111) <= inputs(61);
    layer0_outputs(3112) <= '1';
    layer0_outputs(3113) <= not(inputs(46));
    layer0_outputs(3114) <= not(inputs(120));
    layer0_outputs(3115) <= not(inputs(92));
    layer0_outputs(3116) <= not((inputs(32)) and (inputs(230)));
    layer0_outputs(3117) <= not(inputs(215));
    layer0_outputs(3118) <= (inputs(50)) and not (inputs(36));
    layer0_outputs(3119) <= inputs(77);
    layer0_outputs(3120) <= (inputs(139)) or (inputs(223));
    layer0_outputs(3121) <= not((inputs(133)) or (inputs(164)));
    layer0_outputs(3122) <= inputs(59);
    layer0_outputs(3123) <= '1';
    layer0_outputs(3124) <= not(inputs(45));
    layer0_outputs(3125) <= not((inputs(137)) or (inputs(34)));
    layer0_outputs(3126) <= inputs(100);
    layer0_outputs(3127) <= (inputs(166)) or (inputs(111));
    layer0_outputs(3128) <= inputs(26);
    layer0_outputs(3129) <= '0';
    layer0_outputs(3130) <= not((inputs(33)) xor (inputs(110)));
    layer0_outputs(3131) <= not(inputs(133));
    layer0_outputs(3132) <= not((inputs(255)) or (inputs(236)));
    layer0_outputs(3133) <= '1';
    layer0_outputs(3134) <= not(inputs(117)) or (inputs(10));
    layer0_outputs(3135) <= inputs(23);
    layer0_outputs(3136) <= (inputs(160)) and not (inputs(145));
    layer0_outputs(3137) <= inputs(244);
    layer0_outputs(3138) <= inputs(119);
    layer0_outputs(3139) <= not((inputs(44)) and (inputs(231)));
    layer0_outputs(3140) <= '1';
    layer0_outputs(3141) <= (inputs(106)) xor (inputs(127));
    layer0_outputs(3142) <= not(inputs(152));
    layer0_outputs(3143) <= (inputs(232)) or (inputs(247));
    layer0_outputs(3144) <= not((inputs(182)) xor (inputs(150)));
    layer0_outputs(3145) <= not(inputs(2));
    layer0_outputs(3146) <= (inputs(155)) or (inputs(206));
    layer0_outputs(3147) <= inputs(91);
    layer0_outputs(3148) <= not((inputs(221)) or (inputs(15)));
    layer0_outputs(3149) <= (inputs(201)) and not (inputs(13));
    layer0_outputs(3150) <= (inputs(63)) or (inputs(43));
    layer0_outputs(3151) <= not(inputs(72));
    layer0_outputs(3152) <= (inputs(83)) or (inputs(128));
    layer0_outputs(3153) <= inputs(132);
    layer0_outputs(3154) <= (inputs(244)) or (inputs(116));
    layer0_outputs(3155) <= (inputs(213)) or (inputs(219));
    layer0_outputs(3156) <= not(inputs(60));
    layer0_outputs(3157) <= (inputs(185)) and (inputs(177));
    layer0_outputs(3158) <= not((inputs(218)) xor (inputs(237)));
    layer0_outputs(3159) <= (inputs(198)) or (inputs(164));
    layer0_outputs(3160) <= (inputs(206)) or (inputs(62));
    layer0_outputs(3161) <= '0';
    layer0_outputs(3162) <= not(inputs(248)) or (inputs(146));
    layer0_outputs(3163) <= inputs(226);
    layer0_outputs(3164) <= inputs(230);
    layer0_outputs(3165) <= not((inputs(21)) or (inputs(32)));
    layer0_outputs(3166) <= not(inputs(66)) or (inputs(52));
    layer0_outputs(3167) <= not((inputs(223)) xor (inputs(22)));
    layer0_outputs(3168) <= not((inputs(108)) or (inputs(130)));
    layer0_outputs(3169) <= not((inputs(112)) or (inputs(82)));
    layer0_outputs(3170) <= (inputs(114)) or (inputs(169));
    layer0_outputs(3171) <= not(inputs(74));
    layer0_outputs(3172) <= not(inputs(47)) or (inputs(143));
    layer0_outputs(3173) <= inputs(64);
    layer0_outputs(3174) <= not((inputs(216)) and (inputs(226)));
    layer0_outputs(3175) <= not((inputs(105)) or (inputs(7)));
    layer0_outputs(3176) <= '0';
    layer0_outputs(3177) <= not((inputs(208)) or (inputs(167)));
    layer0_outputs(3178) <= not(inputs(181));
    layer0_outputs(3179) <= (inputs(3)) xor (inputs(101));
    layer0_outputs(3180) <= inputs(21);
    layer0_outputs(3181) <= not(inputs(212));
    layer0_outputs(3182) <= (inputs(179)) and not (inputs(107));
    layer0_outputs(3183) <= (inputs(62)) or (inputs(59));
    layer0_outputs(3184) <= (inputs(182)) or (inputs(5));
    layer0_outputs(3185) <= '1';
    layer0_outputs(3186) <= inputs(165);
    layer0_outputs(3187) <= (inputs(177)) and not (inputs(142));
    layer0_outputs(3188) <= not((inputs(149)) or (inputs(234)));
    layer0_outputs(3189) <= inputs(56);
    layer0_outputs(3190) <= (inputs(214)) and (inputs(214));
    layer0_outputs(3191) <= (inputs(73)) and (inputs(58));
    layer0_outputs(3192) <= inputs(101);
    layer0_outputs(3193) <= inputs(233);
    layer0_outputs(3194) <= not(inputs(32));
    layer0_outputs(3195) <= (inputs(70)) and (inputs(28));
    layer0_outputs(3196) <= not((inputs(199)) or (inputs(192)));
    layer0_outputs(3197) <= not(inputs(86)) or (inputs(1));
    layer0_outputs(3198) <= (inputs(65)) xor (inputs(238));
    layer0_outputs(3199) <= not(inputs(98));
    layer0_outputs(3200) <= (inputs(161)) or (inputs(85));
    layer0_outputs(3201) <= '0';
    layer0_outputs(3202) <= (inputs(114)) and not (inputs(169));
    layer0_outputs(3203) <= not(inputs(83));
    layer0_outputs(3204) <= (inputs(252)) or (inputs(85));
    layer0_outputs(3205) <= inputs(92);
    layer0_outputs(3206) <= not(inputs(122));
    layer0_outputs(3207) <= not(inputs(41)) or (inputs(147));
    layer0_outputs(3208) <= not(inputs(101));
    layer0_outputs(3209) <= (inputs(90)) and not (inputs(248));
    layer0_outputs(3210) <= not(inputs(131));
    layer0_outputs(3211) <= not((inputs(208)) or (inputs(84)));
    layer0_outputs(3212) <= not(inputs(151));
    layer0_outputs(3213) <= (inputs(127)) or (inputs(164));
    layer0_outputs(3214) <= '0';
    layer0_outputs(3215) <= not(inputs(156)) or (inputs(143));
    layer0_outputs(3216) <= not((inputs(70)) xor (inputs(133)));
    layer0_outputs(3217) <= (inputs(243)) and (inputs(174));
    layer0_outputs(3218) <= not(inputs(246));
    layer0_outputs(3219) <= inputs(137);
    layer0_outputs(3220) <= '0';
    layer0_outputs(3221) <= not((inputs(82)) xor (inputs(225)));
    layer0_outputs(3222) <= (inputs(207)) or (inputs(140));
    layer0_outputs(3223) <= inputs(207);
    layer0_outputs(3224) <= not((inputs(231)) or (inputs(143)));
    layer0_outputs(3225) <= (inputs(59)) or (inputs(123));
    layer0_outputs(3226) <= inputs(217);
    layer0_outputs(3227) <= not(inputs(179)) or (inputs(191));
    layer0_outputs(3228) <= (inputs(215)) and (inputs(119));
    layer0_outputs(3229) <= not(inputs(103)) or (inputs(57));
    layer0_outputs(3230) <= inputs(111);
    layer0_outputs(3231) <= not(inputs(22)) or (inputs(84));
    layer0_outputs(3232) <= not(inputs(90));
    layer0_outputs(3233) <= not(inputs(212)) or (inputs(8));
    layer0_outputs(3234) <= not(inputs(223));
    layer0_outputs(3235) <= not((inputs(174)) xor (inputs(2)));
    layer0_outputs(3236) <= not(inputs(3));
    layer0_outputs(3237) <= (inputs(190)) or (inputs(225));
    layer0_outputs(3238) <= (inputs(223)) and (inputs(195));
    layer0_outputs(3239) <= not(inputs(55)) or (inputs(223));
    layer0_outputs(3240) <= (inputs(44)) xor (inputs(34));
    layer0_outputs(3241) <= (inputs(217)) or (inputs(233));
    layer0_outputs(3242) <= (inputs(36)) and (inputs(16));
    layer0_outputs(3243) <= (inputs(84)) or (inputs(64));
    layer0_outputs(3244) <= inputs(165);
    layer0_outputs(3245) <= (inputs(191)) or (inputs(194));
    layer0_outputs(3246) <= not((inputs(183)) and (inputs(7)));
    layer0_outputs(3247) <= (inputs(227)) and not (inputs(172));
    layer0_outputs(3248) <= inputs(131);
    layer0_outputs(3249) <= not(inputs(83)) or (inputs(208));
    layer0_outputs(3250) <= (inputs(253)) xor (inputs(177));
    layer0_outputs(3251) <= inputs(131);
    layer0_outputs(3252) <= not((inputs(247)) and (inputs(54)));
    layer0_outputs(3253) <= '1';
    layer0_outputs(3254) <= (inputs(120)) or (inputs(86));
    layer0_outputs(3255) <= (inputs(20)) xor (inputs(113));
    layer0_outputs(3256) <= inputs(106);
    layer0_outputs(3257) <= not((inputs(158)) or (inputs(230)));
    layer0_outputs(3258) <= inputs(230);
    layer0_outputs(3259) <= (inputs(130)) and (inputs(161));
    layer0_outputs(3260) <= (inputs(123)) xor (inputs(149));
    layer0_outputs(3261) <= (inputs(106)) or (inputs(78));
    layer0_outputs(3262) <= (inputs(18)) or (inputs(155));
    layer0_outputs(3263) <= not(inputs(18));
    layer0_outputs(3264) <= not(inputs(4)) or (inputs(239));
    layer0_outputs(3265) <= not(inputs(71));
    layer0_outputs(3266) <= '1';
    layer0_outputs(3267) <= (inputs(224)) and not (inputs(23));
    layer0_outputs(3268) <= not((inputs(205)) or (inputs(92)));
    layer0_outputs(3269) <= '0';
    layer0_outputs(3270) <= (inputs(10)) xor (inputs(59));
    layer0_outputs(3271) <= (inputs(87)) and (inputs(64));
    layer0_outputs(3272) <= inputs(103);
    layer0_outputs(3273) <= not((inputs(53)) and (inputs(55)));
    layer0_outputs(3274) <= (inputs(77)) xor (inputs(154));
    layer0_outputs(3275) <= (inputs(188)) and not (inputs(48));
    layer0_outputs(3276) <= inputs(15);
    layer0_outputs(3277) <= not((inputs(24)) or (inputs(110)));
    layer0_outputs(3278) <= not((inputs(111)) and (inputs(6)));
    layer0_outputs(3279) <= (inputs(188)) and not (inputs(27));
    layer0_outputs(3280) <= not(inputs(151)) or (inputs(17));
    layer0_outputs(3281) <= (inputs(32)) xor (inputs(80));
    layer0_outputs(3282) <= not(inputs(169));
    layer0_outputs(3283) <= not(inputs(145));
    layer0_outputs(3284) <= inputs(212);
    layer0_outputs(3285) <= (inputs(54)) and (inputs(10));
    layer0_outputs(3286) <= not((inputs(219)) or (inputs(189)));
    layer0_outputs(3287) <= not(inputs(7));
    layer0_outputs(3288) <= (inputs(60)) xor (inputs(30));
    layer0_outputs(3289) <= (inputs(177)) xor (inputs(231));
    layer0_outputs(3290) <= not(inputs(89)) or (inputs(2));
    layer0_outputs(3291) <= (inputs(152)) xor (inputs(146));
    layer0_outputs(3292) <= (inputs(120)) and not (inputs(124));
    layer0_outputs(3293) <= not(inputs(160));
    layer0_outputs(3294) <= not(inputs(123));
    layer0_outputs(3295) <= not(inputs(12)) or (inputs(251));
    layer0_outputs(3296) <= inputs(10);
    layer0_outputs(3297) <= not(inputs(11)) or (inputs(222));
    layer0_outputs(3298) <= not((inputs(48)) or (inputs(225)));
    layer0_outputs(3299) <= (inputs(250)) or (inputs(17));
    layer0_outputs(3300) <= inputs(25);
    layer0_outputs(3301) <= not(inputs(117));
    layer0_outputs(3302) <= inputs(214);
    layer0_outputs(3303) <= not((inputs(147)) xor (inputs(174)));
    layer0_outputs(3304) <= not(inputs(4));
    layer0_outputs(3305) <= inputs(192);
    layer0_outputs(3306) <= not((inputs(89)) or (inputs(157)));
    layer0_outputs(3307) <= not(inputs(186));
    layer0_outputs(3308) <= not(inputs(118)) or (inputs(75));
    layer0_outputs(3309) <= (inputs(100)) or (inputs(253));
    layer0_outputs(3310) <= inputs(98);
    layer0_outputs(3311) <= not(inputs(189));
    layer0_outputs(3312) <= not((inputs(88)) or (inputs(239)));
    layer0_outputs(3313) <= (inputs(3)) and not (inputs(239));
    layer0_outputs(3314) <= inputs(55);
    layer0_outputs(3315) <= not((inputs(210)) xor (inputs(240)));
    layer0_outputs(3316) <= not((inputs(2)) xor (inputs(237)));
    layer0_outputs(3317) <= (inputs(177)) and (inputs(94));
    layer0_outputs(3318) <= inputs(162);
    layer0_outputs(3319) <= (inputs(2)) and not (inputs(91));
    layer0_outputs(3320) <= (inputs(145)) or (inputs(112));
    layer0_outputs(3321) <= not(inputs(189)) or (inputs(92));
    layer0_outputs(3322) <= not(inputs(20));
    layer0_outputs(3323) <= not((inputs(160)) or (inputs(189)));
    layer0_outputs(3324) <= not(inputs(29));
    layer0_outputs(3325) <= not((inputs(203)) or (inputs(239)));
    layer0_outputs(3326) <= (inputs(143)) and not (inputs(119));
    layer0_outputs(3327) <= not(inputs(46)) or (inputs(253));
    layer0_outputs(3328) <= not(inputs(227)) or (inputs(17));
    layer0_outputs(3329) <= (inputs(18)) xor (inputs(250));
    layer0_outputs(3330) <= not(inputs(165));
    layer0_outputs(3331) <= not(inputs(244)) or (inputs(114));
    layer0_outputs(3332) <= not(inputs(179));
    layer0_outputs(3333) <= not(inputs(243));
    layer0_outputs(3334) <= (inputs(8)) or (inputs(156));
    layer0_outputs(3335) <= not(inputs(6)) or (inputs(112));
    layer0_outputs(3336) <= not(inputs(77));
    layer0_outputs(3337) <= not(inputs(176)) or (inputs(0));
    layer0_outputs(3338) <= not(inputs(173)) or (inputs(42));
    layer0_outputs(3339) <= (inputs(169)) and not (inputs(144));
    layer0_outputs(3340) <= not(inputs(198));
    layer0_outputs(3341) <= not(inputs(152));
    layer0_outputs(3342) <= inputs(240);
    layer0_outputs(3343) <= not(inputs(69)) or (inputs(244));
    layer0_outputs(3344) <= '0';
    layer0_outputs(3345) <= not(inputs(100)) or (inputs(149));
    layer0_outputs(3346) <= not(inputs(55));
    layer0_outputs(3347) <= '0';
    layer0_outputs(3348) <= inputs(136);
    layer0_outputs(3349) <= (inputs(26)) and not (inputs(160));
    layer0_outputs(3350) <= not(inputs(70)) or (inputs(143));
    layer0_outputs(3351) <= not(inputs(52));
    layer0_outputs(3352) <= not((inputs(172)) or (inputs(235)));
    layer0_outputs(3353) <= inputs(53);
    layer0_outputs(3354) <= not(inputs(213)) or (inputs(97));
    layer0_outputs(3355) <= not((inputs(129)) or (inputs(67)));
    layer0_outputs(3356) <= not(inputs(229)) or (inputs(237));
    layer0_outputs(3357) <= not((inputs(191)) or (inputs(3)));
    layer0_outputs(3358) <= not(inputs(74)) or (inputs(158));
    layer0_outputs(3359) <= (inputs(167)) and (inputs(59));
    layer0_outputs(3360) <= '0';
    layer0_outputs(3361) <= not(inputs(116));
    layer0_outputs(3362) <= (inputs(252)) xor (inputs(134));
    layer0_outputs(3363) <= not(inputs(145)) or (inputs(34));
    layer0_outputs(3364) <= not(inputs(63));
    layer0_outputs(3365) <= inputs(75);
    layer0_outputs(3366) <= (inputs(137)) xor (inputs(237));
    layer0_outputs(3367) <= not(inputs(98));
    layer0_outputs(3368) <= inputs(247);
    layer0_outputs(3369) <= not((inputs(89)) or (inputs(247)));
    layer0_outputs(3370) <= not(inputs(226));
    layer0_outputs(3371) <= '0';
    layer0_outputs(3372) <= '1';
    layer0_outputs(3373) <= not(inputs(93));
    layer0_outputs(3374) <= (inputs(238)) or (inputs(255));
    layer0_outputs(3375) <= '0';
    layer0_outputs(3376) <= inputs(52);
    layer0_outputs(3377) <= '1';
    layer0_outputs(3378) <= '0';
    layer0_outputs(3379) <= not(inputs(39));
    layer0_outputs(3380) <= '1';
    layer0_outputs(3381) <= not(inputs(148));
    layer0_outputs(3382) <= inputs(105);
    layer0_outputs(3383) <= '1';
    layer0_outputs(3384) <= not(inputs(4));
    layer0_outputs(3385) <= not(inputs(215)) or (inputs(226));
    layer0_outputs(3386) <= inputs(112);
    layer0_outputs(3387) <= (inputs(94)) and not (inputs(200));
    layer0_outputs(3388) <= (inputs(205)) and not (inputs(0));
    layer0_outputs(3389) <= not((inputs(236)) or (inputs(214)));
    layer0_outputs(3390) <= not(inputs(187));
    layer0_outputs(3391) <= not(inputs(149));
    layer0_outputs(3392) <= not(inputs(29));
    layer0_outputs(3393) <= not(inputs(92)) or (inputs(105));
    layer0_outputs(3394) <= '0';
    layer0_outputs(3395) <= not((inputs(122)) and (inputs(14)));
    layer0_outputs(3396) <= (inputs(4)) xor (inputs(69));
    layer0_outputs(3397) <= (inputs(86)) or (inputs(237));
    layer0_outputs(3398) <= (inputs(248)) and not (inputs(222));
    layer0_outputs(3399) <= inputs(9);
    layer0_outputs(3400) <= not((inputs(216)) xor (inputs(183)));
    layer0_outputs(3401) <= (inputs(133)) xor (inputs(197));
    layer0_outputs(3402) <= not((inputs(73)) and (inputs(183)));
    layer0_outputs(3403) <= not((inputs(249)) or (inputs(150)));
    layer0_outputs(3404) <= not(inputs(67));
    layer0_outputs(3405) <= not(inputs(25));
    layer0_outputs(3406) <= '0';
    layer0_outputs(3407) <= (inputs(59)) or (inputs(100));
    layer0_outputs(3408) <= (inputs(216)) and not (inputs(88));
    layer0_outputs(3409) <= not(inputs(192));
    layer0_outputs(3410) <= not(inputs(216));
    layer0_outputs(3411) <= (inputs(187)) or (inputs(60));
    layer0_outputs(3412) <= not(inputs(40));
    layer0_outputs(3413) <= not((inputs(86)) xor (inputs(102)));
    layer0_outputs(3414) <= not(inputs(107)) or (inputs(111));
    layer0_outputs(3415) <= (inputs(46)) or (inputs(234));
    layer0_outputs(3416) <= (inputs(41)) or (inputs(105));
    layer0_outputs(3417) <= (inputs(227)) and not (inputs(180));
    layer0_outputs(3418) <= (inputs(192)) or (inputs(166));
    layer0_outputs(3419) <= inputs(179);
    layer0_outputs(3420) <= (inputs(8)) or (inputs(238));
    layer0_outputs(3421) <= inputs(151);
    layer0_outputs(3422) <= not((inputs(100)) or (inputs(186)));
    layer0_outputs(3423) <= (inputs(2)) or (inputs(93));
    layer0_outputs(3424) <= (inputs(104)) and not (inputs(5));
    layer0_outputs(3425) <= not(inputs(13));
    layer0_outputs(3426) <= inputs(101);
    layer0_outputs(3427) <= '1';
    layer0_outputs(3428) <= not((inputs(138)) or (inputs(186)));
    layer0_outputs(3429) <= (inputs(148)) or (inputs(51));
    layer0_outputs(3430) <= not((inputs(101)) or (inputs(117)));
    layer0_outputs(3431) <= not((inputs(19)) or (inputs(219)));
    layer0_outputs(3432) <= inputs(160);
    layer0_outputs(3433) <= not((inputs(212)) xor (inputs(227)));
    layer0_outputs(3434) <= not((inputs(230)) xor (inputs(191)));
    layer0_outputs(3435) <= (inputs(242)) or (inputs(253));
    layer0_outputs(3436) <= (inputs(194)) and not (inputs(168));
    layer0_outputs(3437) <= inputs(186);
    layer0_outputs(3438) <= not(inputs(248)) or (inputs(61));
    layer0_outputs(3439) <= (inputs(199)) and (inputs(189));
    layer0_outputs(3440) <= not(inputs(24)) or (inputs(132));
    layer0_outputs(3441) <= not(inputs(132)) or (inputs(5));
    layer0_outputs(3442) <= inputs(229);
    layer0_outputs(3443) <= not(inputs(151));
    layer0_outputs(3444) <= not(inputs(156)) or (inputs(29));
    layer0_outputs(3445) <= not(inputs(46)) or (inputs(182));
    layer0_outputs(3446) <= not(inputs(4)) or (inputs(82));
    layer0_outputs(3447) <= (inputs(153)) and not (inputs(28));
    layer0_outputs(3448) <= not(inputs(142));
    layer0_outputs(3449) <= (inputs(239)) or (inputs(223));
    layer0_outputs(3450) <= not(inputs(7));
    layer0_outputs(3451) <= '0';
    layer0_outputs(3452) <= not(inputs(168)) or (inputs(2));
    layer0_outputs(3453) <= not(inputs(35));
    layer0_outputs(3454) <= inputs(126);
    layer0_outputs(3455) <= not(inputs(212));
    layer0_outputs(3456) <= inputs(121);
    layer0_outputs(3457) <= not((inputs(141)) or (inputs(210)));
    layer0_outputs(3458) <= not((inputs(206)) or (inputs(115)));
    layer0_outputs(3459) <= '0';
    layer0_outputs(3460) <= (inputs(230)) or (inputs(169));
    layer0_outputs(3461) <= not((inputs(117)) or (inputs(102)));
    layer0_outputs(3462) <= not(inputs(14));
    layer0_outputs(3463) <= (inputs(190)) or (inputs(158));
    layer0_outputs(3464) <= inputs(104);
    layer0_outputs(3465) <= inputs(25);
    layer0_outputs(3466) <= inputs(253);
    layer0_outputs(3467) <= not((inputs(245)) or (inputs(97)));
    layer0_outputs(3468) <= not((inputs(43)) or (inputs(197)));
    layer0_outputs(3469) <= (inputs(218)) xor (inputs(63));
    layer0_outputs(3470) <= inputs(130);
    layer0_outputs(3471) <= inputs(131);
    layer0_outputs(3472) <= not(inputs(242)) or (inputs(92));
    layer0_outputs(3473) <= inputs(19);
    layer0_outputs(3474) <= not(inputs(183)) or (inputs(253));
    layer0_outputs(3475) <= not(inputs(167)) or (inputs(185));
    layer0_outputs(3476) <= not(inputs(129)) or (inputs(57));
    layer0_outputs(3477) <= not(inputs(193)) or (inputs(173));
    layer0_outputs(3478) <= (inputs(147)) and not (inputs(53));
    layer0_outputs(3479) <= inputs(84);
    layer0_outputs(3480) <= not((inputs(161)) or (inputs(204)));
    layer0_outputs(3481) <= not(inputs(103));
    layer0_outputs(3482) <= (inputs(47)) and (inputs(255));
    layer0_outputs(3483) <= (inputs(40)) and (inputs(166));
    layer0_outputs(3484) <= not((inputs(23)) or (inputs(69)));
    layer0_outputs(3485) <= inputs(98);
    layer0_outputs(3486) <= not((inputs(20)) and (inputs(255)));
    layer0_outputs(3487) <= not(inputs(9));
    layer0_outputs(3488) <= (inputs(191)) and (inputs(8));
    layer0_outputs(3489) <= not(inputs(183)) or (inputs(31));
    layer0_outputs(3490) <= not(inputs(79)) or (inputs(119));
    layer0_outputs(3491) <= inputs(206);
    layer0_outputs(3492) <= (inputs(71)) or (inputs(246));
    layer0_outputs(3493) <= not((inputs(205)) and (inputs(190)));
    layer0_outputs(3494) <= inputs(204);
    layer0_outputs(3495) <= (inputs(52)) and (inputs(157));
    layer0_outputs(3496) <= not((inputs(62)) or (inputs(158)));
    layer0_outputs(3497) <= inputs(245);
    layer0_outputs(3498) <= (inputs(57)) and not (inputs(251));
    layer0_outputs(3499) <= not(inputs(9)) or (inputs(161));
    layer0_outputs(3500) <= (inputs(148)) or (inputs(128));
    layer0_outputs(3501) <= '0';
    layer0_outputs(3502) <= not((inputs(103)) xor (inputs(51)));
    layer0_outputs(3503) <= (inputs(231)) and not (inputs(40));
    layer0_outputs(3504) <= not((inputs(232)) and (inputs(229)));
    layer0_outputs(3505) <= not(inputs(163));
    layer0_outputs(3506) <= not(inputs(255));
    layer0_outputs(3507) <= inputs(143);
    layer0_outputs(3508) <= not(inputs(60)) or (inputs(12));
    layer0_outputs(3509) <= not((inputs(51)) xor (inputs(94)));
    layer0_outputs(3510) <= not((inputs(150)) or (inputs(48)));
    layer0_outputs(3511) <= not((inputs(60)) or (inputs(76)));
    layer0_outputs(3512) <= '0';
    layer0_outputs(3513) <= '0';
    layer0_outputs(3514) <= not((inputs(176)) or (inputs(207)));
    layer0_outputs(3515) <= not((inputs(194)) or (inputs(177)));
    layer0_outputs(3516) <= not(inputs(43));
    layer0_outputs(3517) <= not(inputs(224)) or (inputs(219));
    layer0_outputs(3518) <= (inputs(203)) or (inputs(150));
    layer0_outputs(3519) <= (inputs(88)) and not (inputs(55));
    layer0_outputs(3520) <= '1';
    layer0_outputs(3521) <= '1';
    layer0_outputs(3522) <= not(inputs(189));
    layer0_outputs(3523) <= (inputs(7)) and (inputs(37));
    layer0_outputs(3524) <= not(inputs(49));
    layer0_outputs(3525) <= (inputs(103)) or (inputs(142));
    layer0_outputs(3526) <= not(inputs(235));
    layer0_outputs(3527) <= (inputs(101)) or (inputs(142));
    layer0_outputs(3528) <= not(inputs(25)) or (inputs(169));
    layer0_outputs(3529) <= (inputs(105)) and not (inputs(81));
    layer0_outputs(3530) <= not(inputs(98)) or (inputs(70));
    layer0_outputs(3531) <= not(inputs(184));
    layer0_outputs(3532) <= not(inputs(44)) or (inputs(215));
    layer0_outputs(3533) <= not(inputs(136)) or (inputs(204));
    layer0_outputs(3534) <= (inputs(92)) or (inputs(248));
    layer0_outputs(3535) <= not(inputs(119));
    layer0_outputs(3536) <= not(inputs(23));
    layer0_outputs(3537) <= not(inputs(193));
    layer0_outputs(3538) <= not((inputs(112)) and (inputs(239)));
    layer0_outputs(3539) <= not(inputs(32)) or (inputs(92));
    layer0_outputs(3540) <= (inputs(136)) and not (inputs(138));
    layer0_outputs(3541) <= inputs(117);
    layer0_outputs(3542) <= (inputs(222)) or (inputs(33));
    layer0_outputs(3543) <= not((inputs(254)) and (inputs(162)));
    layer0_outputs(3544) <= (inputs(36)) or (inputs(82));
    layer0_outputs(3545) <= '1';
    layer0_outputs(3546) <= (inputs(23)) and (inputs(27));
    layer0_outputs(3547) <= (inputs(132)) and not (inputs(79));
    layer0_outputs(3548) <= not(inputs(235));
    layer0_outputs(3549) <= not((inputs(236)) and (inputs(235)));
    layer0_outputs(3550) <= (inputs(206)) or (inputs(245));
    layer0_outputs(3551) <= (inputs(193)) or (inputs(41));
    layer0_outputs(3552) <= not((inputs(147)) or (inputs(161)));
    layer0_outputs(3553) <= '0';
    layer0_outputs(3554) <= inputs(162);
    layer0_outputs(3555) <= (inputs(52)) or (inputs(129));
    layer0_outputs(3556) <= not((inputs(86)) or (inputs(193)));
    layer0_outputs(3557) <= not((inputs(142)) xor (inputs(161)));
    layer0_outputs(3558) <= not(inputs(107));
    layer0_outputs(3559) <= not(inputs(184));
    layer0_outputs(3560) <= (inputs(118)) or (inputs(194));
    layer0_outputs(3561) <= (inputs(92)) xor (inputs(72));
    layer0_outputs(3562) <= not(inputs(179));
    layer0_outputs(3563) <= (inputs(205)) xor (inputs(94));
    layer0_outputs(3564) <= not(inputs(7));
    layer0_outputs(3565) <= not((inputs(47)) or (inputs(70)));
    layer0_outputs(3566) <= (inputs(112)) xor (inputs(84));
    layer0_outputs(3567) <= (inputs(200)) and not (inputs(210));
    layer0_outputs(3568) <= not(inputs(160));
    layer0_outputs(3569) <= inputs(30);
    layer0_outputs(3570) <= (inputs(80)) and (inputs(36));
    layer0_outputs(3571) <= not((inputs(62)) or (inputs(242)));
    layer0_outputs(3572) <= (inputs(65)) or (inputs(63));
    layer0_outputs(3573) <= not((inputs(114)) or (inputs(97)));
    layer0_outputs(3574) <= (inputs(240)) or (inputs(198));
    layer0_outputs(3575) <= not((inputs(73)) or (inputs(121)));
    layer0_outputs(3576) <= '1';
    layer0_outputs(3577) <= not(inputs(210));
    layer0_outputs(3578) <= not(inputs(200)) or (inputs(130));
    layer0_outputs(3579) <= (inputs(94)) or (inputs(15));
    layer0_outputs(3580) <= inputs(186);
    layer0_outputs(3581) <= (inputs(189)) and not (inputs(59));
    layer0_outputs(3582) <= (inputs(125)) and not (inputs(182));
    layer0_outputs(3583) <= not(inputs(215)) or (inputs(101));
    layer0_outputs(3584) <= (inputs(59)) and not (inputs(213));
    layer0_outputs(3585) <= not((inputs(153)) or (inputs(236)));
    layer0_outputs(3586) <= not(inputs(245));
    layer0_outputs(3587) <= '1';
    layer0_outputs(3588) <= (inputs(67)) or (inputs(52));
    layer0_outputs(3589) <= (inputs(48)) xor (inputs(103));
    layer0_outputs(3590) <= not((inputs(85)) or (inputs(175)));
    layer0_outputs(3591) <= (inputs(108)) and not (inputs(180));
    layer0_outputs(3592) <= (inputs(237)) and not (inputs(144));
    layer0_outputs(3593) <= '1';
    layer0_outputs(3594) <= not((inputs(39)) and (inputs(123)));
    layer0_outputs(3595) <= inputs(191);
    layer0_outputs(3596) <= inputs(244);
    layer0_outputs(3597) <= (inputs(232)) or (inputs(217));
    layer0_outputs(3598) <= not((inputs(16)) or (inputs(89)));
    layer0_outputs(3599) <= (inputs(163)) and not (inputs(31));
    layer0_outputs(3600) <= (inputs(85)) xor (inputs(113));
    layer0_outputs(3601) <= inputs(211);
    layer0_outputs(3602) <= not(inputs(229)) or (inputs(109));
    layer0_outputs(3603) <= not((inputs(8)) and (inputs(72)));
    layer0_outputs(3604) <= (inputs(175)) or (inputs(210));
    layer0_outputs(3605) <= not(inputs(252)) or (inputs(166));
    layer0_outputs(3606) <= not(inputs(226));
    layer0_outputs(3607) <= not((inputs(157)) or (inputs(229)));
    layer0_outputs(3608) <= not(inputs(146));
    layer0_outputs(3609) <= (inputs(99)) xor (inputs(85));
    layer0_outputs(3610) <= (inputs(6)) and not (inputs(100));
    layer0_outputs(3611) <= inputs(3);
    layer0_outputs(3612) <= (inputs(56)) and not (inputs(102));
    layer0_outputs(3613) <= inputs(48);
    layer0_outputs(3614) <= not(inputs(179));
    layer0_outputs(3615) <= (inputs(26)) and not (inputs(161));
    layer0_outputs(3616) <= not(inputs(28)) or (inputs(199));
    layer0_outputs(3617) <= not((inputs(141)) and (inputs(113)));
    layer0_outputs(3618) <= inputs(23);
    layer0_outputs(3619) <= (inputs(117)) or (inputs(232));
    layer0_outputs(3620) <= (inputs(213)) and not (inputs(240));
    layer0_outputs(3621) <= not((inputs(234)) xor (inputs(106)));
    layer0_outputs(3622) <= not(inputs(121));
    layer0_outputs(3623) <= not(inputs(135));
    layer0_outputs(3624) <= not(inputs(117));
    layer0_outputs(3625) <= inputs(24);
    layer0_outputs(3626) <= inputs(198);
    layer0_outputs(3627) <= not((inputs(199)) or (inputs(192)));
    layer0_outputs(3628) <= inputs(148);
    layer0_outputs(3629) <= not(inputs(204)) or (inputs(114));
    layer0_outputs(3630) <= inputs(142);
    layer0_outputs(3631) <= (inputs(163)) and not (inputs(157));
    layer0_outputs(3632) <= inputs(95);
    layer0_outputs(3633) <= '0';
    layer0_outputs(3634) <= not((inputs(205)) or (inputs(131)));
    layer0_outputs(3635) <= not((inputs(123)) or (inputs(203)));
    layer0_outputs(3636) <= not(inputs(112)) or (inputs(17));
    layer0_outputs(3637) <= not((inputs(33)) xor (inputs(139)));
    layer0_outputs(3638) <= not(inputs(121)) or (inputs(201));
    layer0_outputs(3639) <= not((inputs(234)) xor (inputs(164)));
    layer0_outputs(3640) <= (inputs(74)) and not (inputs(127));
    layer0_outputs(3641) <= (inputs(74)) xor (inputs(42));
    layer0_outputs(3642) <= not((inputs(70)) xor (inputs(12)));
    layer0_outputs(3643) <= (inputs(82)) or (inputs(229));
    layer0_outputs(3644) <= not((inputs(230)) or (inputs(208)));
    layer0_outputs(3645) <= '0';
    layer0_outputs(3646) <= not(inputs(149));
    layer0_outputs(3647) <= inputs(117);
    layer0_outputs(3648) <= not((inputs(101)) or (inputs(29)));
    layer0_outputs(3649) <= (inputs(26)) or (inputs(197));
    layer0_outputs(3650) <= '0';
    layer0_outputs(3651) <= '1';
    layer0_outputs(3652) <= inputs(164);
    layer0_outputs(3653) <= not(inputs(113));
    layer0_outputs(3654) <= '0';
    layer0_outputs(3655) <= inputs(215);
    layer0_outputs(3656) <= not((inputs(98)) and (inputs(242)));
    layer0_outputs(3657) <= inputs(55);
    layer0_outputs(3658) <= inputs(142);
    layer0_outputs(3659) <= not((inputs(188)) or (inputs(223)));
    layer0_outputs(3660) <= (inputs(176)) or (inputs(25));
    layer0_outputs(3661) <= not((inputs(99)) or (inputs(14)));
    layer0_outputs(3662) <= not(inputs(106));
    layer0_outputs(3663) <= '1';
    layer0_outputs(3664) <= not(inputs(9));
    layer0_outputs(3665) <= not((inputs(151)) or (inputs(38)));
    layer0_outputs(3666) <= '1';
    layer0_outputs(3667) <= '0';
    layer0_outputs(3668) <= (inputs(209)) or (inputs(222));
    layer0_outputs(3669) <= (inputs(140)) and not (inputs(169));
    layer0_outputs(3670) <= not(inputs(45)) or (inputs(92));
    layer0_outputs(3671) <= not((inputs(11)) or (inputs(99)));
    layer0_outputs(3672) <= not(inputs(234));
    layer0_outputs(3673) <= not(inputs(217)) or (inputs(113));
    layer0_outputs(3674) <= not((inputs(177)) or (inputs(231)));
    layer0_outputs(3675) <= inputs(158);
    layer0_outputs(3676) <= not((inputs(107)) or (inputs(83)));
    layer0_outputs(3677) <= (inputs(183)) xor (inputs(113));
    layer0_outputs(3678) <= not((inputs(130)) or (inputs(176)));
    layer0_outputs(3679) <= (inputs(111)) or (inputs(141));
    layer0_outputs(3680) <= inputs(93);
    layer0_outputs(3681) <= not(inputs(24));
    layer0_outputs(3682) <= '1';
    layer0_outputs(3683) <= (inputs(27)) and (inputs(242));
    layer0_outputs(3684) <= not(inputs(105)) or (inputs(142));
    layer0_outputs(3685) <= inputs(60);
    layer0_outputs(3686) <= not(inputs(215));
    layer0_outputs(3687) <= not(inputs(134)) or (inputs(19));
    layer0_outputs(3688) <= not(inputs(36)) or (inputs(73));
    layer0_outputs(3689) <= not(inputs(42));
    layer0_outputs(3690) <= (inputs(203)) or (inputs(107));
    layer0_outputs(3691) <= inputs(116);
    layer0_outputs(3692) <= inputs(234);
    layer0_outputs(3693) <= not(inputs(140)) or (inputs(58));
    layer0_outputs(3694) <= not((inputs(221)) xor (inputs(224)));
    layer0_outputs(3695) <= not((inputs(78)) xor (inputs(91)));
    layer0_outputs(3696) <= (inputs(158)) or (inputs(246));
    layer0_outputs(3697) <= not((inputs(34)) or (inputs(192)));
    layer0_outputs(3698) <= inputs(226);
    layer0_outputs(3699) <= not((inputs(188)) or (inputs(24)));
    layer0_outputs(3700) <= inputs(134);
    layer0_outputs(3701) <= '0';
    layer0_outputs(3702) <= (inputs(68)) and not (inputs(222));
    layer0_outputs(3703) <= (inputs(205)) and not (inputs(115));
    layer0_outputs(3704) <= not(inputs(180));
    layer0_outputs(3705) <= (inputs(20)) and not (inputs(93));
    layer0_outputs(3706) <= inputs(58);
    layer0_outputs(3707) <= (inputs(227)) and not (inputs(105));
    layer0_outputs(3708) <= not(inputs(152));
    layer0_outputs(3709) <= not((inputs(193)) or (inputs(240)));
    layer0_outputs(3710) <= '1';
    layer0_outputs(3711) <= (inputs(238)) or (inputs(110));
    layer0_outputs(3712) <= (inputs(164)) xor (inputs(61));
    layer0_outputs(3713) <= not((inputs(204)) or (inputs(157)));
    layer0_outputs(3714) <= inputs(204);
    layer0_outputs(3715) <= (inputs(82)) or (inputs(182));
    layer0_outputs(3716) <= not((inputs(175)) and (inputs(191)));
    layer0_outputs(3717) <= not(inputs(135));
    layer0_outputs(3718) <= (inputs(211)) or (inputs(113));
    layer0_outputs(3719) <= not((inputs(75)) and (inputs(185)));
    layer0_outputs(3720) <= '1';
    layer0_outputs(3721) <= (inputs(9)) and not (inputs(179));
    layer0_outputs(3722) <= (inputs(9)) and (inputs(121));
    layer0_outputs(3723) <= inputs(125);
    layer0_outputs(3724) <= not((inputs(53)) and (inputs(202)));
    layer0_outputs(3725) <= not((inputs(4)) or (inputs(202)));
    layer0_outputs(3726) <= '0';
    layer0_outputs(3727) <= not((inputs(49)) and (inputs(86)));
    layer0_outputs(3728) <= not(inputs(150));
    layer0_outputs(3729) <= inputs(246);
    layer0_outputs(3730) <= (inputs(7)) or (inputs(106));
    layer0_outputs(3731) <= not(inputs(55)) or (inputs(103));
    layer0_outputs(3732) <= '0';
    layer0_outputs(3733) <= (inputs(224)) or (inputs(105));
    layer0_outputs(3734) <= not(inputs(230)) or (inputs(165));
    layer0_outputs(3735) <= inputs(198);
    layer0_outputs(3736) <= not(inputs(246));
    layer0_outputs(3737) <= inputs(18);
    layer0_outputs(3738) <= (inputs(91)) or (inputs(80));
    layer0_outputs(3739) <= not(inputs(231));
    layer0_outputs(3740) <= (inputs(113)) or (inputs(155));
    layer0_outputs(3741) <= inputs(15);
    layer0_outputs(3742) <= not((inputs(192)) or (inputs(31)));
    layer0_outputs(3743) <= (inputs(3)) and (inputs(22));
    layer0_outputs(3744) <= not(inputs(148));
    layer0_outputs(3745) <= (inputs(178)) xor (inputs(53));
    layer0_outputs(3746) <= not(inputs(100)) or (inputs(26));
    layer0_outputs(3747) <= inputs(249);
    layer0_outputs(3748) <= (inputs(22)) and not (inputs(147));
    layer0_outputs(3749) <= not((inputs(130)) or (inputs(193)));
    layer0_outputs(3750) <= not(inputs(141));
    layer0_outputs(3751) <= not((inputs(245)) or (inputs(191)));
    layer0_outputs(3752) <= not(inputs(152));
    layer0_outputs(3753) <= not(inputs(87));
    layer0_outputs(3754) <= (inputs(78)) or (inputs(251));
    layer0_outputs(3755) <= inputs(44);
    layer0_outputs(3756) <= not((inputs(44)) or (inputs(134)));
    layer0_outputs(3757) <= (inputs(29)) or (inputs(149));
    layer0_outputs(3758) <= (inputs(187)) or (inputs(197));
    layer0_outputs(3759) <= not(inputs(238));
    layer0_outputs(3760) <= not((inputs(170)) or (inputs(71)));
    layer0_outputs(3761) <= (inputs(99)) or (inputs(114));
    layer0_outputs(3762) <= not((inputs(152)) xor (inputs(105)));
    layer0_outputs(3763) <= (inputs(34)) and not (inputs(226));
    layer0_outputs(3764) <= (inputs(42)) and not (inputs(203));
    layer0_outputs(3765) <= inputs(126);
    layer0_outputs(3766) <= (inputs(101)) and not (inputs(19));
    layer0_outputs(3767) <= not(inputs(34)) or (inputs(250));
    layer0_outputs(3768) <= (inputs(109)) and (inputs(6));
    layer0_outputs(3769) <= not((inputs(69)) or (inputs(18)));
    layer0_outputs(3770) <= '0';
    layer0_outputs(3771) <= '0';
    layer0_outputs(3772) <= not(inputs(161));
    layer0_outputs(3773) <= '1';
    layer0_outputs(3774) <= (inputs(57)) or (inputs(157));
    layer0_outputs(3775) <= (inputs(190)) and (inputs(73));
    layer0_outputs(3776) <= (inputs(61)) xor (inputs(149));
    layer0_outputs(3777) <= inputs(152);
    layer0_outputs(3778) <= '1';
    layer0_outputs(3779) <= (inputs(219)) or (inputs(205));
    layer0_outputs(3780) <= not(inputs(222));
    layer0_outputs(3781) <= (inputs(60)) xor (inputs(0));
    layer0_outputs(3782) <= '1';
    layer0_outputs(3783) <= (inputs(254)) or (inputs(104));
    layer0_outputs(3784) <= (inputs(17)) and not (inputs(10));
    layer0_outputs(3785) <= not((inputs(175)) or (inputs(227)));
    layer0_outputs(3786) <= not(inputs(212));
    layer0_outputs(3787) <= not((inputs(247)) or (inputs(141)));
    layer0_outputs(3788) <= (inputs(54)) xor (inputs(4));
    layer0_outputs(3789) <= not(inputs(43)) or (inputs(2));
    layer0_outputs(3790) <= inputs(154);
    layer0_outputs(3791) <= inputs(158);
    layer0_outputs(3792) <= not(inputs(71)) or (inputs(223));
    layer0_outputs(3793) <= not((inputs(167)) or (inputs(37)));
    layer0_outputs(3794) <= inputs(227);
    layer0_outputs(3795) <= inputs(59);
    layer0_outputs(3796) <= inputs(88);
    layer0_outputs(3797) <= '1';
    layer0_outputs(3798) <= not((inputs(112)) xor (inputs(44)));
    layer0_outputs(3799) <= (inputs(97)) and not (inputs(153));
    layer0_outputs(3800) <= '1';
    layer0_outputs(3801) <= not(inputs(75));
    layer0_outputs(3802) <= (inputs(167)) and not (inputs(80));
    layer0_outputs(3803) <= '1';
    layer0_outputs(3804) <= not(inputs(133)) or (inputs(254));
    layer0_outputs(3805) <= not(inputs(168));
    layer0_outputs(3806) <= not(inputs(16));
    layer0_outputs(3807) <= inputs(218);
    layer0_outputs(3808) <= '1';
    layer0_outputs(3809) <= '1';
    layer0_outputs(3810) <= not(inputs(25)) or (inputs(113));
    layer0_outputs(3811) <= (inputs(230)) and not (inputs(0));
    layer0_outputs(3812) <= '1';
    layer0_outputs(3813) <= not((inputs(78)) or (inputs(88)));
    layer0_outputs(3814) <= not((inputs(220)) xor (inputs(46)));
    layer0_outputs(3815) <= not(inputs(123)) or (inputs(174));
    layer0_outputs(3816) <= (inputs(228)) or (inputs(18));
    layer0_outputs(3817) <= not(inputs(230));
    layer0_outputs(3818) <= '1';
    layer0_outputs(3819) <= (inputs(148)) or (inputs(184));
    layer0_outputs(3820) <= '1';
    layer0_outputs(3821) <= not(inputs(26));
    layer0_outputs(3822) <= (inputs(35)) or (inputs(213));
    layer0_outputs(3823) <= not(inputs(42));
    layer0_outputs(3824) <= inputs(247);
    layer0_outputs(3825) <= inputs(177);
    layer0_outputs(3826) <= (inputs(242)) and not (inputs(108));
    layer0_outputs(3827) <= not(inputs(86));
    layer0_outputs(3828) <= (inputs(86)) and not (inputs(77));
    layer0_outputs(3829) <= (inputs(113)) or (inputs(82));
    layer0_outputs(3830) <= not(inputs(151));
    layer0_outputs(3831) <= inputs(52);
    layer0_outputs(3832) <= inputs(122);
    layer0_outputs(3833) <= not(inputs(178));
    layer0_outputs(3834) <= not(inputs(171)) or (inputs(151));
    layer0_outputs(3835) <= not((inputs(228)) and (inputs(61)));
    layer0_outputs(3836) <= (inputs(128)) and not (inputs(153));
    layer0_outputs(3837) <= not((inputs(68)) or (inputs(44)));
    layer0_outputs(3838) <= (inputs(45)) or (inputs(94));
    layer0_outputs(3839) <= not((inputs(114)) or (inputs(107)));
    layer0_outputs(3840) <= '0';
    layer0_outputs(3841) <= inputs(195);
    layer0_outputs(3842) <= '0';
    layer0_outputs(3843) <= not((inputs(18)) xor (inputs(109)));
    layer0_outputs(3844) <= not(inputs(214));
    layer0_outputs(3845) <= not(inputs(187));
    layer0_outputs(3846) <= inputs(38);
    layer0_outputs(3847) <= (inputs(102)) or (inputs(146));
    layer0_outputs(3848) <= not(inputs(246));
    layer0_outputs(3849) <= not((inputs(61)) or (inputs(126)));
    layer0_outputs(3850) <= (inputs(222)) and not (inputs(49));
    layer0_outputs(3851) <= inputs(170);
    layer0_outputs(3852) <= (inputs(186)) or (inputs(46));
    layer0_outputs(3853) <= not(inputs(60));
    layer0_outputs(3854) <= '1';
    layer0_outputs(3855) <= not(inputs(81)) or (inputs(124));
    layer0_outputs(3856) <= not((inputs(83)) or (inputs(246)));
    layer0_outputs(3857) <= not((inputs(160)) and (inputs(5)));
    layer0_outputs(3858) <= (inputs(169)) xor (inputs(224));
    layer0_outputs(3859) <= not(inputs(90));
    layer0_outputs(3860) <= not((inputs(255)) or (inputs(166)));
    layer0_outputs(3861) <= inputs(22);
    layer0_outputs(3862) <= not((inputs(163)) or (inputs(236)));
    layer0_outputs(3863) <= not(inputs(120)) or (inputs(119));
    layer0_outputs(3864) <= (inputs(250)) or (inputs(127));
    layer0_outputs(3865) <= (inputs(147)) or (inputs(160));
    layer0_outputs(3866) <= not(inputs(118)) or (inputs(243));
    layer0_outputs(3867) <= (inputs(58)) and not (inputs(145));
    layer0_outputs(3868) <= (inputs(203)) xor (inputs(236));
    layer0_outputs(3869) <= inputs(150);
    layer0_outputs(3870) <= not((inputs(222)) or (inputs(154)));
    layer0_outputs(3871) <= (inputs(81)) and not (inputs(66));
    layer0_outputs(3872) <= not((inputs(143)) or (inputs(234)));
    layer0_outputs(3873) <= not(inputs(93));
    layer0_outputs(3874) <= inputs(59);
    layer0_outputs(3875) <= inputs(89);
    layer0_outputs(3876) <= (inputs(202)) xor (inputs(144));
    layer0_outputs(3877) <= (inputs(24)) xor (inputs(39));
    layer0_outputs(3878) <= not((inputs(164)) or (inputs(148)));
    layer0_outputs(3879) <= (inputs(215)) and not (inputs(246));
    layer0_outputs(3880) <= not(inputs(92));
    layer0_outputs(3881) <= not(inputs(42)) or (inputs(151));
    layer0_outputs(3882) <= not((inputs(58)) or (inputs(142)));
    layer0_outputs(3883) <= not(inputs(246)) or (inputs(17));
    layer0_outputs(3884) <= inputs(82);
    layer0_outputs(3885) <= '0';
    layer0_outputs(3886) <= not(inputs(73));
    layer0_outputs(3887) <= inputs(49);
    layer0_outputs(3888) <= '1';
    layer0_outputs(3889) <= not((inputs(91)) or (inputs(163)));
    layer0_outputs(3890) <= not((inputs(223)) or (inputs(204)));
    layer0_outputs(3891) <= (inputs(244)) or (inputs(156));
    layer0_outputs(3892) <= '1';
    layer0_outputs(3893) <= not((inputs(147)) xor (inputs(118)));
    layer0_outputs(3894) <= inputs(5);
    layer0_outputs(3895) <= not(inputs(159)) or (inputs(47));
    layer0_outputs(3896) <= not((inputs(37)) or (inputs(53)));
    layer0_outputs(3897) <= inputs(163);
    layer0_outputs(3898) <= (inputs(153)) xor (inputs(105));
    layer0_outputs(3899) <= (inputs(203)) and not (inputs(15));
    layer0_outputs(3900) <= (inputs(30)) or (inputs(88));
    layer0_outputs(3901) <= not(inputs(120));
    layer0_outputs(3902) <= '1';
    layer0_outputs(3903) <= not(inputs(64)) or (inputs(0));
    layer0_outputs(3904) <= not(inputs(191));
    layer0_outputs(3905) <= inputs(121);
    layer0_outputs(3906) <= inputs(254);
    layer0_outputs(3907) <= not((inputs(123)) or (inputs(129)));
    layer0_outputs(3908) <= not(inputs(125)) or (inputs(253));
    layer0_outputs(3909) <= not((inputs(188)) xor (inputs(238)));
    layer0_outputs(3910) <= not(inputs(68));
    layer0_outputs(3911) <= not(inputs(52));
    layer0_outputs(3912) <= (inputs(63)) and not (inputs(145));
    layer0_outputs(3913) <= (inputs(41)) and (inputs(22));
    layer0_outputs(3914) <= not(inputs(136)) or (inputs(75));
    layer0_outputs(3915) <= (inputs(229)) and not (inputs(104));
    layer0_outputs(3916) <= inputs(210);
    layer0_outputs(3917) <= inputs(147);
    layer0_outputs(3918) <= (inputs(203)) or (inputs(30));
    layer0_outputs(3919) <= not(inputs(216));
    layer0_outputs(3920) <= not(inputs(87)) or (inputs(235));
    layer0_outputs(3921) <= (inputs(75)) or (inputs(252));
    layer0_outputs(3922) <= (inputs(226)) and not (inputs(109));
    layer0_outputs(3923) <= not((inputs(152)) or (inputs(85)));
    layer0_outputs(3924) <= '0';
    layer0_outputs(3925) <= (inputs(135)) or (inputs(115));
    layer0_outputs(3926) <= not(inputs(229));
    layer0_outputs(3927) <= inputs(231);
    layer0_outputs(3928) <= (inputs(109)) and (inputs(85));
    layer0_outputs(3929) <= (inputs(204)) or (inputs(175));
    layer0_outputs(3930) <= not(inputs(164));
    layer0_outputs(3931) <= not((inputs(88)) and (inputs(137)));
    layer0_outputs(3932) <= not((inputs(110)) and (inputs(199)));
    layer0_outputs(3933) <= inputs(103);
    layer0_outputs(3934) <= (inputs(45)) and not (inputs(226));
    layer0_outputs(3935) <= inputs(120);
    layer0_outputs(3936) <= (inputs(114)) xor (inputs(173));
    layer0_outputs(3937) <= not((inputs(196)) xor (inputs(177)));
    layer0_outputs(3938) <= inputs(201);
    layer0_outputs(3939) <= not(inputs(76));
    layer0_outputs(3940) <= '0';
    layer0_outputs(3941) <= inputs(47);
    layer0_outputs(3942) <= not(inputs(80));
    layer0_outputs(3943) <= not((inputs(65)) and (inputs(176)));
    layer0_outputs(3944) <= (inputs(45)) or (inputs(61));
    layer0_outputs(3945) <= not((inputs(57)) or (inputs(176)));
    layer0_outputs(3946) <= (inputs(210)) or (inputs(183));
    layer0_outputs(3947) <= (inputs(40)) and not (inputs(13));
    layer0_outputs(3948) <= not((inputs(33)) xor (inputs(180)));
    layer0_outputs(3949) <= not((inputs(49)) and (inputs(124)));
    layer0_outputs(3950) <= '1';
    layer0_outputs(3951) <= not(inputs(151));
    layer0_outputs(3952) <= (inputs(6)) or (inputs(127));
    layer0_outputs(3953) <= (inputs(139)) and not (inputs(34));
    layer0_outputs(3954) <= not((inputs(47)) or (inputs(4)));
    layer0_outputs(3955) <= not(inputs(4));
    layer0_outputs(3956) <= inputs(37);
    layer0_outputs(3957) <= (inputs(10)) and not (inputs(153));
    layer0_outputs(3958) <= (inputs(136)) or (inputs(167));
    layer0_outputs(3959) <= not(inputs(73)) or (inputs(131));
    layer0_outputs(3960) <= not((inputs(251)) or (inputs(137)));
    layer0_outputs(3961) <= '0';
    layer0_outputs(3962) <= (inputs(36)) or (inputs(114));
    layer0_outputs(3963) <= not(inputs(237));
    layer0_outputs(3964) <= (inputs(40)) or (inputs(160));
    layer0_outputs(3965) <= not(inputs(227));
    layer0_outputs(3966) <= not(inputs(0));
    layer0_outputs(3967) <= inputs(99);
    layer0_outputs(3968) <= not((inputs(169)) or (inputs(253)));
    layer0_outputs(3969) <= (inputs(151)) and not (inputs(13));
    layer0_outputs(3970) <= not(inputs(207)) or (inputs(56));
    layer0_outputs(3971) <= not((inputs(227)) or (inputs(48)));
    layer0_outputs(3972) <= not((inputs(159)) or (inputs(98)));
    layer0_outputs(3973) <= inputs(49);
    layer0_outputs(3974) <= not(inputs(16));
    layer0_outputs(3975) <= not(inputs(24));
    layer0_outputs(3976) <= (inputs(205)) and not (inputs(39));
    layer0_outputs(3977) <= not((inputs(208)) or (inputs(213)));
    layer0_outputs(3978) <= (inputs(15)) xor (inputs(111));
    layer0_outputs(3979) <= (inputs(211)) or (inputs(227));
    layer0_outputs(3980) <= (inputs(72)) or (inputs(79));
    layer0_outputs(3981) <= (inputs(26)) xor (inputs(148));
    layer0_outputs(3982) <= not(inputs(92));
    layer0_outputs(3983) <= not((inputs(51)) and (inputs(142)));
    layer0_outputs(3984) <= (inputs(83)) or (inputs(69));
    layer0_outputs(3985) <= (inputs(77)) or (inputs(100));
    layer0_outputs(3986) <= not(inputs(147)) or (inputs(29));
    layer0_outputs(3987) <= not(inputs(132));
    layer0_outputs(3988) <= (inputs(213)) and not (inputs(144));
    layer0_outputs(3989) <= not(inputs(214));
    layer0_outputs(3990) <= (inputs(231)) and not (inputs(60));
    layer0_outputs(3991) <= (inputs(247)) xor (inputs(249));
    layer0_outputs(3992) <= not((inputs(105)) or (inputs(135)));
    layer0_outputs(3993) <= (inputs(56)) or (inputs(237));
    layer0_outputs(3994) <= (inputs(16)) and not (inputs(78));
    layer0_outputs(3995) <= not(inputs(25)) or (inputs(99));
    layer0_outputs(3996) <= not((inputs(228)) or (inputs(245)));
    layer0_outputs(3997) <= not(inputs(4));
    layer0_outputs(3998) <= '1';
    layer0_outputs(3999) <= (inputs(246)) and not (inputs(172));
    layer0_outputs(4000) <= not(inputs(60));
    layer0_outputs(4001) <= (inputs(132)) or (inputs(220));
    layer0_outputs(4002) <= not(inputs(12)) or (inputs(109));
    layer0_outputs(4003) <= inputs(224);
    layer0_outputs(4004) <= not(inputs(118));
    layer0_outputs(4005) <= inputs(73);
    layer0_outputs(4006) <= inputs(129);
    layer0_outputs(4007) <= not(inputs(182));
    layer0_outputs(4008) <= (inputs(196)) or (inputs(190));
    layer0_outputs(4009) <= not((inputs(254)) xor (inputs(135)));
    layer0_outputs(4010) <= not((inputs(224)) or (inputs(47)));
    layer0_outputs(4011) <= (inputs(152)) and not (inputs(253));
    layer0_outputs(4012) <= (inputs(133)) and not (inputs(245));
    layer0_outputs(4013) <= inputs(68);
    layer0_outputs(4014) <= (inputs(129)) or (inputs(215));
    layer0_outputs(4015) <= '0';
    layer0_outputs(4016) <= not(inputs(139)) or (inputs(193));
    layer0_outputs(4017) <= not(inputs(255)) or (inputs(171));
    layer0_outputs(4018) <= (inputs(91)) and (inputs(57));
    layer0_outputs(4019) <= not((inputs(204)) xor (inputs(172)));
    layer0_outputs(4020) <= (inputs(111)) xor (inputs(199));
    layer0_outputs(4021) <= not((inputs(49)) or (inputs(99)));
    layer0_outputs(4022) <= (inputs(180)) or (inputs(90));
    layer0_outputs(4023) <= inputs(120);
    layer0_outputs(4024) <= (inputs(163)) or (inputs(22));
    layer0_outputs(4025) <= (inputs(191)) or (inputs(15));
    layer0_outputs(4026) <= not(inputs(108));
    layer0_outputs(4027) <= (inputs(120)) and not (inputs(99));
    layer0_outputs(4028) <= (inputs(233)) or (inputs(225));
    layer0_outputs(4029) <= (inputs(154)) and not (inputs(73));
    layer0_outputs(4030) <= inputs(47);
    layer0_outputs(4031) <= not(inputs(157));
    layer0_outputs(4032) <= (inputs(178)) xor (inputs(37));
    layer0_outputs(4033) <= not(inputs(31));
    layer0_outputs(4034) <= (inputs(109)) or (inputs(67));
    layer0_outputs(4035) <= (inputs(160)) and not (inputs(200));
    layer0_outputs(4036) <= not((inputs(249)) and (inputs(62)));
    layer0_outputs(4037) <= not(inputs(197));
    layer0_outputs(4038) <= (inputs(80)) or (inputs(38));
    layer0_outputs(4039) <= (inputs(216)) and not (inputs(121));
    layer0_outputs(4040) <= not(inputs(201));
    layer0_outputs(4041) <= (inputs(86)) or (inputs(162));
    layer0_outputs(4042) <= inputs(209);
    layer0_outputs(4043) <= (inputs(143)) and (inputs(252));
    layer0_outputs(4044) <= not(inputs(55));
    layer0_outputs(4045) <= not(inputs(225));
    layer0_outputs(4046) <= not(inputs(123));
    layer0_outputs(4047) <= not(inputs(251)) or (inputs(38));
    layer0_outputs(4048) <= not(inputs(221)) or (inputs(249));
    layer0_outputs(4049) <= (inputs(248)) or (inputs(176));
    layer0_outputs(4050) <= (inputs(151)) and not (inputs(180));
    layer0_outputs(4051) <= (inputs(113)) and (inputs(25));
    layer0_outputs(4052) <= (inputs(13)) or (inputs(141));
    layer0_outputs(4053) <= not((inputs(146)) or (inputs(140)));
    layer0_outputs(4054) <= inputs(210);
    layer0_outputs(4055) <= inputs(252);
    layer0_outputs(4056) <= not(inputs(234)) or (inputs(51));
    layer0_outputs(4057) <= inputs(195);
    layer0_outputs(4058) <= not((inputs(189)) or (inputs(204)));
    layer0_outputs(4059) <= '0';
    layer0_outputs(4060) <= '0';
    layer0_outputs(4061) <= inputs(173);
    layer0_outputs(4062) <= not((inputs(184)) or (inputs(44)));
    layer0_outputs(4063) <= not((inputs(72)) and (inputs(35)));
    layer0_outputs(4064) <= not((inputs(66)) or (inputs(64)));
    layer0_outputs(4065) <= inputs(164);
    layer0_outputs(4066) <= not(inputs(147));
    layer0_outputs(4067) <= (inputs(62)) or (inputs(164));
    layer0_outputs(4068) <= (inputs(56)) or (inputs(10));
    layer0_outputs(4069) <= (inputs(164)) or (inputs(98));
    layer0_outputs(4070) <= (inputs(157)) or (inputs(251));
    layer0_outputs(4071) <= inputs(153);
    layer0_outputs(4072) <= '1';
    layer0_outputs(4073) <= '0';
    layer0_outputs(4074) <= not((inputs(220)) or (inputs(160)));
    layer0_outputs(4075) <= not(inputs(73));
    layer0_outputs(4076) <= not(inputs(114));
    layer0_outputs(4077) <= not((inputs(147)) xor (inputs(4)));
    layer0_outputs(4078) <= inputs(134);
    layer0_outputs(4079) <= not(inputs(97)) or (inputs(240));
    layer0_outputs(4080) <= inputs(202);
    layer0_outputs(4081) <= not(inputs(181));
    layer0_outputs(4082) <= not(inputs(18));
    layer0_outputs(4083) <= not((inputs(31)) or (inputs(144)));
    layer0_outputs(4084) <= '0';
    layer0_outputs(4085) <= inputs(122);
    layer0_outputs(4086) <= (inputs(252)) and (inputs(155));
    layer0_outputs(4087) <= not((inputs(13)) xor (inputs(45)));
    layer0_outputs(4088) <= not(inputs(128));
    layer0_outputs(4089) <= not(inputs(201)) or (inputs(97));
    layer0_outputs(4090) <= inputs(3);
    layer0_outputs(4091) <= (inputs(161)) and not (inputs(61));
    layer0_outputs(4092) <= not(inputs(250)) or (inputs(100));
    layer0_outputs(4093) <= inputs(125);
    layer0_outputs(4094) <= not(inputs(34));
    layer0_outputs(4095) <= not(inputs(217));
    layer0_outputs(4096) <= not(inputs(86));
    layer0_outputs(4097) <= '0';
    layer0_outputs(4098) <= (inputs(119)) or (inputs(114));
    layer0_outputs(4099) <= not(inputs(70));
    layer0_outputs(4100) <= not((inputs(7)) or (inputs(203)));
    layer0_outputs(4101) <= '0';
    layer0_outputs(4102) <= not((inputs(239)) or (inputs(210)));
    layer0_outputs(4103) <= '0';
    layer0_outputs(4104) <= (inputs(22)) and (inputs(181));
    layer0_outputs(4105) <= not((inputs(219)) or (inputs(81)));
    layer0_outputs(4106) <= inputs(214);
    layer0_outputs(4107) <= not((inputs(169)) and (inputs(123)));
    layer0_outputs(4108) <= (inputs(91)) or (inputs(13));
    layer0_outputs(4109) <= not(inputs(158));
    layer0_outputs(4110) <= not(inputs(109));
    layer0_outputs(4111) <= (inputs(220)) or (inputs(117));
    layer0_outputs(4112) <= not(inputs(86));
    layer0_outputs(4113) <= not((inputs(183)) or (inputs(224)));
    layer0_outputs(4114) <= (inputs(191)) xor (inputs(188));
    layer0_outputs(4115) <= inputs(201);
    layer0_outputs(4116) <= not((inputs(233)) or (inputs(47)));
    layer0_outputs(4117) <= not(inputs(162)) or (inputs(235));
    layer0_outputs(4118) <= not(inputs(59)) or (inputs(17));
    layer0_outputs(4119) <= inputs(21);
    layer0_outputs(4120) <= not(inputs(178));
    layer0_outputs(4121) <= (inputs(166)) and not (inputs(12));
    layer0_outputs(4122) <= (inputs(231)) and (inputs(228));
    layer0_outputs(4123) <= not(inputs(181));
    layer0_outputs(4124) <= not(inputs(161));
    layer0_outputs(4125) <= (inputs(129)) or (inputs(164));
    layer0_outputs(4126) <= (inputs(79)) and not (inputs(109));
    layer0_outputs(4127) <= not(inputs(120)) or (inputs(207));
    layer0_outputs(4128) <= not(inputs(88)) or (inputs(78));
    layer0_outputs(4129) <= (inputs(239)) or (inputs(177));
    layer0_outputs(4130) <= inputs(231);
    layer0_outputs(4131) <= not((inputs(65)) or (inputs(186)));
    layer0_outputs(4132) <= not((inputs(247)) or (inputs(11)));
    layer0_outputs(4133) <= inputs(17);
    layer0_outputs(4134) <= not(inputs(18)) or (inputs(120));
    layer0_outputs(4135) <= not(inputs(196));
    layer0_outputs(4136) <= inputs(197);
    layer0_outputs(4137) <= not((inputs(156)) or (inputs(88)));
    layer0_outputs(4138) <= not((inputs(171)) or (inputs(85)));
    layer0_outputs(4139) <= not(inputs(120));
    layer0_outputs(4140) <= not(inputs(166)) or (inputs(108));
    layer0_outputs(4141) <= (inputs(95)) and not (inputs(196));
    layer0_outputs(4142) <= not(inputs(44)) or (inputs(236));
    layer0_outputs(4143) <= (inputs(40)) or (inputs(47));
    layer0_outputs(4144) <= (inputs(87)) and not (inputs(207));
    layer0_outputs(4145) <= not((inputs(176)) or (inputs(70)));
    layer0_outputs(4146) <= (inputs(249)) and not (inputs(165));
    layer0_outputs(4147) <= not(inputs(232));
    layer0_outputs(4148) <= (inputs(46)) and not (inputs(223));
    layer0_outputs(4149) <= not(inputs(204));
    layer0_outputs(4150) <= not(inputs(227));
    layer0_outputs(4151) <= not(inputs(180));
    layer0_outputs(4152) <= (inputs(89)) xor (inputs(26));
    layer0_outputs(4153) <= not((inputs(33)) and (inputs(216)));
    layer0_outputs(4154) <= (inputs(91)) or (inputs(178));
    layer0_outputs(4155) <= '1';
    layer0_outputs(4156) <= not(inputs(230)) or (inputs(50));
    layer0_outputs(4157) <= not((inputs(117)) xor (inputs(66)));
    layer0_outputs(4158) <= not(inputs(88)) or (inputs(190));
    layer0_outputs(4159) <= inputs(162);
    layer0_outputs(4160) <= not(inputs(52)) or (inputs(216));
    layer0_outputs(4161) <= (inputs(153)) and not (inputs(44));
    layer0_outputs(4162) <= not((inputs(55)) or (inputs(102)));
    layer0_outputs(4163) <= not(inputs(100)) or (inputs(207));
    layer0_outputs(4164) <= not((inputs(28)) or (inputs(50)));
    layer0_outputs(4165) <= not(inputs(25));
    layer0_outputs(4166) <= not(inputs(204));
    layer0_outputs(4167) <= (inputs(125)) xor (inputs(191));
    layer0_outputs(4168) <= not(inputs(253));
    layer0_outputs(4169) <= inputs(105);
    layer0_outputs(4170) <= not((inputs(26)) xor (inputs(159)));
    layer0_outputs(4171) <= (inputs(115)) and not (inputs(85));
    layer0_outputs(4172) <= (inputs(49)) or (inputs(41));
    layer0_outputs(4173) <= (inputs(135)) and not (inputs(7));
    layer0_outputs(4174) <= not(inputs(166));
    layer0_outputs(4175) <= (inputs(135)) or (inputs(4));
    layer0_outputs(4176) <= not(inputs(184));
    layer0_outputs(4177) <= (inputs(166)) and not (inputs(144));
    layer0_outputs(4178) <= (inputs(141)) xor (inputs(146));
    layer0_outputs(4179) <= not((inputs(250)) xor (inputs(186)));
    layer0_outputs(4180) <= not((inputs(206)) or (inputs(226)));
    layer0_outputs(4181) <= not(inputs(95));
    layer0_outputs(4182) <= not(inputs(135));
    layer0_outputs(4183) <= (inputs(239)) and not (inputs(243));
    layer0_outputs(4184) <= not(inputs(131));
    layer0_outputs(4185) <= not((inputs(96)) or (inputs(144)));
    layer0_outputs(4186) <= not((inputs(95)) and (inputs(132)));
    layer0_outputs(4187) <= not(inputs(43));
    layer0_outputs(4188) <= inputs(233);
    layer0_outputs(4189) <= inputs(122);
    layer0_outputs(4190) <= not(inputs(229));
    layer0_outputs(4191) <= inputs(21);
    layer0_outputs(4192) <= (inputs(109)) or (inputs(6));
    layer0_outputs(4193) <= (inputs(254)) or (inputs(237));
    layer0_outputs(4194) <= not(inputs(86));
    layer0_outputs(4195) <= '0';
    layer0_outputs(4196) <= (inputs(36)) and not (inputs(235));
    layer0_outputs(4197) <= not(inputs(126));
    layer0_outputs(4198) <= inputs(59);
    layer0_outputs(4199) <= not(inputs(117)) or (inputs(255));
    layer0_outputs(4200) <= '0';
    layer0_outputs(4201) <= not(inputs(32));
    layer0_outputs(4202) <= (inputs(100)) or (inputs(13));
    layer0_outputs(4203) <= (inputs(58)) or (inputs(99));
    layer0_outputs(4204) <= not((inputs(69)) xor (inputs(51)));
    layer0_outputs(4205) <= inputs(197);
    layer0_outputs(4206) <= not(inputs(159));
    layer0_outputs(4207) <= (inputs(177)) and not (inputs(78));
    layer0_outputs(4208) <= not((inputs(208)) or (inputs(110)));
    layer0_outputs(4209) <= (inputs(3)) and not (inputs(217));
    layer0_outputs(4210) <= not(inputs(206)) or (inputs(128));
    layer0_outputs(4211) <= not(inputs(56));
    layer0_outputs(4212) <= (inputs(159)) xor (inputs(86));
    layer0_outputs(4213) <= (inputs(163)) or (inputs(176));
    layer0_outputs(4214) <= inputs(52);
    layer0_outputs(4215) <= not(inputs(192)) or (inputs(119));
    layer0_outputs(4216) <= not(inputs(151));
    layer0_outputs(4217) <= '1';
    layer0_outputs(4218) <= (inputs(25)) or (inputs(54));
    layer0_outputs(4219) <= inputs(162);
    layer0_outputs(4220) <= not(inputs(208));
    layer0_outputs(4221) <= not((inputs(110)) or (inputs(60)));
    layer0_outputs(4222) <= not(inputs(238));
    layer0_outputs(4223) <= (inputs(190)) or (inputs(65));
    layer0_outputs(4224) <= not(inputs(85));
    layer0_outputs(4225) <= (inputs(222)) or (inputs(159));
    layer0_outputs(4226) <= (inputs(70)) xor (inputs(82));
    layer0_outputs(4227) <= (inputs(233)) and not (inputs(225));
    layer0_outputs(4228) <= (inputs(35)) xor (inputs(80));
    layer0_outputs(4229) <= not((inputs(177)) or (inputs(9)));
    layer0_outputs(4230) <= not((inputs(152)) or (inputs(102)));
    layer0_outputs(4231) <= inputs(119);
    layer0_outputs(4232) <= inputs(119);
    layer0_outputs(4233) <= not(inputs(79));
    layer0_outputs(4234) <= inputs(197);
    layer0_outputs(4235) <= not((inputs(98)) or (inputs(89)));
    layer0_outputs(4236) <= not(inputs(88));
    layer0_outputs(4237) <= (inputs(23)) xor (inputs(223));
    layer0_outputs(4238) <= not(inputs(93));
    layer0_outputs(4239) <= not(inputs(28));
    layer0_outputs(4240) <= (inputs(20)) and not (inputs(254));
    layer0_outputs(4241) <= inputs(43);
    layer0_outputs(4242) <= inputs(69);
    layer0_outputs(4243) <= (inputs(25)) or (inputs(53));
    layer0_outputs(4244) <= not(inputs(165));
    layer0_outputs(4245) <= not(inputs(153)) or (inputs(209));
    layer0_outputs(4246) <= (inputs(10)) or (inputs(248));
    layer0_outputs(4247) <= '1';
    layer0_outputs(4248) <= inputs(115);
    layer0_outputs(4249) <= (inputs(181)) and not (inputs(192));
    layer0_outputs(4250) <= inputs(63);
    layer0_outputs(4251) <= not(inputs(128));
    layer0_outputs(4252) <= not((inputs(33)) or (inputs(122)));
    layer0_outputs(4253) <= (inputs(214)) and not (inputs(35));
    layer0_outputs(4254) <= (inputs(191)) or (inputs(156));
    layer0_outputs(4255) <= not((inputs(160)) or (inputs(168)));
    layer0_outputs(4256) <= not(inputs(26));
    layer0_outputs(4257) <= inputs(18);
    layer0_outputs(4258) <= inputs(202);
    layer0_outputs(4259) <= (inputs(221)) or (inputs(50));
    layer0_outputs(4260) <= not(inputs(21));
    layer0_outputs(4261) <= inputs(118);
    layer0_outputs(4262) <= not(inputs(235)) or (inputs(173));
    layer0_outputs(4263) <= not(inputs(183));
    layer0_outputs(4264) <= not((inputs(144)) or (inputs(160)));
    layer0_outputs(4265) <= not(inputs(85));
    layer0_outputs(4266) <= not(inputs(209));
    layer0_outputs(4267) <= not(inputs(116)) or (inputs(236));
    layer0_outputs(4268) <= not((inputs(77)) or (inputs(233)));
    layer0_outputs(4269) <= not((inputs(193)) or (inputs(5)));
    layer0_outputs(4270) <= not(inputs(8)) or (inputs(227));
    layer0_outputs(4271) <= not(inputs(204));
    layer0_outputs(4272) <= not(inputs(40));
    layer0_outputs(4273) <= not(inputs(111)) or (inputs(137));
    layer0_outputs(4274) <= not(inputs(115));
    layer0_outputs(4275) <= not(inputs(123));
    layer0_outputs(4276) <= inputs(97);
    layer0_outputs(4277) <= inputs(91);
    layer0_outputs(4278) <= inputs(51);
    layer0_outputs(4279) <= not(inputs(218)) or (inputs(68));
    layer0_outputs(4280) <= not(inputs(102));
    layer0_outputs(4281) <= not((inputs(29)) or (inputs(194)));
    layer0_outputs(4282) <= (inputs(196)) and not (inputs(22));
    layer0_outputs(4283) <= (inputs(118)) and (inputs(71));
    layer0_outputs(4284) <= (inputs(35)) xor (inputs(65));
    layer0_outputs(4285) <= inputs(26);
    layer0_outputs(4286) <= not(inputs(28));
    layer0_outputs(4287) <= not(inputs(38));
    layer0_outputs(4288) <= (inputs(130)) and not (inputs(49));
    layer0_outputs(4289) <= not(inputs(94));
    layer0_outputs(4290) <= not(inputs(231));
    layer0_outputs(4291) <= (inputs(224)) and not (inputs(57));
    layer0_outputs(4292) <= not((inputs(175)) or (inputs(211)));
    layer0_outputs(4293) <= (inputs(144)) and not (inputs(242));
    layer0_outputs(4294) <= not((inputs(239)) xor (inputs(72)));
    layer0_outputs(4295) <= not(inputs(89));
    layer0_outputs(4296) <= not((inputs(97)) xor (inputs(143)));
    layer0_outputs(4297) <= (inputs(215)) and not (inputs(80));
    layer0_outputs(4298) <= not(inputs(21)) or (inputs(176));
    layer0_outputs(4299) <= inputs(72);
    layer0_outputs(4300) <= (inputs(160)) and not (inputs(194));
    layer0_outputs(4301) <= '1';
    layer0_outputs(4302) <= (inputs(226)) or (inputs(26));
    layer0_outputs(4303) <= not(inputs(51)) or (inputs(161));
    layer0_outputs(4304) <= (inputs(84)) and not (inputs(208));
    layer0_outputs(4305) <= not(inputs(212)) or (inputs(241));
    layer0_outputs(4306) <= not((inputs(119)) or (inputs(158)));
    layer0_outputs(4307) <= (inputs(145)) or (inputs(206));
    layer0_outputs(4308) <= inputs(205);
    layer0_outputs(4309) <= inputs(7);
    layer0_outputs(4310) <= inputs(201);
    layer0_outputs(4311) <= (inputs(63)) or (inputs(43));
    layer0_outputs(4312) <= not((inputs(149)) or (inputs(63)));
    layer0_outputs(4313) <= inputs(151);
    layer0_outputs(4314) <= not(inputs(196));
    layer0_outputs(4315) <= inputs(27);
    layer0_outputs(4316) <= inputs(141);
    layer0_outputs(4317) <= inputs(38);
    layer0_outputs(4318) <= (inputs(180)) xor (inputs(28));
    layer0_outputs(4319) <= not(inputs(64));
    layer0_outputs(4320) <= (inputs(128)) and (inputs(239));
    layer0_outputs(4321) <= (inputs(41)) and not (inputs(172));
    layer0_outputs(4322) <= inputs(93);
    layer0_outputs(4323) <= '0';
    layer0_outputs(4324) <= not(inputs(247)) or (inputs(61));
    layer0_outputs(4325) <= not(inputs(208));
    layer0_outputs(4326) <= inputs(187);
    layer0_outputs(4327) <= not(inputs(115)) or (inputs(180));
    layer0_outputs(4328) <= (inputs(153)) and not (inputs(102));
    layer0_outputs(4329) <= not(inputs(98));
    layer0_outputs(4330) <= (inputs(185)) and not (inputs(68));
    layer0_outputs(4331) <= not(inputs(251)) or (inputs(14));
    layer0_outputs(4332) <= inputs(159);
    layer0_outputs(4333) <= inputs(17);
    layer0_outputs(4334) <= (inputs(88)) and not (inputs(42));
    layer0_outputs(4335) <= inputs(106);
    layer0_outputs(4336) <= not(inputs(232));
    layer0_outputs(4337) <= (inputs(32)) and (inputs(51));
    layer0_outputs(4338) <= '1';
    layer0_outputs(4339) <= '0';
    layer0_outputs(4340) <= (inputs(176)) or (inputs(178));
    layer0_outputs(4341) <= not((inputs(130)) xor (inputs(100)));
    layer0_outputs(4342) <= not(inputs(164)) or (inputs(169));
    layer0_outputs(4343) <= not((inputs(16)) or (inputs(182)));
    layer0_outputs(4344) <= inputs(190);
    layer0_outputs(4345) <= not((inputs(195)) xor (inputs(197)));
    layer0_outputs(4346) <= (inputs(202)) and not (inputs(173));
    layer0_outputs(4347) <= not(inputs(2)) or (inputs(254));
    layer0_outputs(4348) <= not(inputs(47));
    layer0_outputs(4349) <= not(inputs(253));
    layer0_outputs(4350) <= inputs(49);
    layer0_outputs(4351) <= not((inputs(43)) and (inputs(231)));
    layer0_outputs(4352) <= not(inputs(247));
    layer0_outputs(4353) <= (inputs(154)) and (inputs(151));
    layer0_outputs(4354) <= not((inputs(111)) or (inputs(255)));
    layer0_outputs(4355) <= not(inputs(166));
    layer0_outputs(4356) <= inputs(147);
    layer0_outputs(4357) <= (inputs(8)) or (inputs(190));
    layer0_outputs(4358) <= not(inputs(85)) or (inputs(17));
    layer0_outputs(4359) <= not(inputs(163));
    layer0_outputs(4360) <= not((inputs(218)) or (inputs(202)));
    layer0_outputs(4361) <= (inputs(49)) or (inputs(232));
    layer0_outputs(4362) <= not((inputs(248)) and (inputs(144)));
    layer0_outputs(4363) <= not((inputs(228)) or (inputs(32)));
    layer0_outputs(4364) <= (inputs(175)) or (inputs(228));
    layer0_outputs(4365) <= inputs(166);
    layer0_outputs(4366) <= (inputs(136)) or (inputs(168));
    layer0_outputs(4367) <= not(inputs(60));
    layer0_outputs(4368) <= not(inputs(69)) or (inputs(92));
    layer0_outputs(4369) <= (inputs(6)) and not (inputs(172));
    layer0_outputs(4370) <= (inputs(35)) and not (inputs(127));
    layer0_outputs(4371) <= (inputs(73)) and not (inputs(52));
    layer0_outputs(4372) <= (inputs(1)) or (inputs(147));
    layer0_outputs(4373) <= not((inputs(194)) xor (inputs(19)));
    layer0_outputs(4374) <= inputs(76);
    layer0_outputs(4375) <= (inputs(5)) and not (inputs(99));
    layer0_outputs(4376) <= (inputs(228)) xor (inputs(2));
    layer0_outputs(4377) <= (inputs(211)) and not (inputs(114));
    layer0_outputs(4378) <= (inputs(91)) or (inputs(229));
    layer0_outputs(4379) <= (inputs(251)) or (inputs(147));
    layer0_outputs(4380) <= not(inputs(43)) or (inputs(201));
    layer0_outputs(4381) <= not((inputs(157)) or (inputs(132)));
    layer0_outputs(4382) <= not(inputs(19)) or (inputs(169));
    layer0_outputs(4383) <= '1';
    layer0_outputs(4384) <= inputs(100);
    layer0_outputs(4385) <= inputs(178);
    layer0_outputs(4386) <= not(inputs(128)) or (inputs(192));
    layer0_outputs(4387) <= not(inputs(81));
    layer0_outputs(4388) <= inputs(163);
    layer0_outputs(4389) <= (inputs(131)) xor (inputs(17));
    layer0_outputs(4390) <= inputs(171);
    layer0_outputs(4391) <= not(inputs(26));
    layer0_outputs(4392) <= not(inputs(46)) or (inputs(97));
    layer0_outputs(4393) <= (inputs(67)) or (inputs(185));
    layer0_outputs(4394) <= not((inputs(252)) xor (inputs(203)));
    layer0_outputs(4395) <= inputs(183);
    layer0_outputs(4396) <= (inputs(184)) or (inputs(197));
    layer0_outputs(4397) <= inputs(226);
    layer0_outputs(4398) <= not(inputs(230));
    layer0_outputs(4399) <= not(inputs(167));
    layer0_outputs(4400) <= not((inputs(58)) or (inputs(167)));
    layer0_outputs(4401) <= not((inputs(123)) or (inputs(95)));
    layer0_outputs(4402) <= inputs(151);
    layer0_outputs(4403) <= not(inputs(196)) or (inputs(175));
    layer0_outputs(4404) <= not((inputs(42)) and (inputs(249)));
    layer0_outputs(4405) <= not(inputs(249));
    layer0_outputs(4406) <= inputs(79);
    layer0_outputs(4407) <= inputs(50);
    layer0_outputs(4408) <= not((inputs(119)) or (inputs(97)));
    layer0_outputs(4409) <= not((inputs(155)) or (inputs(60)));
    layer0_outputs(4410) <= not(inputs(163));
    layer0_outputs(4411) <= inputs(21);
    layer0_outputs(4412) <= '0';
    layer0_outputs(4413) <= not(inputs(27));
    layer0_outputs(4414) <= (inputs(90)) and (inputs(225));
    layer0_outputs(4415) <= inputs(101);
    layer0_outputs(4416) <= (inputs(27)) or (inputs(167));
    layer0_outputs(4417) <= not(inputs(78));
    layer0_outputs(4418) <= (inputs(23)) or (inputs(51));
    layer0_outputs(4419) <= not((inputs(230)) and (inputs(171)));
    layer0_outputs(4420) <= (inputs(196)) and (inputs(37));
    layer0_outputs(4421) <= not((inputs(89)) or (inputs(35)));
    layer0_outputs(4422) <= inputs(202);
    layer0_outputs(4423) <= not(inputs(102)) or (inputs(150));
    layer0_outputs(4424) <= (inputs(19)) and (inputs(145));
    layer0_outputs(4425) <= '0';
    layer0_outputs(4426) <= (inputs(162)) or (inputs(85));
    layer0_outputs(4427) <= (inputs(43)) and not (inputs(13));
    layer0_outputs(4428) <= inputs(27);
    layer0_outputs(4429) <= not((inputs(46)) or (inputs(60)));
    layer0_outputs(4430) <= not((inputs(148)) xor (inputs(230)));
    layer0_outputs(4431) <= not((inputs(86)) or (inputs(101)));
    layer0_outputs(4432) <= not((inputs(184)) or (inputs(213)));
    layer0_outputs(4433) <= '1';
    layer0_outputs(4434) <= (inputs(19)) or (inputs(33));
    layer0_outputs(4435) <= not((inputs(254)) and (inputs(13)));
    layer0_outputs(4436) <= not((inputs(248)) xor (inputs(231)));
    layer0_outputs(4437) <= not((inputs(207)) or (inputs(108)));
    layer0_outputs(4438) <= not(inputs(72));
    layer0_outputs(4439) <= not(inputs(114)) or (inputs(238));
    layer0_outputs(4440) <= (inputs(188)) and not (inputs(101));
    layer0_outputs(4441) <= inputs(12);
    layer0_outputs(4442) <= inputs(135);
    layer0_outputs(4443) <= (inputs(50)) and (inputs(114));
    layer0_outputs(4444) <= (inputs(149)) and not (inputs(194));
    layer0_outputs(4445) <= (inputs(181)) and (inputs(0));
    layer0_outputs(4446) <= not(inputs(69)) or (inputs(30));
    layer0_outputs(4447) <= not((inputs(151)) or (inputs(119)));
    layer0_outputs(4448) <= not(inputs(136)) or (inputs(192));
    layer0_outputs(4449) <= (inputs(166)) or (inputs(133));
    layer0_outputs(4450) <= not(inputs(218));
    layer0_outputs(4451) <= (inputs(75)) and not (inputs(208));
    layer0_outputs(4452) <= '0';
    layer0_outputs(4453) <= not((inputs(2)) or (inputs(124)));
    layer0_outputs(4454) <= (inputs(57)) or (inputs(180));
    layer0_outputs(4455) <= not(inputs(167)) or (inputs(135));
    layer0_outputs(4456) <= inputs(237);
    layer0_outputs(4457) <= (inputs(37)) or (inputs(206));
    layer0_outputs(4458) <= not(inputs(126)) or (inputs(241));
    layer0_outputs(4459) <= (inputs(27)) or (inputs(86));
    layer0_outputs(4460) <= inputs(137);
    layer0_outputs(4461) <= not((inputs(207)) or (inputs(172)));
    layer0_outputs(4462) <= (inputs(178)) or (inputs(130));
    layer0_outputs(4463) <= not(inputs(107));
    layer0_outputs(4464) <= not(inputs(50));
    layer0_outputs(4465) <= not(inputs(138)) or (inputs(78));
    layer0_outputs(4466) <= inputs(73);
    layer0_outputs(4467) <= not(inputs(156));
    layer0_outputs(4468) <= inputs(216);
    layer0_outputs(4469) <= (inputs(107)) or (inputs(103));
    layer0_outputs(4470) <= not((inputs(187)) or (inputs(222)));
    layer0_outputs(4471) <= not((inputs(229)) and (inputs(180)));
    layer0_outputs(4472) <= not(inputs(165)) or (inputs(171));
    layer0_outputs(4473) <= not((inputs(44)) or (inputs(251)));
    layer0_outputs(4474) <= inputs(183);
    layer0_outputs(4475) <= (inputs(138)) or (inputs(109));
    layer0_outputs(4476) <= not(inputs(153));
    layer0_outputs(4477) <= inputs(92);
    layer0_outputs(4478) <= not(inputs(220)) or (inputs(22));
    layer0_outputs(4479) <= not((inputs(37)) or (inputs(108)));
    layer0_outputs(4480) <= not(inputs(147)) or (inputs(184));
    layer0_outputs(4481) <= not(inputs(194));
    layer0_outputs(4482) <= (inputs(155)) and not (inputs(81));
    layer0_outputs(4483) <= not(inputs(75)) or (inputs(113));
    layer0_outputs(4484) <= inputs(4);
    layer0_outputs(4485) <= not((inputs(162)) xor (inputs(143)));
    layer0_outputs(4486) <= inputs(56);
    layer0_outputs(4487) <= not(inputs(64)) or (inputs(179));
    layer0_outputs(4488) <= (inputs(141)) or (inputs(240));
    layer0_outputs(4489) <= (inputs(168)) and not (inputs(171));
    layer0_outputs(4490) <= (inputs(43)) and not (inputs(146));
    layer0_outputs(4491) <= not(inputs(152));
    layer0_outputs(4492) <= (inputs(152)) and not (inputs(191));
    layer0_outputs(4493) <= not(inputs(126));
    layer0_outputs(4494) <= not(inputs(153));
    layer0_outputs(4495) <= inputs(243);
    layer0_outputs(4496) <= inputs(10);
    layer0_outputs(4497) <= not((inputs(21)) or (inputs(47)));
    layer0_outputs(4498) <= not((inputs(46)) or (inputs(12)));
    layer0_outputs(4499) <= '0';
    layer0_outputs(4500) <= not(inputs(80));
    layer0_outputs(4501) <= not(inputs(229));
    layer0_outputs(4502) <= inputs(75);
    layer0_outputs(4503) <= inputs(134);
    layer0_outputs(4504) <= (inputs(14)) xor (inputs(31));
    layer0_outputs(4505) <= (inputs(105)) xor (inputs(136));
    layer0_outputs(4506) <= not(inputs(43)) or (inputs(188));
    layer0_outputs(4507) <= not((inputs(59)) or (inputs(127)));
    layer0_outputs(4508) <= not(inputs(142)) or (inputs(0));
    layer0_outputs(4509) <= inputs(102);
    layer0_outputs(4510) <= (inputs(245)) or (inputs(26));
    layer0_outputs(4511) <= (inputs(22)) xor (inputs(244));
    layer0_outputs(4512) <= (inputs(46)) and not (inputs(53));
    layer0_outputs(4513) <= (inputs(60)) xor (inputs(28));
    layer0_outputs(4514) <= not((inputs(198)) and (inputs(111)));
    layer0_outputs(4515) <= not(inputs(165));
    layer0_outputs(4516) <= not((inputs(39)) and (inputs(210)));
    layer0_outputs(4517) <= not(inputs(19)) or (inputs(82));
    layer0_outputs(4518) <= not(inputs(109));
    layer0_outputs(4519) <= (inputs(57)) or (inputs(91));
    layer0_outputs(4520) <= not(inputs(68));
    layer0_outputs(4521) <= (inputs(108)) and not (inputs(6));
    layer0_outputs(4522) <= not((inputs(168)) or (inputs(68)));
    layer0_outputs(4523) <= not(inputs(147));
    layer0_outputs(4524) <= not((inputs(110)) or (inputs(125)));
    layer0_outputs(4525) <= inputs(115);
    layer0_outputs(4526) <= not((inputs(171)) or (inputs(211)));
    layer0_outputs(4527) <= (inputs(208)) or (inputs(57));
    layer0_outputs(4528) <= not((inputs(250)) or (inputs(116)));
    layer0_outputs(4529) <= (inputs(34)) and not (inputs(240));
    layer0_outputs(4530) <= inputs(199);
    layer0_outputs(4531) <= not(inputs(186));
    layer0_outputs(4532) <= not(inputs(248));
    layer0_outputs(4533) <= (inputs(152)) or (inputs(197));
    layer0_outputs(4534) <= (inputs(7)) and not (inputs(154));
    layer0_outputs(4535) <= not((inputs(30)) or (inputs(90)));
    layer0_outputs(4536) <= not((inputs(255)) or (inputs(8)));
    layer0_outputs(4537) <= not(inputs(56)) or (inputs(236));
    layer0_outputs(4538) <= inputs(207);
    layer0_outputs(4539) <= not((inputs(217)) or (inputs(212)));
    layer0_outputs(4540) <= '0';
    layer0_outputs(4541) <= (inputs(182)) and not (inputs(31));
    layer0_outputs(4542) <= inputs(209);
    layer0_outputs(4543) <= not(inputs(233));
    layer0_outputs(4544) <= (inputs(187)) and (inputs(185));
    layer0_outputs(4545) <= not(inputs(82)) or (inputs(8));
    layer0_outputs(4546) <= (inputs(152)) or (inputs(254));
    layer0_outputs(4547) <= not(inputs(91)) or (inputs(176));
    layer0_outputs(4548) <= not(inputs(123));
    layer0_outputs(4549) <= not((inputs(3)) and (inputs(57)));
    layer0_outputs(4550) <= not(inputs(178));
    layer0_outputs(4551) <= (inputs(71)) xor (inputs(43));
    layer0_outputs(4552) <= (inputs(50)) or (inputs(123));
    layer0_outputs(4553) <= '0';
    layer0_outputs(4554) <= (inputs(206)) xor (inputs(50));
    layer0_outputs(4555) <= not(inputs(197));
    layer0_outputs(4556) <= inputs(66);
    layer0_outputs(4557) <= not(inputs(212));
    layer0_outputs(4558) <= not(inputs(220)) or (inputs(248));
    layer0_outputs(4559) <= inputs(254);
    layer0_outputs(4560) <= not(inputs(37));
    layer0_outputs(4561) <= inputs(129);
    layer0_outputs(4562) <= inputs(227);
    layer0_outputs(4563) <= not(inputs(244));
    layer0_outputs(4564) <= not((inputs(73)) xor (inputs(12)));
    layer0_outputs(4565) <= not((inputs(90)) or (inputs(126)));
    layer0_outputs(4566) <= not((inputs(42)) or (inputs(28)));
    layer0_outputs(4567) <= not((inputs(225)) or (inputs(104)));
    layer0_outputs(4568) <= not(inputs(156));
    layer0_outputs(4569) <= not((inputs(128)) or (inputs(250)));
    layer0_outputs(4570) <= not((inputs(238)) or (inputs(86)));
    layer0_outputs(4571) <= (inputs(228)) and not (inputs(111));
    layer0_outputs(4572) <= (inputs(147)) or (inputs(207));
    layer0_outputs(4573) <= (inputs(133)) xor (inputs(34));
    layer0_outputs(4574) <= not((inputs(228)) or (inputs(54)));
    layer0_outputs(4575) <= not((inputs(167)) or (inputs(105)));
    layer0_outputs(4576) <= not((inputs(13)) and (inputs(195)));
    layer0_outputs(4577) <= not(inputs(201)) or (inputs(185));
    layer0_outputs(4578) <= '0';
    layer0_outputs(4579) <= not((inputs(140)) or (inputs(125)));
    layer0_outputs(4580) <= (inputs(217)) and not (inputs(70));
    layer0_outputs(4581) <= not((inputs(122)) or (inputs(120)));
    layer0_outputs(4582) <= inputs(67);
    layer0_outputs(4583) <= not((inputs(175)) or (inputs(95)));
    layer0_outputs(4584) <= not(inputs(99));
    layer0_outputs(4585) <= not(inputs(213));
    layer0_outputs(4586) <= not(inputs(39));
    layer0_outputs(4587) <= not(inputs(229));
    layer0_outputs(4588) <= (inputs(36)) or (inputs(137));
    layer0_outputs(4589) <= not((inputs(143)) or (inputs(204)));
    layer0_outputs(4590) <= (inputs(121)) or (inputs(106));
    layer0_outputs(4591) <= '1';
    layer0_outputs(4592) <= inputs(22);
    layer0_outputs(4593) <= not((inputs(175)) or (inputs(189)));
    layer0_outputs(4594) <= (inputs(6)) or (inputs(124));
    layer0_outputs(4595) <= (inputs(86)) and not (inputs(33));
    layer0_outputs(4596) <= inputs(234);
    layer0_outputs(4597) <= (inputs(229)) and not (inputs(122));
    layer0_outputs(4598) <= (inputs(63)) or (inputs(159));
    layer0_outputs(4599) <= not(inputs(202));
    layer0_outputs(4600) <= inputs(6);
    layer0_outputs(4601) <= inputs(69);
    layer0_outputs(4602) <= inputs(174);
    layer0_outputs(4603) <= (inputs(152)) or (inputs(96));
    layer0_outputs(4604) <= not(inputs(213)) or (inputs(88));
    layer0_outputs(4605) <= (inputs(95)) or (inputs(195));
    layer0_outputs(4606) <= not(inputs(231));
    layer0_outputs(4607) <= (inputs(63)) xor (inputs(26));
    layer0_outputs(4608) <= (inputs(146)) or (inputs(146));
    layer0_outputs(4609) <= not(inputs(39));
    layer0_outputs(4610) <= not(inputs(211)) or (inputs(95));
    layer0_outputs(4611) <= '0';
    layer0_outputs(4612) <= not(inputs(76));
    layer0_outputs(4613) <= inputs(110);
    layer0_outputs(4614) <= (inputs(193)) xor (inputs(73));
    layer0_outputs(4615) <= not(inputs(115)) or (inputs(238));
    layer0_outputs(4616) <= inputs(128);
    layer0_outputs(4617) <= not(inputs(226));
    layer0_outputs(4618) <= (inputs(74)) and not (inputs(171));
    layer0_outputs(4619) <= (inputs(111)) or (inputs(86));
    layer0_outputs(4620) <= '0';
    layer0_outputs(4621) <= not(inputs(151));
    layer0_outputs(4622) <= inputs(252);
    layer0_outputs(4623) <= (inputs(34)) and (inputs(83));
    layer0_outputs(4624) <= (inputs(6)) and not (inputs(205));
    layer0_outputs(4625) <= '0';
    layer0_outputs(4626) <= not(inputs(147)) or (inputs(244));
    layer0_outputs(4627) <= (inputs(44)) or (inputs(155));
    layer0_outputs(4628) <= '0';
    layer0_outputs(4629) <= not(inputs(92));
    layer0_outputs(4630) <= '0';
    layer0_outputs(4631) <= (inputs(48)) or (inputs(238));
    layer0_outputs(4632) <= not(inputs(184));
    layer0_outputs(4633) <= not(inputs(238)) or (inputs(249));
    layer0_outputs(4634) <= not(inputs(166));
    layer0_outputs(4635) <= not(inputs(127)) or (inputs(240));
    layer0_outputs(4636) <= not(inputs(24));
    layer0_outputs(4637) <= not(inputs(111));
    layer0_outputs(4638) <= inputs(46);
    layer0_outputs(4639) <= (inputs(15)) xor (inputs(202));
    layer0_outputs(4640) <= not(inputs(236)) or (inputs(241));
    layer0_outputs(4641) <= (inputs(103)) or (inputs(102));
    layer0_outputs(4642) <= (inputs(227)) and not (inputs(67));
    layer0_outputs(4643) <= (inputs(212)) and not (inputs(58));
    layer0_outputs(4644) <= inputs(63);
    layer0_outputs(4645) <= not((inputs(196)) or (inputs(82)));
    layer0_outputs(4646) <= inputs(233);
    layer0_outputs(4647) <= not((inputs(76)) xor (inputs(96)));
    layer0_outputs(4648) <= not(inputs(59)) or (inputs(130));
    layer0_outputs(4649) <= not(inputs(228));
    layer0_outputs(4650) <= (inputs(153)) and not (inputs(7));
    layer0_outputs(4651) <= inputs(130);
    layer0_outputs(4652) <= not((inputs(131)) or (inputs(234)));
    layer0_outputs(4653) <= not(inputs(196));
    layer0_outputs(4654) <= inputs(121);
    layer0_outputs(4655) <= not((inputs(22)) and (inputs(10)));
    layer0_outputs(4656) <= (inputs(101)) and not (inputs(18));
    layer0_outputs(4657) <= not(inputs(230));
    layer0_outputs(4658) <= not(inputs(102)) or (inputs(207));
    layer0_outputs(4659) <= (inputs(150)) or (inputs(168));
    layer0_outputs(4660) <= not(inputs(4));
    layer0_outputs(4661) <= (inputs(22)) and not (inputs(203));
    layer0_outputs(4662) <= (inputs(38)) and not (inputs(31));
    layer0_outputs(4663) <= not((inputs(80)) or (inputs(168)));
    layer0_outputs(4664) <= (inputs(124)) and not (inputs(211));
    layer0_outputs(4665) <= not(inputs(128));
    layer0_outputs(4666) <= not(inputs(157)) or (inputs(184));
    layer0_outputs(4667) <= (inputs(22)) and not (inputs(102));
    layer0_outputs(4668) <= not(inputs(22));
    layer0_outputs(4669) <= (inputs(165)) and not (inputs(47));
    layer0_outputs(4670) <= not((inputs(49)) or (inputs(33)));
    layer0_outputs(4671) <= not((inputs(185)) and (inputs(125)));
    layer0_outputs(4672) <= (inputs(61)) and (inputs(50));
    layer0_outputs(4673) <= not(inputs(245)) or (inputs(121));
    layer0_outputs(4674) <= not((inputs(243)) xor (inputs(34)));
    layer0_outputs(4675) <= '0';
    layer0_outputs(4676) <= not((inputs(62)) or (inputs(56)));
    layer0_outputs(4677) <= not(inputs(78));
    layer0_outputs(4678) <= not(inputs(119)) or (inputs(193));
    layer0_outputs(4679) <= (inputs(37)) and not (inputs(144));
    layer0_outputs(4680) <= not((inputs(158)) or (inputs(27)));
    layer0_outputs(4681) <= (inputs(197)) or (inputs(125));
    layer0_outputs(4682) <= inputs(124);
    layer0_outputs(4683) <= not((inputs(172)) or (inputs(107)));
    layer0_outputs(4684) <= not((inputs(192)) or (inputs(230)));
    layer0_outputs(4685) <= (inputs(189)) or (inputs(51));
    layer0_outputs(4686) <= '0';
    layer0_outputs(4687) <= '1';
    layer0_outputs(4688) <= not((inputs(190)) or (inputs(62)));
    layer0_outputs(4689) <= inputs(160);
    layer0_outputs(4690) <= not((inputs(104)) or (inputs(51)));
    layer0_outputs(4691) <= not((inputs(15)) and (inputs(94)));
    layer0_outputs(4692) <= not(inputs(166)) or (inputs(172));
    layer0_outputs(4693) <= not(inputs(194));
    layer0_outputs(4694) <= (inputs(196)) xor (inputs(225));
    layer0_outputs(4695) <= (inputs(58)) or (inputs(78));
    layer0_outputs(4696) <= inputs(120);
    layer0_outputs(4697) <= inputs(193);
    layer0_outputs(4698) <= (inputs(174)) or (inputs(56));
    layer0_outputs(4699) <= inputs(85);
    layer0_outputs(4700) <= '0';
    layer0_outputs(4701) <= not(inputs(196)) or (inputs(23));
    layer0_outputs(4702) <= not((inputs(15)) or (inputs(178)));
    layer0_outputs(4703) <= (inputs(110)) or (inputs(134));
    layer0_outputs(4704) <= inputs(21);
    layer0_outputs(4705) <= (inputs(90)) or (inputs(122));
    layer0_outputs(4706) <= not(inputs(91)) or (inputs(253));
    layer0_outputs(4707) <= inputs(210);
    layer0_outputs(4708) <= not(inputs(143));
    layer0_outputs(4709) <= (inputs(237)) or (inputs(180));
    layer0_outputs(4710) <= '0';
    layer0_outputs(4711) <= inputs(179);
    layer0_outputs(4712) <= not(inputs(94));
    layer0_outputs(4713) <= not(inputs(155));
    layer0_outputs(4714) <= (inputs(79)) and (inputs(105));
    layer0_outputs(4715) <= (inputs(194)) and not (inputs(64));
    layer0_outputs(4716) <= (inputs(141)) and not (inputs(17));
    layer0_outputs(4717) <= not((inputs(216)) or (inputs(118)));
    layer0_outputs(4718) <= not(inputs(133));
    layer0_outputs(4719) <= (inputs(32)) and not (inputs(234));
    layer0_outputs(4720) <= inputs(146);
    layer0_outputs(4721) <= (inputs(106)) and not (inputs(55));
    layer0_outputs(4722) <= '0';
    layer0_outputs(4723) <= (inputs(0)) or (inputs(33));
    layer0_outputs(4724) <= not(inputs(24));
    layer0_outputs(4725) <= not((inputs(46)) or (inputs(163)));
    layer0_outputs(4726) <= not((inputs(116)) or (inputs(117)));
    layer0_outputs(4727) <= not(inputs(42)) or (inputs(167));
    layer0_outputs(4728) <= not((inputs(94)) xor (inputs(135)));
    layer0_outputs(4729) <= '0';
    layer0_outputs(4730) <= inputs(10);
    layer0_outputs(4731) <= (inputs(29)) and (inputs(240));
    layer0_outputs(4732) <= not(inputs(103)) or (inputs(182));
    layer0_outputs(4733) <= (inputs(172)) or (inputs(236));
    layer0_outputs(4734) <= not(inputs(44)) or (inputs(103));
    layer0_outputs(4735) <= not(inputs(114));
    layer0_outputs(4736) <= inputs(69);
    layer0_outputs(4737) <= inputs(43);
    layer0_outputs(4738) <= not((inputs(59)) and (inputs(206)));
    layer0_outputs(4739) <= (inputs(99)) and not (inputs(207));
    layer0_outputs(4740) <= (inputs(72)) and not (inputs(96));
    layer0_outputs(4741) <= not((inputs(63)) or (inputs(19)));
    layer0_outputs(4742) <= not(inputs(210)) or (inputs(56));
    layer0_outputs(4743) <= (inputs(181)) and not (inputs(146));
    layer0_outputs(4744) <= '0';
    layer0_outputs(4745) <= not((inputs(152)) and (inputs(179)));
    layer0_outputs(4746) <= inputs(132);
    layer0_outputs(4747) <= inputs(37);
    layer0_outputs(4748) <= '1';
    layer0_outputs(4749) <= '0';
    layer0_outputs(4750) <= (inputs(128)) and not (inputs(1));
    layer0_outputs(4751) <= not(inputs(25));
    layer0_outputs(4752) <= inputs(145);
    layer0_outputs(4753) <= not(inputs(118)) or (inputs(6));
    layer0_outputs(4754) <= inputs(129);
    layer0_outputs(4755) <= not(inputs(24));
    layer0_outputs(4756) <= inputs(138);
    layer0_outputs(4757) <= not((inputs(149)) xor (inputs(102)));
    layer0_outputs(4758) <= (inputs(134)) or (inputs(152));
    layer0_outputs(4759) <= (inputs(77)) and not (inputs(2));
    layer0_outputs(4760) <= (inputs(177)) or (inputs(121));
    layer0_outputs(4761) <= (inputs(128)) and not (inputs(96));
    layer0_outputs(4762) <= not(inputs(2)) or (inputs(244));
    layer0_outputs(4763) <= (inputs(98)) and not (inputs(48));
    layer0_outputs(4764) <= (inputs(23)) and (inputs(25));
    layer0_outputs(4765) <= not(inputs(167)) or (inputs(99));
    layer0_outputs(4766) <= (inputs(178)) and not (inputs(71));
    layer0_outputs(4767) <= not(inputs(153));
    layer0_outputs(4768) <= not((inputs(165)) or (inputs(165)));
    layer0_outputs(4769) <= not((inputs(164)) xor (inputs(143)));
    layer0_outputs(4770) <= (inputs(56)) and not (inputs(167));
    layer0_outputs(4771) <= inputs(127);
    layer0_outputs(4772) <= (inputs(112)) and not (inputs(250));
    layer0_outputs(4773) <= not(inputs(29)) or (inputs(34));
    layer0_outputs(4774) <= inputs(25);
    layer0_outputs(4775) <= not((inputs(116)) or (inputs(167)));
    layer0_outputs(4776) <= (inputs(107)) and not (inputs(198));
    layer0_outputs(4777) <= not(inputs(8)) or (inputs(97));
    layer0_outputs(4778) <= not(inputs(231));
    layer0_outputs(4779) <= inputs(64);
    layer0_outputs(4780) <= (inputs(229)) or (inputs(34));
    layer0_outputs(4781) <= not(inputs(157));
    layer0_outputs(4782) <= (inputs(231)) and not (inputs(252));
    layer0_outputs(4783) <= not(inputs(168));
    layer0_outputs(4784) <= inputs(40);
    layer0_outputs(4785) <= not(inputs(164)) or (inputs(247));
    layer0_outputs(4786) <= not((inputs(132)) and (inputs(97)));
    layer0_outputs(4787) <= (inputs(45)) and not (inputs(217));
    layer0_outputs(4788) <= not(inputs(102));
    layer0_outputs(4789) <= not(inputs(171));
    layer0_outputs(4790) <= '0';
    layer0_outputs(4791) <= not((inputs(43)) or (inputs(63)));
    layer0_outputs(4792) <= not((inputs(103)) or (inputs(136)));
    layer0_outputs(4793) <= '1';
    layer0_outputs(4794) <= not(inputs(255)) or (inputs(235));
    layer0_outputs(4795) <= not(inputs(163)) or (inputs(10));
    layer0_outputs(4796) <= '1';
    layer0_outputs(4797) <= not((inputs(20)) or (inputs(179)));
    layer0_outputs(4798) <= (inputs(16)) or (inputs(123));
    layer0_outputs(4799) <= not((inputs(43)) or (inputs(154)));
    layer0_outputs(4800) <= (inputs(31)) and not (inputs(203));
    layer0_outputs(4801) <= inputs(231);
    layer0_outputs(4802) <= not(inputs(174)) or (inputs(97));
    layer0_outputs(4803) <= not(inputs(151)) or (inputs(224));
    layer0_outputs(4804) <= (inputs(119)) and not (inputs(204));
    layer0_outputs(4805) <= not(inputs(69)) or (inputs(127));
    layer0_outputs(4806) <= not(inputs(51));
    layer0_outputs(4807) <= (inputs(75)) or (inputs(49));
    layer0_outputs(4808) <= not((inputs(51)) and (inputs(55)));
    layer0_outputs(4809) <= inputs(210);
    layer0_outputs(4810) <= not(inputs(85)) or (inputs(79));
    layer0_outputs(4811) <= inputs(63);
    layer0_outputs(4812) <= inputs(127);
    layer0_outputs(4813) <= not((inputs(3)) or (inputs(218)));
    layer0_outputs(4814) <= (inputs(172)) xor (inputs(231));
    layer0_outputs(4815) <= '1';
    layer0_outputs(4816) <= inputs(84);
    layer0_outputs(4817) <= not((inputs(96)) xor (inputs(71)));
    layer0_outputs(4818) <= '0';
    layer0_outputs(4819) <= inputs(81);
    layer0_outputs(4820) <= not((inputs(88)) or (inputs(219)));
    layer0_outputs(4821) <= (inputs(0)) and (inputs(62));
    layer0_outputs(4822) <= not(inputs(209));
    layer0_outputs(4823) <= inputs(84);
    layer0_outputs(4824) <= (inputs(150)) and not (inputs(15));
    layer0_outputs(4825) <= '0';
    layer0_outputs(4826) <= (inputs(79)) or (inputs(72));
    layer0_outputs(4827) <= not(inputs(243));
    layer0_outputs(4828) <= not(inputs(97));
    layer0_outputs(4829) <= not((inputs(232)) and (inputs(173)));
    layer0_outputs(4830) <= (inputs(236)) and not (inputs(205));
    layer0_outputs(4831) <= (inputs(192)) or (inputs(199));
    layer0_outputs(4832) <= (inputs(238)) and (inputs(210));
    layer0_outputs(4833) <= not((inputs(16)) or (inputs(194)));
    layer0_outputs(4834) <= not((inputs(69)) or (inputs(148)));
    layer0_outputs(4835) <= inputs(180);
    layer0_outputs(4836) <= not(inputs(133)) or (inputs(142));
    layer0_outputs(4837) <= not(inputs(123));
    layer0_outputs(4838) <= inputs(247);
    layer0_outputs(4839) <= '1';
    layer0_outputs(4840) <= not((inputs(154)) xor (inputs(64)));
    layer0_outputs(4841) <= inputs(137);
    layer0_outputs(4842) <= inputs(178);
    layer0_outputs(4843) <= (inputs(183)) or (inputs(129));
    layer0_outputs(4844) <= not((inputs(34)) or (inputs(134)));
    layer0_outputs(4845) <= not(inputs(182));
    layer0_outputs(4846) <= inputs(17);
    layer0_outputs(4847) <= (inputs(28)) and not (inputs(158));
    layer0_outputs(4848) <= (inputs(159)) or (inputs(158));
    layer0_outputs(4849) <= not(inputs(250));
    layer0_outputs(4850) <= '0';
    layer0_outputs(4851) <= not((inputs(145)) or (inputs(20)));
    layer0_outputs(4852) <= (inputs(67)) and not (inputs(48));
    layer0_outputs(4853) <= inputs(82);
    layer0_outputs(4854) <= not(inputs(16)) or (inputs(230));
    layer0_outputs(4855) <= not(inputs(22));
    layer0_outputs(4856) <= (inputs(176)) and not (inputs(142));
    layer0_outputs(4857) <= (inputs(62)) and not (inputs(74));
    layer0_outputs(4858) <= (inputs(48)) xor (inputs(211));
    layer0_outputs(4859) <= not((inputs(241)) or (inputs(150)));
    layer0_outputs(4860) <= not(inputs(233));
    layer0_outputs(4861) <= not(inputs(22)) or (inputs(158));
    layer0_outputs(4862) <= inputs(1);
    layer0_outputs(4863) <= not((inputs(171)) or (inputs(30)));
    layer0_outputs(4864) <= inputs(130);
    layer0_outputs(4865) <= not(inputs(36));
    layer0_outputs(4866) <= not(inputs(56)) or (inputs(6));
    layer0_outputs(4867) <= not(inputs(74));
    layer0_outputs(4868) <= (inputs(104)) and not (inputs(98));
    layer0_outputs(4869) <= inputs(7);
    layer0_outputs(4870) <= inputs(214);
    layer0_outputs(4871) <= (inputs(30)) and not (inputs(89));
    layer0_outputs(4872) <= (inputs(209)) or (inputs(38));
    layer0_outputs(4873) <= not((inputs(117)) or (inputs(15)));
    layer0_outputs(4874) <= inputs(104);
    layer0_outputs(4875) <= inputs(189);
    layer0_outputs(4876) <= inputs(62);
    layer0_outputs(4877) <= inputs(14);
    layer0_outputs(4878) <= not(inputs(107)) or (inputs(215));
    layer0_outputs(4879) <= (inputs(101)) and (inputs(27));
    layer0_outputs(4880) <= not(inputs(150)) or (inputs(37));
    layer0_outputs(4881) <= (inputs(116)) xor (inputs(20));
    layer0_outputs(4882) <= not(inputs(139));
    layer0_outputs(4883) <= inputs(168);
    layer0_outputs(4884) <= not((inputs(246)) or (inputs(210)));
    layer0_outputs(4885) <= (inputs(250)) or (inputs(235));
    layer0_outputs(4886) <= inputs(15);
    layer0_outputs(4887) <= '1';
    layer0_outputs(4888) <= not((inputs(180)) xor (inputs(242)));
    layer0_outputs(4889) <= (inputs(0)) and not (inputs(41));
    layer0_outputs(4890) <= (inputs(100)) and not (inputs(140));
    layer0_outputs(4891) <= (inputs(126)) and (inputs(71));
    layer0_outputs(4892) <= '1';
    layer0_outputs(4893) <= not((inputs(178)) or (inputs(111)));
    layer0_outputs(4894) <= not((inputs(20)) or (inputs(99)));
    layer0_outputs(4895) <= (inputs(154)) and not (inputs(31));
    layer0_outputs(4896) <= (inputs(252)) or (inputs(196));
    layer0_outputs(4897) <= not(inputs(24));
    layer0_outputs(4898) <= not(inputs(135));
    layer0_outputs(4899) <= not((inputs(38)) or (inputs(96)));
    layer0_outputs(4900) <= not(inputs(115));
    layer0_outputs(4901) <= not(inputs(90));
    layer0_outputs(4902) <= inputs(40);
    layer0_outputs(4903) <= '0';
    layer0_outputs(4904) <= not(inputs(164));
    layer0_outputs(4905) <= '1';
    layer0_outputs(4906) <= (inputs(161)) or (inputs(110));
    layer0_outputs(4907) <= (inputs(120)) or (inputs(144));
    layer0_outputs(4908) <= (inputs(115)) and not (inputs(170));
    layer0_outputs(4909) <= inputs(144);
    layer0_outputs(4910) <= inputs(227);
    layer0_outputs(4911) <= not((inputs(104)) and (inputs(132)));
    layer0_outputs(4912) <= not(inputs(10));
    layer0_outputs(4913) <= inputs(144);
    layer0_outputs(4914) <= (inputs(173)) and not (inputs(124));
    layer0_outputs(4915) <= inputs(168);
    layer0_outputs(4916) <= not(inputs(128));
    layer0_outputs(4917) <= inputs(94);
    layer0_outputs(4918) <= (inputs(245)) and (inputs(79));
    layer0_outputs(4919) <= inputs(89);
    layer0_outputs(4920) <= not(inputs(91));
    layer0_outputs(4921) <= not(inputs(189));
    layer0_outputs(4922) <= (inputs(52)) or (inputs(53));
    layer0_outputs(4923) <= not(inputs(132)) or (inputs(177));
    layer0_outputs(4924) <= inputs(183);
    layer0_outputs(4925) <= not((inputs(51)) or (inputs(244)));
    layer0_outputs(4926) <= '1';
    layer0_outputs(4927) <= (inputs(78)) and not (inputs(223));
    layer0_outputs(4928) <= (inputs(190)) xor (inputs(95));
    layer0_outputs(4929) <= (inputs(245)) and not (inputs(126));
    layer0_outputs(4930) <= not(inputs(5));
    layer0_outputs(4931) <= not(inputs(231));
    layer0_outputs(4932) <= not(inputs(208));
    layer0_outputs(4933) <= inputs(1);
    layer0_outputs(4934) <= (inputs(233)) and not (inputs(145));
    layer0_outputs(4935) <= (inputs(59)) and not (inputs(188));
    layer0_outputs(4936) <= (inputs(186)) or (inputs(64));
    layer0_outputs(4937) <= inputs(73);
    layer0_outputs(4938) <= inputs(138);
    layer0_outputs(4939) <= not(inputs(224)) or (inputs(126));
    layer0_outputs(4940) <= not(inputs(172));
    layer0_outputs(4941) <= not(inputs(75));
    layer0_outputs(4942) <= inputs(233);
    layer0_outputs(4943) <= inputs(168);
    layer0_outputs(4944) <= (inputs(151)) and not (inputs(71));
    layer0_outputs(4945) <= inputs(213);
    layer0_outputs(4946) <= not(inputs(116));
    layer0_outputs(4947) <= (inputs(47)) and not (inputs(126));
    layer0_outputs(4948) <= (inputs(33)) or (inputs(176));
    layer0_outputs(4949) <= not((inputs(164)) or (inputs(192)));
    layer0_outputs(4950) <= not((inputs(33)) or (inputs(232)));
    layer0_outputs(4951) <= not(inputs(148));
    layer0_outputs(4952) <= (inputs(13)) and (inputs(111));
    layer0_outputs(4953) <= (inputs(92)) xor (inputs(255));
    layer0_outputs(4954) <= (inputs(158)) or (inputs(34));
    layer0_outputs(4955) <= inputs(180);
    layer0_outputs(4956) <= not(inputs(221));
    layer0_outputs(4957) <= (inputs(179)) xor (inputs(30));
    layer0_outputs(4958) <= not(inputs(35));
    layer0_outputs(4959) <= not(inputs(153));
    layer0_outputs(4960) <= (inputs(203)) or (inputs(17));
    layer0_outputs(4961) <= inputs(45);
    layer0_outputs(4962) <= (inputs(190)) and not (inputs(157));
    layer0_outputs(4963) <= (inputs(236)) and not (inputs(170));
    layer0_outputs(4964) <= (inputs(215)) xor (inputs(248));
    layer0_outputs(4965) <= not((inputs(48)) or (inputs(135)));
    layer0_outputs(4966) <= not((inputs(29)) or (inputs(181)));
    layer0_outputs(4967) <= (inputs(213)) or (inputs(229));
    layer0_outputs(4968) <= inputs(215);
    layer0_outputs(4969) <= not(inputs(213));
    layer0_outputs(4970) <= (inputs(5)) and not (inputs(14));
    layer0_outputs(4971) <= (inputs(67)) xor (inputs(224));
    layer0_outputs(4972) <= inputs(21);
    layer0_outputs(4973) <= (inputs(228)) or (inputs(222));
    layer0_outputs(4974) <= not(inputs(54)) or (inputs(9));
    layer0_outputs(4975) <= (inputs(72)) xor (inputs(23));
    layer0_outputs(4976) <= not(inputs(46));
    layer0_outputs(4977) <= not(inputs(77)) or (inputs(237));
    layer0_outputs(4978) <= not(inputs(151));
    layer0_outputs(4979) <= inputs(6);
    layer0_outputs(4980) <= '1';
    layer0_outputs(4981) <= (inputs(38)) and not (inputs(158));
    layer0_outputs(4982) <= not(inputs(223));
    layer0_outputs(4983) <= (inputs(12)) and not (inputs(151));
    layer0_outputs(4984) <= not((inputs(149)) or (inputs(188)));
    layer0_outputs(4985) <= inputs(248);
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= (inputs(48)) xor (inputs(116));
    layer0_outputs(4988) <= '0';
    layer0_outputs(4989) <= not(inputs(203));
    layer0_outputs(4990) <= inputs(196);
    layer0_outputs(4991) <= (inputs(238)) or (inputs(137));
    layer0_outputs(4992) <= '1';
    layer0_outputs(4993) <= not((inputs(3)) or (inputs(5)));
    layer0_outputs(4994) <= (inputs(124)) and not (inputs(183));
    layer0_outputs(4995) <= not(inputs(24));
    layer0_outputs(4996) <= not(inputs(1));
    layer0_outputs(4997) <= not(inputs(70)) or (inputs(251));
    layer0_outputs(4998) <= (inputs(156)) or (inputs(138));
    layer0_outputs(4999) <= not((inputs(225)) or (inputs(232)));
    layer0_outputs(5000) <= not(inputs(252));
    layer0_outputs(5001) <= inputs(146);
    layer0_outputs(5002) <= not(inputs(131));
    layer0_outputs(5003) <= inputs(62);
    layer0_outputs(5004) <= '0';
    layer0_outputs(5005) <= inputs(138);
    layer0_outputs(5006) <= not(inputs(0));
    layer0_outputs(5007) <= not(inputs(89));
    layer0_outputs(5008) <= not((inputs(84)) and (inputs(226)));
    layer0_outputs(5009) <= not(inputs(54)) or (inputs(232));
    layer0_outputs(5010) <= inputs(136);
    layer0_outputs(5011) <= (inputs(25)) or (inputs(2));
    layer0_outputs(5012) <= '1';
    layer0_outputs(5013) <= (inputs(224)) xor (inputs(153));
    layer0_outputs(5014) <= not((inputs(84)) or (inputs(68)));
    layer0_outputs(5015) <= not(inputs(40)) or (inputs(239));
    layer0_outputs(5016) <= not(inputs(159)) or (inputs(126));
    layer0_outputs(5017) <= inputs(133);
    layer0_outputs(5018) <= (inputs(49)) or (inputs(2));
    layer0_outputs(5019) <= inputs(23);
    layer0_outputs(5020) <= inputs(134);
    layer0_outputs(5021) <= not(inputs(24));
    layer0_outputs(5022) <= (inputs(62)) and not (inputs(247));
    layer0_outputs(5023) <= (inputs(16)) xor (inputs(64));
    layer0_outputs(5024) <= not(inputs(99));
    layer0_outputs(5025) <= (inputs(198)) and not (inputs(54));
    layer0_outputs(5026) <= (inputs(186)) xor (inputs(83));
    layer0_outputs(5027) <= (inputs(93)) or (inputs(50));
    layer0_outputs(5028) <= not(inputs(39));
    layer0_outputs(5029) <= not((inputs(101)) or (inputs(94)));
    layer0_outputs(5030) <= not((inputs(175)) and (inputs(146)));
    layer0_outputs(5031) <= inputs(245);
    layer0_outputs(5032) <= (inputs(51)) and (inputs(118));
    layer0_outputs(5033) <= not((inputs(194)) or (inputs(191)));
    layer0_outputs(5034) <= inputs(243);
    layer0_outputs(5035) <= not((inputs(14)) xor (inputs(160)));
    layer0_outputs(5036) <= (inputs(106)) and not (inputs(5));
    layer0_outputs(5037) <= not(inputs(101)) or (inputs(216));
    layer0_outputs(5038) <= (inputs(180)) xor (inputs(32));
    layer0_outputs(5039) <= not((inputs(41)) xor (inputs(105)));
    layer0_outputs(5040) <= not(inputs(32));
    layer0_outputs(5041) <= not(inputs(194));
    layer0_outputs(5042) <= inputs(149);
    layer0_outputs(5043) <= not((inputs(169)) or (inputs(98)));
    layer0_outputs(5044) <= not((inputs(96)) and (inputs(147)));
    layer0_outputs(5045) <= (inputs(19)) or (inputs(253));
    layer0_outputs(5046) <= not((inputs(55)) and (inputs(112)));
    layer0_outputs(5047) <= not((inputs(242)) and (inputs(176)));
    layer0_outputs(5048) <= (inputs(220)) and not (inputs(156));
    layer0_outputs(5049) <= (inputs(114)) and not (inputs(239));
    layer0_outputs(5050) <= inputs(184);
    layer0_outputs(5051) <= inputs(86);
    layer0_outputs(5052) <= not((inputs(2)) or (inputs(68)));
    layer0_outputs(5053) <= (inputs(222)) and not (inputs(129));
    layer0_outputs(5054) <= (inputs(3)) and not (inputs(255));
    layer0_outputs(5055) <= not((inputs(209)) or (inputs(188)));
    layer0_outputs(5056) <= inputs(209);
    layer0_outputs(5057) <= (inputs(252)) and not (inputs(212));
    layer0_outputs(5058) <= inputs(179);
    layer0_outputs(5059) <= not((inputs(204)) xor (inputs(68)));
    layer0_outputs(5060) <= (inputs(90)) xor (inputs(106));
    layer0_outputs(5061) <= (inputs(137)) and not (inputs(223));
    layer0_outputs(5062) <= not((inputs(188)) or (inputs(149)));
    layer0_outputs(5063) <= not(inputs(68));
    layer0_outputs(5064) <= inputs(149);
    layer0_outputs(5065) <= (inputs(103)) and not (inputs(14));
    layer0_outputs(5066) <= not(inputs(99));
    layer0_outputs(5067) <= inputs(114);
    layer0_outputs(5068) <= inputs(135);
    layer0_outputs(5069) <= not(inputs(162));
    layer0_outputs(5070) <= '0';
    layer0_outputs(5071) <= (inputs(136)) and not (inputs(77));
    layer0_outputs(5072) <= not((inputs(146)) or (inputs(223)));
    layer0_outputs(5073) <= inputs(126);
    layer0_outputs(5074) <= not(inputs(122)) or (inputs(233));
    layer0_outputs(5075) <= '0';
    layer0_outputs(5076) <= not((inputs(212)) xor (inputs(181)));
    layer0_outputs(5077) <= (inputs(119)) or (inputs(125));
    layer0_outputs(5078) <= not((inputs(79)) or (inputs(4)));
    layer0_outputs(5079) <= not(inputs(107)) or (inputs(87));
    layer0_outputs(5080) <= inputs(136);
    layer0_outputs(5081) <= not(inputs(38));
    layer0_outputs(5082) <= not((inputs(47)) xor (inputs(184)));
    layer0_outputs(5083) <= (inputs(132)) xor (inputs(101));
    layer0_outputs(5084) <= not(inputs(41)) or (inputs(80));
    layer0_outputs(5085) <= not(inputs(150));
    layer0_outputs(5086) <= not(inputs(111)) or (inputs(42));
    layer0_outputs(5087) <= not((inputs(32)) xor (inputs(167)));
    layer0_outputs(5088) <= not(inputs(136)) or (inputs(194));
    layer0_outputs(5089) <= '1';
    layer0_outputs(5090) <= inputs(213);
    layer0_outputs(5091) <= (inputs(14)) or (inputs(109));
    layer0_outputs(5092) <= (inputs(35)) and not (inputs(70));
    layer0_outputs(5093) <= not((inputs(25)) or (inputs(34)));
    layer0_outputs(5094) <= (inputs(121)) or (inputs(104));
    layer0_outputs(5095) <= (inputs(38)) and (inputs(104));
    layer0_outputs(5096) <= (inputs(221)) or (inputs(99));
    layer0_outputs(5097) <= '0';
    layer0_outputs(5098) <= inputs(98);
    layer0_outputs(5099) <= not((inputs(203)) xor (inputs(16)));
    layer0_outputs(5100) <= not(inputs(233)) or (inputs(110));
    layer0_outputs(5101) <= not((inputs(92)) or (inputs(125)));
    layer0_outputs(5102) <= not(inputs(185));
    layer0_outputs(5103) <= inputs(130);
    layer0_outputs(5104) <= '0';
    layer0_outputs(5105) <= not((inputs(212)) or (inputs(112)));
    layer0_outputs(5106) <= (inputs(72)) and (inputs(119));
    layer0_outputs(5107) <= not((inputs(60)) or (inputs(19)));
    layer0_outputs(5108) <= inputs(245);
    layer0_outputs(5109) <= inputs(75);
    layer0_outputs(5110) <= not((inputs(189)) or (inputs(89)));
    layer0_outputs(5111) <= (inputs(202)) or (inputs(180));
    layer0_outputs(5112) <= inputs(96);
    layer0_outputs(5113) <= '1';
    layer0_outputs(5114) <= '1';
    layer0_outputs(5115) <= (inputs(223)) or (inputs(56));
    layer0_outputs(5116) <= inputs(116);
    layer0_outputs(5117) <= (inputs(46)) and not (inputs(62));
    layer0_outputs(5118) <= not(inputs(248)) or (inputs(32));
    layer0_outputs(5119) <= (inputs(69)) or (inputs(48));
    layer1_outputs(0) <= (layer0_outputs(4186)) and not (layer0_outputs(2688));
    layer1_outputs(1) <= not(layer0_outputs(2583));
    layer1_outputs(2) <= not((layer0_outputs(1448)) and (layer0_outputs(4929)));
    layer1_outputs(3) <= not((layer0_outputs(1728)) or (layer0_outputs(2709)));
    layer1_outputs(4) <= '1';
    layer1_outputs(5) <= not(layer0_outputs(1595)) or (layer0_outputs(174));
    layer1_outputs(6) <= layer0_outputs(39);
    layer1_outputs(7) <= not((layer0_outputs(3960)) and (layer0_outputs(4605)));
    layer1_outputs(8) <= not((layer0_outputs(2237)) or (layer0_outputs(4163)));
    layer1_outputs(9) <= (layer0_outputs(3662)) and not (layer0_outputs(4190));
    layer1_outputs(10) <= layer0_outputs(414);
    layer1_outputs(11) <= layer0_outputs(761);
    layer1_outputs(12) <= (layer0_outputs(1119)) and (layer0_outputs(3794));
    layer1_outputs(13) <= '0';
    layer1_outputs(14) <= not(layer0_outputs(2148));
    layer1_outputs(15) <= (layer0_outputs(1308)) and not (layer0_outputs(4761));
    layer1_outputs(16) <= (layer0_outputs(3413)) or (layer0_outputs(2752));
    layer1_outputs(17) <= layer0_outputs(4360);
    layer1_outputs(18) <= not((layer0_outputs(545)) or (layer0_outputs(4534)));
    layer1_outputs(19) <= (layer0_outputs(2991)) or (layer0_outputs(4050));
    layer1_outputs(20) <= not(layer0_outputs(3556));
    layer1_outputs(21) <= not(layer0_outputs(3975));
    layer1_outputs(22) <= not(layer0_outputs(230));
    layer1_outputs(23) <= (layer0_outputs(5023)) or (layer0_outputs(2309));
    layer1_outputs(24) <= not(layer0_outputs(213));
    layer1_outputs(25) <= not(layer0_outputs(805));
    layer1_outputs(26) <= not((layer0_outputs(2825)) xor (layer0_outputs(5020)));
    layer1_outputs(27) <= '1';
    layer1_outputs(28) <= (layer0_outputs(897)) or (layer0_outputs(2145));
    layer1_outputs(29) <= not(layer0_outputs(4763));
    layer1_outputs(30) <= layer0_outputs(1304);
    layer1_outputs(31) <= not(layer0_outputs(2297));
    layer1_outputs(32) <= not(layer0_outputs(580));
    layer1_outputs(33) <= (layer0_outputs(3387)) and not (layer0_outputs(564));
    layer1_outputs(34) <= not(layer0_outputs(3789));
    layer1_outputs(35) <= layer0_outputs(176);
    layer1_outputs(36) <= layer0_outputs(3061);
    layer1_outputs(37) <= not(layer0_outputs(1746));
    layer1_outputs(38) <= (layer0_outputs(4604)) and not (layer0_outputs(2767));
    layer1_outputs(39) <= not(layer0_outputs(1222));
    layer1_outputs(40) <= (layer0_outputs(3087)) or (layer0_outputs(2521));
    layer1_outputs(41) <= (layer0_outputs(344)) or (layer0_outputs(1812));
    layer1_outputs(42) <= not(layer0_outputs(3146));
    layer1_outputs(43) <= '1';
    layer1_outputs(44) <= not(layer0_outputs(3750));
    layer1_outputs(45) <= (layer0_outputs(825)) and (layer0_outputs(3377));
    layer1_outputs(46) <= not((layer0_outputs(544)) or (layer0_outputs(1122)));
    layer1_outputs(47) <= not(layer0_outputs(2288)) or (layer0_outputs(1719));
    layer1_outputs(48) <= not(layer0_outputs(1030)) or (layer0_outputs(1868));
    layer1_outputs(49) <= not(layer0_outputs(1765));
    layer1_outputs(50) <= not(layer0_outputs(1066)) or (layer0_outputs(3715));
    layer1_outputs(51) <= (layer0_outputs(4820)) and (layer0_outputs(236));
    layer1_outputs(52) <= layer0_outputs(1456);
    layer1_outputs(53) <= (layer0_outputs(2649)) xor (layer0_outputs(418));
    layer1_outputs(54) <= layer0_outputs(3098);
    layer1_outputs(55) <= (layer0_outputs(2142)) or (layer0_outputs(4825));
    layer1_outputs(56) <= layer0_outputs(315);
    layer1_outputs(57) <= (layer0_outputs(2188)) and (layer0_outputs(3104));
    layer1_outputs(58) <= layer0_outputs(2269);
    layer1_outputs(59) <= (layer0_outputs(1821)) and (layer0_outputs(2181));
    layer1_outputs(60) <= not(layer0_outputs(4937));
    layer1_outputs(61) <= layer0_outputs(2606);
    layer1_outputs(62) <= layer0_outputs(3606);
    layer1_outputs(63) <= not(layer0_outputs(4287));
    layer1_outputs(64) <= layer0_outputs(4038);
    layer1_outputs(65) <= (layer0_outputs(766)) and (layer0_outputs(2900));
    layer1_outputs(66) <= (layer0_outputs(1852)) and not (layer0_outputs(2408));
    layer1_outputs(67) <= not((layer0_outputs(3673)) or (layer0_outputs(3989)));
    layer1_outputs(68) <= (layer0_outputs(2448)) xor (layer0_outputs(777));
    layer1_outputs(69) <= not(layer0_outputs(2571)) or (layer0_outputs(3699));
    layer1_outputs(70) <= layer0_outputs(407);
    layer1_outputs(71) <= layer0_outputs(2585);
    layer1_outputs(72) <= layer0_outputs(3);
    layer1_outputs(73) <= (layer0_outputs(24)) and not (layer0_outputs(34));
    layer1_outputs(74) <= layer0_outputs(150);
    layer1_outputs(75) <= (layer0_outputs(4713)) and not (layer0_outputs(56));
    layer1_outputs(76) <= layer0_outputs(4829);
    layer1_outputs(77) <= layer0_outputs(423);
    layer1_outputs(78) <= not(layer0_outputs(1306)) or (layer0_outputs(2684));
    layer1_outputs(79) <= (layer0_outputs(3029)) and not (layer0_outputs(2775));
    layer1_outputs(80) <= (layer0_outputs(2597)) or (layer0_outputs(1371));
    layer1_outputs(81) <= not(layer0_outputs(3845)) or (layer0_outputs(3492));
    layer1_outputs(82) <= (layer0_outputs(3004)) and not (layer0_outputs(2440));
    layer1_outputs(83) <= layer0_outputs(3234);
    layer1_outputs(84) <= (layer0_outputs(1345)) or (layer0_outputs(4378));
    layer1_outputs(85) <= '1';
    layer1_outputs(86) <= not(layer0_outputs(531));
    layer1_outputs(87) <= layer0_outputs(2222);
    layer1_outputs(88) <= not((layer0_outputs(4327)) and (layer0_outputs(4500)));
    layer1_outputs(89) <= layer0_outputs(58);
    layer1_outputs(90) <= (layer0_outputs(312)) and (layer0_outputs(191));
    layer1_outputs(91) <= not(layer0_outputs(4364));
    layer1_outputs(92) <= not(layer0_outputs(2502));
    layer1_outputs(93) <= (layer0_outputs(3754)) or (layer0_outputs(1180));
    layer1_outputs(94) <= layer0_outputs(3684);
    layer1_outputs(95) <= not(layer0_outputs(445));
    layer1_outputs(96) <= not((layer0_outputs(2296)) or (layer0_outputs(4672)));
    layer1_outputs(97) <= (layer0_outputs(4968)) and not (layer0_outputs(878));
    layer1_outputs(98) <= (layer0_outputs(2832)) and not (layer0_outputs(2685));
    layer1_outputs(99) <= not(layer0_outputs(1077));
    layer1_outputs(100) <= (layer0_outputs(3457)) and not (layer0_outputs(2664));
    layer1_outputs(101) <= not(layer0_outputs(3502));
    layer1_outputs(102) <= (layer0_outputs(2276)) and not (layer0_outputs(4237));
    layer1_outputs(103) <= not(layer0_outputs(3927));
    layer1_outputs(104) <= (layer0_outputs(567)) and not (layer0_outputs(167));
    layer1_outputs(105) <= not((layer0_outputs(3544)) or (layer0_outputs(5117)));
    layer1_outputs(106) <= layer0_outputs(3288);
    layer1_outputs(107) <= '0';
    layer1_outputs(108) <= (layer0_outputs(5046)) xor (layer0_outputs(805));
    layer1_outputs(109) <= not(layer0_outputs(1922));
    layer1_outputs(110) <= layer0_outputs(4324);
    layer1_outputs(111) <= '1';
    layer1_outputs(112) <= (layer0_outputs(2134)) and not (layer0_outputs(2862));
    layer1_outputs(113) <= '1';
    layer1_outputs(114) <= not((layer0_outputs(3950)) and (layer0_outputs(441)));
    layer1_outputs(115) <= (layer0_outputs(2574)) and (layer0_outputs(3964));
    layer1_outputs(116) <= not((layer0_outputs(67)) or (layer0_outputs(28)));
    layer1_outputs(117) <= layer0_outputs(2708);
    layer1_outputs(118) <= layer0_outputs(2515);
    layer1_outputs(119) <= not(layer0_outputs(3155)) or (layer0_outputs(2506));
    layer1_outputs(120) <= not(layer0_outputs(3679)) or (layer0_outputs(4434));
    layer1_outputs(121) <= layer0_outputs(2802);
    layer1_outputs(122) <= layer0_outputs(2221);
    layer1_outputs(123) <= not(layer0_outputs(168));
    layer1_outputs(124) <= '0';
    layer1_outputs(125) <= layer0_outputs(2863);
    layer1_outputs(126) <= (layer0_outputs(2836)) and not (layer0_outputs(3251));
    layer1_outputs(127) <= not(layer0_outputs(1424));
    layer1_outputs(128) <= not((layer0_outputs(2719)) and (layer0_outputs(210)));
    layer1_outputs(129) <= '1';
    layer1_outputs(130) <= not((layer0_outputs(1279)) or (layer0_outputs(4073)));
    layer1_outputs(131) <= (layer0_outputs(2771)) and (layer0_outputs(713));
    layer1_outputs(132) <= '1';
    layer1_outputs(133) <= layer0_outputs(747);
    layer1_outputs(134) <= layer0_outputs(2817);
    layer1_outputs(135) <= (layer0_outputs(147)) or (layer0_outputs(904));
    layer1_outputs(136) <= layer0_outputs(4286);
    layer1_outputs(137) <= not(layer0_outputs(4434));
    layer1_outputs(138) <= not(layer0_outputs(846)) or (layer0_outputs(3821));
    layer1_outputs(139) <= (layer0_outputs(2965)) xor (layer0_outputs(55));
    layer1_outputs(140) <= (layer0_outputs(3783)) and not (layer0_outputs(1845));
    layer1_outputs(141) <= not((layer0_outputs(2070)) and (layer0_outputs(3187)));
    layer1_outputs(142) <= layer0_outputs(4026);
    layer1_outputs(143) <= '1';
    layer1_outputs(144) <= not((layer0_outputs(156)) and (layer0_outputs(840)));
    layer1_outputs(145) <= (layer0_outputs(1352)) and not (layer0_outputs(508));
    layer1_outputs(146) <= (layer0_outputs(2136)) and not (layer0_outputs(1310));
    layer1_outputs(147) <= (layer0_outputs(170)) and (layer0_outputs(2262));
    layer1_outputs(148) <= not(layer0_outputs(3109)) or (layer0_outputs(2647));
    layer1_outputs(149) <= not(layer0_outputs(2274));
    layer1_outputs(150) <= not(layer0_outputs(1958));
    layer1_outputs(151) <= not(layer0_outputs(1021));
    layer1_outputs(152) <= (layer0_outputs(2855)) and not (layer0_outputs(4856));
    layer1_outputs(153) <= not(layer0_outputs(5008));
    layer1_outputs(154) <= layer0_outputs(2623);
    layer1_outputs(155) <= not(layer0_outputs(853));
    layer1_outputs(156) <= not(layer0_outputs(4927));
    layer1_outputs(157) <= (layer0_outputs(715)) and not (layer0_outputs(2801));
    layer1_outputs(158) <= not(layer0_outputs(1926)) or (layer0_outputs(1770));
    layer1_outputs(159) <= layer0_outputs(4448);
    layer1_outputs(160) <= not(layer0_outputs(1347)) or (layer0_outputs(3652));
    layer1_outputs(161) <= not((layer0_outputs(2933)) and (layer0_outputs(2285)));
    layer1_outputs(162) <= not(layer0_outputs(3121));
    layer1_outputs(163) <= layer0_outputs(250);
    layer1_outputs(164) <= (layer0_outputs(4851)) and (layer0_outputs(4607));
    layer1_outputs(165) <= not(layer0_outputs(4558));
    layer1_outputs(166) <= (layer0_outputs(2093)) or (layer0_outputs(1169));
    layer1_outputs(167) <= (layer0_outputs(94)) and not (layer0_outputs(2278));
    layer1_outputs(168) <= not(layer0_outputs(1976));
    layer1_outputs(169) <= (layer0_outputs(4635)) and not (layer0_outputs(2872));
    layer1_outputs(170) <= not((layer0_outputs(812)) xor (layer0_outputs(581)));
    layer1_outputs(171) <= layer0_outputs(5058);
    layer1_outputs(172) <= not(layer0_outputs(3682)) or (layer0_outputs(663));
    layer1_outputs(173) <= not(layer0_outputs(3220)) or (layer0_outputs(287));
    layer1_outputs(174) <= not(layer0_outputs(2071));
    layer1_outputs(175) <= not((layer0_outputs(2303)) or (layer0_outputs(916)));
    layer1_outputs(176) <= layer0_outputs(2292);
    layer1_outputs(177) <= not(layer0_outputs(2231)) or (layer0_outputs(563));
    layer1_outputs(178) <= layer0_outputs(4752);
    layer1_outputs(179) <= not(layer0_outputs(1508));
    layer1_outputs(180) <= not(layer0_outputs(2497));
    layer1_outputs(181) <= layer0_outputs(4279);
    layer1_outputs(182) <= not((layer0_outputs(3946)) and (layer0_outputs(4713)));
    layer1_outputs(183) <= '1';
    layer1_outputs(184) <= (layer0_outputs(735)) or (layer0_outputs(752));
    layer1_outputs(185) <= layer0_outputs(2156);
    layer1_outputs(186) <= layer0_outputs(1627);
    layer1_outputs(187) <= (layer0_outputs(1711)) and not (layer0_outputs(879));
    layer1_outputs(188) <= not(layer0_outputs(800));
    layer1_outputs(189) <= (layer0_outputs(4029)) and (layer0_outputs(2985));
    layer1_outputs(190) <= not(layer0_outputs(1292));
    layer1_outputs(191) <= (layer0_outputs(4562)) xor (layer0_outputs(2412));
    layer1_outputs(192) <= not((layer0_outputs(1146)) and (layer0_outputs(3040)));
    layer1_outputs(193) <= not(layer0_outputs(579));
    layer1_outputs(194) <= not(layer0_outputs(2919));
    layer1_outputs(195) <= not(layer0_outputs(74)) or (layer0_outputs(80));
    layer1_outputs(196) <= layer0_outputs(1563);
    layer1_outputs(197) <= not(layer0_outputs(2356)) or (layer0_outputs(3766));
    layer1_outputs(198) <= layer0_outputs(1630);
    layer1_outputs(199) <= not(layer0_outputs(2963)) or (layer0_outputs(325));
    layer1_outputs(200) <= layer0_outputs(2994);
    layer1_outputs(201) <= not(layer0_outputs(3489));
    layer1_outputs(202) <= not((layer0_outputs(2384)) or (layer0_outputs(1737)));
    layer1_outputs(203) <= layer0_outputs(3370);
    layer1_outputs(204) <= (layer0_outputs(2901)) and not (layer0_outputs(4491));
    layer1_outputs(205) <= (layer0_outputs(4688)) and (layer0_outputs(4351));
    layer1_outputs(206) <= (layer0_outputs(4472)) or (layer0_outputs(3818));
    layer1_outputs(207) <= layer0_outputs(1067);
    layer1_outputs(208) <= not(layer0_outputs(3612));
    layer1_outputs(209) <= not(layer0_outputs(3286)) or (layer0_outputs(1027));
    layer1_outputs(210) <= (layer0_outputs(2951)) and not (layer0_outputs(1330));
    layer1_outputs(211) <= (layer0_outputs(4833)) and not (layer0_outputs(1219));
    layer1_outputs(212) <= layer0_outputs(1057);
    layer1_outputs(213) <= (layer0_outputs(3788)) or (layer0_outputs(949));
    layer1_outputs(214) <= not(layer0_outputs(4629));
    layer1_outputs(215) <= not((layer0_outputs(1933)) or (layer0_outputs(2556)));
    layer1_outputs(216) <= not(layer0_outputs(3058));
    layer1_outputs(217) <= (layer0_outputs(4105)) and not (layer0_outputs(2912));
    layer1_outputs(218) <= layer0_outputs(3208);
    layer1_outputs(219) <= '1';
    layer1_outputs(220) <= '0';
    layer1_outputs(221) <= not((layer0_outputs(4793)) and (layer0_outputs(1048)));
    layer1_outputs(222) <= layer0_outputs(1393);
    layer1_outputs(223) <= '0';
    layer1_outputs(224) <= not(layer0_outputs(2117));
    layer1_outputs(225) <= not(layer0_outputs(1571)) or (layer0_outputs(2179));
    layer1_outputs(226) <= not(layer0_outputs(882));
    layer1_outputs(227) <= layer0_outputs(1977);
    layer1_outputs(228) <= not(layer0_outputs(23));
    layer1_outputs(229) <= (layer0_outputs(2619)) xor (layer0_outputs(3302));
    layer1_outputs(230) <= not(layer0_outputs(5063));
    layer1_outputs(231) <= not((layer0_outputs(1729)) xor (layer0_outputs(1742)));
    layer1_outputs(232) <= (layer0_outputs(202)) or (layer0_outputs(2310));
    layer1_outputs(233) <= layer0_outputs(1492);
    layer1_outputs(234) <= not(layer0_outputs(1726)) or (layer0_outputs(1465));
    layer1_outputs(235) <= (layer0_outputs(4234)) and not (layer0_outputs(3561));
    layer1_outputs(236) <= not(layer0_outputs(2926)) or (layer0_outputs(3450));
    layer1_outputs(237) <= layer0_outputs(2245);
    layer1_outputs(238) <= layer0_outputs(1786);
    layer1_outputs(239) <= (layer0_outputs(3955)) and not (layer0_outputs(952));
    layer1_outputs(240) <= (layer0_outputs(4411)) or (layer0_outputs(1664));
    layer1_outputs(241) <= not(layer0_outputs(1991));
    layer1_outputs(242) <= not((layer0_outputs(3697)) and (layer0_outputs(290)));
    layer1_outputs(243) <= (layer0_outputs(375)) and (layer0_outputs(601));
    layer1_outputs(244) <= not((layer0_outputs(4665)) and (layer0_outputs(4345)));
    layer1_outputs(245) <= not((layer0_outputs(518)) and (layer0_outputs(4739)));
    layer1_outputs(246) <= (layer0_outputs(713)) and (layer0_outputs(2425));
    layer1_outputs(247) <= not(layer0_outputs(994)) or (layer0_outputs(402));
    layer1_outputs(248) <= (layer0_outputs(319)) and not (layer0_outputs(1543));
    layer1_outputs(249) <= not(layer0_outputs(396));
    layer1_outputs(250) <= not(layer0_outputs(1968)) or (layer0_outputs(3099));
    layer1_outputs(251) <= layer0_outputs(1046);
    layer1_outputs(252) <= not(layer0_outputs(82));
    layer1_outputs(253) <= (layer0_outputs(2325)) and (layer0_outputs(2486));
    layer1_outputs(254) <= not(layer0_outputs(1716));
    layer1_outputs(255) <= '0';
    layer1_outputs(256) <= not(layer0_outputs(1951));
    layer1_outputs(257) <= not(layer0_outputs(5100));
    layer1_outputs(258) <= (layer0_outputs(3699)) or (layer0_outputs(126));
    layer1_outputs(259) <= not(layer0_outputs(2050));
    layer1_outputs(260) <= not(layer0_outputs(1504)) or (layer0_outputs(2637));
    layer1_outputs(261) <= not(layer0_outputs(1485));
    layer1_outputs(262) <= '1';
    layer1_outputs(263) <= (layer0_outputs(4423)) and not (layer0_outputs(3985));
    layer1_outputs(264) <= layer0_outputs(372);
    layer1_outputs(265) <= layer0_outputs(1505);
    layer1_outputs(266) <= (layer0_outputs(3446)) or (layer0_outputs(4521));
    layer1_outputs(267) <= not(layer0_outputs(1490)) or (layer0_outputs(135));
    layer1_outputs(268) <= (layer0_outputs(2895)) and (layer0_outputs(121));
    layer1_outputs(269) <= (layer0_outputs(128)) and not (layer0_outputs(300));
    layer1_outputs(270) <= not(layer0_outputs(4048));
    layer1_outputs(271) <= not((layer0_outputs(1004)) and (layer0_outputs(1397)));
    layer1_outputs(272) <= not(layer0_outputs(2888)) or (layer0_outputs(2802));
    layer1_outputs(273) <= not(layer0_outputs(1141));
    layer1_outputs(274) <= '0';
    layer1_outputs(275) <= not(layer0_outputs(1582));
    layer1_outputs(276) <= not(layer0_outputs(3098)) or (layer0_outputs(3284));
    layer1_outputs(277) <= not((layer0_outputs(703)) xor (layer0_outputs(996)));
    layer1_outputs(278) <= not((layer0_outputs(2251)) and (layer0_outputs(2601)));
    layer1_outputs(279) <= not(layer0_outputs(44));
    layer1_outputs(280) <= not(layer0_outputs(3017));
    layer1_outputs(281) <= layer0_outputs(1636);
    layer1_outputs(282) <= (layer0_outputs(1128)) or (layer0_outputs(1050));
    layer1_outputs(283) <= (layer0_outputs(73)) and not (layer0_outputs(2609));
    layer1_outputs(284) <= not((layer0_outputs(5106)) and (layer0_outputs(1642)));
    layer1_outputs(285) <= '1';
    layer1_outputs(286) <= layer0_outputs(757);
    layer1_outputs(287) <= layer0_outputs(3653);
    layer1_outputs(288) <= layer0_outputs(1489);
    layer1_outputs(289) <= layer0_outputs(4841);
    layer1_outputs(290) <= not(layer0_outputs(4760));
    layer1_outputs(291) <= '1';
    layer1_outputs(292) <= not(layer0_outputs(2765));
    layer1_outputs(293) <= not(layer0_outputs(17)) or (layer0_outputs(1442));
    layer1_outputs(294) <= not(layer0_outputs(3438)) or (layer0_outputs(884));
    layer1_outputs(295) <= '0';
    layer1_outputs(296) <= layer0_outputs(4022);
    layer1_outputs(297) <= not(layer0_outputs(2630));
    layer1_outputs(298) <= not((layer0_outputs(2187)) or (layer0_outputs(2402)));
    layer1_outputs(299) <= (layer0_outputs(4860)) and (layer0_outputs(4471));
    layer1_outputs(300) <= '0';
    layer1_outputs(301) <= layer0_outputs(4042);
    layer1_outputs(302) <= (layer0_outputs(3222)) and not (layer0_outputs(604));
    layer1_outputs(303) <= (layer0_outputs(3775)) or (layer0_outputs(1629));
    layer1_outputs(304) <= layer0_outputs(1863);
    layer1_outputs(305) <= (layer0_outputs(2657)) and not (layer0_outputs(4070));
    layer1_outputs(306) <= layer0_outputs(9);
    layer1_outputs(307) <= not(layer0_outputs(4897));
    layer1_outputs(308) <= (layer0_outputs(2522)) xor (layer0_outputs(4228));
    layer1_outputs(309) <= not(layer0_outputs(2650));
    layer1_outputs(310) <= layer0_outputs(3434);
    layer1_outputs(311) <= not(layer0_outputs(4981));
    layer1_outputs(312) <= (layer0_outputs(1980)) and (layer0_outputs(1590));
    layer1_outputs(313) <= not(layer0_outputs(2366));
    layer1_outputs(314) <= not(layer0_outputs(1593)) or (layer0_outputs(2682));
    layer1_outputs(315) <= not(layer0_outputs(4595));
    layer1_outputs(316) <= not(layer0_outputs(2383)) or (layer0_outputs(1920));
    layer1_outputs(317) <= layer0_outputs(627);
    layer1_outputs(318) <= (layer0_outputs(1470)) and not (layer0_outputs(5064));
    layer1_outputs(319) <= (layer0_outputs(1405)) and (layer0_outputs(2876));
    layer1_outputs(320) <= (layer0_outputs(3139)) xor (layer0_outputs(945));
    layer1_outputs(321) <= not(layer0_outputs(696));
    layer1_outputs(322) <= (layer0_outputs(4940)) and not (layer0_outputs(2167));
    layer1_outputs(323) <= not((layer0_outputs(228)) and (layer0_outputs(958)));
    layer1_outputs(324) <= layer0_outputs(1158);
    layer1_outputs(325) <= layer0_outputs(4123);
    layer1_outputs(326) <= not(layer0_outputs(3320));
    layer1_outputs(327) <= layer0_outputs(836);
    layer1_outputs(328) <= not(layer0_outputs(32)) or (layer0_outputs(505));
    layer1_outputs(329) <= not((layer0_outputs(783)) or (layer0_outputs(677)));
    layer1_outputs(330) <= (layer0_outputs(2402)) and not (layer0_outputs(4565));
    layer1_outputs(331) <= layer0_outputs(4276);
    layer1_outputs(332) <= (layer0_outputs(2942)) xor (layer0_outputs(1519));
    layer1_outputs(333) <= layer0_outputs(3239);
    layer1_outputs(334) <= layer0_outputs(2816);
    layer1_outputs(335) <= layer0_outputs(4236);
    layer1_outputs(336) <= (layer0_outputs(3696)) and (layer0_outputs(1054));
    layer1_outputs(337) <= not((layer0_outputs(1643)) or (layer0_outputs(2988)));
    layer1_outputs(338) <= not(layer0_outputs(2364)) or (layer0_outputs(3607));
    layer1_outputs(339) <= layer0_outputs(1312);
    layer1_outputs(340) <= not(layer0_outputs(427)) or (layer0_outputs(2449));
    layer1_outputs(341) <= (layer0_outputs(1782)) and not (layer0_outputs(3751));
    layer1_outputs(342) <= layer0_outputs(4008);
    layer1_outputs(343) <= not(layer0_outputs(3116)) or (layer0_outputs(3149));
    layer1_outputs(344) <= (layer0_outputs(9)) and (layer0_outputs(3218));
    layer1_outputs(345) <= layer0_outputs(5031);
    layer1_outputs(346) <= (layer0_outputs(1847)) and not (layer0_outputs(883));
    layer1_outputs(347) <= not(layer0_outputs(3930));
    layer1_outputs(348) <= not((layer0_outputs(4309)) or (layer0_outputs(720)));
    layer1_outputs(349) <= not(layer0_outputs(4279));
    layer1_outputs(350) <= layer0_outputs(2720);
    layer1_outputs(351) <= not(layer0_outputs(4657));
    layer1_outputs(352) <= not(layer0_outputs(4763)) or (layer0_outputs(4798));
    layer1_outputs(353) <= layer0_outputs(435);
    layer1_outputs(354) <= not(layer0_outputs(4026)) or (layer0_outputs(5054));
    layer1_outputs(355) <= layer0_outputs(1949);
    layer1_outputs(356) <= '1';
    layer1_outputs(357) <= not((layer0_outputs(2482)) and (layer0_outputs(3137)));
    layer1_outputs(358) <= layer0_outputs(2499);
    layer1_outputs(359) <= (layer0_outputs(3120)) xor (layer0_outputs(154));
    layer1_outputs(360) <= not(layer0_outputs(1009));
    layer1_outputs(361) <= not(layer0_outputs(2041));
    layer1_outputs(362) <= not(layer0_outputs(492));
    layer1_outputs(363) <= (layer0_outputs(4401)) and not (layer0_outputs(1213));
    layer1_outputs(364) <= (layer0_outputs(4094)) and not (layer0_outputs(5039));
    layer1_outputs(365) <= not((layer0_outputs(5052)) and (layer0_outputs(2876)));
    layer1_outputs(366) <= (layer0_outputs(3827)) and (layer0_outputs(5019));
    layer1_outputs(367) <= not((layer0_outputs(4888)) and (layer0_outputs(4405)));
    layer1_outputs(368) <= layer0_outputs(1185);
    layer1_outputs(369) <= layer0_outputs(222);
    layer1_outputs(370) <= (layer0_outputs(4503)) and not (layer0_outputs(2838));
    layer1_outputs(371) <= layer0_outputs(4197);
    layer1_outputs(372) <= layer0_outputs(3373);
    layer1_outputs(373) <= not(layer0_outputs(3623));
    layer1_outputs(374) <= layer0_outputs(700);
    layer1_outputs(375) <= layer0_outputs(349);
    layer1_outputs(376) <= layer0_outputs(1209);
    layer1_outputs(377) <= '1';
    layer1_outputs(378) <= (layer0_outputs(1999)) or (layer0_outputs(392));
    layer1_outputs(379) <= layer0_outputs(1016);
    layer1_outputs(380) <= not(layer0_outputs(4386)) or (layer0_outputs(1217));
    layer1_outputs(381) <= (layer0_outputs(3030)) and (layer0_outputs(1864));
    layer1_outputs(382) <= layer0_outputs(3466);
    layer1_outputs(383) <= not(layer0_outputs(2609));
    layer1_outputs(384) <= layer0_outputs(1380);
    layer1_outputs(385) <= (layer0_outputs(3716)) xor (layer0_outputs(753));
    layer1_outputs(386) <= (layer0_outputs(632)) and (layer0_outputs(3742));
    layer1_outputs(387) <= not((layer0_outputs(1045)) or (layer0_outputs(4251)));
    layer1_outputs(388) <= not(layer0_outputs(3422)) or (layer0_outputs(14));
    layer1_outputs(389) <= not(layer0_outputs(2132)) or (layer0_outputs(4623));
    layer1_outputs(390) <= layer0_outputs(543);
    layer1_outputs(391) <= layer0_outputs(1312);
    layer1_outputs(392) <= layer0_outputs(2874);
    layer1_outputs(393) <= layer0_outputs(3388);
    layer1_outputs(394) <= layer0_outputs(1231);
    layer1_outputs(395) <= not((layer0_outputs(3425)) xor (layer0_outputs(796)));
    layer1_outputs(396) <= not((layer0_outputs(3695)) and (layer0_outputs(3133)));
    layer1_outputs(397) <= (layer0_outputs(353)) or (layer0_outputs(1430));
    layer1_outputs(398) <= (layer0_outputs(204)) and not (layer0_outputs(72));
    layer1_outputs(399) <= layer0_outputs(640);
    layer1_outputs(400) <= (layer0_outputs(3515)) and not (layer0_outputs(1717));
    layer1_outputs(401) <= layer0_outputs(1226);
    layer1_outputs(402) <= (layer0_outputs(4814)) and not (layer0_outputs(1547));
    layer1_outputs(403) <= layer0_outputs(2859);
    layer1_outputs(404) <= not(layer0_outputs(4331)) or (layer0_outputs(4835));
    layer1_outputs(405) <= not(layer0_outputs(4417));
    layer1_outputs(406) <= '0';
    layer1_outputs(407) <= (layer0_outputs(3338)) and (layer0_outputs(3311));
    layer1_outputs(408) <= layer0_outputs(3566);
    layer1_outputs(409) <= (layer0_outputs(2675)) xor (layer0_outputs(2938));
    layer1_outputs(410) <= (layer0_outputs(5077)) and (layer0_outputs(986));
    layer1_outputs(411) <= (layer0_outputs(4048)) and not (layer0_outputs(1970));
    layer1_outputs(412) <= (layer0_outputs(4838)) and (layer0_outputs(4855));
    layer1_outputs(413) <= not(layer0_outputs(2357)) or (layer0_outputs(422));
    layer1_outputs(414) <= not((layer0_outputs(4288)) xor (layer0_outputs(3787)));
    layer1_outputs(415) <= not(layer0_outputs(1400));
    layer1_outputs(416) <= (layer0_outputs(4325)) and not (layer0_outputs(3626));
    layer1_outputs(417) <= layer0_outputs(4728);
    layer1_outputs(418) <= not((layer0_outputs(1538)) or (layer0_outputs(178)));
    layer1_outputs(419) <= '1';
    layer1_outputs(420) <= not(layer0_outputs(3956)) or (layer0_outputs(2432));
    layer1_outputs(421) <= not((layer0_outputs(4706)) and (layer0_outputs(1435)));
    layer1_outputs(422) <= not((layer0_outputs(1911)) or (layer0_outputs(4861)));
    layer1_outputs(423) <= layer0_outputs(758);
    layer1_outputs(424) <= not((layer0_outputs(3010)) xor (layer0_outputs(4992)));
    layer1_outputs(425) <= layer0_outputs(4951);
    layer1_outputs(426) <= not(layer0_outputs(4411));
    layer1_outputs(427) <= (layer0_outputs(3490)) or (layer0_outputs(2413));
    layer1_outputs(428) <= not(layer0_outputs(3037)) or (layer0_outputs(258));
    layer1_outputs(429) <= not((layer0_outputs(2960)) and (layer0_outputs(4683)));
    layer1_outputs(430) <= layer0_outputs(2858);
    layer1_outputs(431) <= not(layer0_outputs(4587)) or (layer0_outputs(3053));
    layer1_outputs(432) <= not(layer0_outputs(2579)) or (layer0_outputs(2907));
    layer1_outputs(433) <= not(layer0_outputs(3671));
    layer1_outputs(434) <= (layer0_outputs(939)) xor (layer0_outputs(1075));
    layer1_outputs(435) <= layer0_outputs(2620);
    layer1_outputs(436) <= not(layer0_outputs(4461));
    layer1_outputs(437) <= (layer0_outputs(1385)) and not (layer0_outputs(2556));
    layer1_outputs(438) <= not(layer0_outputs(662)) or (layer0_outputs(2910));
    layer1_outputs(439) <= (layer0_outputs(190)) and (layer0_outputs(3800));
    layer1_outputs(440) <= not(layer0_outputs(2102));
    layer1_outputs(441) <= (layer0_outputs(3129)) and (layer0_outputs(3726));
    layer1_outputs(442) <= layer0_outputs(942);
    layer1_outputs(443) <= (layer0_outputs(4290)) and not (layer0_outputs(470));
    layer1_outputs(444) <= not(layer0_outputs(1169)) or (layer0_outputs(2422));
    layer1_outputs(445) <= not(layer0_outputs(3220)) or (layer0_outputs(3252));
    layer1_outputs(446) <= not((layer0_outputs(2623)) or (layer0_outputs(2287)));
    layer1_outputs(447) <= not(layer0_outputs(3399));
    layer1_outputs(448) <= not((layer0_outputs(4212)) or (layer0_outputs(424)));
    layer1_outputs(449) <= not(layer0_outputs(1596)) or (layer0_outputs(1806));
    layer1_outputs(450) <= (layer0_outputs(1321)) and not (layer0_outputs(899));
    layer1_outputs(451) <= (layer0_outputs(998)) and not (layer0_outputs(3600));
    layer1_outputs(452) <= not(layer0_outputs(3909)) or (layer0_outputs(1796));
    layer1_outputs(453) <= layer0_outputs(2200);
    layer1_outputs(454) <= (layer0_outputs(1346)) and not (layer0_outputs(428));
    layer1_outputs(455) <= '1';
    layer1_outputs(456) <= not(layer0_outputs(689)) or (layer0_outputs(4442));
    layer1_outputs(457) <= not(layer0_outputs(4110));
    layer1_outputs(458) <= not(layer0_outputs(1628));
    layer1_outputs(459) <= not(layer0_outputs(1223));
    layer1_outputs(460) <= not((layer0_outputs(1280)) and (layer0_outputs(2571)));
    layer1_outputs(461) <= (layer0_outputs(1423)) and (layer0_outputs(530));
    layer1_outputs(462) <= '1';
    layer1_outputs(463) <= not(layer0_outputs(2783)) or (layer0_outputs(4452));
    layer1_outputs(464) <= not(layer0_outputs(84));
    layer1_outputs(465) <= not(layer0_outputs(311));
    layer1_outputs(466) <= not((layer0_outputs(2171)) or (layer0_outputs(673)));
    layer1_outputs(467) <= (layer0_outputs(1195)) or (layer0_outputs(3852));
    layer1_outputs(468) <= '1';
    layer1_outputs(469) <= not((layer0_outputs(1979)) and (layer0_outputs(1804)));
    layer1_outputs(470) <= layer0_outputs(3976);
    layer1_outputs(471) <= '0';
    layer1_outputs(472) <= layer0_outputs(1182);
    layer1_outputs(473) <= not(layer0_outputs(4174));
    layer1_outputs(474) <= not((layer0_outputs(3072)) or (layer0_outputs(1861)));
    layer1_outputs(475) <= not((layer0_outputs(3619)) or (layer0_outputs(4229)));
    layer1_outputs(476) <= (layer0_outputs(4429)) or (layer0_outputs(1776));
    layer1_outputs(477) <= not((layer0_outputs(526)) xor (layer0_outputs(2371)));
    layer1_outputs(478) <= layer0_outputs(1101);
    layer1_outputs(479) <= not(layer0_outputs(520));
    layer1_outputs(480) <= layer0_outputs(1362);
    layer1_outputs(481) <= layer0_outputs(1728);
    layer1_outputs(482) <= (layer0_outputs(2255)) and not (layer0_outputs(5018));
    layer1_outputs(483) <= not((layer0_outputs(3823)) xor (layer0_outputs(1539)));
    layer1_outputs(484) <= not(layer0_outputs(1142)) or (layer0_outputs(4012));
    layer1_outputs(485) <= '0';
    layer1_outputs(486) <= (layer0_outputs(3333)) and not (layer0_outputs(4267));
    layer1_outputs(487) <= (layer0_outputs(2466)) xor (layer0_outputs(2893));
    layer1_outputs(488) <= layer0_outputs(4787);
    layer1_outputs(489) <= not((layer0_outputs(1306)) or (layer0_outputs(4853)));
    layer1_outputs(490) <= not(layer0_outputs(1165));
    layer1_outputs(491) <= layer0_outputs(4907);
    layer1_outputs(492) <= not(layer0_outputs(4394)) or (layer0_outputs(454));
    layer1_outputs(493) <= layer0_outputs(2256);
    layer1_outputs(494) <= not(layer0_outputs(2186));
    layer1_outputs(495) <= '1';
    layer1_outputs(496) <= (layer0_outputs(4208)) or (layer0_outputs(4291));
    layer1_outputs(497) <= not((layer0_outputs(585)) and (layer0_outputs(2960)));
    layer1_outputs(498) <= layer0_outputs(2978);
    layer1_outputs(499) <= not(layer0_outputs(2507));
    layer1_outputs(500) <= not(layer0_outputs(2018));
    layer1_outputs(501) <= not((layer0_outputs(2033)) xor (layer0_outputs(3068)));
    layer1_outputs(502) <= not(layer0_outputs(1982)) or (layer0_outputs(1453));
    layer1_outputs(503) <= not(layer0_outputs(4586));
    layer1_outputs(504) <= not(layer0_outputs(784));
    layer1_outputs(505) <= not(layer0_outputs(4128));
    layer1_outputs(506) <= (layer0_outputs(3935)) and not (layer0_outputs(3572));
    layer1_outputs(507) <= not((layer0_outputs(4973)) xor (layer0_outputs(2967)));
    layer1_outputs(508) <= '0';
    layer1_outputs(509) <= not(layer0_outputs(2041)) or (layer0_outputs(2237));
    layer1_outputs(510) <= (layer0_outputs(2924)) and not (layer0_outputs(1955));
    layer1_outputs(511) <= not(layer0_outputs(2214));
    layer1_outputs(512) <= (layer0_outputs(3853)) and not (layer0_outputs(3989));
    layer1_outputs(513) <= not(layer0_outputs(3829));
    layer1_outputs(514) <= not(layer0_outputs(359));
    layer1_outputs(515) <= (layer0_outputs(3647)) and not (layer0_outputs(1664));
    layer1_outputs(516) <= (layer0_outputs(4472)) and not (layer0_outputs(2992));
    layer1_outputs(517) <= not(layer0_outputs(1785));
    layer1_outputs(518) <= (layer0_outputs(2584)) or (layer0_outputs(1316));
    layer1_outputs(519) <= not((layer0_outputs(3049)) or (layer0_outputs(4377)));
    layer1_outputs(520) <= layer0_outputs(1467);
    layer1_outputs(521) <= not((layer0_outputs(4098)) and (layer0_outputs(848)));
    layer1_outputs(522) <= (layer0_outputs(4601)) xor (layer0_outputs(2655));
    layer1_outputs(523) <= layer0_outputs(1879);
    layer1_outputs(524) <= not((layer0_outputs(4685)) xor (layer0_outputs(1252)));
    layer1_outputs(525) <= not((layer0_outputs(871)) and (layer0_outputs(4482)));
    layer1_outputs(526) <= not(layer0_outputs(947)) or (layer0_outputs(1292));
    layer1_outputs(527) <= not(layer0_outputs(4363)) or (layer0_outputs(2751));
    layer1_outputs(528) <= (layer0_outputs(1514)) or (layer0_outputs(503));
    layer1_outputs(529) <= not(layer0_outputs(3753)) or (layer0_outputs(447));
    layer1_outputs(530) <= not((layer0_outputs(3267)) or (layer0_outputs(2759)));
    layer1_outputs(531) <= '0';
    layer1_outputs(532) <= (layer0_outputs(5024)) and (layer0_outputs(3949));
    layer1_outputs(533) <= not(layer0_outputs(3645));
    layer1_outputs(534) <= not(layer0_outputs(2123));
    layer1_outputs(535) <= not(layer0_outputs(3200));
    layer1_outputs(536) <= '1';
    layer1_outputs(537) <= (layer0_outputs(4817)) or (layer0_outputs(4957));
    layer1_outputs(538) <= not((layer0_outputs(534)) and (layer0_outputs(3397)));
    layer1_outputs(539) <= '1';
    layer1_outputs(540) <= not((layer0_outputs(3332)) and (layer0_outputs(1623)));
    layer1_outputs(541) <= not(layer0_outputs(3189)) or (layer0_outputs(4333));
    layer1_outputs(542) <= layer0_outputs(2625);
    layer1_outputs(543) <= not(layer0_outputs(3883));
    layer1_outputs(544) <= not((layer0_outputs(737)) xor (layer0_outputs(4086)));
    layer1_outputs(545) <= not((layer0_outputs(1408)) xor (layer0_outputs(1115)));
    layer1_outputs(546) <= not((layer0_outputs(2180)) or (layer0_outputs(3824)));
    layer1_outputs(547) <= layer0_outputs(3877);
    layer1_outputs(548) <= not(layer0_outputs(2806)) or (layer0_outputs(4716));
    layer1_outputs(549) <= layer0_outputs(2698);
    layer1_outputs(550) <= (layer0_outputs(1015)) xor (layer0_outputs(931));
    layer1_outputs(551) <= not(layer0_outputs(3535));
    layer1_outputs(552) <= (layer0_outputs(2340)) or (layer0_outputs(519));
    layer1_outputs(553) <= not(layer0_outputs(4694));
    layer1_outputs(554) <= not(layer0_outputs(1331));
    layer1_outputs(555) <= layer0_outputs(772);
    layer1_outputs(556) <= (layer0_outputs(3606)) and not (layer0_outputs(3182));
    layer1_outputs(557) <= not(layer0_outputs(4418));
    layer1_outputs(558) <= not(layer0_outputs(3709)) or (layer0_outputs(3314));
    layer1_outputs(559) <= not(layer0_outputs(438));
    layer1_outputs(560) <= not(layer0_outputs(809));
    layer1_outputs(561) <= (layer0_outputs(3126)) or (layer0_outputs(4525));
    layer1_outputs(562) <= (layer0_outputs(120)) and not (layer0_outputs(4963));
    layer1_outputs(563) <= not((layer0_outputs(1188)) and (layer0_outputs(2289)));
    layer1_outputs(564) <= not(layer0_outputs(274));
    layer1_outputs(565) <= not((layer0_outputs(2738)) and (layer0_outputs(1204)));
    layer1_outputs(566) <= layer0_outputs(769);
    layer1_outputs(567) <= layer0_outputs(2621);
    layer1_outputs(568) <= not(layer0_outputs(5082)) or (layer0_outputs(4532));
    layer1_outputs(569) <= not((layer0_outputs(4040)) or (layer0_outputs(4605)));
    layer1_outputs(570) <= not(layer0_outputs(3832));
    layer1_outputs(571) <= '0';
    layer1_outputs(572) <= layer0_outputs(4238);
    layer1_outputs(573) <= layer0_outputs(4294);
    layer1_outputs(574) <= not(layer0_outputs(4923)) or (layer0_outputs(2150));
    layer1_outputs(575) <= not(layer0_outputs(2540)) or (layer0_outputs(4581));
    layer1_outputs(576) <= layer0_outputs(4791);
    layer1_outputs(577) <= (layer0_outputs(4157)) and not (layer0_outputs(2188));
    layer1_outputs(578) <= (layer0_outputs(3698)) and not (layer0_outputs(3703));
    layer1_outputs(579) <= not(layer0_outputs(4468)) or (layer0_outputs(1729));
    layer1_outputs(580) <= not(layer0_outputs(787)) or (layer0_outputs(2841));
    layer1_outputs(581) <= not((layer0_outputs(232)) and (layer0_outputs(2945)));
    layer1_outputs(582) <= not(layer0_outputs(3474)) or (layer0_outputs(395));
    layer1_outputs(583) <= not(layer0_outputs(1732));
    layer1_outputs(584) <= (layer0_outputs(2016)) and not (layer0_outputs(3508));
    layer1_outputs(585) <= not((layer0_outputs(242)) and (layer0_outputs(941)));
    layer1_outputs(586) <= not(layer0_outputs(3549)) or (layer0_outputs(603));
    layer1_outputs(587) <= (layer0_outputs(1293)) or (layer0_outputs(4615));
    layer1_outputs(588) <= not(layer0_outputs(3328));
    layer1_outputs(589) <= not(layer0_outputs(572));
    layer1_outputs(590) <= (layer0_outputs(3283)) and not (layer0_outputs(4064));
    layer1_outputs(591) <= '0';
    layer1_outputs(592) <= not(layer0_outputs(3869)) or (layer0_outputs(4002));
    layer1_outputs(593) <= (layer0_outputs(4719)) or (layer0_outputs(4999));
    layer1_outputs(594) <= (layer0_outputs(2605)) and not (layer0_outputs(3598));
    layer1_outputs(595) <= (layer0_outputs(3406)) and (layer0_outputs(3230));
    layer1_outputs(596) <= (layer0_outputs(2835)) and (layer0_outputs(4172));
    layer1_outputs(597) <= not((layer0_outputs(5078)) and (layer0_outputs(4421)));
    layer1_outputs(598) <= (layer0_outputs(2056)) and not (layer0_outputs(1674));
    layer1_outputs(599) <= not((layer0_outputs(3792)) and (layer0_outputs(1632)));
    layer1_outputs(600) <= layer0_outputs(1297);
    layer1_outputs(601) <= layer0_outputs(5049);
    layer1_outputs(602) <= not(layer0_outputs(1024));
    layer1_outputs(603) <= not(layer0_outputs(892));
    layer1_outputs(604) <= layer0_outputs(5109);
    layer1_outputs(605) <= not(layer0_outputs(1153)) or (layer0_outputs(1944));
    layer1_outputs(606) <= not(layer0_outputs(1597)) or (layer0_outputs(3318));
    layer1_outputs(607) <= (layer0_outputs(4598)) and not (layer0_outputs(3016));
    layer1_outputs(608) <= '0';
    layer1_outputs(609) <= '0';
    layer1_outputs(610) <= (layer0_outputs(3768)) and not (layer0_outputs(1076));
    layer1_outputs(611) <= not(layer0_outputs(4816));
    layer1_outputs(612) <= not((layer0_outputs(14)) or (layer0_outputs(4270)));
    layer1_outputs(613) <= '1';
    layer1_outputs(614) <= not(layer0_outputs(1858)) or (layer0_outputs(499));
    layer1_outputs(615) <= not((layer0_outputs(1219)) or (layer0_outputs(2873)));
    layer1_outputs(616) <= (layer0_outputs(1802)) or (layer0_outputs(4013));
    layer1_outputs(617) <= not(layer0_outputs(3619)) or (layer0_outputs(794));
    layer1_outputs(618) <= not(layer0_outputs(875));
    layer1_outputs(619) <= layer0_outputs(286);
    layer1_outputs(620) <= not((layer0_outputs(977)) and (layer0_outputs(3292)));
    layer1_outputs(621) <= not(layer0_outputs(776));
    layer1_outputs(622) <= not((layer0_outputs(1405)) and (layer0_outputs(2065)));
    layer1_outputs(623) <= not((layer0_outputs(952)) and (layer0_outputs(4384)));
    layer1_outputs(624) <= layer0_outputs(4285);
    layer1_outputs(625) <= layer0_outputs(4112);
    layer1_outputs(626) <= not(layer0_outputs(1706)) or (layer0_outputs(3523));
    layer1_outputs(627) <= layer0_outputs(2569);
    layer1_outputs(628) <= layer0_outputs(2881);
    layer1_outputs(629) <= layer0_outputs(3841);
    layer1_outputs(630) <= not(layer0_outputs(4738)) or (layer0_outputs(2654));
    layer1_outputs(631) <= '1';
    layer1_outputs(632) <= not((layer0_outputs(1052)) or (layer0_outputs(2226)));
    layer1_outputs(633) <= not((layer0_outputs(2391)) and (layer0_outputs(4173)));
    layer1_outputs(634) <= (layer0_outputs(4904)) and (layer0_outputs(1922));
    layer1_outputs(635) <= not((layer0_outputs(2045)) xor (layer0_outputs(3092)));
    layer1_outputs(636) <= not(layer0_outputs(2714));
    layer1_outputs(637) <= not(layer0_outputs(137));
    layer1_outputs(638) <= not(layer0_outputs(1631)) or (layer0_outputs(3798));
    layer1_outputs(639) <= '1';
    layer1_outputs(640) <= not(layer0_outputs(4680));
    layer1_outputs(641) <= (layer0_outputs(385)) or (layer0_outputs(5088));
    layer1_outputs(642) <= (layer0_outputs(2377)) or (layer0_outputs(1640));
    layer1_outputs(643) <= layer0_outputs(651);
    layer1_outputs(644) <= (layer0_outputs(1787)) and (layer0_outputs(3110));
    layer1_outputs(645) <= not(layer0_outputs(4621));
    layer1_outputs(646) <= not(layer0_outputs(2135));
    layer1_outputs(647) <= layer0_outputs(4785);
    layer1_outputs(648) <= not(layer0_outputs(724)) or (layer0_outputs(427));
    layer1_outputs(649) <= (layer0_outputs(1684)) and not (layer0_outputs(3142));
    layer1_outputs(650) <= layer0_outputs(299);
    layer1_outputs(651) <= not(layer0_outputs(2820)) or (layer0_outputs(2126));
    layer1_outputs(652) <= (layer0_outputs(1037)) xor (layer0_outputs(1074));
    layer1_outputs(653) <= (layer0_outputs(4872)) or (layer0_outputs(4422));
    layer1_outputs(654) <= (layer0_outputs(1547)) and not (layer0_outputs(1273));
    layer1_outputs(655) <= (layer0_outputs(1515)) and (layer0_outputs(5016));
    layer1_outputs(656) <= not(layer0_outputs(921));
    layer1_outputs(657) <= layer0_outputs(5056);
    layer1_outputs(658) <= (layer0_outputs(705)) and not (layer0_outputs(4956));
    layer1_outputs(659) <= (layer0_outputs(4400)) or (layer0_outputs(481));
    layer1_outputs(660) <= (layer0_outputs(3685)) or (layer0_outputs(2407));
    layer1_outputs(661) <= layer0_outputs(112);
    layer1_outputs(662) <= '1';
    layer1_outputs(663) <= layer0_outputs(4780);
    layer1_outputs(664) <= not(layer0_outputs(3995));
    layer1_outputs(665) <= (layer0_outputs(4451)) and (layer0_outputs(4742));
    layer1_outputs(666) <= (layer0_outputs(2733)) and not (layer0_outputs(4991));
    layer1_outputs(667) <= not(layer0_outputs(3332));
    layer1_outputs(668) <= not((layer0_outputs(4464)) and (layer0_outputs(3774)));
    layer1_outputs(669) <= layer0_outputs(2917);
    layer1_outputs(670) <= not(layer0_outputs(2339));
    layer1_outputs(671) <= not(layer0_outputs(4574));
    layer1_outputs(672) <= not(layer0_outputs(585)) or (layer0_outputs(1890));
    layer1_outputs(673) <= not(layer0_outputs(3245)) or (layer0_outputs(326));
    layer1_outputs(674) <= not(layer0_outputs(226)) or (layer0_outputs(4006));
    layer1_outputs(675) <= layer0_outputs(3535);
    layer1_outputs(676) <= layer0_outputs(2794);
    layer1_outputs(677) <= not(layer0_outputs(1705));
    layer1_outputs(678) <= (layer0_outputs(4438)) xor (layer0_outputs(4828));
    layer1_outputs(679) <= (layer0_outputs(3803)) and not (layer0_outputs(4733));
    layer1_outputs(680) <= layer0_outputs(642);
    layer1_outputs(681) <= layer0_outputs(74);
    layer1_outputs(682) <= (layer0_outputs(1179)) xor (layer0_outputs(2125));
    layer1_outputs(683) <= not(layer0_outputs(4379)) or (layer0_outputs(4366));
    layer1_outputs(684) <= not(layer0_outputs(4344));
    layer1_outputs(685) <= not((layer0_outputs(2899)) or (layer0_outputs(874)));
    layer1_outputs(686) <= not((layer0_outputs(1378)) and (layer0_outputs(959)));
    layer1_outputs(687) <= (layer0_outputs(4816)) and (layer0_outputs(2477));
    layer1_outputs(688) <= not((layer0_outputs(4775)) and (layer0_outputs(3901)));
    layer1_outputs(689) <= not((layer0_outputs(1848)) and (layer0_outputs(3350)));
    layer1_outputs(690) <= not(layer0_outputs(1310));
    layer1_outputs(691) <= (layer0_outputs(2881)) or (layer0_outputs(4961));
    layer1_outputs(692) <= layer0_outputs(4360);
    layer1_outputs(693) <= not((layer0_outputs(198)) and (layer0_outputs(231)));
    layer1_outputs(694) <= (layer0_outputs(507)) or (layer0_outputs(132));
    layer1_outputs(695) <= not(layer0_outputs(2052));
    layer1_outputs(696) <= not(layer0_outputs(1396));
    layer1_outputs(697) <= not((layer0_outputs(3095)) or (layer0_outputs(4501)));
    layer1_outputs(698) <= not(layer0_outputs(877)) or (layer0_outputs(5025));
    layer1_outputs(699) <= not(layer0_outputs(3948)) or (layer0_outputs(2659));
    layer1_outputs(700) <= '1';
    layer1_outputs(701) <= (layer0_outputs(1510)) and not (layer0_outputs(4370));
    layer1_outputs(702) <= layer0_outputs(4426);
    layer1_outputs(703) <= not(layer0_outputs(4523)) or (layer0_outputs(4836));
    layer1_outputs(704) <= not(layer0_outputs(3588));
    layer1_outputs(705) <= not(layer0_outputs(2204)) or (layer0_outputs(1651));
    layer1_outputs(706) <= not(layer0_outputs(3951)) or (layer0_outputs(563));
    layer1_outputs(707) <= (layer0_outputs(1136)) and not (layer0_outputs(1381));
    layer1_outputs(708) <= not(layer0_outputs(3574));
    layer1_outputs(709) <= not(layer0_outputs(1887));
    layer1_outputs(710) <= not((layer0_outputs(3327)) and (layer0_outputs(2447)));
    layer1_outputs(711) <= layer0_outputs(1554);
    layer1_outputs(712) <= layer0_outputs(1983);
    layer1_outputs(713) <= (layer0_outputs(3398)) and not (layer0_outputs(4145));
    layer1_outputs(714) <= layer0_outputs(4866);
    layer1_outputs(715) <= not(layer0_outputs(2172));
    layer1_outputs(716) <= not((layer0_outputs(4907)) and (layer0_outputs(4118)));
    layer1_outputs(717) <= layer0_outputs(1519);
    layer1_outputs(718) <= layer0_outputs(1910);
    layer1_outputs(719) <= '1';
    layer1_outputs(720) <= (layer0_outputs(793)) xor (layer0_outputs(2964));
    layer1_outputs(721) <= not((layer0_outputs(3826)) or (layer0_outputs(2855)));
    layer1_outputs(722) <= not(layer0_outputs(3051));
    layer1_outputs(723) <= not(layer0_outputs(2271)) or (layer0_outputs(1236));
    layer1_outputs(724) <= not(layer0_outputs(958));
    layer1_outputs(725) <= not(layer0_outputs(1939));
    layer1_outputs(726) <= (layer0_outputs(157)) and (layer0_outputs(4505));
    layer1_outputs(727) <= layer0_outputs(618);
    layer1_outputs(728) <= layer0_outputs(1992);
    layer1_outputs(729) <= not(layer0_outputs(867));
    layer1_outputs(730) <= (layer0_outputs(986)) and (layer0_outputs(3551));
    layer1_outputs(731) <= not(layer0_outputs(3064));
    layer1_outputs(732) <= not(layer0_outputs(2983));
    layer1_outputs(733) <= (layer0_outputs(4917)) and (layer0_outputs(4268));
    layer1_outputs(734) <= layer0_outputs(4462);
    layer1_outputs(735) <= not(layer0_outputs(3971));
    layer1_outputs(736) <= (layer0_outputs(2631)) and not (layer0_outputs(4616));
    layer1_outputs(737) <= not(layer0_outputs(2716));
    layer1_outputs(738) <= (layer0_outputs(3736)) and (layer0_outputs(3477));
    layer1_outputs(739) <= (layer0_outputs(1821)) and not (layer0_outputs(1575));
    layer1_outputs(740) <= not(layer0_outputs(4485));
    layer1_outputs(741) <= not(layer0_outputs(1978)) or (layer0_outputs(5053));
    layer1_outputs(742) <= not(layer0_outputs(133));
    layer1_outputs(743) <= layer0_outputs(3404);
    layer1_outputs(744) <= layer0_outputs(4042);
    layer1_outputs(745) <= not(layer0_outputs(1763));
    layer1_outputs(746) <= not((layer0_outputs(2078)) or (layer0_outputs(144)));
    layer1_outputs(747) <= not(layer0_outputs(2723)) or (layer0_outputs(3351));
    layer1_outputs(748) <= (layer0_outputs(2375)) or (layer0_outputs(3266));
    layer1_outputs(749) <= not(layer0_outputs(2249)) or (layer0_outputs(529));
    layer1_outputs(750) <= (layer0_outputs(125)) or (layer0_outputs(2004));
    layer1_outputs(751) <= layer0_outputs(2280);
    layer1_outputs(752) <= (layer0_outputs(4188)) and not (layer0_outputs(2595));
    layer1_outputs(753) <= not(layer0_outputs(2277));
    layer1_outputs(754) <= not(layer0_outputs(4391));
    layer1_outputs(755) <= not(layer0_outputs(4366));
    layer1_outputs(756) <= not(layer0_outputs(517));
    layer1_outputs(757) <= layer0_outputs(3634);
    layer1_outputs(758) <= (layer0_outputs(879)) and not (layer0_outputs(1221));
    layer1_outputs(759) <= layer0_outputs(2213);
    layer1_outputs(760) <= not(layer0_outputs(4464));
    layer1_outputs(761) <= not(layer0_outputs(4337)) or (layer0_outputs(35));
    layer1_outputs(762) <= (layer0_outputs(2544)) and not (layer0_outputs(1775));
    layer1_outputs(763) <= (layer0_outputs(135)) and not (layer0_outputs(205));
    layer1_outputs(764) <= not(layer0_outputs(573)) or (layer0_outputs(3170));
    layer1_outputs(765) <= (layer0_outputs(5013)) and (layer0_outputs(2984));
    layer1_outputs(766) <= not(layer0_outputs(4226));
    layer1_outputs(767) <= layer0_outputs(1384);
    layer1_outputs(768) <= not(layer0_outputs(2456)) or (layer0_outputs(1117));
    layer1_outputs(769) <= not(layer0_outputs(2122));
    layer1_outputs(770) <= (layer0_outputs(4087)) and not (layer0_outputs(4723));
    layer1_outputs(771) <= not(layer0_outputs(1838));
    layer1_outputs(772) <= not(layer0_outputs(4506)) or (layer0_outputs(437));
    layer1_outputs(773) <= '0';
    layer1_outputs(774) <= (layer0_outputs(189)) or (layer0_outputs(4223));
    layer1_outputs(775) <= (layer0_outputs(4430)) and not (layer0_outputs(4746));
    layer1_outputs(776) <= not(layer0_outputs(788));
    layer1_outputs(777) <= not(layer0_outputs(3104));
    layer1_outputs(778) <= '1';
    layer1_outputs(779) <= layer0_outputs(3971);
    layer1_outputs(780) <= not((layer0_outputs(760)) or (layer0_outputs(4174)));
    layer1_outputs(781) <= layer0_outputs(1104);
    layer1_outputs(782) <= '1';
    layer1_outputs(783) <= not(layer0_outputs(2573));
    layer1_outputs(784) <= layer0_outputs(3658);
    layer1_outputs(785) <= not((layer0_outputs(183)) or (layer0_outputs(710)));
    layer1_outputs(786) <= not((layer0_outputs(2108)) and (layer0_outputs(4129)));
    layer1_outputs(787) <= not(layer0_outputs(3839));
    layer1_outputs(788) <= not(layer0_outputs(2707));
    layer1_outputs(789) <= not(layer0_outputs(2064));
    layer1_outputs(790) <= layer0_outputs(2218);
    layer1_outputs(791) <= layer0_outputs(3858);
    layer1_outputs(792) <= not(layer0_outputs(1057)) or (layer0_outputs(3182));
    layer1_outputs(793) <= layer0_outputs(4117);
    layer1_outputs(794) <= (layer0_outputs(5076)) and not (layer0_outputs(4390));
    layer1_outputs(795) <= not((layer0_outputs(910)) and (layer0_outputs(1525)));
    layer1_outputs(796) <= not(layer0_outputs(756)) or (layer0_outputs(1672));
    layer1_outputs(797) <= (layer0_outputs(4876)) or (layer0_outputs(687));
    layer1_outputs(798) <= not((layer0_outputs(629)) or (layer0_outputs(3470)));
    layer1_outputs(799) <= '1';
    layer1_outputs(800) <= layer0_outputs(2619);
    layer1_outputs(801) <= layer0_outputs(5110);
    layer1_outputs(802) <= not(layer0_outputs(3206)) or (layer0_outputs(1109));
    layer1_outputs(803) <= (layer0_outputs(938)) or (layer0_outputs(2147));
    layer1_outputs(804) <= not((layer0_outputs(223)) and (layer0_outputs(1031)));
    layer1_outputs(805) <= not(layer0_outputs(2652)) or (layer0_outputs(2880));
    layer1_outputs(806) <= not(layer0_outputs(2161)) or (layer0_outputs(2185));
    layer1_outputs(807) <= layer0_outputs(3046);
    layer1_outputs(808) <= not(layer0_outputs(1403));
    layer1_outputs(809) <= (layer0_outputs(1464)) and not (layer0_outputs(1875));
    layer1_outputs(810) <= not(layer0_outputs(310)) or (layer0_outputs(2238));
    layer1_outputs(811) <= not(layer0_outputs(3770));
    layer1_outputs(812) <= not(layer0_outputs(4577)) or (layer0_outputs(792));
    layer1_outputs(813) <= (layer0_outputs(2374)) or (layer0_outputs(1442));
    layer1_outputs(814) <= (layer0_outputs(3136)) and (layer0_outputs(974));
    layer1_outputs(815) <= layer0_outputs(3318);
    layer1_outputs(816) <= (layer0_outputs(4343)) and not (layer0_outputs(4559));
    layer1_outputs(817) <= not((layer0_outputs(1776)) and (layer0_outputs(4702)));
    layer1_outputs(818) <= (layer0_outputs(1145)) or (layer0_outputs(1118));
    layer1_outputs(819) <= (layer0_outputs(604)) or (layer0_outputs(2718));
    layer1_outputs(820) <= not(layer0_outputs(3257)) or (layer0_outputs(281));
    layer1_outputs(821) <= layer0_outputs(5024);
    layer1_outputs(822) <= not(layer0_outputs(4404));
    layer1_outputs(823) <= (layer0_outputs(4926)) or (layer0_outputs(1527));
    layer1_outputs(824) <= layer0_outputs(2150);
    layer1_outputs(825) <= not(layer0_outputs(3116)) or (layer0_outputs(1934));
    layer1_outputs(826) <= (layer0_outputs(4752)) or (layer0_outputs(4023));
    layer1_outputs(827) <= (layer0_outputs(523)) and not (layer0_outputs(873));
    layer1_outputs(828) <= (layer0_outputs(4270)) or (layer0_outputs(4312));
    layer1_outputs(829) <= '1';
    layer1_outputs(830) <= not(layer0_outputs(1650));
    layer1_outputs(831) <= not(layer0_outputs(716));
    layer1_outputs(832) <= layer0_outputs(2860);
    layer1_outputs(833) <= (layer0_outputs(3395)) and not (layer0_outputs(4528));
    layer1_outputs(834) <= not((layer0_outputs(801)) or (layer0_outputs(2087)));
    layer1_outputs(835) <= layer0_outputs(3461);
    layer1_outputs(836) <= '0';
    layer1_outputs(837) <= not(layer0_outputs(1271)) or (layer0_outputs(4886));
    layer1_outputs(838) <= (layer0_outputs(3505)) and (layer0_outputs(378));
    layer1_outputs(839) <= (layer0_outputs(2773)) or (layer0_outputs(1569));
    layer1_outputs(840) <= layer0_outputs(3358);
    layer1_outputs(841) <= (layer0_outputs(3354)) or (layer0_outputs(1475));
    layer1_outputs(842) <= (layer0_outputs(68)) and not (layer0_outputs(52));
    layer1_outputs(843) <= not((layer0_outputs(657)) xor (layer0_outputs(3136)));
    layer1_outputs(844) <= not(layer0_outputs(5078));
    layer1_outputs(845) <= '1';
    layer1_outputs(846) <= not(layer0_outputs(590));
    layer1_outputs(847) <= not((layer0_outputs(3236)) or (layer0_outputs(239)));
    layer1_outputs(848) <= not((layer0_outputs(2427)) or (layer0_outputs(852)));
    layer1_outputs(849) <= (layer0_outputs(1771)) and not (layer0_outputs(2281));
    layer1_outputs(850) <= not((layer0_outputs(2225)) or (layer0_outputs(3774)));
    layer1_outputs(851) <= layer0_outputs(1103);
    layer1_outputs(852) <= layer0_outputs(3143);
    layer1_outputs(853) <= (layer0_outputs(3107)) or (layer0_outputs(698));
    layer1_outputs(854) <= not((layer0_outputs(3777)) or (layer0_outputs(4501)));
    layer1_outputs(855) <= not((layer0_outputs(978)) and (layer0_outputs(3615)));
    layer1_outputs(856) <= (layer0_outputs(43)) or (layer0_outputs(794));
    layer1_outputs(857) <= not((layer0_outputs(1994)) or (layer0_outputs(3137)));
    layer1_outputs(858) <= not(layer0_outputs(2353)) or (layer0_outputs(1583));
    layer1_outputs(859) <= not((layer0_outputs(3067)) and (layer0_outputs(782)));
    layer1_outputs(860) <= (layer0_outputs(368)) and (layer0_outputs(1227));
    layer1_outputs(861) <= not((layer0_outputs(4387)) or (layer0_outputs(4794)));
    layer1_outputs(862) <= (layer0_outputs(2558)) and not (layer0_outputs(3796));
    layer1_outputs(863) <= layer0_outputs(52);
    layer1_outputs(864) <= not(layer0_outputs(1924));
    layer1_outputs(865) <= not(layer0_outputs(954)) or (layer0_outputs(4633));
    layer1_outputs(866) <= (layer0_outputs(1635)) and (layer0_outputs(2032));
    layer1_outputs(867) <= not((layer0_outputs(3813)) and (layer0_outputs(180)));
    layer1_outputs(868) <= '0';
    layer1_outputs(869) <= not(layer0_outputs(4707));
    layer1_outputs(870) <= (layer0_outputs(4079)) and not (layer0_outputs(1677));
    layer1_outputs(871) <= '1';
    layer1_outputs(872) <= not(layer0_outputs(1749));
    layer1_outputs(873) <= not(layer0_outputs(1476));
    layer1_outputs(874) <= not((layer0_outputs(341)) or (layer0_outputs(1633)));
    layer1_outputs(875) <= not((layer0_outputs(2370)) or (layer0_outputs(1497)));
    layer1_outputs(876) <= not(layer0_outputs(184)) or (layer0_outputs(3665));
    layer1_outputs(877) <= (layer0_outputs(824)) and (layer0_outputs(4136));
    layer1_outputs(878) <= not(layer0_outputs(3827));
    layer1_outputs(879) <= not(layer0_outputs(1638)) or (layer0_outputs(303));
    layer1_outputs(880) <= not(layer0_outputs(4547));
    layer1_outputs(881) <= (layer0_outputs(981)) and (layer0_outputs(4050));
    layer1_outputs(882) <= not(layer0_outputs(2356));
    layer1_outputs(883) <= layer0_outputs(3917);
    layer1_outputs(884) <= (layer0_outputs(3731)) and (layer0_outputs(4912));
    layer1_outputs(885) <= not(layer0_outputs(4410));
    layer1_outputs(886) <= not((layer0_outputs(4610)) and (layer0_outputs(2112)));
    layer1_outputs(887) <= not(layer0_outputs(3591)) or (layer0_outputs(697));
    layer1_outputs(888) <= layer0_outputs(2153);
    layer1_outputs(889) <= not(layer0_outputs(2541));
    layer1_outputs(890) <= not(layer0_outputs(3044));
    layer1_outputs(891) <= (layer0_outputs(4762)) and (layer0_outputs(4924));
    layer1_outputs(892) <= (layer0_outputs(4306)) and not (layer0_outputs(4334));
    layer1_outputs(893) <= not(layer0_outputs(1715)) or (layer0_outputs(4389));
    layer1_outputs(894) <= not(layer0_outputs(2210)) or (layer0_outputs(4979));
    layer1_outputs(895) <= not((layer0_outputs(2366)) or (layer0_outputs(3910)));
    layer1_outputs(896) <= not(layer0_outputs(3913));
    layer1_outputs(897) <= not(layer0_outputs(640));
    layer1_outputs(898) <= layer0_outputs(787);
    layer1_outputs(899) <= not(layer0_outputs(3132));
    layer1_outputs(900) <= not(layer0_outputs(1637));
    layer1_outputs(901) <= not(layer0_outputs(2149)) or (layer0_outputs(3237));
    layer1_outputs(902) <= not((layer0_outputs(4740)) and (layer0_outputs(1851)));
    layer1_outputs(903) <= (layer0_outputs(912)) and not (layer0_outputs(523));
    layer1_outputs(904) <= (layer0_outputs(764)) or (layer0_outputs(1234));
    layer1_outputs(905) <= not(layer0_outputs(1700));
    layer1_outputs(906) <= not(layer0_outputs(2939));
    layer1_outputs(907) <= (layer0_outputs(2244)) or (layer0_outputs(1314));
    layer1_outputs(908) <= not(layer0_outputs(3506)) or (layer0_outputs(4396));
    layer1_outputs(909) <= not((layer0_outputs(4692)) xor (layer0_outputs(2601)));
    layer1_outputs(910) <= not(layer0_outputs(4900));
    layer1_outputs(911) <= not((layer0_outputs(158)) and (layer0_outputs(750)));
    layer1_outputs(912) <= not(layer0_outputs(113));
    layer1_outputs(913) <= not(layer0_outputs(808));
    layer1_outputs(914) <= layer0_outputs(4080);
    layer1_outputs(915) <= not(layer0_outputs(1477)) or (layer0_outputs(198));
    layer1_outputs(916) <= (layer0_outputs(2628)) and not (layer0_outputs(3435));
    layer1_outputs(917) <= not((layer0_outputs(1996)) and (layer0_outputs(4496)));
    layer1_outputs(918) <= (layer0_outputs(732)) and not (layer0_outputs(844));
    layer1_outputs(919) <= (layer0_outputs(1698)) and not (layer0_outputs(820));
    layer1_outputs(920) <= not(layer0_outputs(4899));
    layer1_outputs(921) <= not((layer0_outputs(2454)) xor (layer0_outputs(1854)));
    layer1_outputs(922) <= not(layer0_outputs(1701));
    layer1_outputs(923) <= not(layer0_outputs(854));
    layer1_outputs(924) <= not(layer0_outputs(4958));
    layer1_outputs(925) <= not((layer0_outputs(2154)) or (layer0_outputs(4143)));
    layer1_outputs(926) <= (layer0_outputs(821)) xor (layer0_outputs(4269));
    layer1_outputs(927) <= not((layer0_outputs(3262)) and (layer0_outputs(1902)));
    layer1_outputs(928) <= not((layer0_outputs(387)) and (layer0_outputs(3363)));
    layer1_outputs(929) <= not(layer0_outputs(1982));
    layer1_outputs(930) <= not((layer0_outputs(683)) or (layer0_outputs(4969)));
    layer1_outputs(931) <= (layer0_outputs(1340)) and (layer0_outputs(3541));
    layer1_outputs(932) <= layer0_outputs(2405);
    layer1_outputs(933) <= not(layer0_outputs(3984));
    layer1_outputs(934) <= not((layer0_outputs(3382)) xor (layer0_outputs(3267)));
    layer1_outputs(935) <= not(layer0_outputs(1656)) or (layer0_outputs(2240));
    layer1_outputs(936) <= (layer0_outputs(4637)) and not (layer0_outputs(4322));
    layer1_outputs(937) <= not(layer0_outputs(4576));
    layer1_outputs(938) <= (layer0_outputs(3346)) xor (layer0_outputs(4608));
    layer1_outputs(939) <= (layer0_outputs(3570)) or (layer0_outputs(3344));
    layer1_outputs(940) <= '1';
    layer1_outputs(941) <= not(layer0_outputs(2128));
    layer1_outputs(942) <= not((layer0_outputs(2608)) or (layer0_outputs(1947)));
    layer1_outputs(943) <= not(layer0_outputs(3427)) or (layer0_outputs(1228));
    layer1_outputs(944) <= not(layer0_outputs(3756));
    layer1_outputs(945) <= not(layer0_outputs(1945)) or (layer0_outputs(3927));
    layer1_outputs(946) <= not(layer0_outputs(2660)) or (layer0_outputs(4754));
    layer1_outputs(947) <= not((layer0_outputs(4171)) and (layer0_outputs(4357)));
    layer1_outputs(948) <= not(layer0_outputs(2612));
    layer1_outputs(949) <= not((layer0_outputs(4168)) and (layer0_outputs(647)));
    layer1_outputs(950) <= (layer0_outputs(2690)) or (layer0_outputs(4676));
    layer1_outputs(951) <= layer0_outputs(3264);
    layer1_outputs(952) <= (layer0_outputs(3811)) and (layer0_outputs(4115));
    layer1_outputs(953) <= not((layer0_outputs(1927)) and (layer0_outputs(4273)));
    layer1_outputs(954) <= layer0_outputs(2223);
    layer1_outputs(955) <= not(layer0_outputs(3919)) or (layer0_outputs(5081));
    layer1_outputs(956) <= not((layer0_outputs(832)) or (layer0_outputs(2947)));
    layer1_outputs(957) <= not(layer0_outputs(1097));
    layer1_outputs(958) <= (layer0_outputs(2715)) and (layer0_outputs(2220));
    layer1_outputs(959) <= not((layer0_outputs(891)) or (layer0_outputs(3566)));
    layer1_outputs(960) <= (layer0_outputs(784)) and (layer0_outputs(1454));
    layer1_outputs(961) <= '1';
    layer1_outputs(962) <= layer0_outputs(1939);
    layer1_outputs(963) <= not(layer0_outputs(346)) or (layer0_outputs(2144));
    layer1_outputs(964) <= layer0_outputs(116);
    layer1_outputs(965) <= (layer0_outputs(3076)) xor (layer0_outputs(2562));
    layer1_outputs(966) <= layer0_outputs(4308);
    layer1_outputs(967) <= not(layer0_outputs(2692));
    layer1_outputs(968) <= not(layer0_outputs(1126));
    layer1_outputs(969) <= (layer0_outputs(3277)) and (layer0_outputs(2892));
    layer1_outputs(970) <= (layer0_outputs(1028)) and not (layer0_outputs(5093));
    layer1_outputs(971) <= layer0_outputs(660);
    layer1_outputs(972) <= (layer0_outputs(4240)) and not (layer0_outputs(1584));
    layer1_outputs(973) <= not(layer0_outputs(3997));
    layer1_outputs(974) <= not(layer0_outputs(3361)) or (layer0_outputs(566));
    layer1_outputs(975) <= (layer0_outputs(4799)) or (layer0_outputs(1499));
    layer1_outputs(976) <= not(layer0_outputs(2092));
    layer1_outputs(977) <= (layer0_outputs(3086)) or (layer0_outputs(1008));
    layer1_outputs(978) <= not((layer0_outputs(2360)) or (layer0_outputs(1653)));
    layer1_outputs(979) <= '0';
    layer1_outputs(980) <= (layer0_outputs(4531)) xor (layer0_outputs(3540));
    layer1_outputs(981) <= layer0_outputs(1650);
    layer1_outputs(982) <= layer0_outputs(2911);
    layer1_outputs(983) <= not(layer0_outputs(2448));
    layer1_outputs(984) <= not((layer0_outputs(2193)) or (layer0_outputs(3769)));
    layer1_outputs(985) <= (layer0_outputs(1103)) or (layer0_outputs(3483));
    layer1_outputs(986) <= (layer0_outputs(2778)) and not (layer0_outputs(1594));
    layer1_outputs(987) <= layer0_outputs(1357);
    layer1_outputs(988) <= (layer0_outputs(3065)) and not (layer0_outputs(4789));
    layer1_outputs(989) <= (layer0_outputs(714)) and (layer0_outputs(4620));
    layer1_outputs(990) <= not((layer0_outputs(3705)) or (layer0_outputs(1635)));
    layer1_outputs(991) <= (layer0_outputs(2447)) and (layer0_outputs(2437));
    layer1_outputs(992) <= (layer0_outputs(3764)) and not (layer0_outputs(1429));
    layer1_outputs(993) <= (layer0_outputs(4268)) and not (layer0_outputs(2361));
    layer1_outputs(994) <= not(layer0_outputs(1072));
    layer1_outputs(995) <= not((layer0_outputs(1088)) and (layer0_outputs(1750)));
    layer1_outputs(996) <= not((layer0_outputs(1722)) or (layer0_outputs(4374)));
    layer1_outputs(997) <= (layer0_outputs(177)) and not (layer0_outputs(3781));
    layer1_outputs(998) <= not(layer0_outputs(2079));
    layer1_outputs(999) <= not(layer0_outputs(2094));
    layer1_outputs(1000) <= not(layer0_outputs(1129));
    layer1_outputs(1001) <= not((layer0_outputs(2127)) or (layer0_outputs(4211)));
    layer1_outputs(1002) <= layer0_outputs(2534);
    layer1_outputs(1003) <= not((layer0_outputs(3433)) and (layer0_outputs(347)));
    layer1_outputs(1004) <= layer0_outputs(2240);
    layer1_outputs(1005) <= '1';
    layer1_outputs(1006) <= (layer0_outputs(3705)) or (layer0_outputs(3585));
    layer1_outputs(1007) <= not(layer0_outputs(1090)) or (layer0_outputs(4819));
    layer1_outputs(1008) <= (layer0_outputs(1742)) and not (layer0_outputs(3448));
    layer1_outputs(1009) <= layer0_outputs(209);
    layer1_outputs(1010) <= not(layer0_outputs(5033));
    layer1_outputs(1011) <= not(layer0_outputs(816));
    layer1_outputs(1012) <= layer0_outputs(1784);
    layer1_outputs(1013) <= layer0_outputs(2921);
    layer1_outputs(1014) <= not((layer0_outputs(277)) or (layer0_outputs(2922)));
    layer1_outputs(1015) <= not((layer0_outputs(1244)) or (layer0_outputs(2906)));
    layer1_outputs(1016) <= layer0_outputs(3174);
    layer1_outputs(1017) <= not(layer0_outputs(2539));
    layer1_outputs(1018) <= not(layer0_outputs(4970));
    layer1_outputs(1019) <= not(layer0_outputs(3845));
    layer1_outputs(1020) <= not((layer0_outputs(2860)) xor (layer0_outputs(4905)));
    layer1_outputs(1021) <= (layer0_outputs(959)) xor (layer0_outputs(4559));
    layer1_outputs(1022) <= not(layer0_outputs(2570));
    layer1_outputs(1023) <= not(layer0_outputs(846));
    layer1_outputs(1024) <= (layer0_outputs(4222)) and not (layer0_outputs(3631));
    layer1_outputs(1025) <= not(layer0_outputs(2707)) or (layer0_outputs(2170));
    layer1_outputs(1026) <= layer0_outputs(2263);
    layer1_outputs(1027) <= not(layer0_outputs(2330)) or (layer0_outputs(4144));
    layer1_outputs(1028) <= not(layer0_outputs(929)) or (layer0_outputs(3468));
    layer1_outputs(1029) <= not(layer0_outputs(4005));
    layer1_outputs(1030) <= layer0_outputs(5036);
    layer1_outputs(1031) <= layer0_outputs(3103);
    layer1_outputs(1032) <= layer0_outputs(5013);
    layer1_outputs(1033) <= layer0_outputs(2904);
    layer1_outputs(1034) <= (layer0_outputs(5016)) or (layer0_outputs(484));
    layer1_outputs(1035) <= (layer0_outputs(4921)) or (layer0_outputs(310));
    layer1_outputs(1036) <= not(layer0_outputs(3685));
    layer1_outputs(1037) <= not(layer0_outputs(2501));
    layer1_outputs(1038) <= layer0_outputs(252);
    layer1_outputs(1039) <= '1';
    layer1_outputs(1040) <= (layer0_outputs(811)) or (layer0_outputs(4497));
    layer1_outputs(1041) <= not(layer0_outputs(4147)) or (layer0_outputs(648));
    layer1_outputs(1042) <= not(layer0_outputs(3473));
    layer1_outputs(1043) <= not((layer0_outputs(1166)) or (layer0_outputs(3422)));
    layer1_outputs(1044) <= not((layer0_outputs(1298)) or (layer0_outputs(4663)));
    layer1_outputs(1045) <= not(layer0_outputs(483));
    layer1_outputs(1046) <= (layer0_outputs(3761)) xor (layer0_outputs(4001));
    layer1_outputs(1047) <= not((layer0_outputs(679)) or (layer0_outputs(1369)));
    layer1_outputs(1048) <= (layer0_outputs(1216)) xor (layer0_outputs(454));
    layer1_outputs(1049) <= (layer0_outputs(2043)) and (layer0_outputs(1670));
    layer1_outputs(1050) <= not((layer0_outputs(354)) and (layer0_outputs(3739)));
    layer1_outputs(1051) <= (layer0_outputs(2509)) and not (layer0_outputs(2726));
    layer1_outputs(1052) <= layer0_outputs(65);
    layer1_outputs(1053) <= not(layer0_outputs(3467));
    layer1_outputs(1054) <= not(layer0_outputs(4739));
    layer1_outputs(1055) <= (layer0_outputs(4132)) or (layer0_outputs(278));
    layer1_outputs(1056) <= (layer0_outputs(1194)) and (layer0_outputs(2948));
    layer1_outputs(1057) <= not((layer0_outputs(3731)) and (layer0_outputs(4663)));
    layer1_outputs(1058) <= '0';
    layer1_outputs(1059) <= not(layer0_outputs(2224));
    layer1_outputs(1060) <= layer0_outputs(3482);
    layer1_outputs(1061) <= not(layer0_outputs(1770)) or (layer0_outputs(1992));
    layer1_outputs(1062) <= not(layer0_outputs(3674));
    layer1_outputs(1063) <= '0';
    layer1_outputs(1064) <= not(layer0_outputs(4358));
    layer1_outputs(1065) <= not(layer0_outputs(3933));
    layer1_outputs(1066) <= layer0_outputs(1249);
    layer1_outputs(1067) <= not(layer0_outputs(257)) or (layer0_outputs(3066));
    layer1_outputs(1068) <= not(layer0_outputs(4603)) or (layer0_outputs(843));
    layer1_outputs(1069) <= not(layer0_outputs(708)) or (layer0_outputs(656));
    layer1_outputs(1070) <= not(layer0_outputs(3646)) or (layer0_outputs(769));
    layer1_outputs(1071) <= layer0_outputs(1450);
    layer1_outputs(1072) <= (layer0_outputs(4208)) and (layer0_outputs(2005));
    layer1_outputs(1073) <= (layer0_outputs(2388)) or (layer0_outputs(2760));
    layer1_outputs(1074) <= layer0_outputs(2505);
    layer1_outputs(1075) <= (layer0_outputs(4461)) and not (layer0_outputs(3003));
    layer1_outputs(1076) <= (layer0_outputs(1376)) and (layer0_outputs(2590));
    layer1_outputs(1077) <= not(layer0_outputs(1587));
    layer1_outputs(1078) <= not(layer0_outputs(4075));
    layer1_outputs(1079) <= not(layer0_outputs(3880));
    layer1_outputs(1080) <= layer0_outputs(3714);
    layer1_outputs(1081) <= not(layer0_outputs(1275)) or (layer0_outputs(1829));
    layer1_outputs(1082) <= '1';
    layer1_outputs(1083) <= not(layer0_outputs(2885)) or (layer0_outputs(4305));
    layer1_outputs(1084) <= '1';
    layer1_outputs(1085) <= (layer0_outputs(4628)) and (layer0_outputs(3740));
    layer1_outputs(1086) <= (layer0_outputs(3290)) and not (layer0_outputs(3279));
    layer1_outputs(1087) <= (layer0_outputs(2487)) and not (layer0_outputs(3069));
    layer1_outputs(1088) <= (layer0_outputs(3612)) or (layer0_outputs(2959));
    layer1_outputs(1089) <= (layer0_outputs(3348)) and not (layer0_outputs(3765));
    layer1_outputs(1090) <= layer0_outputs(4397);
    layer1_outputs(1091) <= layer0_outputs(1344);
    layer1_outputs(1092) <= not(layer0_outputs(4689)) or (layer0_outputs(4678));
    layer1_outputs(1093) <= layer0_outputs(2281);
    layer1_outputs(1094) <= layer0_outputs(1873);
    layer1_outputs(1095) <= not(layer0_outputs(4758));
    layer1_outputs(1096) <= '0';
    layer1_outputs(1097) <= (layer0_outputs(2255)) and not (layer0_outputs(2987));
    layer1_outputs(1098) <= not(layer0_outputs(4594));
    layer1_outputs(1099) <= layer0_outputs(1121);
    layer1_outputs(1100) <= not(layer0_outputs(599)) or (layer0_outputs(2701));
    layer1_outputs(1101) <= (layer0_outputs(403)) and not (layer0_outputs(4233));
    layer1_outputs(1102) <= not(layer0_outputs(490)) or (layer0_outputs(504));
    layer1_outputs(1103) <= (layer0_outputs(328)) and not (layer0_outputs(2301));
    layer1_outputs(1104) <= (layer0_outputs(3303)) and (layer0_outputs(223));
    layer1_outputs(1105) <= layer0_outputs(2241);
    layer1_outputs(1106) <= not((layer0_outputs(1603)) and (layer0_outputs(2055)));
    layer1_outputs(1107) <= not((layer0_outputs(4573)) or (layer0_outputs(4125)));
    layer1_outputs(1108) <= not(layer0_outputs(1123)) or (layer0_outputs(1960));
    layer1_outputs(1109) <= (layer0_outputs(2737)) and not (layer0_outputs(917));
    layer1_outputs(1110) <= (layer0_outputs(2611)) and not (layer0_outputs(2594));
    layer1_outputs(1111) <= layer0_outputs(2345);
    layer1_outputs(1112) <= (layer0_outputs(1150)) xor (layer0_outputs(124));
    layer1_outputs(1113) <= layer0_outputs(1692);
    layer1_outputs(1114) <= (layer0_outputs(1269)) or (layer0_outputs(3715));
    layer1_outputs(1115) <= (layer0_outputs(2409)) and (layer0_outputs(2011));
    layer1_outputs(1116) <= not(layer0_outputs(2756));
    layer1_outputs(1117) <= not(layer0_outputs(3229)) or (layer0_outputs(1307));
    layer1_outputs(1118) <= (layer0_outputs(318)) or (layer0_outputs(830));
    layer1_outputs(1119) <= not((layer0_outputs(80)) or (layer0_outputs(2581)));
    layer1_outputs(1120) <= (layer0_outputs(50)) and not (layer0_outputs(4740));
    layer1_outputs(1121) <= (layer0_outputs(4785)) and not (layer0_outputs(1688));
    layer1_outputs(1122) <= not(layer0_outputs(737));
    layer1_outputs(1123) <= layer0_outputs(772);
    layer1_outputs(1124) <= not(layer0_outputs(712)) or (layer0_outputs(3300));
    layer1_outputs(1125) <= not(layer0_outputs(3625));
    layer1_outputs(1126) <= (layer0_outputs(1783)) or (layer0_outputs(4771));
    layer1_outputs(1127) <= (layer0_outputs(4469)) and not (layer0_outputs(3208));
    layer1_outputs(1128) <= not(layer0_outputs(351)) or (layer0_outputs(4872));
    layer1_outputs(1129) <= not((layer0_outputs(2575)) and (layer0_outputs(2533)));
    layer1_outputs(1130) <= not(layer0_outputs(4889)) or (layer0_outputs(2895));
    layer1_outputs(1131) <= (layer0_outputs(3020)) or (layer0_outputs(3016));
    layer1_outputs(1132) <= (layer0_outputs(2813)) and not (layer0_outputs(79));
    layer1_outputs(1133) <= not(layer0_outputs(4134)) or (layer0_outputs(96));
    layer1_outputs(1134) <= '0';
    layer1_outputs(1135) <= (layer0_outputs(2805)) and not (layer0_outputs(2412));
    layer1_outputs(1136) <= layer0_outputs(4204);
    layer1_outputs(1137) <= (layer0_outputs(881)) and (layer0_outputs(4591));
    layer1_outputs(1138) <= not(layer0_outputs(4053));
    layer1_outputs(1139) <= (layer0_outputs(1548)) and not (layer0_outputs(4848));
    layer1_outputs(1140) <= (layer0_outputs(4592)) and (layer0_outputs(4571));
    layer1_outputs(1141) <= not(layer0_outputs(4179));
    layer1_outputs(1142) <= layer0_outputs(239);
    layer1_outputs(1143) <= layer0_outputs(372);
    layer1_outputs(1144) <= not(layer0_outputs(4646));
    layer1_outputs(1145) <= layer0_outputs(1777);
    layer1_outputs(1146) <= layer0_outputs(2323);
    layer1_outputs(1147) <= layer0_outputs(4019);
    layer1_outputs(1148) <= not((layer0_outputs(468)) or (layer0_outputs(4085)));
    layer1_outputs(1149) <= not(layer0_outputs(4930)) or (layer0_outputs(1539));
    layer1_outputs(1150) <= not(layer0_outputs(591));
    layer1_outputs(1151) <= not((layer0_outputs(4881)) and (layer0_outputs(1903)));
    layer1_outputs(1152) <= (layer0_outputs(2526)) or (layer0_outputs(196));
    layer1_outputs(1153) <= layer0_outputs(2076);
    layer1_outputs(1154) <= not(layer0_outputs(3469));
    layer1_outputs(1155) <= not(layer0_outputs(3922)) or (layer0_outputs(2949));
    layer1_outputs(1156) <= layer0_outputs(2698);
    layer1_outputs(1157) <= not((layer0_outputs(3257)) and (layer0_outputs(4950)));
    layer1_outputs(1158) <= layer0_outputs(2919);
    layer1_outputs(1159) <= (layer0_outputs(3883)) and (layer0_outputs(3224));
    layer1_outputs(1160) <= layer0_outputs(270);
    layer1_outputs(1161) <= not((layer0_outputs(1697)) or (layer0_outputs(4132)));
    layer1_outputs(1162) <= (layer0_outputs(1891)) and not (layer0_outputs(3694));
    layer1_outputs(1163) <= not(layer0_outputs(4542));
    layer1_outputs(1164) <= not((layer0_outputs(1912)) xor (layer0_outputs(5107)));
    layer1_outputs(1165) <= '1';
    layer1_outputs(1166) <= layer0_outputs(4274);
    layer1_outputs(1167) <= not(layer0_outputs(4197));
    layer1_outputs(1168) <= not(layer0_outputs(3851));
    layer1_outputs(1169) <= not(layer0_outputs(4982)) or (layer0_outputs(2069));
    layer1_outputs(1170) <= layer0_outputs(717);
    layer1_outputs(1171) <= layer0_outputs(3630);
    layer1_outputs(1172) <= not(layer0_outputs(2324)) or (layer0_outputs(2952));
    layer1_outputs(1173) <= not(layer0_outputs(1542)) or (layer0_outputs(4143));
    layer1_outputs(1174) <= not(layer0_outputs(2438));
    layer1_outputs(1175) <= layer0_outputs(3510);
    layer1_outputs(1176) <= not(layer0_outputs(4837)) or (layer0_outputs(4922));
    layer1_outputs(1177) <= not(layer0_outputs(2983));
    layer1_outputs(1178) <= not(layer0_outputs(4365));
    layer1_outputs(1179) <= (layer0_outputs(2076)) and not (layer0_outputs(211));
    layer1_outputs(1180) <= not(layer0_outputs(2660));
    layer1_outputs(1181) <= (layer0_outputs(4112)) and (layer0_outputs(376));
    layer1_outputs(1182) <= not(layer0_outputs(2693)) or (layer0_outputs(4904));
    layer1_outputs(1183) <= not((layer0_outputs(4631)) or (layer0_outputs(3255)));
    layer1_outputs(1184) <= (layer0_outputs(4936)) and not (layer0_outputs(455));
    layer1_outputs(1185) <= (layer0_outputs(2928)) or (layer0_outputs(3723));
    layer1_outputs(1186) <= not(layer0_outputs(2946));
    layer1_outputs(1187) <= layer0_outputs(4153);
    layer1_outputs(1188) <= layer0_outputs(2520);
    layer1_outputs(1189) <= not((layer0_outputs(4004)) and (layer0_outputs(4046)));
    layer1_outputs(1190) <= (layer0_outputs(4492)) and not (layer0_outputs(2031));
    layer1_outputs(1191) <= not(layer0_outputs(1521)) or (layer0_outputs(3458));
    layer1_outputs(1192) <= not(layer0_outputs(1765));
    layer1_outputs(1193) <= not((layer0_outputs(3101)) and (layer0_outputs(6)));
    layer1_outputs(1194) <= layer0_outputs(1069);
    layer1_outputs(1195) <= not(layer0_outputs(2139));
    layer1_outputs(1196) <= '1';
    layer1_outputs(1197) <= not(layer0_outputs(4830));
    layer1_outputs(1198) <= (layer0_outputs(2349)) or (layer0_outputs(4510));
    layer1_outputs(1199) <= '0';
    layer1_outputs(1200) <= not(layer0_outputs(2058)) or (layer0_outputs(4729));
    layer1_outputs(1201) <= '1';
    layer1_outputs(1202) <= layer0_outputs(3944);
    layer1_outputs(1203) <= not((layer0_outputs(1752)) and (layer0_outputs(3543)));
    layer1_outputs(1204) <= layer0_outputs(3114);
    layer1_outputs(1205) <= not(layer0_outputs(4272)) or (layer0_outputs(2490));
    layer1_outputs(1206) <= layer0_outputs(2811);
    layer1_outputs(1207) <= '0';
    layer1_outputs(1208) <= not(layer0_outputs(4380)) or (layer0_outputs(1849));
    layer1_outputs(1209) <= not(layer0_outputs(1426));
    layer1_outputs(1210) <= layer0_outputs(960);
    layer1_outputs(1211) <= not((layer0_outputs(1727)) and (layer0_outputs(2270)));
    layer1_outputs(1212) <= not((layer0_outputs(3521)) and (layer0_outputs(3097)));
    layer1_outputs(1213) <= not((layer0_outputs(3897)) and (layer0_outputs(5028)));
    layer1_outputs(1214) <= not((layer0_outputs(3001)) or (layer0_outputs(940)));
    layer1_outputs(1215) <= (layer0_outputs(2023)) and (layer0_outputs(1759));
    layer1_outputs(1216) <= not(layer0_outputs(4730)) or (layer0_outputs(2337));
    layer1_outputs(1217) <= not(layer0_outputs(3655));
    layer1_outputs(1218) <= (layer0_outputs(2118)) and not (layer0_outputs(249));
    layer1_outputs(1219) <= not((layer0_outputs(4673)) and (layer0_outputs(2512)));
    layer1_outputs(1220) <= not((layer0_outputs(4726)) xor (layer0_outputs(1258)));
    layer1_outputs(1221) <= (layer0_outputs(566)) and (layer0_outputs(5061));
    layer1_outputs(1222) <= (layer0_outputs(684)) and (layer0_outputs(5042));
    layer1_outputs(1223) <= layer0_outputs(3251);
    layer1_outputs(1224) <= (layer0_outputs(4116)) and (layer0_outputs(5080));
    layer1_outputs(1225) <= not(layer0_outputs(2677)) or (layer0_outputs(1249));
    layer1_outputs(1226) <= not(layer0_outputs(176));
    layer1_outputs(1227) <= (layer0_outputs(3590)) and not (layer0_outputs(3058));
    layer1_outputs(1228) <= not(layer0_outputs(3292)) or (layer0_outputs(4059));
    layer1_outputs(1229) <= not(layer0_outputs(2295));
    layer1_outputs(1230) <= not(layer0_outputs(1757)) or (layer0_outputs(626));
    layer1_outputs(1231) <= not((layer0_outputs(2976)) or (layer0_outputs(3746)));
    layer1_outputs(1232) <= (layer0_outputs(1356)) and not (layer0_outputs(4813));
    layer1_outputs(1233) <= layer0_outputs(1645);
    layer1_outputs(1234) <= layer0_outputs(4603);
    layer1_outputs(1235) <= not(layer0_outputs(3784)) or (layer0_outputs(3822));
    layer1_outputs(1236) <= not(layer0_outputs(876));
    layer1_outputs(1237) <= (layer0_outputs(4189)) and not (layer0_outputs(152));
    layer1_outputs(1238) <= '1';
    layer1_outputs(1239) <= (layer0_outputs(5059)) or (layer0_outputs(4216));
    layer1_outputs(1240) <= not(layer0_outputs(103)) or (layer0_outputs(810));
    layer1_outputs(1241) <= not(layer0_outputs(851)) or (layer0_outputs(1175));
    layer1_outputs(1242) <= layer0_outputs(2886);
    layer1_outputs(1243) <= not(layer0_outputs(1972)) or (layer0_outputs(3966));
    layer1_outputs(1244) <= not(layer0_outputs(2747));
    layer1_outputs(1245) <= not(layer0_outputs(548));
    layer1_outputs(1246) <= not(layer0_outputs(473)) or (layer0_outputs(954));
    layer1_outputs(1247) <= not(layer0_outputs(4355));
    layer1_outputs(1248) <= not(layer0_outputs(414)) or (layer0_outputs(1403));
    layer1_outputs(1249) <= layer0_outputs(3154);
    layer1_outputs(1250) <= layer0_outputs(1322);
    layer1_outputs(1251) <= (layer0_outputs(2868)) and not (layer0_outputs(138));
    layer1_outputs(1252) <= layer0_outputs(3734);
    layer1_outputs(1253) <= not(layer0_outputs(69)) or (layer0_outputs(1458));
    layer1_outputs(1254) <= layer0_outputs(1064);
    layer1_outputs(1255) <= '0';
    layer1_outputs(1256) <= not((layer0_outputs(4346)) and (layer0_outputs(112)));
    layer1_outputs(1257) <= (layer0_outputs(4504)) or (layer0_outputs(2336));
    layer1_outputs(1258) <= not((layer0_outputs(1658)) and (layer0_outputs(1997)));
    layer1_outputs(1259) <= (layer0_outputs(2818)) and not (layer0_outputs(4575));
    layer1_outputs(1260) <= not(layer0_outputs(615));
    layer1_outputs(1261) <= layer0_outputs(3580);
    layer1_outputs(1262) <= not(layer0_outputs(219));
    layer1_outputs(1263) <= '0';
    layer1_outputs(1264) <= layer0_outputs(4248);
    layer1_outputs(1265) <= layer0_outputs(4097);
    layer1_outputs(1266) <= not(layer0_outputs(1473)) or (layer0_outputs(1168));
    layer1_outputs(1267) <= '1';
    layer1_outputs(1268) <= layer0_outputs(4646);
    layer1_outputs(1269) <= (layer0_outputs(492)) and (layer0_outputs(3296));
    layer1_outputs(1270) <= (layer0_outputs(283)) and (layer0_outputs(804));
    layer1_outputs(1271) <= '0';
    layer1_outputs(1272) <= not(layer0_outputs(478));
    layer1_outputs(1273) <= not(layer0_outputs(3704)) or (layer0_outputs(3735));
    layer1_outputs(1274) <= not(layer0_outputs(2372)) or (layer0_outputs(2894));
    layer1_outputs(1275) <= (layer0_outputs(974)) and not (layer0_outputs(1152));
    layer1_outputs(1276) <= not(layer0_outputs(2368));
    layer1_outputs(1277) <= not(layer0_outputs(4444));
    layer1_outputs(1278) <= not((layer0_outputs(4516)) and (layer0_outputs(1938)));
    layer1_outputs(1279) <= (layer0_outputs(4547)) and (layer0_outputs(463));
    layer1_outputs(1280) <= layer0_outputs(333);
    layer1_outputs(1281) <= not(layer0_outputs(3107));
    layer1_outputs(1282) <= (layer0_outputs(1339)) and not (layer0_outputs(3906));
    layer1_outputs(1283) <= not(layer0_outputs(1807));
    layer1_outputs(1284) <= layer0_outputs(4813);
    layer1_outputs(1285) <= not((layer0_outputs(2418)) xor (layer0_outputs(2847)));
    layer1_outputs(1286) <= not(layer0_outputs(127)) or (layer0_outputs(214));
    layer1_outputs(1287) <= layer0_outputs(3221);
    layer1_outputs(1288) <= (layer0_outputs(628)) and (layer0_outputs(3886));
    layer1_outputs(1289) <= (layer0_outputs(2497)) and (layer0_outputs(2583));
    layer1_outputs(1290) <= not(layer0_outputs(1188));
    layer1_outputs(1291) <= layer0_outputs(3832);
    layer1_outputs(1292) <= (layer0_outputs(3829)) or (layer0_outputs(3717));
    layer1_outputs(1293) <= '0';
    layer1_outputs(1294) <= (layer0_outputs(4412)) xor (layer0_outputs(2877));
    layer1_outputs(1295) <= not(layer0_outputs(3804)) or (layer0_outputs(4146));
    layer1_outputs(1296) <= (layer0_outputs(2826)) and (layer0_outputs(1056));
    layer1_outputs(1297) <= not(layer0_outputs(2662));
    layer1_outputs(1298) <= (layer0_outputs(680)) xor (layer0_outputs(4145));
    layer1_outputs(1299) <= not(layer0_outputs(4966));
    layer1_outputs(1300) <= '0';
    layer1_outputs(1301) <= not((layer0_outputs(4823)) and (layer0_outputs(928)));
    layer1_outputs(1302) <= layer0_outputs(2599);
    layer1_outputs(1303) <= not(layer0_outputs(2025)) or (layer0_outputs(3134));
    layer1_outputs(1304) <= not((layer0_outputs(3613)) or (layer0_outputs(1723)));
    layer1_outputs(1305) <= (layer0_outputs(4787)) or (layer0_outputs(2190));
    layer1_outputs(1306) <= '0';
    layer1_outputs(1307) <= (layer0_outputs(4220)) and (layer0_outputs(1313));
    layer1_outputs(1308) <= (layer0_outputs(4135)) and not (layer0_outputs(1178));
    layer1_outputs(1309) <= not(layer0_outputs(631)) or (layer0_outputs(3691));
    layer1_outputs(1310) <= (layer0_outputs(203)) and not (layer0_outputs(1895));
    layer1_outputs(1311) <= not(layer0_outputs(1029));
    layer1_outputs(1312) <= not(layer0_outputs(464));
    layer1_outputs(1313) <= (layer0_outputs(2594)) xor (layer0_outputs(902));
    layer1_outputs(1314) <= (layer0_outputs(308)) and not (layer0_outputs(215));
    layer1_outputs(1315) <= (layer0_outputs(2243)) and not (layer0_outputs(3957));
    layer1_outputs(1316) <= (layer0_outputs(2073)) or (layer0_outputs(4178));
    layer1_outputs(1317) <= not(layer0_outputs(4266));
    layer1_outputs(1318) <= layer0_outputs(3305);
    layer1_outputs(1319) <= layer0_outputs(4123);
    layer1_outputs(1320) <= not(layer0_outputs(3432)) or (layer0_outputs(722));
    layer1_outputs(1321) <= not((layer0_outputs(4533)) or (layer0_outputs(1859)));
    layer1_outputs(1322) <= layer0_outputs(1715);
    layer1_outputs(1323) <= not(layer0_outputs(4058));
    layer1_outputs(1324) <= not(layer0_outputs(2528));
    layer1_outputs(1325) <= not((layer0_outputs(5017)) and (layer0_outputs(1342)));
    layer1_outputs(1326) <= not(layer0_outputs(278)) or (layer0_outputs(1341));
    layer1_outputs(1327) <= not((layer0_outputs(683)) and (layer0_outputs(661)));
    layer1_outputs(1328) <= (layer0_outputs(3179)) or (layer0_outputs(382));
    layer1_outputs(1329) <= not(layer0_outputs(3802));
    layer1_outputs(1330) <= layer0_outputs(1957);
    layer1_outputs(1331) <= not(layer0_outputs(4655)) or (layer0_outputs(56));
    layer1_outputs(1332) <= not(layer0_outputs(218)) or (layer0_outputs(4169));
    layer1_outputs(1333) <= layer0_outputs(2582);
    layer1_outputs(1334) <= (layer0_outputs(868)) and not (layer0_outputs(1530));
    layer1_outputs(1335) <= (layer0_outputs(2666)) and not (layer0_outputs(3908));
    layer1_outputs(1336) <= layer0_outputs(2482);
    layer1_outputs(1337) <= not(layer0_outputs(4792));
    layer1_outputs(1338) <= not((layer0_outputs(107)) and (layer0_outputs(2869)));
    layer1_outputs(1339) <= not(layer0_outputs(3349));
    layer1_outputs(1340) <= layer0_outputs(4714);
    layer1_outputs(1341) <= not(layer0_outputs(739));
    layer1_outputs(1342) <= not(layer0_outputs(4660)) or (layer0_outputs(4140));
    layer1_outputs(1343) <= not(layer0_outputs(4557));
    layer1_outputs(1344) <= not((layer0_outputs(1262)) xor (layer0_outputs(1898)));
    layer1_outputs(1345) <= layer0_outputs(4119);
    layer1_outputs(1346) <= not(layer0_outputs(4607));
    layer1_outputs(1347) <= not(layer0_outputs(1159));
    layer1_outputs(1348) <= not(layer0_outputs(4848));
    layer1_outputs(1349) <= (layer0_outputs(2484)) and (layer0_outputs(2433));
    layer1_outputs(1350) <= (layer0_outputs(1866)) xor (layer0_outputs(4626));
    layer1_outputs(1351) <= (layer0_outputs(1004)) xor (layer0_outputs(4207));
    layer1_outputs(1352) <= not(layer0_outputs(3881));
    layer1_outputs(1353) <= (layer0_outputs(4299)) and not (layer0_outputs(2797));
    layer1_outputs(1354) <= not((layer0_outputs(2283)) or (layer0_outputs(2239)));
    layer1_outputs(1355) <= not(layer0_outputs(3898));
    layer1_outputs(1356) <= not((layer0_outputs(1238)) and (layer0_outputs(229)));
    layer1_outputs(1357) <= (layer0_outputs(4959)) and (layer0_outputs(4252));
    layer1_outputs(1358) <= (layer0_outputs(2242)) and not (layer0_outputs(3985));
    layer1_outputs(1359) <= not(layer0_outputs(3536)) or (layer0_outputs(54));
    layer1_outputs(1360) <= (layer0_outputs(2182)) and (layer0_outputs(2627));
    layer1_outputs(1361) <= layer0_outputs(3336);
    layer1_outputs(1362) <= not((layer0_outputs(282)) or (layer0_outputs(1183)));
    layer1_outputs(1363) <= not(layer0_outputs(3145)) or (layer0_outputs(2887));
    layer1_outputs(1364) <= layer0_outputs(2385);
    layer1_outputs(1365) <= layer0_outputs(2811);
    layer1_outputs(1366) <= (layer0_outputs(4548)) and not (layer0_outputs(2884));
    layer1_outputs(1367) <= '0';
    layer1_outputs(1368) <= (layer0_outputs(3785)) or (layer0_outputs(1291));
    layer1_outputs(1369) <= not(layer0_outputs(3433));
    layer1_outputs(1370) <= not(layer0_outputs(2658)) or (layer0_outputs(4831));
    layer1_outputs(1371) <= (layer0_outputs(964)) xor (layer0_outputs(5069));
    layer1_outputs(1372) <= (layer0_outputs(1779)) and not (layer0_outputs(3916));
    layer1_outputs(1373) <= layer0_outputs(3336);
    layer1_outputs(1374) <= (layer0_outputs(3862)) and (layer0_outputs(450));
    layer1_outputs(1375) <= (layer0_outputs(2457)) and not (layer0_outputs(4133));
    layer1_outputs(1376) <= not(layer0_outputs(1838)) or (layer0_outputs(245));
    layer1_outputs(1377) <= layer0_outputs(3458);
    layer1_outputs(1378) <= not(layer0_outputs(3684));
    layer1_outputs(1379) <= layer0_outputs(1082);
    layer1_outputs(1380) <= not((layer0_outputs(4198)) and (layer0_outputs(4314)));
    layer1_outputs(1381) <= (layer0_outputs(4065)) and (layer0_outputs(2112));
    layer1_outputs(1382) <= (layer0_outputs(6)) and not (layer0_outputs(575));
    layer1_outputs(1383) <= not(layer0_outputs(998));
    layer1_outputs(1384) <= layer0_outputs(3584);
    layer1_outputs(1385) <= not((layer0_outputs(456)) xor (layer0_outputs(1713)));
    layer1_outputs(1386) <= not((layer0_outputs(3122)) xor (layer0_outputs(322)));
    layer1_outputs(1387) <= layer0_outputs(2965);
    layer1_outputs(1388) <= layer0_outputs(2678);
    layer1_outputs(1389) <= not(layer0_outputs(3099));
    layer1_outputs(1390) <= not(layer0_outputs(2487)) or (layer0_outputs(291));
    layer1_outputs(1391) <= (layer0_outputs(1568)) and (layer0_outputs(2745));
    layer1_outputs(1392) <= not(layer0_outputs(2468)) or (layer0_outputs(1166));
    layer1_outputs(1393) <= (layer0_outputs(91)) and (layer0_outputs(3150));
    layer1_outputs(1394) <= not((layer0_outputs(4724)) and (layer0_outputs(3866)));
    layer1_outputs(1395) <= layer0_outputs(1724);
    layer1_outputs(1396) <= not(layer0_outputs(3402)) or (layer0_outputs(3761));
    layer1_outputs(1397) <= not(layer0_outputs(2665));
    layer1_outputs(1398) <= (layer0_outputs(3062)) and not (layer0_outputs(2704));
    layer1_outputs(1399) <= not(layer0_outputs(2297)) or (layer0_outputs(4350));
    layer1_outputs(1400) <= (layer0_outputs(4645)) and not (layer0_outputs(3641));
    layer1_outputs(1401) <= not((layer0_outputs(583)) or (layer0_outputs(2890)));
    layer1_outputs(1402) <= layer0_outputs(390);
    layer1_outputs(1403) <= not(layer0_outputs(2761));
    layer1_outputs(1404) <= not(layer0_outputs(1053)) or (layer0_outputs(5001));
    layer1_outputs(1405) <= not((layer0_outputs(29)) xor (layer0_outputs(2639)));
    layer1_outputs(1406) <= (layer0_outputs(3124)) and not (layer0_outputs(4704));
    layer1_outputs(1407) <= not((layer0_outputs(4176)) and (layer0_outputs(358)));
    layer1_outputs(1408) <= not(layer0_outputs(4778));
    layer1_outputs(1409) <= (layer0_outputs(4743)) and not (layer0_outputs(2600));
    layer1_outputs(1410) <= layer0_outputs(3261);
    layer1_outputs(1411) <= not(layer0_outputs(4383));
    layer1_outputs(1412) <= not(layer0_outputs(5037)) or (layer0_outputs(289));
    layer1_outputs(1413) <= layer0_outputs(751);
    layer1_outputs(1414) <= layer0_outputs(78);
    layer1_outputs(1415) <= layer0_outputs(2848);
    layer1_outputs(1416) <= (layer0_outputs(3762)) and (layer0_outputs(758));
    layer1_outputs(1417) <= not(layer0_outputs(4305));
    layer1_outputs(1418) <= (layer0_outputs(309)) and (layer0_outputs(2486));
    layer1_outputs(1419) <= not((layer0_outputs(3595)) or (layer0_outputs(108)));
    layer1_outputs(1420) <= not((layer0_outputs(4757)) or (layer0_outputs(1126)));
    layer1_outputs(1421) <= (layer0_outputs(2382)) or (layer0_outputs(1735));
    layer1_outputs(1422) <= not(layer0_outputs(594));
    layer1_outputs(1423) <= (layer0_outputs(450)) and not (layer0_outputs(3283));
    layer1_outputs(1424) <= not(layer0_outputs(4202));
    layer1_outputs(1425) <= '0';
    layer1_outputs(1426) <= layer0_outputs(643);
    layer1_outputs(1427) <= not(layer0_outputs(3783));
    layer1_outputs(1428) <= (layer0_outputs(4045)) and not (layer0_outputs(448));
    layer1_outputs(1429) <= not(layer0_outputs(340));
    layer1_outputs(1430) <= layer0_outputs(3562);
    layer1_outputs(1431) <= not((layer0_outputs(2731)) xor (layer0_outputs(3412)));
    layer1_outputs(1432) <= (layer0_outputs(182)) and (layer0_outputs(3113));
    layer1_outputs(1433) <= layer0_outputs(3411);
    layer1_outputs(1434) <= not((layer0_outputs(2185)) xor (layer0_outputs(1158)));
    layer1_outputs(1435) <= (layer0_outputs(1167)) and not (layer0_outputs(3904));
    layer1_outputs(1436) <= not(layer0_outputs(3114));
    layer1_outputs(1437) <= layer0_outputs(635);
    layer1_outputs(1438) <= not(layer0_outputs(185));
    layer1_outputs(1439) <= not(layer0_outputs(4551));
    layer1_outputs(1440) <= layer0_outputs(1858);
    layer1_outputs(1441) <= (layer0_outputs(104)) or (layer0_outputs(129));
    layer1_outputs(1442) <= layer0_outputs(1074);
    layer1_outputs(1443) <= not(layer0_outputs(3547));
    layer1_outputs(1444) <= not(layer0_outputs(425));
    layer1_outputs(1445) <= (layer0_outputs(1428)) and (layer0_outputs(2832));
    layer1_outputs(1446) <= not(layer0_outputs(2560)) or (layer0_outputs(106));
    layer1_outputs(1447) <= (layer0_outputs(2355)) and not (layer0_outputs(1165));
    layer1_outputs(1448) <= not((layer0_outputs(2137)) and (layer0_outputs(2861)));
    layer1_outputs(1449) <= not(layer0_outputs(2928));
    layer1_outputs(1450) <= not(layer0_outputs(400));
    layer1_outputs(1451) <= not(layer0_outputs(4783));
    layer1_outputs(1452) <= (layer0_outputs(4455)) and not (layer0_outputs(4998));
    layer1_outputs(1453) <= layer0_outputs(4224);
    layer1_outputs(1454) <= (layer0_outputs(2765)) or (layer0_outputs(2555));
    layer1_outputs(1455) <= (layer0_outputs(267)) and not (layer0_outputs(1517));
    layer1_outputs(1456) <= (layer0_outputs(509)) xor (layer0_outputs(2649));
    layer1_outputs(1457) <= not(layer0_outputs(3434)) or (layer0_outputs(494));
    layer1_outputs(1458) <= (layer0_outputs(759)) or (layer0_outputs(4449));
    layer1_outputs(1459) <= not(layer0_outputs(304)) or (layer0_outputs(420));
    layer1_outputs(1460) <= layer0_outputs(5072);
    layer1_outputs(1461) <= not(layer0_outputs(4761));
    layer1_outputs(1462) <= not(layer0_outputs(3181));
    layer1_outputs(1463) <= not(layer0_outputs(3708));
    layer1_outputs(1464) <= not(layer0_outputs(404));
    layer1_outputs(1465) <= layer0_outputs(3856);
    layer1_outputs(1466) <= not((layer0_outputs(4302)) xor (layer0_outputs(2927)));
    layer1_outputs(1467) <= (layer0_outputs(4479)) and not (layer0_outputs(2067));
    layer1_outputs(1468) <= not((layer0_outputs(3875)) or (layer0_outputs(4868)));
    layer1_outputs(1469) <= not(layer0_outputs(1624));
    layer1_outputs(1470) <= '1';
    layer1_outputs(1471) <= (layer0_outputs(65)) or (layer0_outputs(485));
    layer1_outputs(1472) <= not(layer0_outputs(1429));
    layer1_outputs(1473) <= not((layer0_outputs(3698)) and (layer0_outputs(1837)));
    layer1_outputs(1474) <= layer0_outputs(2776);
    layer1_outputs(1475) <= (layer0_outputs(2224)) and not (layer0_outputs(610));
    layer1_outputs(1476) <= not((layer0_outputs(0)) and (layer0_outputs(2768)));
    layer1_outputs(1477) <= not(layer0_outputs(4935));
    layer1_outputs(1478) <= not(layer0_outputs(2362));
    layer1_outputs(1479) <= layer0_outputs(3523);
    layer1_outputs(1480) <= not((layer0_outputs(1404)) and (layer0_outputs(291)));
    layer1_outputs(1481) <= (layer0_outputs(3804)) and not (layer0_outputs(809));
    layer1_outputs(1482) <= layer0_outputs(4140);
    layer1_outputs(1483) <= not(layer0_outputs(1517));
    layer1_outputs(1484) <= not((layer0_outputs(342)) and (layer0_outputs(1553)));
    layer1_outputs(1485) <= not(layer0_outputs(602));
    layer1_outputs(1486) <= not((layer0_outputs(3310)) xor (layer0_outputs(2002)));
    layer1_outputs(1487) <= layer0_outputs(2640);
    layer1_outputs(1488) <= layer0_outputs(4089);
    layer1_outputs(1489) <= layer0_outputs(4606);
    layer1_outputs(1490) <= not(layer0_outputs(4841));
    layer1_outputs(1491) <= (layer0_outputs(4987)) or (layer0_outputs(940));
    layer1_outputs(1492) <= layer0_outputs(1865);
    layer1_outputs(1493) <= (layer0_outputs(3306)) or (layer0_outputs(4278));
    layer1_outputs(1494) <= not(layer0_outputs(2164));
    layer1_outputs(1495) <= (layer0_outputs(2774)) or (layer0_outputs(412));
    layer1_outputs(1496) <= not((layer0_outputs(877)) and (layer0_outputs(1347)));
    layer1_outputs(1497) <= layer0_outputs(1857);
    layer1_outputs(1498) <= not(layer0_outputs(2982));
    layer1_outputs(1499) <= not(layer0_outputs(3529));
    layer1_outputs(1500) <= not(layer0_outputs(5095)) or (layer0_outputs(1935));
    layer1_outputs(1501) <= '0';
    layer1_outputs(1502) <= (layer0_outputs(2197)) and (layer0_outputs(4595));
    layer1_outputs(1503) <= not((layer0_outputs(1505)) or (layer0_outputs(760)));
    layer1_outputs(1504) <= not(layer0_outputs(217)) or (layer0_outputs(5038));
    layer1_outputs(1505) <= not((layer0_outputs(4661)) or (layer0_outputs(3763)));
    layer1_outputs(1506) <= not(layer0_outputs(3356));
    layer1_outputs(1507) <= '0';
    layer1_outputs(1508) <= (layer0_outputs(2903)) and not (layer0_outputs(3280));
    layer1_outputs(1509) <= '0';
    layer1_outputs(1510) <= not((layer0_outputs(2310)) or (layer0_outputs(3138)));
    layer1_outputs(1511) <= '1';
    layer1_outputs(1512) <= (layer0_outputs(3240)) or (layer0_outputs(3690));
    layer1_outputs(1513) <= '0';
    layer1_outputs(1514) <= (layer0_outputs(1023)) and not (layer0_outputs(4489));
    layer1_outputs(1515) <= not((layer0_outputs(3055)) and (layer0_outputs(4564)));
    layer1_outputs(1516) <= not((layer0_outputs(2130)) xor (layer0_outputs(2568)));
    layer1_outputs(1517) <= (layer0_outputs(2536)) or (layer0_outputs(4032));
    layer1_outputs(1518) <= (layer0_outputs(4780)) or (layer0_outputs(898));
    layer1_outputs(1519) <= not(layer0_outputs(5067));
    layer1_outputs(1520) <= not(layer0_outputs(5101)) or (layer0_outputs(2887));
    layer1_outputs(1521) <= (layer0_outputs(4847)) and not (layer0_outputs(917));
    layer1_outputs(1522) <= (layer0_outputs(4169)) and (layer0_outputs(4232));
    layer1_outputs(1523) <= layer0_outputs(4617);
    layer1_outputs(1524) <= (layer0_outputs(4106)) or (layer0_outputs(2734));
    layer1_outputs(1525) <= layer0_outputs(4769);
    layer1_outputs(1526) <= (layer0_outputs(2362)) and not (layer0_outputs(1150));
    layer1_outputs(1527) <= not((layer0_outputs(3594)) and (layer0_outputs(4420)));
    layer1_outputs(1528) <= not(layer0_outputs(1516)) or (layer0_outputs(2071));
    layer1_outputs(1529) <= not((layer0_outputs(142)) or (layer0_outputs(1445)));
    layer1_outputs(1530) <= not(layer0_outputs(3868));
    layer1_outputs(1531) <= not(layer0_outputs(3232));
    layer1_outputs(1532) <= (layer0_outputs(1789)) and (layer0_outputs(4587));
    layer1_outputs(1533) <= (layer0_outputs(973)) xor (layer0_outputs(1016));
    layer1_outputs(1534) <= not(layer0_outputs(1801)) or (layer0_outputs(1224));
    layer1_outputs(1535) <= (layer0_outputs(602)) and not (layer0_outputs(1990));
    layer1_outputs(1536) <= layer0_outputs(16);
    layer1_outputs(1537) <= '1';
    layer1_outputs(1538) <= not((layer0_outputs(880)) or (layer0_outputs(105)));
    layer1_outputs(1539) <= not(layer0_outputs(3111)) or (layer0_outputs(1731));
    layer1_outputs(1540) <= (layer0_outputs(1702)) and not (layer0_outputs(1305));
    layer1_outputs(1541) <= (layer0_outputs(1478)) and not (layer0_outputs(671));
    layer1_outputs(1542) <= not(layer0_outputs(4658));
    layer1_outputs(1543) <= '0';
    layer1_outputs(1544) <= layer0_outputs(4868);
    layer1_outputs(1545) <= layer0_outputs(2994);
    layer1_outputs(1546) <= not(layer0_outputs(2214));
    layer1_outputs(1547) <= not((layer0_outputs(4701)) or (layer0_outputs(1148)));
    layer1_outputs(1548) <= not(layer0_outputs(3299)) or (layer0_outputs(1843));
    layer1_outputs(1549) <= not(layer0_outputs(3837)) or (layer0_outputs(4103));
    layer1_outputs(1550) <= layer0_outputs(4600);
    layer1_outputs(1551) <= (layer0_outputs(3352)) and (layer0_outputs(2901));
    layer1_outputs(1552) <= (layer0_outputs(3331)) or (layer0_outputs(4774));
    layer1_outputs(1553) <= layer0_outputs(4429);
    layer1_outputs(1554) <= not(layer0_outputs(1144));
    layer1_outputs(1555) <= layer0_outputs(3864);
    layer1_outputs(1556) <= not((layer0_outputs(4035)) or (layer0_outputs(2500)));
    layer1_outputs(1557) <= not(layer0_outputs(1803)) or (layer0_outputs(4833));
    layer1_outputs(1558) <= layer0_outputs(4037);
    layer1_outputs(1559) <= not(layer0_outputs(2668)) or (layer0_outputs(1276));
    layer1_outputs(1560) <= (layer0_outputs(889)) or (layer0_outputs(1839));
    layer1_outputs(1561) <= not(layer0_outputs(598)) or (layer0_outputs(2142));
    layer1_outputs(1562) <= layer0_outputs(5044);
    layer1_outputs(1563) <= not(layer0_outputs(2103));
    layer1_outputs(1564) <= layer0_outputs(117);
    layer1_outputs(1565) <= not((layer0_outputs(503)) and (layer0_outputs(660)));
    layer1_outputs(1566) <= not(layer0_outputs(3706));
    layer1_outputs(1567) <= layer0_outputs(906);
    layer1_outputs(1568) <= layer0_outputs(2952);
    layer1_outputs(1569) <= layer0_outputs(3813);
    layer1_outputs(1570) <= not(layer0_outputs(1550));
    layer1_outputs(1571) <= layer0_outputs(3315);
    layer1_outputs(1572) <= not(layer0_outputs(4352));
    layer1_outputs(1573) <= not(layer0_outputs(2302)) or (layer0_outputs(3412));
    layer1_outputs(1574) <= (layer0_outputs(3429)) and not (layer0_outputs(1436));
    layer1_outputs(1575) <= not(layer0_outputs(1176));
    layer1_outputs(1576) <= not(layer0_outputs(3130)) or (layer0_outputs(2028));
    layer1_outputs(1577) <= layer0_outputs(5014);
    layer1_outputs(1578) <= layer0_outputs(3522);
    layer1_outputs(1579) <= not(layer0_outputs(3873)) or (layer0_outputs(664));
    layer1_outputs(1580) <= not((layer0_outputs(2552)) or (layer0_outputs(4318)));
    layer1_outputs(1581) <= layer0_outputs(753);
    layer1_outputs(1582) <= layer0_outputs(1258);
    layer1_outputs(1583) <= (layer0_outputs(4691)) and not (layer0_outputs(1348));
    layer1_outputs(1584) <= (layer0_outputs(726)) or (layer0_outputs(2477));
    layer1_outputs(1585) <= layer0_outputs(2036);
    layer1_outputs(1586) <= (layer0_outputs(1333)) and not (layer0_outputs(87));
    layer1_outputs(1587) <= layer0_outputs(5059);
    layer1_outputs(1588) <= not(layer0_outputs(1700)) or (layer0_outputs(1598));
    layer1_outputs(1589) <= not(layer0_outputs(4018));
    layer1_outputs(1590) <= layer0_outputs(1590);
    layer1_outputs(1591) <= not(layer0_outputs(1573)) or (layer0_outputs(599));
    layer1_outputs(1592) <= not((layer0_outputs(762)) and (layer0_outputs(3728)));
    layer1_outputs(1593) <= not(layer0_outputs(3475));
    layer1_outputs(1594) <= layer0_outputs(3862);
    layer1_outputs(1595) <= (layer0_outputs(4945)) or (layer0_outputs(4948));
    layer1_outputs(1596) <= (layer0_outputs(1274)) and (layer0_outputs(220));
    layer1_outputs(1597) <= (layer0_outputs(889)) xor (layer0_outputs(899));
    layer1_outputs(1598) <= not(layer0_outputs(4031));
    layer1_outputs(1599) <= not((layer0_outputs(2713)) or (layer0_outputs(4629)));
    layer1_outputs(1600) <= not(layer0_outputs(3060));
    layer1_outputs(1601) <= layer0_outputs(4515);
    layer1_outputs(1602) <= layer0_outputs(1705);
    layer1_outputs(1603) <= layer0_outputs(4057);
    layer1_outputs(1604) <= layer0_outputs(4690);
    layer1_outputs(1605) <= not((layer0_outputs(4125)) or (layer0_outputs(4867)));
    layer1_outputs(1606) <= (layer0_outputs(1070)) or (layer0_outputs(110));
    layer1_outputs(1607) <= not(layer0_outputs(2417));
    layer1_outputs(1608) <= layer0_outputs(2990);
    layer1_outputs(1609) <= (layer0_outputs(411)) and not (layer0_outputs(181));
    layer1_outputs(1610) <= (layer0_outputs(3309)) and (layer0_outputs(319));
    layer1_outputs(1611) <= '0';
    layer1_outputs(1612) <= not((layer0_outputs(5025)) or (layer0_outputs(2696)));
    layer1_outputs(1613) <= layer0_outputs(2828);
    layer1_outputs(1614) <= not(layer0_outputs(2635));
    layer1_outputs(1615) <= (layer0_outputs(396)) or (layer0_outputs(217));
    layer1_outputs(1616) <= not((layer0_outputs(2209)) xor (layer0_outputs(1253)));
    layer1_outputs(1617) <= not(layer0_outputs(961));
    layer1_outputs(1618) <= not((layer0_outputs(4912)) or (layer0_outputs(700)));
    layer1_outputs(1619) <= not(layer0_outputs(4998)) or (layer0_outputs(3596));
    layer1_outputs(1620) <= not(layer0_outputs(2809));
    layer1_outputs(1621) <= not(layer0_outputs(411));
    layer1_outputs(1622) <= (layer0_outputs(1833)) or (layer0_outputs(715));
    layer1_outputs(1623) <= (layer0_outputs(3794)) or (layer0_outputs(5101));
    layer1_outputs(1624) <= (layer0_outputs(3951)) and not (layer0_outputs(5001));
    layer1_outputs(1625) <= '1';
    layer1_outputs(1626) <= not(layer0_outputs(3089)) or (layer0_outputs(4539));
    layer1_outputs(1627) <= not(layer0_outputs(3416));
    layer1_outputs(1628) <= not((layer0_outputs(2648)) and (layer0_outputs(3625)));
    layer1_outputs(1629) <= (layer0_outputs(3994)) or (layer0_outputs(3575));
    layer1_outputs(1630) <= layer0_outputs(3160);
    layer1_outputs(1631) <= (layer0_outputs(1850)) and not (layer0_outputs(2746));
    layer1_outputs(1632) <= (layer0_outputs(2231)) or (layer0_outputs(5084));
    layer1_outputs(1633) <= not((layer0_outputs(651)) or (layer0_outputs(151)));
    layer1_outputs(1634) <= not(layer0_outputs(1152));
    layer1_outputs(1635) <= not(layer0_outputs(394)) or (layer0_outputs(920));
    layer1_outputs(1636) <= (layer0_outputs(1789)) xor (layer0_outputs(2069));
    layer1_outputs(1637) <= (layer0_outputs(3503)) or (layer0_outputs(676));
    layer1_outputs(1638) <= not((layer0_outputs(814)) and (layer0_outputs(2279)));
    layer1_outputs(1639) <= not((layer0_outputs(2598)) and (layer0_outputs(3530)));
    layer1_outputs(1640) <= not(layer0_outputs(1224));
    layer1_outputs(1641) <= (layer0_outputs(578)) and (layer0_outputs(844));
    layer1_outputs(1642) <= layer0_outputs(3670);
    layer1_outputs(1643) <= layer0_outputs(177);
    layer1_outputs(1644) <= layer0_outputs(3729);
    layer1_outputs(1645) <= (layer0_outputs(2493)) and not (layer0_outputs(2434));
    layer1_outputs(1646) <= '1';
    layer1_outputs(1647) <= not(layer0_outputs(4886)) or (layer0_outputs(2342));
    layer1_outputs(1648) <= layer0_outputs(3086);
    layer1_outputs(1649) <= (layer0_outputs(3674)) and not (layer0_outputs(1437));
    layer1_outputs(1650) <= layer0_outputs(2154);
    layer1_outputs(1651) <= layer0_outputs(3400);
    layer1_outputs(1652) <= not(layer0_outputs(2852));
    layer1_outputs(1653) <= not(layer0_outputs(2192));
    layer1_outputs(1654) <= not(layer0_outputs(1009)) or (layer0_outputs(4193));
    layer1_outputs(1655) <= not((layer0_outputs(3940)) or (layer0_outputs(2047)));
    layer1_outputs(1656) <= (layer0_outputs(366)) and (layer0_outputs(3574));
    layer1_outputs(1657) <= not(layer0_outputs(2316)) or (layer0_outputs(4034));
    layer1_outputs(1658) <= not((layer0_outputs(3896)) and (layer0_outputs(1546)));
    layer1_outputs(1659) <= layer0_outputs(2277);
    layer1_outputs(1660) <= not(layer0_outputs(2161));
    layer1_outputs(1661) <= not(layer0_outputs(1896));
    layer1_outputs(1662) <= layer0_outputs(79);
    layer1_outputs(1663) <= (layer0_outputs(4444)) xor (layer0_outputs(457));
    layer1_outputs(1664) <= not(layer0_outputs(1605));
    layer1_outputs(1665) <= not(layer0_outputs(944)) or (layer0_outputs(162));
    layer1_outputs(1666) <= (layer0_outputs(4613)) and (layer0_outputs(4333));
    layer1_outputs(1667) <= not(layer0_outputs(4239)) or (layer0_outputs(2937));
    layer1_outputs(1668) <= not(layer0_outputs(3778)) or (layer0_outputs(3545));
    layer1_outputs(1669) <= not(layer0_outputs(2739));
    layer1_outputs(1670) <= layer0_outputs(3838);
    layer1_outputs(1671) <= not((layer0_outputs(719)) or (layer0_outputs(2169)));
    layer1_outputs(1672) <= layer0_outputs(528);
    layer1_outputs(1673) <= not(layer0_outputs(2971));
    layer1_outputs(1674) <= not(layer0_outputs(3184));
    layer1_outputs(1675) <= (layer0_outputs(1000)) or (layer0_outputs(4223));
    layer1_outputs(1676) <= not((layer0_outputs(2939)) or (layer0_outputs(40)));
    layer1_outputs(1677) <= not(layer0_outputs(4425)) or (layer0_outputs(1995));
    layer1_outputs(1678) <= layer0_outputs(41);
    layer1_outputs(1679) <= layer0_outputs(4558);
    layer1_outputs(1680) <= not(layer0_outputs(2644)) or (layer0_outputs(4588));
    layer1_outputs(1681) <= layer0_outputs(5010);
    layer1_outputs(1682) <= (layer0_outputs(1744)) or (layer0_outputs(302));
    layer1_outputs(1683) <= (layer0_outputs(1693)) and not (layer0_outputs(3038));
    layer1_outputs(1684) <= '0';
    layer1_outputs(1685) <= layer0_outputs(3496);
    layer1_outputs(1686) <= (layer0_outputs(4056)) or (layer0_outputs(139));
    layer1_outputs(1687) <= not((layer0_outputs(2781)) or (layer0_outputs(3603)));
    layer1_outputs(1688) <= not(layer0_outputs(2518)) or (layer0_outputs(3463));
    layer1_outputs(1689) <= layer0_outputs(1111);
    layer1_outputs(1690) <= '0';
    layer1_outputs(1691) <= (layer0_outputs(3298)) and (layer0_outputs(101));
    layer1_outputs(1692) <= '0';
    layer1_outputs(1693) <= not((layer0_outputs(2503)) xor (layer0_outputs(643)));
    layer1_outputs(1694) <= (layer0_outputs(4545)) and not (layer0_outputs(1425));
    layer1_outputs(1695) <= not(layer0_outputs(3791));
    layer1_outputs(1696) <= (layer0_outputs(404)) and not (layer0_outputs(3604));
    layer1_outputs(1697) <= (layer0_outputs(2431)) or (layer0_outputs(4246));
    layer1_outputs(1698) <= not((layer0_outputs(48)) xor (layer0_outputs(243)));
    layer1_outputs(1699) <= layer0_outputs(3668);
    layer1_outputs(1700) <= layer0_outputs(3751);
    layer1_outputs(1701) <= not(layer0_outputs(2580));
    layer1_outputs(1702) <= not(layer0_outputs(2735));
    layer1_outputs(1703) <= not(layer0_outputs(1326));
    layer1_outputs(1704) <= layer0_outputs(2515);
    layer1_outputs(1705) <= (layer0_outputs(2419)) and not (layer0_outputs(3368));
    layer1_outputs(1706) <= not(layer0_outputs(4002)) or (layer0_outputs(3090));
    layer1_outputs(1707) <= not((layer0_outputs(3929)) xor (layer0_outputs(4188)));
    layer1_outputs(1708) <= not(layer0_outputs(3510));
    layer1_outputs(1709) <= not((layer0_outputs(4410)) and (layer0_outputs(4512)));
    layer1_outputs(1710) <= layer0_outputs(4481);
    layer1_outputs(1711) <= layer0_outputs(1225);
    layer1_outputs(1712) <= not(layer0_outputs(1387));
    layer1_outputs(1713) <= layer0_outputs(1399);
    layer1_outputs(1714) <= (layer0_outputs(1950)) and (layer0_outputs(1666));
    layer1_outputs(1715) <= (layer0_outputs(4783)) and not (layer0_outputs(4953));
    layer1_outputs(1716) <= not(layer0_outputs(4709));
    layer1_outputs(1717) <= not(layer0_outputs(1574));
    layer1_outputs(1718) <= not((layer0_outputs(4090)) or (layer0_outputs(4678)));
    layer1_outputs(1719) <= (layer0_outputs(529)) and (layer0_outputs(2804));
    layer1_outputs(1720) <= layer0_outputs(2558);
    layer1_outputs(1721) <= (layer0_outputs(434)) and (layer0_outputs(1524));
    layer1_outputs(1722) <= not(layer0_outputs(3485));
    layer1_outputs(1723) <= not(layer0_outputs(4100)) or (layer0_outputs(1740));
    layer1_outputs(1724) <= not(layer0_outputs(4075));
    layer1_outputs(1725) <= (layer0_outputs(221)) and (layer0_outputs(4709));
    layer1_outputs(1726) <= not((layer0_outputs(2780)) xor (layer0_outputs(1840)));
    layer1_outputs(1727) <= not(layer0_outputs(288));
    layer1_outputs(1728) <= not((layer0_outputs(3122)) or (layer0_outputs(1189)));
    layer1_outputs(1729) <= '1';
    layer1_outputs(1730) <= (layer0_outputs(467)) and not (layer0_outputs(4264));
    layer1_outputs(1731) <= not(layer0_outputs(227));
    layer1_outputs(1732) <= (layer0_outputs(2970)) and (layer0_outputs(4522));
    layer1_outputs(1733) <= layer0_outputs(839);
    layer1_outputs(1734) <= '0';
    layer1_outputs(1735) <= not(layer0_outputs(3840)) or (layer0_outputs(2668));
    layer1_outputs(1736) <= not(layer0_outputs(1379)) or (layer0_outputs(4356));
    layer1_outputs(1737) <= (layer0_outputs(1812)) and not (layer0_outputs(4351));
    layer1_outputs(1738) <= (layer0_outputs(2274)) xor (layer0_outputs(116));
    layer1_outputs(1739) <= (layer0_outputs(580)) and not (layer0_outputs(500));
    layer1_outputs(1740) <= not(layer0_outputs(2221)) or (layer0_outputs(1387));
    layer1_outputs(1741) <= layer0_outputs(4385);
    layer1_outputs(1742) <= not((layer0_outputs(3946)) or (layer0_outputs(562)));
    layer1_outputs(1743) <= (layer0_outputs(1708)) and not (layer0_outputs(4340));
    layer1_outputs(1744) <= not(layer0_outputs(4199));
    layer1_outputs(1745) <= '1';
    layer1_outputs(1746) <= not(layer0_outputs(1701));
    layer1_outputs(1747) <= not((layer0_outputs(633)) and (layer0_outputs(4971)));
    layer1_outputs(1748) <= layer0_outputs(442);
    layer1_outputs(1749) <= (layer0_outputs(3218)) and not (layer0_outputs(4505));
    layer1_outputs(1750) <= not(layer0_outputs(232)) or (layer0_outputs(1540));
    layer1_outputs(1751) <= not(layer0_outputs(3744)) or (layer0_outputs(63));
    layer1_outputs(1752) <= layer0_outputs(4542);
    layer1_outputs(1753) <= not(layer0_outputs(1831));
    layer1_outputs(1754) <= not(layer0_outputs(1018));
    layer1_outputs(1755) <= not(layer0_outputs(3905));
    layer1_outputs(1756) <= (layer0_outputs(2107)) and not (layer0_outputs(1865));
    layer1_outputs(1757) <= (layer0_outputs(3974)) xor (layer0_outputs(4696));
    layer1_outputs(1758) <= not(layer0_outputs(5112));
    layer1_outputs(1759) <= (layer0_outputs(579)) and (layer0_outputs(4511));
    layer1_outputs(1760) <= not(layer0_outputs(513));
    layer1_outputs(1761) <= (layer0_outputs(4659)) and not (layer0_outputs(171));
    layer1_outputs(1762) <= layer0_outputs(5035);
    layer1_outputs(1763) <= (layer0_outputs(3035)) xor (layer0_outputs(2152));
    layer1_outputs(1764) <= (layer0_outputs(2444)) and (layer0_outputs(206));
    layer1_outputs(1765) <= (layer0_outputs(1007)) and (layer0_outputs(1562));
    layer1_outputs(1766) <= '1';
    layer1_outputs(1767) <= (layer0_outputs(2974)) xor (layer0_outputs(4612));
    layer1_outputs(1768) <= not((layer0_outputs(1907)) and (layer0_outputs(1871)));
    layer1_outputs(1769) <= not(layer0_outputs(2908)) or (layer0_outputs(415));
    layer1_outputs(1770) <= not(layer0_outputs(1607)) or (layer0_outputs(475));
    layer1_outputs(1771) <= not(layer0_outputs(510)) or (layer0_outputs(3622));
    layer1_outputs(1772) <= '0';
    layer1_outputs(1773) <= layer0_outputs(3190);
    layer1_outputs(1774) <= not(layer0_outputs(2195));
    layer1_outputs(1775) <= layer0_outputs(1561);
    layer1_outputs(1776) <= not(layer0_outputs(3890)) or (layer0_outputs(2037));
    layer1_outputs(1777) <= (layer0_outputs(4647)) and not (layer0_outputs(577));
    layer1_outputs(1778) <= not((layer0_outputs(1319)) xor (layer0_outputs(2702)));
    layer1_outputs(1779) <= not((layer0_outputs(3012)) or (layer0_outputs(3576)));
    layer1_outputs(1780) <= (layer0_outputs(1767)) xor (layer0_outputs(3527));
    layer1_outputs(1781) <= '1';
    layer1_outputs(1782) <= not((layer0_outputs(2335)) or (layer0_outputs(3337)));
    layer1_outputs(1783) <= layer0_outputs(4293);
    layer1_outputs(1784) <= layer0_outputs(3196);
    layer1_outputs(1785) <= layer0_outputs(306);
    layer1_outputs(1786) <= layer0_outputs(2316);
    layer1_outputs(1787) <= not((layer0_outputs(4297)) and (layer0_outputs(2429)));
    layer1_outputs(1788) <= layer0_outputs(4840);
    layer1_outputs(1789) <= not(layer0_outputs(1927));
    layer1_outputs(1790) <= not(layer0_outputs(3968));
    layer1_outputs(1791) <= (layer0_outputs(3407)) xor (layer0_outputs(4701));
    layer1_outputs(1792) <= layer0_outputs(4835);
    layer1_outputs(1793) <= layer0_outputs(1390);
    layer1_outputs(1794) <= not(layer0_outputs(4384));
    layer1_outputs(1795) <= (layer0_outputs(1867)) and not (layer0_outputs(2545));
    layer1_outputs(1796) <= not((layer0_outputs(1419)) or (layer0_outputs(1662)));
    layer1_outputs(1797) <= not(layer0_outputs(2539));
    layer1_outputs(1798) <= (layer0_outputs(3575)) and (layer0_outputs(3663));
    layer1_outputs(1799) <= (layer0_outputs(2652)) and (layer0_outputs(1820));
    layer1_outputs(1800) <= not(layer0_outputs(2260)) or (layer0_outputs(3559));
    layer1_outputs(1801) <= not((layer0_outputs(4438)) xor (layer0_outputs(4041)));
    layer1_outputs(1802) <= not((layer0_outputs(1181)) or (layer0_outputs(160)));
    layer1_outputs(1803) <= not(layer0_outputs(1604));
    layer1_outputs(1804) <= '1';
    layer1_outputs(1805) <= not(layer0_outputs(5029));
    layer1_outputs(1806) <= not(layer0_outputs(4227));
    layer1_outputs(1807) <= (layer0_outputs(432)) xor (layer0_outputs(2123));
    layer1_outputs(1808) <= (layer0_outputs(3509)) and (layer0_outputs(692));
    layer1_outputs(1809) <= (layer0_outputs(4972)) or (layer0_outputs(3416));
    layer1_outputs(1810) <= (layer0_outputs(2909)) xor (layer0_outputs(2097));
    layer1_outputs(1811) <= not(layer0_outputs(911));
    layer1_outputs(1812) <= (layer0_outputs(2347)) or (layer0_outputs(2906));
    layer1_outputs(1813) <= (layer0_outputs(4699)) or (layer0_outputs(2870));
    layer1_outputs(1814) <= not(layer0_outputs(4345)) or (layer0_outputs(1981));
    layer1_outputs(1815) <= not(layer0_outputs(3507));
    layer1_outputs(1816) <= (layer0_outputs(4266)) and not (layer0_outputs(3560));
    layer1_outputs(1817) <= (layer0_outputs(2070)) and not (layer0_outputs(1491));
    layer1_outputs(1818) <= layer0_outputs(3675);
    layer1_outputs(1819) <= (layer0_outputs(729)) or (layer0_outputs(1846));
    layer1_outputs(1820) <= layer0_outputs(3779);
    layer1_outputs(1821) <= layer0_outputs(685);
    layer1_outputs(1822) <= (layer0_outputs(2535)) or (layer0_outputs(1355));
    layer1_outputs(1823) <= not(layer0_outputs(1324));
    layer1_outputs(1824) <= not(layer0_outputs(3361));
    layer1_outputs(1825) <= not(layer0_outputs(4271));
    layer1_outputs(1826) <= not(layer0_outputs(4649)) or (layer0_outputs(3846));
    layer1_outputs(1827) <= not(layer0_outputs(3592));
    layer1_outputs(1828) <= layer0_outputs(4142);
    layer1_outputs(1829) <= not(layer0_outputs(4797)) or (layer0_outputs(2998));
    layer1_outputs(1830) <= (layer0_outputs(2615)) and (layer0_outputs(2537));
    layer1_outputs(1831) <= not((layer0_outputs(4440)) or (layer0_outputs(332)));
    layer1_outputs(1832) <= not((layer0_outputs(1182)) and (layer0_outputs(2861)));
    layer1_outputs(1833) <= layer0_outputs(3152);
    layer1_outputs(1834) <= not(layer0_outputs(4246));
    layer1_outputs(1835) <= layer0_outputs(4483);
    layer1_outputs(1836) <= (layer0_outputs(4893)) and not (layer0_outputs(4408));
    layer1_outputs(1837) <= not(layer0_outputs(4213));
    layer1_outputs(1838) <= not(layer0_outputs(1686));
    layer1_outputs(1839) <= not(layer0_outputs(3680));
    layer1_outputs(1840) <= not(layer0_outputs(214));
    layer1_outputs(1841) <= (layer0_outputs(2651)) and not (layer0_outputs(615));
    layer1_outputs(1842) <= (layer0_outputs(2085)) and not (layer0_outputs(4092));
    layer1_outputs(1843) <= (layer0_outputs(4250)) and (layer0_outputs(1586));
    layer1_outputs(1844) <= layer0_outputs(22);
    layer1_outputs(1845) <= not((layer0_outputs(3023)) and (layer0_outputs(3988)));
    layer1_outputs(1846) <= (layer0_outputs(4745)) and (layer0_outputs(5087));
    layer1_outputs(1847) <= (layer0_outputs(2785)) or (layer0_outputs(1588));
    layer1_outputs(1848) <= layer0_outputs(2450);
    layer1_outputs(1849) <= (layer0_outputs(4550)) and not (layer0_outputs(1100));
    layer1_outputs(1850) <= not((layer0_outputs(3937)) and (layer0_outputs(2143)));
    layer1_outputs(1851) <= not(layer0_outputs(4910)) or (layer0_outputs(119));
    layer1_outputs(1852) <= (layer0_outputs(3314)) or (layer0_outputs(1349));
    layer1_outputs(1853) <= not(layer0_outputs(4019));
    layer1_outputs(1854) <= not(layer0_outputs(4032));
    layer1_outputs(1855) <= (layer0_outputs(3242)) or (layer0_outputs(1694));
    layer1_outputs(1856) <= (layer0_outputs(4287)) and not (layer0_outputs(1072));
    layer1_outputs(1857) <= not(layer0_outputs(1479)) or (layer0_outputs(3613));
    layer1_outputs(1858) <= not(layer0_outputs(951));
    layer1_outputs(1859) <= not((layer0_outputs(1644)) or (layer0_outputs(2273)));
    layer1_outputs(1860) <= not(layer0_outputs(2073));
    layer1_outputs(1861) <= not(layer0_outputs(555));
    layer1_outputs(1862) <= (layer0_outputs(3494)) and not (layer0_outputs(2087));
    layer1_outputs(1863) <= not(layer0_outputs(2822));
    layer1_outputs(1864) <= layer0_outputs(3367);
    layer1_outputs(1865) <= not(layer0_outputs(1340));
    layer1_outputs(1866) <= not(layer0_outputs(1695));
    layer1_outputs(1867) <= layer0_outputs(4397);
    layer1_outputs(1868) <= layer0_outputs(1415);
    layer1_outputs(1869) <= layer0_outputs(1371);
    layer1_outputs(1870) <= not((layer0_outputs(2113)) or (layer0_outputs(4141)));
    layer1_outputs(1871) <= not((layer0_outputs(4488)) xor (layer0_outputs(3173)));
    layer1_outputs(1872) <= (layer0_outputs(12)) and not (layer0_outputs(601));
    layer1_outputs(1873) <= not(layer0_outputs(1303));
    layer1_outputs(1874) <= not((layer0_outputs(93)) and (layer0_outputs(1936)));
    layer1_outputs(1875) <= not(layer0_outputs(2687));
    layer1_outputs(1876) <= not(layer0_outputs(3465));
    layer1_outputs(1877) <= not(layer0_outputs(3386));
    layer1_outputs(1878) <= not(layer0_outputs(3135)) or (layer0_outputs(1612));
    layer1_outputs(1879) <= layer0_outputs(3234);
    layer1_outputs(1880) <= not(layer0_outputs(3850));
    layer1_outputs(1881) <= (layer0_outputs(3233)) and not (layer0_outputs(3597));
    layer1_outputs(1882) <= not(layer0_outputs(4590));
    layer1_outputs(1883) <= not(layer0_outputs(1206)) or (layer0_outputs(4022));
    layer1_outputs(1884) <= layer0_outputs(4503);
    layer1_outputs(1885) <= (layer0_outputs(2080)) and not (layer0_outputs(4430));
    layer1_outputs(1886) <= (layer0_outputs(4458)) and not (layer0_outputs(3489));
    layer1_outputs(1887) <= not(layer0_outputs(3886)) or (layer0_outputs(2369));
    layer1_outputs(1888) <= not((layer0_outputs(4118)) and (layer0_outputs(1852)));
    layer1_outputs(1889) <= layer0_outputs(1503);
    layer1_outputs(1890) <= '0';
    layer1_outputs(1891) <= layer0_outputs(1136);
    layer1_outputs(1892) <= not(layer0_outputs(2530)) or (layer0_outputs(285));
    layer1_outputs(1893) <= '0';
    layer1_outputs(1894) <= not(layer0_outputs(3094));
    layer1_outputs(1895) <= (layer0_outputs(3672)) and not (layer0_outputs(196));
    layer1_outputs(1896) <= not(layer0_outputs(2424)) or (layer0_outputs(3289));
    layer1_outputs(1897) <= not(layer0_outputs(302)) or (layer0_outputs(4332));
    layer1_outputs(1898) <= not(layer0_outputs(3901));
    layer1_outputs(1899) <= (layer0_outputs(3881)) and not (layer0_outputs(4506));
    layer1_outputs(1900) <= not(layer0_outputs(892));
    layer1_outputs(1901) <= not(layer0_outputs(570));
    layer1_outputs(1902) <= not(layer0_outputs(1337));
    layer1_outputs(1903) <= not((layer0_outputs(1309)) xor (layer0_outputs(3082)));
    layer1_outputs(1904) <= not(layer0_outputs(1413)) or (layer0_outputs(361));
    layer1_outputs(1905) <= not(layer0_outputs(507));
    layer1_outputs(1906) <= not(layer0_outputs(3152));
    layer1_outputs(1907) <= layer0_outputs(3156);
    layer1_outputs(1908) <= not(layer0_outputs(2247));
    layer1_outputs(1909) <= not(layer0_outputs(2709));
    layer1_outputs(1910) <= (layer0_outputs(201)) and (layer0_outputs(765));
    layer1_outputs(1911) <= (layer0_outputs(666)) or (layer0_outputs(617));
    layer1_outputs(1912) <= (layer0_outputs(2322)) and not (layer0_outputs(3638));
    layer1_outputs(1913) <= layer0_outputs(1411);
    layer1_outputs(1914) <= (layer0_outputs(4790)) and (layer0_outputs(1559));
    layer1_outputs(1915) <= not((layer0_outputs(3480)) and (layer0_outputs(2080)));
    layer1_outputs(1916) <= layer0_outputs(2433);
    layer1_outputs(1917) <= (layer0_outputs(3978)) and not (layer0_outputs(3540));
    layer1_outputs(1918) <= (layer0_outputs(4812)) or (layer0_outputs(1063));
    layer1_outputs(1919) <= '0';
    layer1_outputs(1920) <= (layer0_outputs(4412)) and (layer0_outputs(3709));
    layer1_outputs(1921) <= not(layer0_outputs(1533));
    layer1_outputs(1922) <= '0';
    layer1_outputs(1923) <= (layer0_outputs(4920)) and (layer0_outputs(2365));
    layer1_outputs(1924) <= not(layer0_outputs(5026));
    layer1_outputs(1925) <= (layer0_outputs(4258)) and (layer0_outputs(3440));
    layer1_outputs(1926) <= not(layer0_outputs(1255));
    layer1_outputs(1927) <= not(layer0_outputs(95));
    layer1_outputs(1928) <= layer0_outputs(3579);
    layer1_outputs(1929) <= not(layer0_outputs(4182));
    layer1_outputs(1930) <= (layer0_outputs(304)) and not (layer0_outputs(3223));
    layer1_outputs(1931) <= not(layer0_outputs(4156));
    layer1_outputs(1932) <= not(layer0_outputs(4203));
    layer1_outputs(1933) <= layer0_outputs(2724);
    layer1_outputs(1934) <= not(layer0_outputs(1584)) or (layer0_outputs(3276));
    layer1_outputs(1935) <= not(layer0_outputs(350));
    layer1_outputs(1936) <= '0';
    layer1_outputs(1937) <= (layer0_outputs(7)) or (layer0_outputs(1079));
    layer1_outputs(1938) <= layer0_outputs(4016);
    layer1_outputs(1939) <= not(layer0_outputs(184));
    layer1_outputs(1940) <= not(layer0_outputs(331));
    layer1_outputs(1941) <= not(layer0_outputs(4431)) or (layer0_outputs(2215));
    layer1_outputs(1942) <= not(layer0_outputs(3260));
    layer1_outputs(1943) <= (layer0_outputs(930)) and (layer0_outputs(3573));
    layer1_outputs(1944) <= layer0_outputs(4382);
    layer1_outputs(1945) <= (layer0_outputs(1916)) and not (layer0_outputs(1296));
    layer1_outputs(1946) <= (layer0_outputs(2388)) and (layer0_outputs(3487));
    layer1_outputs(1947) <= (layer0_outputs(3621)) and not (layer0_outputs(3847));
    layer1_outputs(1948) <= not(layer0_outputs(4773)) or (layer0_outputs(2305));
    layer1_outputs(1949) <= not((layer0_outputs(495)) and (layer0_outputs(2742)));
    layer1_outputs(1950) <= layer0_outputs(3165);
    layer1_outputs(1951) <= not(layer0_outputs(455)) or (layer0_outputs(147));
    layer1_outputs(1952) <= layer0_outputs(1413);
    layer1_outputs(1953) <= (layer0_outputs(3999)) and (layer0_outputs(3531));
    layer1_outputs(1954) <= not((layer0_outputs(926)) xor (layer0_outputs(4165)));
    layer1_outputs(1955) <= not(layer0_outputs(199));
    layer1_outputs(1956) <= layer0_outputs(4071);
    layer1_outputs(1957) <= not(layer0_outputs(4550)) or (layer0_outputs(3742));
    layer1_outputs(1958) <= not(layer0_outputs(166)) or (layer0_outputs(2163));
    layer1_outputs(1959) <= not(layer0_outputs(4802)) or (layer0_outputs(872));
    layer1_outputs(1960) <= not(layer0_outputs(3043));
    layer1_outputs(1961) <= (layer0_outputs(4513)) and not (layer0_outputs(2466));
    layer1_outputs(1962) <= not(layer0_outputs(498));
    layer1_outputs(1963) <= not(layer0_outputs(307));
    layer1_outputs(1964) <= (layer0_outputs(4235)) or (layer0_outputs(1095));
    layer1_outputs(1965) <= (layer0_outputs(2915)) and (layer0_outputs(315));
    layer1_outputs(1966) <= (layer0_outputs(2854)) and (layer0_outputs(740));
    layer1_outputs(1967) <= not((layer0_outputs(2428)) xor (layer0_outputs(1542)));
    layer1_outputs(1968) <= not(layer0_outputs(1617)) or (layer0_outputs(1085));
    layer1_outputs(1969) <= not((layer0_outputs(3970)) and (layer0_outputs(2969)));
    layer1_outputs(1970) <= not(layer0_outputs(4919)) or (layer0_outputs(4521));
    layer1_outputs(1971) <= '0';
    layer1_outputs(1972) <= layer0_outputs(4852);
    layer1_outputs(1973) <= not(layer0_outputs(5028));
    layer1_outputs(1974) <= not((layer0_outputs(3707)) or (layer0_outputs(3807)));
    layer1_outputs(1975) <= not((layer0_outputs(2337)) xor (layer0_outputs(53)));
    layer1_outputs(1976) <= (layer0_outputs(780)) and not (layer0_outputs(918));
    layer1_outputs(1977) <= not(layer0_outputs(4272));
    layer1_outputs(1978) <= (layer0_outputs(2584)) or (layer0_outputs(1435));
    layer1_outputs(1979) <= '0';
    layer1_outputs(1980) <= not(layer0_outputs(2229));
    layer1_outputs(1981) <= not((layer0_outputs(3091)) xor (layer0_outputs(4784)));
    layer1_outputs(1982) <= (layer0_outputs(4602)) and (layer0_outputs(2768));
    layer1_outputs(1983) <= layer0_outputs(509);
    layer1_outputs(1984) <= (layer0_outputs(365)) and (layer0_outputs(4767));
    layer1_outputs(1985) <= not(layer0_outputs(480));
    layer1_outputs(1986) <= not((layer0_outputs(2380)) or (layer0_outputs(745)));
    layer1_outputs(1987) <= (layer0_outputs(1361)) and (layer0_outputs(3900));
    layer1_outputs(1988) <= layer0_outputs(1040);
    layer1_outputs(1989) <= not(layer0_outputs(4163)) or (layer0_outputs(963));
    layer1_outputs(1990) <= (layer0_outputs(2891)) and (layer0_outputs(3306));
    layer1_outputs(1991) <= layer0_outputs(1550);
    layer1_outputs(1992) <= not((layer0_outputs(1273)) and (layer0_outputs(614)));
    layer1_outputs(1993) <= (layer0_outputs(2808)) or (layer0_outputs(3192));
    layer1_outputs(1994) <= not(layer0_outputs(1490));
    layer1_outputs(1995) <= layer0_outputs(834);
    layer1_outputs(1996) <= not(layer0_outputs(1991));
    layer1_outputs(1997) <= (layer0_outputs(895)) and (layer0_outputs(4189));
    layer1_outputs(1998) <= (layer0_outputs(35)) or (layer0_outputs(356));
    layer1_outputs(1999) <= not(layer0_outputs(1786)) or (layer0_outputs(3191));
    layer1_outputs(2000) <= not(layer0_outputs(603)) or (layer0_outputs(4421));
    layer1_outputs(2001) <= not(layer0_outputs(1841));
    layer1_outputs(2002) <= not(layer0_outputs(5116)) or (layer0_outputs(2490));
    layer1_outputs(2003) <= not(layer0_outputs(1575)) or (layer0_outputs(1618));
    layer1_outputs(2004) <= not(layer0_outputs(1665)) or (layer0_outputs(2929));
    layer1_outputs(2005) <= not((layer0_outputs(4454)) or (layer0_outputs(3230)));
    layer1_outputs(2006) <= not(layer0_outputs(1463)) or (layer0_outputs(466));
    layer1_outputs(2007) <= '1';
    layer1_outputs(2008) <= not(layer0_outputs(3565)) or (layer0_outputs(2350));
    layer1_outputs(2009) <= layer0_outputs(1501);
    layer1_outputs(2010) <= layer0_outputs(1791);
    layer1_outputs(2011) <= (layer0_outputs(2414)) and (layer0_outputs(4161));
    layer1_outputs(2012) <= (layer0_outputs(2125)) xor (layer0_outputs(338));
    layer1_outputs(2013) <= not(layer0_outputs(1383));
    layer1_outputs(2014) <= not(layer0_outputs(551));
    layer1_outputs(2015) <= (layer0_outputs(1391)) and (layer0_outputs(326));
    layer1_outputs(2016) <= layer0_outputs(2641);
    layer1_outputs(2017) <= (layer0_outputs(1455)) and (layer0_outputs(1215));
    layer1_outputs(2018) <= '0';
    layer1_outputs(2019) <= not(layer0_outputs(92));
    layer1_outputs(2020) <= (layer0_outputs(4919)) and not (layer0_outputs(487));
    layer1_outputs(2021) <= not(layer0_outputs(4281)) or (layer0_outputs(2631));
    layer1_outputs(2022) <= not(layer0_outputs(4642));
    layer1_outputs(2023) <= layer0_outputs(4697);
    layer1_outputs(2024) <= '1';
    layer1_outputs(2025) <= layer0_outputs(967);
    layer1_outputs(2026) <= layer0_outputs(3020);
    layer1_outputs(2027) <= layer0_outputs(3811);
    layer1_outputs(2028) <= not(layer0_outputs(4543)) or (layer0_outputs(4689));
    layer1_outputs(2029) <= not((layer0_outputs(841)) or (layer0_outputs(99)));
    layer1_outputs(2030) <= (layer0_outputs(173)) or (layer0_outputs(3473));
    layer1_outputs(2031) <= not(layer0_outputs(4526)) or (layer0_outputs(3329));
    layer1_outputs(2032) <= layer0_outputs(255);
    layer1_outputs(2033) <= not((layer0_outputs(2138)) and (layer0_outputs(4127)));
    layer1_outputs(2034) <= not((layer0_outputs(4818)) xor (layer0_outputs(4177)));
    layer1_outputs(2035) <= (layer0_outputs(4218)) and not (layer0_outputs(1841));
    layer1_outputs(2036) <= not((layer0_outputs(3341)) or (layer0_outputs(1225)));
    layer1_outputs(2037) <= not(layer0_outputs(36));
    layer1_outputs(2038) <= not((layer0_outputs(3227)) and (layer0_outputs(1200)));
    layer1_outputs(2039) <= (layer0_outputs(3925)) or (layer0_outputs(799));
    layer1_outputs(2040) <= (layer0_outputs(3425)) or (layer0_outputs(5048));
    layer1_outputs(2041) <= (layer0_outputs(4571)) and not (layer0_outputs(1932));
    layer1_outputs(2042) <= not(layer0_outputs(3151)) or (layer0_outputs(2792));
    layer1_outputs(2043) <= (layer0_outputs(4082)) and not (layer0_outputs(4172));
    layer1_outputs(2044) <= (layer0_outputs(194)) and not (layer0_outputs(1342));
    layer1_outputs(2045) <= '0';
    layer1_outputs(2046) <= not((layer0_outputs(2248)) and (layer0_outputs(301)));
    layer1_outputs(2047) <= not(layer0_outputs(5035));
    layer1_outputs(2048) <= not(layer0_outputs(1973));
    layer1_outputs(2049) <= not(layer0_outputs(4237));
    layer1_outputs(2050) <= (layer0_outputs(2111)) and (layer0_outputs(1317));
    layer1_outputs(2051) <= (layer0_outputs(2378)) and not (layer0_outputs(1932));
    layer1_outputs(2052) <= (layer0_outputs(3863)) and (layer0_outputs(2503));
    layer1_outputs(2053) <= layer0_outputs(1313);
    layer1_outputs(2054) <= not(layer0_outputs(4377));
    layer1_outputs(2055) <= not((layer0_outputs(5119)) and (layer0_outputs(2159)));
    layer1_outputs(2056) <= (layer0_outputs(3036)) and not (layer0_outputs(3611));
    layer1_outputs(2057) <= (layer0_outputs(2734)) xor (layer0_outputs(1438));
    layer1_outputs(2058) <= not((layer0_outputs(3484)) or (layer0_outputs(38)));
    layer1_outputs(2059) <= not(layer0_outputs(3867)) or (layer0_outputs(3981));
    layer1_outputs(2060) <= not(layer0_outputs(3389));
    layer1_outputs(2061) <= layer0_outputs(3231);
    layer1_outputs(2062) <= (layer0_outputs(3885)) and (layer0_outputs(2567));
    layer1_outputs(2063) <= (layer0_outputs(4676)) and (layer0_outputs(3713));
    layer1_outputs(2064) <= not(layer0_outputs(578)) or (layer0_outputs(3018));
    layer1_outputs(2065) <= (layer0_outputs(3258)) or (layer0_outputs(4899));
    layer1_outputs(2066) <= not(layer0_outputs(3998)) or (layer0_outputs(808));
    layer1_outputs(2067) <= not(layer0_outputs(2304)) or (layer0_outputs(4786));
    layer1_outputs(2068) <= layer0_outputs(2338);
    layer1_outputs(2069) <= not(layer0_outputs(1914));
    layer1_outputs(2070) <= (layer0_outputs(5022)) and not (layer0_outputs(2955));
    layer1_outputs(2071) <= layer0_outputs(3614);
    layer1_outputs(2072) <= (layer0_outputs(2175)) or (layer0_outputs(2859));
    layer1_outputs(2073) <= not(layer0_outputs(1232));
    layer1_outputs(2074) <= (layer0_outputs(789)) and not (layer0_outputs(4866));
    layer1_outputs(2075) <= not(layer0_outputs(3571)) or (layer0_outputs(1760));
    layer1_outputs(2076) <= (layer0_outputs(3819)) and not (layer0_outputs(2891));
    layer1_outputs(2077) <= not(layer0_outputs(3249));
    layer1_outputs(2078) <= not(layer0_outputs(3126));
    layer1_outputs(2079) <= not(layer0_outputs(1338)) or (layer0_outputs(711));
    layer1_outputs(2080) <= (layer0_outputs(2262)) and not (layer0_outputs(1658));
    layer1_outputs(2081) <= layer0_outputs(3802);
    layer1_outputs(2082) <= not(layer0_outputs(670));
    layer1_outputs(2083) <= not(layer0_outputs(4748)) or (layer0_outputs(863));
    layer1_outputs(2084) <= (layer0_outputs(2795)) and (layer0_outputs(1381));
    layer1_outputs(2085) <= not(layer0_outputs(920));
    layer1_outputs(2086) <= not(layer0_outputs(2031)) or (layer0_outputs(2973));
    layer1_outputs(2087) <= not(layer0_outputs(2476));
    layer1_outputs(2088) <= not(layer0_outputs(1256));
    layer1_outputs(2089) <= not(layer0_outputs(4240));
    layer1_outputs(2090) <= not(layer0_outputs(4509));
    layer1_outputs(2091) <= (layer0_outputs(3141)) or (layer0_outputs(4541));
    layer1_outputs(2092) <= not((layer0_outputs(3565)) xor (layer0_outputs(3952)));
    layer1_outputs(2093) <= not(layer0_outputs(5055)) or (layer0_outputs(1824));
    layer1_outputs(2094) <= (layer0_outputs(1457)) and not (layer0_outputs(3720));
    layer1_outputs(2095) <= '1';
    layer1_outputs(2096) <= not(layer0_outputs(4949)) or (layer0_outputs(3938));
    layer1_outputs(2097) <= not((layer0_outputs(3542)) or (layer0_outputs(4418)));
    layer1_outputs(2098) <= not(layer0_outputs(1909)) or (layer0_outputs(1967));
    layer1_outputs(2099) <= layer0_outputs(461);
    layer1_outputs(2100) <= (layer0_outputs(3192)) and (layer0_outputs(91));
    layer1_outputs(2101) <= (layer0_outputs(1192)) and (layer0_outputs(4930));
    layer1_outputs(2102) <= not(layer0_outputs(1309)) or (layer0_outputs(2461));
    layer1_outputs(2103) <= not(layer0_outputs(734)) or (layer0_outputs(514));
    layer1_outputs(2104) <= not((layer0_outputs(30)) and (layer0_outputs(3428)));
    layer1_outputs(2105) <= (layer0_outputs(1068)) and not (layer0_outputs(2024));
    layer1_outputs(2106) <= (layer0_outputs(4941)) or (layer0_outputs(1469));
    layer1_outputs(2107) <= (layer0_outputs(4296)) and (layer0_outputs(2864));
    layer1_outputs(2108) <= (layer0_outputs(4552)) and (layer0_outputs(833));
    layer1_outputs(2109) <= not(layer0_outputs(3668)) or (layer0_outputs(4104));
    layer1_outputs(2110) <= not(layer0_outputs(102));
    layer1_outputs(2111) <= layer0_outputs(2951);
    layer1_outputs(2112) <= layer0_outputs(2381);
    layer1_outputs(2113) <= not(layer0_outputs(1478));
    layer1_outputs(2114) <= not(layer0_outputs(281));
    layer1_outputs(2115) <= (layer0_outputs(4859)) and not (layer0_outputs(3972));
    layer1_outputs(2116) <= layer0_outputs(3563);
    layer1_outputs(2117) <= (layer0_outputs(4997)) and not (layer0_outputs(4651));
    layer1_outputs(2118) <= not((layer0_outputs(2496)) xor (layer0_outputs(3420)));
    layer1_outputs(2119) <= (layer0_outputs(722)) and (layer0_outputs(359));
    layer1_outputs(2120) <= layer0_outputs(759);
    layer1_outputs(2121) <= (layer0_outputs(270)) and not (layer0_outputs(2935));
    layer1_outputs(2122) <= not((layer0_outputs(1647)) or (layer0_outputs(449)));
    layer1_outputs(2123) <= (layer0_outputs(1594)) xor (layer0_outputs(2331));
    layer1_outputs(2124) <= not((layer0_outputs(3132)) xor (layer0_outputs(1206)));
    layer1_outputs(2125) <= not(layer0_outputs(2465));
    layer1_outputs(2126) <= (layer0_outputs(2426)) and not (layer0_outputs(3719));
    layer1_outputs(2127) <= (layer0_outputs(2324)) and (layer0_outputs(2035));
    layer1_outputs(2128) <= (layer0_outputs(1065)) and (layer0_outputs(1913));
    layer1_outputs(2129) <= not(layer0_outputs(2714));
    layer1_outputs(2130) <= layer0_outputs(4388);
    layer1_outputs(2131) <= '0';
    layer1_outputs(2132) <= not(layer0_outputs(2856));
    layer1_outputs(2133) <= (layer0_outputs(614)) xor (layer0_outputs(1581));
    layer1_outputs(2134) <= not(layer0_outputs(3447)) or (layer0_outputs(2591));
    layer1_outputs(2135) <= (layer0_outputs(2682)) or (layer0_outputs(3450));
    layer1_outputs(2136) <= not(layer0_outputs(870)) or (layer0_outputs(3964));
    layer1_outputs(2137) <= not(layer0_outputs(1703));
    layer1_outputs(2138) <= not(layer0_outputs(4721)) or (layer0_outputs(831));
    layer1_outputs(2139) <= layer0_outputs(4069);
    layer1_outputs(2140) <= not((layer0_outputs(1106)) and (layer0_outputs(1659)));
    layer1_outputs(2141) <= layer0_outputs(565);
    layer1_outputs(2142) <= (layer0_outputs(13)) or (layer0_outputs(1694));
    layer1_outputs(2143) <= layer0_outputs(3486);
    layer1_outputs(2144) <= '0';
    layer1_outputs(2145) <= not(layer0_outputs(4076));
    layer1_outputs(2146) <= (layer0_outputs(4573)) or (layer0_outputs(64));
    layer1_outputs(2147) <= layer0_outputs(1739);
    layer1_outputs(2148) <= (layer0_outputs(2958)) or (layer0_outputs(4732));
    layer1_outputs(2149) <= not(layer0_outputs(2610));
    layer1_outputs(2150) <= layer0_outputs(3920);
    layer1_outputs(2151) <= layer0_outputs(3891);
    layer1_outputs(2152) <= not(layer0_outputs(4579));
    layer1_outputs(2153) <= not(layer0_outputs(1374));
    layer1_outputs(2154) <= not((layer0_outputs(2099)) or (layer0_outputs(2762)));
    layer1_outputs(2155) <= layer0_outputs(3598);
    layer1_outputs(2156) <= not((layer0_outputs(2830)) xor (layer0_outputs(3054)));
    layer1_outputs(2157) <= not(layer0_outputs(1235)) or (layer0_outputs(2736));
    layer1_outputs(2158) <= not((layer0_outputs(338)) or (layer0_outputs(1096)));
    layer1_outputs(2159) <= not(layer0_outputs(4580));
    layer1_outputs(2160) <= layer0_outputs(3005);
    layer1_outputs(2161) <= (layer0_outputs(5079)) and not (layer0_outputs(1159));
    layer1_outputs(2162) <= (layer0_outputs(925)) and (layer0_outputs(2866));
    layer1_outputs(2163) <= layer0_outputs(688);
    layer1_outputs(2164) <= (layer0_outputs(1248)) or (layer0_outputs(2110));
    layer1_outputs(2165) <= '0';
    layer1_outputs(2166) <= (layer0_outputs(4181)) and not (layer0_outputs(3456));
    layer1_outputs(2167) <= (layer0_outputs(245)) xor (layer0_outputs(5079));
    layer1_outputs(2168) <= layer0_outputs(1142);
    layer1_outputs(2169) <= (layer0_outputs(3629)) and not (layer0_outputs(495));
    layer1_outputs(2170) <= (layer0_outputs(2758)) and (layer0_outputs(1762));
    layer1_outputs(2171) <= (layer0_outputs(1015)) and not (layer0_outputs(3070));
    layer1_outputs(2172) <= '0';
    layer1_outputs(2173) <= not(layer0_outputs(268));
    layer1_outputs(2174) <= not(layer0_outputs(1359));
    layer1_outputs(2175) <= not(layer0_outputs(4403));
    layer1_outputs(2176) <= not(layer0_outputs(3629)) or (layer0_outputs(1077));
    layer1_outputs(2177) <= layer0_outputs(903);
    layer1_outputs(2178) <= not(layer0_outputs(257));
    layer1_outputs(2179) <= (layer0_outputs(1589)) and not (layer0_outputs(311));
    layer1_outputs(2180) <= '0';
    layer1_outputs(2181) <= not((layer0_outputs(1012)) or (layer0_outputs(3733)));
    layer1_outputs(2182) <= (layer0_outputs(1745)) and not (layer0_outputs(3285));
    layer1_outputs(2183) <= (layer0_outputs(5002)) and not (layer0_outputs(1839));
    layer1_outputs(2184) <= layer0_outputs(3472);
    layer1_outputs(2185) <= not(layer0_outputs(5043));
    layer1_outputs(2186) <= not(layer0_outputs(856)) or (layer0_outputs(247));
    layer1_outputs(2187) <= not(layer0_outputs(502)) or (layer0_outputs(4902));
    layer1_outputs(2188) <= (layer0_outputs(1200)) and (layer0_outputs(199));
    layer1_outputs(2189) <= not(layer0_outputs(4176));
    layer1_outputs(2190) <= (layer0_outputs(1017)) and not (layer0_outputs(1329));
    layer1_outputs(2191) <= (layer0_outputs(3671)) and not (layer0_outputs(2671));
    layer1_outputs(2192) <= not(layer0_outputs(3442));
    layer1_outputs(2193) <= not(layer0_outputs(2211));
    layer1_outputs(2194) <= layer0_outputs(2519);
    layer1_outputs(2195) <= layer0_outputs(1560);
    layer1_outputs(2196) <= not(layer0_outputs(4311)) or (layer0_outputs(4275));
    layer1_outputs(2197) <= not((layer0_outputs(2578)) and (layer0_outputs(3414)));
    layer1_outputs(2198) <= not((layer0_outputs(192)) or (layer0_outputs(4616)));
    layer1_outputs(2199) <= '1';
    layer1_outputs(2200) <= (layer0_outputs(3367)) and not (layer0_outputs(2075));
    layer1_outputs(2201) <= not(layer0_outputs(795)) or (layer0_outputs(4478));
    layer1_outputs(2202) <= not(layer0_outputs(251));
    layer1_outputs(2203) <= not(layer0_outputs(2284)) or (layer0_outputs(2845));
    layer1_outputs(2204) <= not(layer0_outputs(3211));
    layer1_outputs(2205) <= (layer0_outputs(616)) and not (layer0_outputs(3272));
    layer1_outputs(2206) <= not(layer0_outputs(1666));
    layer1_outputs(2207) <= not(layer0_outputs(4768));
    layer1_outputs(2208) <= (layer0_outputs(1923)) and not (layer0_outputs(402));
    layer1_outputs(2209) <= not(layer0_outputs(608));
    layer1_outputs(2210) <= layer0_outputs(3640);
    layer1_outputs(2211) <= layer0_outputs(4967);
    layer1_outputs(2212) <= not(layer0_outputs(5065));
    layer1_outputs(2213) <= (layer0_outputs(4530)) and not (layer0_outputs(681));
    layer1_outputs(2214) <= not((layer0_outputs(2104)) and (layer0_outputs(2758)));
    layer1_outputs(2215) <= not(layer0_outputs(280)) or (layer0_outputs(493));
    layer1_outputs(2216) <= not(layer0_outputs(1801));
    layer1_outputs(2217) <= (layer0_outputs(1161)) and (layer0_outputs(3747));
    layer1_outputs(2218) <= (layer0_outputs(2189)) and (layer0_outputs(1093));
    layer1_outputs(2219) <= not((layer0_outputs(3940)) and (layer0_outputs(4456)));
    layer1_outputs(2220) <= '0';
    layer1_outputs(2221) <= layer0_outputs(4193);
    layer1_outputs(2222) <= (layer0_outputs(1380)) and (layer0_outputs(2877));
    layer1_outputs(2223) <= not(layer0_outputs(475));
    layer1_outputs(2224) <= not(layer0_outputs(3589));
    layer1_outputs(2225) <= (layer0_outputs(2390)) and (layer0_outputs(1984));
    layer1_outputs(2226) <= (layer0_outputs(3894)) or (layer0_outputs(3664));
    layer1_outputs(2227) <= not(layer0_outputs(1854)) or (layer0_outputs(4162));
    layer1_outputs(2228) <= not((layer0_outputs(4877)) or (layer0_outputs(3080)));
    layer1_outputs(2229) <= (layer0_outputs(1622)) and not (layer0_outputs(3140));
    layer1_outputs(2230) <= layer0_outputs(2282);
    layer1_outputs(2231) <= (layer0_outputs(3254)) and (layer0_outputs(4099));
    layer1_outputs(2232) <= layer0_outputs(4361);
    layer1_outputs(2233) <= not((layer0_outputs(568)) xor (layer0_outputs(1755)));
    layer1_outputs(2234) <= (layer0_outputs(1198)) xor (layer0_outputs(1147));
    layer1_outputs(2235) <= not(layer0_outputs(2048));
    layer1_outputs(2236) <= not(layer0_outputs(3374)) or (layer0_outputs(2387));
    layer1_outputs(2237) <= not(layer0_outputs(593));
    layer1_outputs(2238) <= layer0_outputs(4178);
    layer1_outputs(2239) <= not((layer0_outputs(3228)) or (layer0_outputs(3271)));
    layer1_outputs(2240) <= (layer0_outputs(1394)) and not (layer0_outputs(201));
    layer1_outputs(2241) <= not(layer0_outputs(3516));
    layer1_outputs(2242) <= not((layer0_outputs(3461)) or (layer0_outputs(4344)));
    layer1_outputs(2243) <= layer0_outputs(1213);
    layer1_outputs(2244) <= not(layer0_outputs(1035)) or (layer0_outputs(3529));
    layer1_outputs(2245) <= layer0_outputs(1655);
    layer1_outputs(2246) <= (layer0_outputs(472)) and (layer0_outputs(2151));
    layer1_outputs(2247) <= not(layer0_outputs(4102));
    layer1_outputs(2248) <= not(layer0_outputs(1321)) or (layer0_outputs(4671));
    layer1_outputs(2249) <= layer0_outputs(3748);
    layer1_outputs(2250) <= not(layer0_outputs(2205)) or (layer0_outputs(435));
    layer1_outputs(2251) <= not((layer0_outputs(518)) xor (layer0_outputs(1247)));
    layer1_outputs(2252) <= (layer0_outputs(3233)) or (layer0_outputs(2889));
    layer1_outputs(2253) <= not(layer0_outputs(3358)) or (layer0_outputs(2913));
    layer1_outputs(2254) <= (layer0_outputs(3073)) and (layer0_outputs(3730));
    layer1_outputs(2255) <= (layer0_outputs(3045)) and not (layer0_outputs(613));
    layer1_outputs(2256) <= not((layer0_outputs(3084)) or (layer0_outputs(3626)));
    layer1_outputs(2257) <= not(layer0_outputs(531));
    layer1_outputs(2258) <= not((layer0_outputs(3713)) and (layer0_outputs(3912)));
    layer1_outputs(2259) <= layer0_outputs(2773);
    layer1_outputs(2260) <= not((layer0_outputs(1804)) and (layer0_outputs(157)));
    layer1_outputs(2261) <= layer0_outputs(259);
    layer1_outputs(2262) <= not(layer0_outputs(4850)) or (layer0_outputs(4186));
    layer1_outputs(2263) <= (layer0_outputs(2336)) and (layer0_outputs(685));
    layer1_outputs(2264) <= '1';
    layer1_outputs(2265) <= (layer0_outputs(3896)) or (layer0_outputs(4864));
    layer1_outputs(2266) <= not(layer0_outputs(4082)) or (layer0_outputs(1907));
    layer1_outputs(2267) <= not(layer0_outputs(2421));
    layer1_outputs(2268) <= not(layer0_outputs(4807)) or (layer0_outputs(2725));
    layer1_outputs(2269) <= '0';
    layer1_outputs(2270) <= layer0_outputs(3681);
    layer1_outputs(2271) <= not(layer0_outputs(1543));
    layer1_outputs(2272) <= (layer0_outputs(561)) or (layer0_outputs(2145));
    layer1_outputs(2273) <= layer0_outputs(1557);
    layer1_outputs(2274) <= not(layer0_outputs(0)) or (layer0_outputs(4035));
    layer1_outputs(2275) <= (layer0_outputs(2504)) and (layer0_outputs(3953));
    layer1_outputs(2276) <= layer0_outputs(1644);
    layer1_outputs(2277) <= (layer0_outputs(4850)) or (layer0_outputs(4651));
    layer1_outputs(2278) <= not((layer0_outputs(4527)) or (layer0_outputs(3841)));
    layer1_outputs(2279) <= '0';
    layer1_outputs(2280) <= layer0_outputs(3284);
    layer1_outputs(2281) <= '0';
    layer1_outputs(2282) <= (layer0_outputs(600)) xor (layer0_outputs(4467));
    layer1_outputs(2283) <= not(layer0_outputs(2735)) or (layer0_outputs(3844));
    layer1_outputs(2284) <= not((layer0_outputs(5052)) xor (layer0_outputs(1)));
    layer1_outputs(2285) <= (layer0_outputs(4548)) or (layer0_outputs(305));
    layer1_outputs(2286) <= (layer0_outputs(3380)) and (layer0_outputs(1349));
    layer1_outputs(2287) <= layer0_outputs(1325);
    layer1_outputs(2288) <= not(layer0_outputs(2936)) or (layer0_outputs(3526));
    layer1_outputs(2289) <= layer0_outputs(2544);
    layer1_outputs(2290) <= not(layer0_outputs(3191));
    layer1_outputs(2291) <= (layer0_outputs(598)) and (layer0_outputs(2003));
    layer1_outputs(2292) <= not(layer0_outputs(4465)) or (layer0_outputs(3917));
    layer1_outputs(2293) <= not(layer0_outputs(2972));
    layer1_outputs(2294) <= not(layer0_outputs(1252));
    layer1_outputs(2295) <= not((layer0_outputs(1416)) xor (layer0_outputs(3914)));
    layer1_outputs(2296) <= '0';
    layer1_outputs(2297) <= (layer0_outputs(2435)) and (layer0_outputs(2808));
    layer1_outputs(2298) <= not(layer0_outputs(705));
    layer1_outputs(2299) <= (layer0_outputs(1899)) xor (layer0_outputs(2689));
    layer1_outputs(2300) <= layer0_outputs(3219);
    layer1_outputs(2301) <= not(layer0_outputs(3106)) or (layer0_outputs(244));
    layer1_outputs(2302) <= not((layer0_outputs(3265)) xor (layer0_outputs(2453)));
    layer1_outputs(2303) <= (layer0_outputs(1061)) and (layer0_outputs(4413));
    layer1_outputs(2304) <= not(layer0_outputs(2523)) or (layer0_outputs(3053));
    layer1_outputs(2305) <= not((layer0_outputs(595)) and (layer0_outputs(1934)));
    layer1_outputs(2306) <= not(layer0_outputs(7));
    layer1_outputs(2307) <= (layer0_outputs(1747)) and not (layer0_outputs(1712));
    layer1_outputs(2308) <= not(layer0_outputs(3737));
    layer1_outputs(2309) <= not((layer0_outputs(2883)) or (layer0_outputs(2166)));
    layer1_outputs(2310) <= not(layer0_outputs(169));
    layer1_outputs(2311) <= not((layer0_outputs(647)) and (layer0_outputs(1498)));
    layer1_outputs(2312) <= layer0_outputs(4093);
    layer1_outputs(2313) <= not(layer0_outputs(1089));
    layer1_outputs(2314) <= layer0_outputs(497);
    layer1_outputs(2315) <= layer0_outputs(4451);
    layer1_outputs(2316) <= (layer0_outputs(1452)) and (layer0_outputs(2819));
    layer1_outputs(2317) <= not(layer0_outputs(2685));
    layer1_outputs(2318) <= layer0_outputs(1167);
    layer1_outputs(2319) <= layer0_outputs(835);
    layer1_outputs(2320) <= not(layer0_outputs(1637));
    layer1_outputs(2321) <= not((layer0_outputs(3226)) or (layer0_outputs(407)));
    layer1_outputs(2322) <= not(layer0_outputs(5071)) or (layer0_outputs(3022));
    layer1_outputs(2323) <= layer0_outputs(2165);
    layer1_outputs(2324) <= (layer0_outputs(3688)) or (layer0_outputs(3806));
    layer1_outputs(2325) <= (layer0_outputs(4135)) and (layer0_outputs(3057));
    layer1_outputs(2326) <= not(layer0_outputs(4693));
    layer1_outputs(2327) <= not((layer0_outputs(4148)) or (layer0_outputs(953)));
    layer1_outputs(2328) <= (layer0_outputs(3753)) and not (layer0_outputs(2003));
    layer1_outputs(2329) <= not((layer0_outputs(3263)) and (layer0_outputs(4427)));
    layer1_outputs(2330) <= not(layer0_outputs(1156));
    layer1_outputs(2331) <= '1';
    layer1_outputs(2332) <= not(layer0_outputs(4206)) or (layer0_outputs(3409));
    layer1_outputs(2333) <= (layer0_outputs(2564)) and not (layer0_outputs(5034));
    layer1_outputs(2334) <= layer0_outputs(2320);
    layer1_outputs(2335) <= layer0_outputs(4694);
    layer1_outputs(2336) <= '1';
    layer1_outputs(2337) <= (layer0_outputs(3238)) and not (layer0_outputs(4045));
    layer1_outputs(2338) <= not(layer0_outputs(2847));
    layer1_outputs(2339) <= not(layer0_outputs(3312)) or (layer0_outputs(813));
    layer1_outputs(2340) <= not((layer0_outputs(587)) xor (layer0_outputs(2916)));
    layer1_outputs(2341) <= not(layer0_outputs(714)) or (layer0_outputs(1461));
    layer1_outputs(2342) <= layer0_outputs(4579);
    layer1_outputs(2343) <= not((layer0_outputs(2445)) and (layer0_outputs(2101)));
    layer1_outputs(2344) <= (layer0_outputs(3307)) or (layer0_outputs(4460));
    layer1_outputs(2345) <= not(layer0_outputs(1795)) or (layer0_outputs(3078));
    layer1_outputs(2346) <= not((layer0_outputs(205)) or (layer0_outputs(479)));
    layer1_outputs(2347) <= layer0_outputs(1964);
    layer1_outputs(2348) <= not(layer0_outputs(431));
    layer1_outputs(2349) <= not(layer0_outputs(2252));
    layer1_outputs(2350) <= '0';
    layer1_outputs(2351) <= not(layer0_outputs(1711));
    layer1_outputs(2352) <= not(layer0_outputs(2632));
    layer1_outputs(2353) <= not(layer0_outputs(3828));
    layer1_outputs(2354) <= layer0_outputs(5087);
    layer1_outputs(2355) <= not((layer0_outputs(2363)) xor (layer0_outputs(3379)));
    layer1_outputs(2356) <= not((layer0_outputs(1746)) and (layer0_outputs(389)));
    layer1_outputs(2357) <= not((layer0_outputs(468)) or (layer0_outputs(1178)));
    layer1_outputs(2358) <= not(layer0_outputs(4486));
    layer1_outputs(2359) <= layer0_outputs(4883);
    layer1_outputs(2360) <= layer0_outputs(2766);
    layer1_outputs(2361) <= (layer0_outputs(3161)) and not (layer0_outputs(4185));
    layer1_outputs(2362) <= not(layer0_outputs(2977));
    layer1_outputs(2363) <= (layer0_outputs(3749)) or (layer0_outputs(3365));
    layer1_outputs(2364) <= not((layer0_outputs(1608)) and (layer0_outputs(4334)));
    layer1_outputs(2365) <= not(layer0_outputs(4737));
    layer1_outputs(2366) <= '1';
    layer1_outputs(2367) <= not(layer0_outputs(4308)) or (layer0_outputs(421));
    layer1_outputs(2368) <= not(layer0_outputs(1293));
    layer1_outputs(2369) <= (layer0_outputs(3235)) or (layer0_outputs(249));
    layer1_outputs(2370) <= layer0_outputs(2834);
    layer1_outputs(2371) <= not((layer0_outputs(2298)) or (layer0_outputs(4284)));
    layer1_outputs(2372) <= not(layer0_outputs(3213));
    layer1_outputs(2373) <= not(layer0_outputs(1275));
    layer1_outputs(2374) <= (layer0_outputs(2850)) and not (layer0_outputs(145));
    layer1_outputs(2375) <= (layer0_outputs(283)) or (layer0_outputs(2411));
    layer1_outputs(2376) <= layer0_outputs(2344);
    layer1_outputs(2377) <= not(layer0_outputs(4557));
    layer1_outputs(2378) <= layer0_outputs(1554);
    layer1_outputs(2379) <= (layer0_outputs(2521)) and not (layer0_outputs(934));
    layer1_outputs(2380) <= (layer0_outputs(4692)) xor (layer0_outputs(143));
    layer1_outputs(2381) <= not(layer0_outputs(3497));
    layer1_outputs(2382) <= '1';
    layer1_outputs(2383) <= (layer0_outputs(4233)) and (layer0_outputs(2810));
    layer1_outputs(2384) <= (layer0_outputs(4825)) and not (layer0_outputs(1549));
    layer1_outputs(2385) <= layer0_outputs(1763);
    layer1_outputs(2386) <= not((layer0_outputs(4374)) or (layer0_outputs(4183)));
    layer1_outputs(2387) <= not((layer0_outputs(3546)) or (layer0_outputs(277)));
    layer1_outputs(2388) <= layer0_outputs(3074);
    layer1_outputs(2389) <= not((layer0_outputs(2190)) xor (layer0_outputs(4632)));
    layer1_outputs(2390) <= not(layer0_outputs(1750));
    layer1_outputs(2391) <= layer0_outputs(2572);
    layer1_outputs(2392) <= (layer0_outputs(1859)) xor (layer0_outputs(860));
    layer1_outputs(2393) <= not((layer0_outputs(2932)) and (layer0_outputs(636)));
    layer1_outputs(2394) <= layer0_outputs(3564);
    layer1_outputs(2395) <= not((layer0_outputs(4388)) or (layer0_outputs(4440)));
    layer1_outputs(2396) <= not((layer0_outputs(320)) or (layer0_outputs(2043)));
    layer1_outputs(2397) <= not(layer0_outputs(2136)) or (layer0_outputs(821));
    layer1_outputs(2398) <= layer0_outputs(1976);
    layer1_outputs(2399) <= not(layer0_outputs(4205));
    layer1_outputs(2400) <= not((layer0_outputs(5069)) xor (layer0_outputs(2359)));
    layer1_outputs(2401) <= not((layer0_outputs(2541)) and (layer0_outputs(946)));
    layer1_outputs(2402) <= (layer0_outputs(4609)) and not (layer0_outputs(3021));
    layer1_outputs(2403) <= (layer0_outputs(779)) and not (layer0_outputs(4622));
    layer1_outputs(2404) <= not((layer0_outputs(3608)) and (layer0_outputs(4471)));
    layer1_outputs(2405) <= (layer0_outputs(4729)) or (layer0_outputs(2238));
    layer1_outputs(2406) <= not(layer0_outputs(3352));
    layer1_outputs(2407) <= (layer0_outputs(4358)) and not (layer0_outputs(5112));
    layer1_outputs(2408) <= '1';
    layer1_outputs(2409) <= (layer0_outputs(5000)) and (layer0_outputs(4167));
    layer1_outputs(2410) <= not(layer0_outputs(2759));
    layer1_outputs(2411) <= layer0_outputs(1097);
    layer1_outputs(2412) <= '1';
    layer1_outputs(2413) <= (layer0_outputs(2160)) and not (layer0_outputs(4914));
    layer1_outputs(2414) <= not(layer0_outputs(306));
    layer1_outputs(2415) <= layer0_outputs(4999);
    layer1_outputs(2416) <= not(layer0_outputs(1602)) or (layer0_outputs(896));
    layer1_outputs(2417) <= not(layer0_outputs(1541)) or (layer0_outputs(3834));
    layer1_outputs(2418) <= (layer0_outputs(4556)) or (layer0_outputs(1886));
    layer1_outputs(2419) <= (layer0_outputs(4801)) and not (layer0_outputs(4555));
    layer1_outputs(2420) <= layer0_outputs(3729);
    layer1_outputs(2421) <= '1';
    layer1_outputs(2422) <= not((layer0_outputs(4965)) xor (layer0_outputs(1748)));
    layer1_outputs(2423) <= not(layer0_outputs(3014)) or (layer0_outputs(3632));
    layer1_outputs(2424) <= not(layer0_outputs(2233)) or (layer0_outputs(3958));
    layer1_outputs(2425) <= not(layer0_outputs(1351));
    layer1_outputs(2426) <= not(layer0_outputs(3430)) or (layer0_outputs(3334));
    layer1_outputs(2427) <= not(layer0_outputs(3175));
    layer1_outputs(2428) <= (layer0_outputs(4227)) and not (layer0_outputs(2997));
    layer1_outputs(2429) <= layer0_outputs(3079);
    layer1_outputs(2430) <= layer0_outputs(3203);
    layer1_outputs(2431) <= (layer0_outputs(3342)) or (layer0_outputs(3700));
    layer1_outputs(2432) <= '0';
    layer1_outputs(2433) <= layer0_outputs(3476);
    layer1_outputs(2434) <= not(layer0_outputs(2519)) or (layer0_outputs(3187));
    layer1_outputs(2435) <= not((layer0_outputs(2993)) or (layer0_outputs(1327)));
    layer1_outputs(2436) <= (layer0_outputs(512)) and (layer0_outputs(2981));
    layer1_outputs(2437) <= (layer0_outputs(352)) and not (layer0_outputs(2651));
    layer1_outputs(2438) <= not((layer0_outputs(4822)) and (layer0_outputs(1013)));
    layer1_outputs(2439) <= not(layer0_outputs(1409)) or (layer0_outputs(4675));
    layer1_outputs(2440) <= not(layer0_outputs(3558));
    layer1_outputs(2441) <= '1';
    layer1_outputs(2442) <= not(layer0_outputs(1532));
    layer1_outputs(2443) <= '0';
    layer1_outputs(2444) <= layer0_outputs(3913);
    layer1_outputs(2445) <= not(layer0_outputs(1495)) or (layer0_outputs(4258));
    layer1_outputs(2446) <= (layer0_outputs(3511)) and (layer0_outputs(1138));
    layer1_outputs(2447) <= (layer0_outputs(4263)) and not (layer0_outputs(155));
    layer1_outputs(2448) <= not((layer0_outputs(4263)) and (layer0_outputs(2492)));
    layer1_outputs(2449) <= layer0_outputs(2358);
    layer1_outputs(2450) <= layer0_outputs(2848);
    layer1_outputs(2451) <= (layer0_outputs(2741)) and not (layer0_outputs(2566));
    layer1_outputs(2452) <= (layer0_outputs(3075)) or (layer0_outputs(3770));
    layer1_outputs(2453) <= layer0_outputs(4221);
    layer1_outputs(2454) <= not((layer0_outputs(4037)) or (layer0_outputs(1842)));
    layer1_outputs(2455) <= (layer0_outputs(1947)) and not (layer0_outputs(4679));
    layer1_outputs(2456) <= (layer0_outputs(1929)) or (layer0_outputs(3887));
    layer1_outputs(2457) <= (layer0_outputs(2931)) and not (layer0_outputs(4480));
    layer1_outputs(2458) <= layer0_outputs(5084);
    layer1_outputs(2459) <= layer0_outputs(61);
    layer1_outputs(2460) <= not((layer0_outputs(4733)) and (layer0_outputs(4079)));
    layer1_outputs(2461) <= layer0_outputs(1265);
    layer1_outputs(2462) <= not(layer0_outputs(3738)) or (layer0_outputs(3562));
    layer1_outputs(2463) <= not(layer0_outputs(4636));
    layer1_outputs(2464) <= not((layer0_outputs(947)) or (layer0_outputs(1323)));
    layer1_outputs(2465) <= not(layer0_outputs(576));
    layer1_outputs(2466) <= not((layer0_outputs(2252)) or (layer0_outputs(3755)));
    layer1_outputs(2467) <= layer0_outputs(3889);
    layer1_outputs(2468) <= (layer0_outputs(4326)) and (layer0_outputs(3398));
    layer1_outputs(2469) <= not((layer0_outputs(1674)) and (layer0_outputs(919)));
    layer1_outputs(2470) <= layer0_outputs(792);
    layer1_outputs(2471) <= not(layer0_outputs(4715));
    layer1_outputs(2472) <= layer0_outputs(3614);
    layer1_outputs(2473) <= (layer0_outputs(1279)) or (layer0_outputs(506));
    layer1_outputs(2474) <= not(layer0_outputs(2896)) or (layer0_outputs(4888));
    layer1_outputs(2475) <= not(layer0_outputs(1326)) or (layer0_outputs(3722));
    layer1_outputs(2476) <= not(layer0_outputs(1444));
    layer1_outputs(2477) <= not(layer0_outputs(2401));
    layer1_outputs(2478) <= (layer0_outputs(1747)) or (layer0_outputs(4395));
    layer1_outputs(2479) <= '1';
    layer1_outputs(2480) <= not(layer0_outputs(2200)) or (layer0_outputs(3810));
    layer1_outputs(2481) <= '0';
    layer1_outputs(2482) <= not((layer0_outputs(1245)) and (layer0_outputs(4362)));
    layer1_outputs(2483) <= layer0_outputs(2559);
    layer1_outputs(2484) <= not(layer0_outputs(2770)) or (layer0_outputs(4181));
    layer1_outputs(2485) <= not((layer0_outputs(1619)) and (layer0_outputs(3791)));
    layer1_outputs(2486) <= not(layer0_outputs(638)) or (layer0_outputs(4818));
    layer1_outputs(2487) <= layer0_outputs(3511);
    layer1_outputs(2488) <= not((layer0_outputs(4014)) and (layer0_outputs(25)));
    layer1_outputs(2489) <= layer0_outputs(476);
    layer1_outputs(2490) <= (layer0_outputs(1601)) and not (layer0_outputs(2646));
    layer1_outputs(2491) <= layer0_outputs(3695);
    layer1_outputs(2492) <= '1';
    layer1_outputs(2493) <= layer0_outputs(1576);
    layer1_outputs(2494) <= not((layer0_outputs(451)) or (layer0_outputs(2382)));
    layer1_outputs(2495) <= not((layer0_outputs(4932)) and (layer0_outputs(446)));
    layer1_outputs(2496) <= '0';
    layer1_outputs(2497) <= '1';
    layer1_outputs(2498) <= not((layer0_outputs(866)) xor (layer0_outputs(873)));
    layer1_outputs(2499) <= not(layer0_outputs(2613)) or (layer0_outputs(3039));
    layer1_outputs(2500) <= not(layer0_outputs(2246)) or (layer0_outputs(1725));
    layer1_outputs(2501) <= (layer0_outputs(1427)) or (layer0_outputs(2100));
    layer1_outputs(2502) <= layer0_outputs(4894);
    layer1_outputs(2503) <= not(layer0_outputs(2635)) or (layer0_outputs(4685));
    layer1_outputs(2504) <= (layer0_outputs(3323)) and not (layer0_outputs(3196));
    layer1_outputs(2505) <= layer0_outputs(2780);
    layer1_outputs(2506) <= not(layer0_outputs(2101));
    layer1_outputs(2507) <= (layer0_outputs(2611)) and not (layer0_outputs(961));
    layer1_outputs(2508) <= not(layer0_outputs(4011)) or (layer0_outputs(861));
    layer1_outputs(2509) <= (layer0_outputs(3720)) xor (layer0_outputs(654));
    layer1_outputs(2510) <= layer0_outputs(4051);
    layer1_outputs(2511) <= layer0_outputs(3170);
    layer1_outputs(2512) <= layer0_outputs(4364);
    layer1_outputs(2513) <= (layer0_outputs(323)) and (layer0_outputs(2204));
    layer1_outputs(2514) <= layer0_outputs(4365);
    layer1_outputs(2515) <= layer0_outputs(272);
    layer1_outputs(2516) <= (layer0_outputs(2311)) and not (layer0_outputs(1829));
    layer1_outputs(2517) <= (layer0_outputs(1173)) and not (layer0_outputs(1288));
    layer1_outputs(2518) <= not((layer0_outputs(478)) xor (layer0_outputs(4003)));
    layer1_outputs(2519) <= not((layer0_outputs(3779)) and (layer0_outputs(3399)));
    layer1_outputs(2520) <= layer0_outputs(611);
    layer1_outputs(2521) <= not((layer0_outputs(1471)) or (layer0_outputs(1697)));
    layer1_outputs(2522) <= '1';
    layer1_outputs(2523) <= not((layer0_outputs(957)) or (layer0_outputs(349)));
    layer1_outputs(2524) <= (layer0_outputs(950)) and not (layer0_outputs(4329));
    layer1_outputs(2525) <= (layer0_outputs(4165)) xor (layer0_outputs(2462));
    layer1_outputs(2526) <= not(layer0_outputs(4114));
    layer1_outputs(2527) <= '1';
    layer1_outputs(2528) <= not(layer0_outputs(2800)) or (layer0_outputs(3542));
    layer1_outputs(2529) <= not(layer0_outputs(3322)) or (layer0_outputs(3111));
    layer1_outputs(2530) <= not(layer0_outputs(1717)) or (layer0_outputs(4979));
    layer1_outputs(2531) <= layer0_outputs(4078);
    layer1_outputs(2532) <= not((layer0_outputs(332)) and (layer0_outputs(309)));
    layer1_outputs(2533) <= layer0_outputs(1529);
    layer1_outputs(2534) <= not((layer0_outputs(2149)) and (layer0_outputs(4401)));
    layer1_outputs(2535) <= (layer0_outputs(4184)) xor (layer0_outputs(783));
    layer1_outputs(2536) <= (layer0_outputs(2564)) and (layer0_outputs(573));
    layer1_outputs(2537) <= not(layer0_outputs(4684));
    layer1_outputs(2538) <= (layer0_outputs(3721)) and (layer0_outputs(4932));
    layer1_outputs(2539) <= not(layer0_outputs(2483));
    layer1_outputs(2540) <= not(layer0_outputs(803));
    layer1_outputs(2541) <= (layer0_outputs(853)) and (layer0_outputs(4433));
    layer1_outputs(2542) <= layer0_outputs(134);
    layer1_outputs(2543) <= not(layer0_outputs(290));
    layer1_outputs(2544) <= '0';
    layer1_outputs(2545) <= (layer0_outputs(1330)) and (layer0_outputs(4087));
    layer1_outputs(2546) <= (layer0_outputs(4666)) or (layer0_outputs(3637));
    layer1_outputs(2547) <= not((layer0_outputs(97)) xor (layer0_outputs(1513)));
    layer1_outputs(2548) <= (layer0_outputs(4487)) and not (layer0_outputs(2040));
    layer1_outputs(2549) <= not((layer0_outputs(4034)) or (layer0_outputs(1278)));
    layer1_outputs(2550) <= not(layer0_outputs(2947)) or (layer0_outputs(4522));
    layer1_outputs(2551) <= not((layer0_outputs(3123)) or (layer0_outputs(1197)));
    layer1_outputs(2552) <= not(layer0_outputs(3953)) or (layer0_outputs(4796));
    layer1_outputs(2553) <= not(layer0_outputs(4920)) or (layer0_outputs(1741));
    layer1_outputs(2554) <= not(layer0_outputs(4328));
    layer1_outputs(2555) <= '1';
    layer1_outputs(2556) <= not((layer0_outputs(2846)) or (layer0_outputs(4088)));
    layer1_outputs(2557) <= not((layer0_outputs(2851)) or (layer0_outputs(938)));
    layer1_outputs(2558) <= (layer0_outputs(894)) and (layer0_outputs(117));
    layer1_outputs(2559) <= not(layer0_outputs(3687));
    layer1_outputs(2560) <= layer0_outputs(2034);
    layer1_outputs(2561) <= not(layer0_outputs(1567));
    layer1_outputs(2562) <= (layer0_outputs(459)) and not (layer0_outputs(2349));
    layer1_outputs(2563) <= (layer0_outputs(2105)) or (layer0_outputs(1141));
    layer1_outputs(2564) <= (layer0_outputs(1137)) and not (layer0_outputs(274));
    layer1_outputs(2565) <= not(layer0_outputs(828));
    layer1_outputs(2566) <= '0';
    layer1_outputs(2567) <= layer0_outputs(261);
    layer1_outputs(2568) <= not(layer0_outputs(2304));
    layer1_outputs(2569) <= not((layer0_outputs(1454)) and (layer0_outputs(1430)));
    layer1_outputs(2570) <= not(layer0_outputs(916));
    layer1_outputs(2571) <= layer0_outputs(4880);
    layer1_outputs(2572) <= '0';
    layer1_outputs(2573) <= not((layer0_outputs(669)) and (layer0_outputs(1559)));
    layer1_outputs(2574) <= not(layer0_outputs(1609)) or (layer0_outputs(3102));
    layer1_outputs(2575) <= not((layer0_outputs(4975)) and (layer0_outputs(4518)));
    layer1_outputs(2576) <= not((layer0_outputs(2146)) xor (layer0_outputs(533)));
    layer1_outputs(2577) <= (layer0_outputs(4538)) or (layer0_outputs(1373));
    layer1_outputs(2578) <= (layer0_outputs(1011)) and not (layer0_outputs(2775));
    layer1_outputs(2579) <= '1';
    layer1_outputs(2580) <= not((layer0_outputs(4606)) and (layer0_outputs(1175)));
    layer1_outputs(2581) <= not(layer0_outputs(1203)) or (layer0_outputs(2459));
    layer1_outputs(2582) <= (layer0_outputs(756)) and (layer0_outputs(2184));
    layer1_outputs(2583) <= (layer0_outputs(3346)) xor (layer0_outputs(3947));
    layer1_outputs(2584) <= (layer0_outputs(3939)) or (layer0_outputs(4391));
    layer1_outputs(2585) <= not(layer0_outputs(2614));
    layer1_outputs(2586) <= not(layer0_outputs(1099));
    layer1_outputs(2587) <= (layer0_outputs(2272)) and not (layer0_outputs(2962));
    layer1_outputs(2588) <= (layer0_outputs(3782)) and (layer0_outputs(2084));
    layer1_outputs(2589) <= not((layer0_outputs(918)) or (layer0_outputs(2989)));
    layer1_outputs(2590) <= not((layer0_outputs(3869)) and (layer0_outputs(1295)));
    layer1_outputs(2591) <= not(layer0_outputs(2223));
    layer1_outputs(2592) <= not((layer0_outputs(3487)) or (layer0_outputs(2697)));
    layer1_outputs(2593) <= not(layer0_outputs(2227));
    layer1_outputs(2594) <= not((layer0_outputs(4926)) and (layer0_outputs(4419)));
    layer1_outputs(2595) <= layer0_outputs(3117);
    layer1_outputs(2596) <= (layer0_outputs(556)) or (layer0_outputs(105));
    layer1_outputs(2597) <= (layer0_outputs(380)) xor (layer0_outputs(94));
    layer1_outputs(2598) <= not(layer0_outputs(1678));
    layer1_outputs(2599) <= not(layer0_outputs(2394));
    layer1_outputs(2600) <= not((layer0_outputs(4201)) and (layer0_outputs(4130)));
    layer1_outputs(2601) <= not(layer0_outputs(47));
    layer1_outputs(2602) <= layer0_outputs(1171);
    layer1_outputs(2603) <= not(layer0_outputs(27));
    layer1_outputs(2604) <= (layer0_outputs(3764)) and not (layer0_outputs(740));
    layer1_outputs(2605) <= not(layer0_outputs(4782));
    layer1_outputs(2606) <= layer0_outputs(791);
    layer1_outputs(2607) <= not(layer0_outputs(3179));
    layer1_outputs(2608) <= not(layer0_outputs(2365));
    layer1_outputs(2609) <= not(layer0_outputs(4482));
    layer1_outputs(2610) <= not(layer0_outputs(3291)) or (layer0_outputs(4664));
    layer1_outputs(2611) <= not(layer0_outputs(3915));
    layer1_outputs(2612) <= not((layer0_outputs(3250)) or (layer0_outputs(4623)));
    layer1_outputs(2613) <= layer0_outputs(4030);
    layer1_outputs(2614) <= (layer0_outputs(2740)) and not (layer0_outputs(2831));
    layer1_outputs(2615) <= layer0_outputs(1752);
    layer1_outputs(2616) <= not(layer0_outputs(4527));
    layer1_outputs(2617) <= not(layer0_outputs(3763)) or (layer0_outputs(931));
    layer1_outputs(2618) <= not((layer0_outputs(5054)) and (layer0_outputs(2455)));
    layer1_outputs(2619) <= layer0_outputs(2038);
    layer1_outputs(2620) <= '1';
    layer1_outputs(2621) <= (layer0_outputs(2332)) and not (layer0_outputs(1660));
    layer1_outputs(2622) <= not(layer0_outputs(2542));
    layer1_outputs(2623) <= not(layer0_outputs(4768));
    layer1_outputs(2624) <= (layer0_outputs(4300)) and (layer0_outputs(1774));
    layer1_outputs(2625) <= not(layer0_outputs(1754)) or (layer0_outputs(2420));
    layer1_outputs(2626) <= layer0_outputs(4863);
    layer1_outputs(2627) <= not(layer0_outputs(3308)) or (layer0_outputs(1449));
    layer1_outputs(2628) <= not(layer0_outputs(716)) or (layer0_outputs(5021));
    layer1_outputs(2629) <= not(layer0_outputs(649));
    layer1_outputs(2630) <= (layer0_outputs(2102)) xor (layer0_outputs(4021));
    layer1_outputs(2631) <= '1';
    layer1_outputs(2632) <= not((layer0_outputs(3902)) or (layer0_outputs(3278)));
    layer1_outputs(2633) <= not(layer0_outputs(3865));
    layer1_outputs(2634) <= (layer0_outputs(1451)) and not (layer0_outputs(4583));
    layer1_outputs(2635) <= not(layer0_outputs(3077)) or (layer0_outputs(210));
    layer1_outputs(2636) <= (layer0_outputs(2398)) and (layer0_outputs(1738));
    layer1_outputs(2637) <= (layer0_outputs(1227)) xor (layer0_outputs(160));
    layer1_outputs(2638) <= not(layer0_outputs(4708));
    layer1_outputs(2639) <= not(layer0_outputs(2052));
    layer1_outputs(2640) <= not(layer0_outputs(2953)) or (layer0_outputs(1649));
    layer1_outputs(2641) <= not(layer0_outputs(4705)) or (layer0_outputs(3478));
    layer1_outputs(2642) <= (layer0_outputs(1464)) and not (layer0_outputs(1209));
    layer1_outputs(2643) <= '0';
    layer1_outputs(2644) <= (layer0_outputs(1751)) or (layer0_outputs(2749));
    layer1_outputs(2645) <= not(layer0_outputs(3097));
    layer1_outputs(2646) <= not(layer0_outputs(1905)) or (layer0_outputs(2788));
    layer1_outputs(2647) <= not(layer0_outputs(1713));
    layer1_outputs(2648) <= (layer0_outputs(5108)) and (layer0_outputs(1945));
    layer1_outputs(2649) <= not(layer0_outputs(900)) or (layer0_outputs(4995));
    layer1_outputs(2650) <= not((layer0_outputs(3333)) and (layer0_outputs(3215)));
    layer1_outputs(2651) <= layer0_outputs(1173);
    layer1_outputs(2652) <= layer0_outputs(4001);
    layer1_outputs(2653) <= '1';
    layer1_outputs(2654) <= layer0_outputs(1446);
    layer1_outputs(2655) <= layer0_outputs(1218);
    layer1_outputs(2656) <= (layer0_outputs(4788)) and not (layer0_outputs(2911));
    layer1_outputs(2657) <= not(layer0_outputs(3666)) or (layer0_outputs(778));
    layer1_outputs(2658) <= layer0_outputs(586);
    layer1_outputs(2659) <= not(layer0_outputs(4086));
    layer1_outputs(2660) <= not((layer0_outputs(1401)) and (layer0_outputs(4776)));
    layer1_outputs(2661) <= not(layer0_outputs(259));
    layer1_outputs(2662) <= '0';
    layer1_outputs(2663) <= not(layer0_outputs(3323)) or (layer0_outputs(5045));
    layer1_outputs(2664) <= not(layer0_outputs(1679));
    layer1_outputs(2665) <= not((layer0_outputs(4672)) or (layer0_outputs(725)));
    layer1_outputs(2666) <= not((layer0_outputs(4940)) xor (layer0_outputs(4989)));
    layer1_outputs(2667) <= not(layer0_outputs(665));
    layer1_outputs(2668) <= not(layer0_outputs(816)) or (layer0_outputs(4648));
    layer1_outputs(2669) <= layer0_outputs(4698);
    layer1_outputs(2670) <= not(layer0_outputs(2000));
    layer1_outputs(2671) <= not(layer0_outputs(1959)) or (layer0_outputs(2543));
    layer1_outputs(2672) <= not(layer0_outputs(1421)) or (layer0_outputs(1425));
    layer1_outputs(2673) <= not(layer0_outputs(907));
    layer1_outputs(2674) <= not((layer0_outputs(4554)) and (layer0_outputs(1567)));
    layer1_outputs(2675) <= layer0_outputs(3403);
    layer1_outputs(2676) <= (layer0_outputs(2014)) and not (layer0_outputs(3339));
    layer1_outputs(2677) <= (layer0_outputs(3893)) and not (layer0_outputs(5049));
    layer1_outputs(2678) <= layer0_outputs(3609);
    layer1_outputs(2679) <= not(layer0_outputs(318)) or (layer0_outputs(1266));
    layer1_outputs(2680) <= layer0_outputs(1242);
    layer1_outputs(2681) <= (layer0_outputs(1264)) and not (layer0_outputs(66));
    layer1_outputs(2682) <= (layer0_outputs(2658)) and (layer0_outputs(1572));
    layer1_outputs(2683) <= not(layer0_outputs(3048));
    layer1_outputs(2684) <= not(layer0_outputs(4597)) or (layer0_outputs(659));
    layer1_outputs(2685) <= (layer0_outputs(4120)) and (layer0_outputs(1210));
    layer1_outputs(2686) <= (layer0_outputs(460)) and not (layer0_outputs(2417));
    layer1_outputs(2687) <= layer0_outputs(1236);
    layer1_outputs(2688) <= not((layer0_outputs(4151)) or (layer0_outputs(118)));
    layer1_outputs(2689) <= '1';
    layer1_outputs(2690) <= (layer0_outputs(3801)) or (layer0_outputs(398));
    layer1_outputs(2691) <= not((layer0_outputs(4972)) or (layer0_outputs(2909)));
    layer1_outputs(2692) <= layer0_outputs(4159);
    layer1_outputs(2693) <= (layer0_outputs(3961)) and (layer0_outputs(3878));
    layer1_outputs(2694) <= (layer0_outputs(4428)) and not (layer0_outputs(3658));
    layer1_outputs(2695) <= not(layer0_outputs(4));
    layer1_outputs(2696) <= (layer0_outputs(1874)) or (layer0_outputs(1394));
    layer1_outputs(2697) <= (layer0_outputs(2953)) and not (layer0_outputs(5105));
    layer1_outputs(2698) <= (layer0_outputs(845)) and not (layer0_outputs(733));
    layer1_outputs(2699) <= not((layer0_outputs(337)) or (layer0_outputs(1059)));
    layer1_outputs(2700) <= (layer0_outputs(2627)) or (layer0_outputs(141));
    layer1_outputs(2701) <= not(layer0_outputs(4296));
    layer1_outputs(2702) <= (layer0_outputs(1198)) or (layer0_outputs(2346));
    layer1_outputs(2703) <= layer0_outputs(4119);
    layer1_outputs(2704) <= (layer0_outputs(33)) or (layer0_outputs(4484));
    layer1_outputs(2705) <= layer0_outputs(730);
    layer1_outputs(2706) <= not(layer0_outputs(3503));
    layer1_outputs(2707) <= not(layer0_outputs(1392));
    layer1_outputs(2708) <= layer0_outputs(3530);
    layer1_outputs(2709) <= (layer0_outputs(2198)) and not (layer0_outputs(2506));
    layer1_outputs(2710) <= not(layer0_outputs(2576));
    layer1_outputs(2711) <= (layer0_outputs(731)) and (layer0_outputs(2547));
    layer1_outputs(2712) <= not(layer0_outputs(1862));
    layer1_outputs(2713) <= layer0_outputs(2872);
    layer1_outputs(2714) <= layer0_outputs(4024);
    layer1_outputs(2715) <= not((layer0_outputs(869)) and (layer0_outputs(2958)));
    layer1_outputs(2716) <= (layer0_outputs(3172)) and not (layer0_outputs(2977));
    layer1_outputs(2717) <= not(layer0_outputs(2670));
    layer1_outputs(2718) <= not(layer0_outputs(3649)) or (layer0_outputs(3700));
    layer1_outputs(2719) <= not(layer0_outputs(1534)) or (layer0_outputs(827));
    layer1_outputs(2720) <= (layer0_outputs(2526)) xor (layer0_outputs(3219));
    layer1_outputs(2721) <= not((layer0_outputs(1487)) xor (layer0_outputs(2851)));
    layer1_outputs(2722) <= layer0_outputs(1842);
    layer1_outputs(2723) <= not(layer0_outputs(4104));
    layer1_outputs(2724) <= (layer0_outputs(3861)) and (layer0_outputs(950));
    layer1_outputs(2725) <= '1';
    layer1_outputs(2726) <= not(layer0_outputs(154)) or (layer0_outputs(4108));
    layer1_outputs(2727) <= not(layer0_outputs(1535));
    layer1_outputs(2728) <= (layer0_outputs(4996)) and (layer0_outputs(4409));
    layer1_outputs(2729) <= (layer0_outputs(2732)) or (layer0_outputs(159));
    layer1_outputs(2730) <= not((layer0_outputs(5017)) xor (layer0_outputs(1300)));
    layer1_outputs(2731) <= not((layer0_outputs(2329)) and (layer0_outputs(142)));
    layer1_outputs(2732) <= layer0_outputs(3504);
    layer1_outputs(2733) <= layer0_outputs(2400);
    layer1_outputs(2734) <= (layer0_outputs(3861)) and not (layer0_outputs(1556));
    layer1_outputs(2735) <= (layer0_outputs(3762)) and (layer0_outputs(77));
    layer1_outputs(2736) <= (layer0_outputs(1873)) or (layer0_outputs(2409));
    layer1_outputs(2737) <= not(layer0_outputs(3194)) or (layer0_outputs(4784));
    layer1_outputs(2738) <= not(layer0_outputs(4009));
    layer1_outputs(2739) <= layer0_outputs(4667);
    layer1_outputs(2740) <= layer0_outputs(2854);
    layer1_outputs(2741) <= (layer0_outputs(384)) and (layer0_outputs(395));
    layer1_outputs(2742) <= layer0_outputs(1900);
    layer1_outputs(2743) <= (layer0_outputs(3178)) and (layer0_outputs(4149));
    layer1_outputs(2744) <= layer0_outputs(5102);
    layer1_outputs(2745) <= layer0_outputs(2678);
    layer1_outputs(2746) <= not(layer0_outputs(476));
    layer1_outputs(2747) <= not((layer0_outputs(4481)) or (layer0_outputs(5004)));
    layer1_outputs(2748) <= not(layer0_outputs(3281));
    layer1_outputs(2749) <= layer0_outputs(4280);
    layer1_outputs(2750) <= not(layer0_outputs(2634)) or (layer0_outputs(2995));
    layer1_outputs(2751) <= (layer0_outputs(2993)) and not (layer0_outputs(170));
    layer1_outputs(2752) <= (layer0_outputs(4330)) xor (layer0_outputs(3840));
    layer1_outputs(2753) <= not((layer0_outputs(44)) or (layer0_outputs(521)));
    layer1_outputs(2754) <= layer0_outputs(5066);
    layer1_outputs(2755) <= '1';
    layer1_outputs(2756) <= (layer0_outputs(2961)) and not (layer0_outputs(2314));
    layer1_outputs(2757) <= '0';
    layer1_outputs(2758) <= layer0_outputs(3021);
    layer1_outputs(2759) <= not((layer0_outputs(2987)) xor (layer0_outputs(1943)));
    layer1_outputs(2760) <= not(layer0_outputs(515));
    layer1_outputs(2761) <= not(layer0_outputs(3100)) or (layer0_outputs(2625));
    layer1_outputs(2762) <= not(layer0_outputs(2138));
    layer1_outputs(2763) <= not(layer0_outputs(2563)) or (layer0_outputs(2931));
    layer1_outputs(2764) <= (layer0_outputs(256)) and (layer0_outputs(2222));
    layer1_outputs(2765) <= not((layer0_outputs(1395)) and (layer0_outputs(885)));
    layer1_outputs(2766) <= layer0_outputs(3942);
    layer1_outputs(2767) <= (layer0_outputs(1805)) and not (layer0_outputs(4245));
    layer1_outputs(2768) <= layer0_outputs(1942);
    layer1_outputs(2769) <= layer0_outputs(921);
    layer1_outputs(2770) <= not(layer0_outputs(4906));
    layer1_outputs(2771) <= (layer0_outputs(596)) and (layer0_outputs(3995));
    layer1_outputs(2772) <= layer0_outputs(5074);
    layer1_outputs(2773) <= '1';
    layer1_outputs(2774) <= '0';
    layer1_outputs(2775) <= not(layer0_outputs(649)) or (layer0_outputs(4161));
    layer1_outputs(2776) <= not((layer0_outputs(2484)) xor (layer0_outputs(1845)));
    layer1_outputs(2777) <= layer0_outputs(3644);
    layer1_outputs(2778) <= not(layer0_outputs(4398)) or (layer0_outputs(1222));
    layer1_outputs(2779) <= (layer0_outputs(4969)) and not (layer0_outputs(1815));
    layer1_outputs(2780) <= not(layer0_outputs(2513));
    layer1_outputs(2781) <= (layer0_outputs(4337)) and not (layer0_outputs(4994));
    layer1_outputs(2782) <= not(layer0_outputs(884));
    layer1_outputs(2783) <= not(layer0_outputs(4965));
    layer1_outputs(2784) <= not((layer0_outputs(1023)) and (layer0_outputs(3343)));
    layer1_outputs(2785) <= (layer0_outputs(1135)) or (layer0_outputs(1120));
    layer1_outputs(2786) <= (layer0_outputs(4859)) and (layer0_outputs(4662));
    layer1_outputs(2787) <= not(layer0_outputs(4619));
    layer1_outputs(2788) <= layer0_outputs(1221);
    layer1_outputs(2789) <= layer0_outputs(3959);
    layer1_outputs(2790) <= not(layer0_outputs(943)) or (layer0_outputs(3768));
    layer1_outputs(2791) <= not(layer0_outputs(4490));
    layer1_outputs(2792) <= not((layer0_outputs(1089)) and (layer0_outputs(2408)));
    layer1_outputs(2793) <= layer0_outputs(3465);
    layer1_outputs(2794) <= (layer0_outputs(363)) and not (layer0_outputs(1531));
    layer1_outputs(2795) <= (layer0_outputs(1391)) and not (layer0_outputs(2968));
    layer1_outputs(2796) <= not(layer0_outputs(5088)) or (layer0_outputs(2638));
    layer1_outputs(2797) <= (layer0_outputs(3216)) or (layer0_outputs(1720));
    layer1_outputs(2798) <= layer0_outputs(2114);
    layer1_outputs(2799) <= (layer0_outputs(972)) xor (layer0_outputs(977));
    layer1_outputs(2800) <= not(layer0_outputs(4650));
    layer1_outputs(2801) <= not(layer0_outputs(1005)) or (layer0_outputs(1282));
    layer1_outputs(2802) <= not(layer0_outputs(471));
    layer1_outputs(2803) <= not(layer0_outputs(4158));
    layer1_outputs(2804) <= not((layer0_outputs(3795)) and (layer0_outputs(3096)));
    layer1_outputs(2805) <= (layer0_outputs(4640)) and (layer0_outputs(2089));
    layer1_outputs(2806) <= not(layer0_outputs(3806));
    layer1_outputs(2807) <= (layer0_outputs(1769)) and (layer0_outputs(5002));
    layer1_outputs(2808) <= layer0_outputs(4009);
    layer1_outputs(2809) <= layer0_outputs(4832);
    layer1_outputs(2810) <= not(layer0_outputs(519));
    layer1_outputs(2811) <= layer0_outputs(1540);
    layer1_outputs(2812) <= not(layer0_outputs(4403));
    layer1_outputs(2813) <= (layer0_outputs(4332)) xor (layer0_outputs(262));
    layer1_outputs(2814) <= '0';
    layer1_outputs(2815) <= (layer0_outputs(5009)) or (layer0_outputs(172));
    layer1_outputs(2816) <= not((layer0_outputs(2934)) and (layer0_outputs(1592)));
    layer1_outputs(2817) <= (layer0_outputs(4117)) and not (layer0_outputs(2046));
    layer1_outputs(2818) <= layer0_outputs(1565);
    layer1_outputs(2819) <= (layer0_outputs(2878)) and (layer0_outputs(1095));
    layer1_outputs(2820) <= not(layer0_outputs(2413));
    layer1_outputs(2821) <= (layer0_outputs(976)) and (layer0_outputs(1132));
    layer1_outputs(2822) <= not((layer0_outputs(1220)) xor (layer0_outputs(686)));
    layer1_outputs(2823) <= (layer0_outputs(3127)) and (layer0_outputs(1290));
    layer1_outputs(2824) <= not(layer0_outputs(3936));
    layer1_outputs(2825) <= (layer0_outputs(3443)) and not (layer0_outputs(3362));
    layer1_outputs(2826) <= (layer0_outputs(4913)) and (layer0_outputs(1163));
    layer1_outputs(2827) <= not(layer0_outputs(4244)) or (layer0_outputs(4475));
    layer1_outputs(2828) <= layer0_outputs(3484);
    layer1_outputs(2829) <= not((layer0_outputs(3235)) and (layer0_outputs(3316)));
    layer1_outputs(2830) <= not((layer0_outputs(4638)) and (layer0_outputs(1790)));
    layer1_outputs(2831) <= not(layer0_outputs(983));
    layer1_outputs(2832) <= (layer0_outputs(2203)) and not (layer0_outputs(2596));
    layer1_outputs(2833) <= not(layer0_outputs(4099));
    layer1_outputs(2834) <= layer0_outputs(3611);
    layer1_outputs(2835) <= (layer0_outputs(2199)) and (layer0_outputs(2364));
    layer1_outputs(2836) <= (layer0_outputs(294)) and not (layer0_outputs(2936));
    layer1_outputs(2837) <= layer0_outputs(3897);
    layer1_outputs(2838) <= (layer0_outputs(3833)) and (layer0_outputs(4480));
    layer1_outputs(2839) <= (layer0_outputs(4865)) xor (layer0_outputs(2191));
    layer1_outputs(2840) <= layer0_outputs(4677);
    layer1_outputs(2841) <= not(layer0_outputs(4053));
    layer1_outputs(2842) <= not(layer0_outputs(4327));
    layer1_outputs(2843) <= (layer0_outputs(388)) and not (layer0_outputs(5085));
    layer1_outputs(2844) <= (layer0_outputs(4192)) or (layer0_outputs(2432));
    layer1_outputs(2845) <= (layer0_outputs(3169)) and (layer0_outputs(4253));
    layer1_outputs(2846) <= not((layer0_outputs(4982)) and (layer0_outputs(2285)));
    layer1_outputs(2847) <= '1';
    layer1_outputs(2848) <= layer0_outputs(1472);
    layer1_outputs(2849) <= not(layer0_outputs(1272)) or (layer0_outputs(499));
    layer1_outputs(2850) <= (layer0_outputs(567)) and not (layer0_outputs(4896));
    layer1_outputs(2851) <= '1';
    layer1_outputs(2852) <= not(layer0_outputs(2460)) or (layer0_outputs(4753));
    layer1_outputs(2853) <= (layer0_outputs(527)) and (layer0_outputs(2327));
    layer1_outputs(2854) <= not((layer0_outputs(968)) and (layer0_outputs(3661)));
    layer1_outputs(2855) <= not(layer0_outputs(4743));
    layer1_outputs(2856) <= (layer0_outputs(4966)) and not (layer0_outputs(93));
    layer1_outputs(2857) <= layer0_outputs(4735);
    layer1_outputs(2858) <= not(layer0_outputs(4232)) or (layer0_outputs(3319));
    layer1_outputs(2859) <= not(layer0_outputs(2774));
    layer1_outputs(2860) <= not(layer0_outputs(2517));
    layer1_outputs(2861) <= not(layer0_outputs(2393));
    layer1_outputs(2862) <= not(layer0_outputs(305)) or (layer0_outputs(2843));
    layer1_outputs(2863) <= layer0_outputs(4684);
    layer1_outputs(2864) <= layer0_outputs(1915);
    layer1_outputs(2865) <= '0';
    layer1_outputs(2866) <= (layer0_outputs(1483)) xor (layer0_outputs(3973));
    layer1_outputs(2867) <= not(layer0_outputs(59)) or (layer0_outputs(2436));
    layer1_outputs(2868) <= layer0_outputs(3037);
    layer1_outputs(2869) <= (layer0_outputs(3024)) and not (layer0_outputs(103));
    layer1_outputs(2870) <= not(layer0_outputs(1509));
    layer1_outputs(2871) <= (layer0_outputs(279)) and not (layer0_outputs(3426));
    layer1_outputs(2872) <= (layer0_outputs(3303)) xor (layer0_outputs(234));
    layer1_outputs(2873) <= not(layer0_outputs(3183));
    layer1_outputs(2874) <= not((layer0_outputs(4795)) and (layer0_outputs(4918)));
    layer1_outputs(2875) <= not((layer0_outputs(733)) or (layer0_outputs(4081)));
    layer1_outputs(2876) <= (layer0_outputs(2415)) and not (layer0_outputs(5096));
    layer1_outputs(2877) <= (layer0_outputs(2663)) and not (layer0_outputs(4052));
    layer1_outputs(2878) <= not(layer0_outputs(1962)) or (layer0_outputs(2095));
    layer1_outputs(2879) <= (layer0_outputs(1775)) and not (layer0_outputs(2202));
    layer1_outputs(2880) <= (layer0_outputs(5111)) and (layer0_outputs(2842));
    layer1_outputs(2881) <= '1';
    layer1_outputs(2882) <= not(layer0_outputs(4200));
    layer1_outputs(2883) <= layer0_outputs(3414);
    layer1_outputs(2884) <= layer0_outputs(2049);
    layer1_outputs(2885) <= not(layer0_outputs(3401));
    layer1_outputs(2886) <= layer0_outputs(2629);
    layer1_outputs(2887) <= layer0_outputs(2283);
    layer1_outputs(2888) <= (layer0_outputs(4280)) and (layer0_outputs(3573));
    layer1_outputs(2889) <= layer0_outputs(979);
    layer1_outputs(2890) <= not(layer0_outputs(4479));
    layer1_outputs(2891) <= not((layer0_outputs(1772)) and (layer0_outputs(4474)));
    layer1_outputs(2892) <= not(layer0_outputs(2329));
    layer1_outputs(2893) <= (layer0_outputs(2144)) xor (layer0_outputs(4863));
    layer1_outputs(2894) <= (layer0_outputs(2639)) and not (layer0_outputs(3451));
    layer1_outputs(2895) <= '1';
    layer1_outputs(2896) <= (layer0_outputs(1794)) or (layer0_outputs(3692));
    layer1_outputs(2897) <= layer0_outputs(4159);
    layer1_outputs(2898) <= (layer0_outputs(3993)) or (layer0_outputs(2140));
    layer1_outputs(2899) <= layer0_outputs(1114);
    layer1_outputs(2900) <= layer0_outputs(927);
    layer1_outputs(2901) <= not(layer0_outputs(4523));
    layer1_outputs(2902) <= not((layer0_outputs(1314)) and (layer0_outputs(4509)));
    layer1_outputs(2903) <= layer0_outputs(581);
    layer1_outputs(2904) <= not((layer0_outputs(4453)) xor (layer0_outputs(2694)));
    layer1_outputs(2905) <= '1';
    layer1_outputs(2906) <= not((layer0_outputs(48)) or (layer0_outputs(3243)));
    layer1_outputs(2907) <= (layer0_outputs(4661)) and (layer0_outputs(4470));
    layer1_outputs(2908) <= (layer0_outputs(2585)) and not (layer0_outputs(4254));
    layer1_outputs(2909) <= layer0_outputs(1466);
    layer1_outputs(2910) <= layer0_outputs(330);
    layer1_outputs(2911) <= (layer0_outputs(2516)) or (layer0_outputs(3687));
    layer1_outputs(2912) <= layer0_outputs(23);
    layer1_outputs(2913) <= '0';
    layer1_outputs(2914) <= not(layer0_outputs(75)) or (layer0_outputs(1881));
    layer1_outputs(2915) <= (layer0_outputs(1094)) or (layer0_outputs(3776));
    layer1_outputs(2916) <= (layer0_outputs(4485)) and not (layer0_outputs(4072));
    layer1_outputs(2917) <= layer0_outputs(1287);
    layer1_outputs(2918) <= not(layer0_outputs(764));
    layer1_outputs(2919) <= layer0_outputs(993);
    layer1_outputs(2920) <= '0';
    layer1_outputs(2921) <= not((layer0_outputs(3594)) and (layer0_outputs(1186)));
    layer1_outputs(2922) <= not(layer0_outputs(3552));
    layer1_outputs(2923) <= layer0_outputs(4695);
    layer1_outputs(2924) <= layer0_outputs(3374);
    layer1_outputs(2925) <= not(layer0_outputs(3185)) or (layer0_outputs(3552));
    layer1_outputs(2926) <= (layer0_outputs(1969)) and not (layer0_outputs(817));
    layer1_outputs(2927) <= layer0_outputs(1596);
    layer1_outputs(2928) <= (layer0_outputs(3954)) and (layer0_outputs(1299));
    layer1_outputs(2929) <= (layer0_outputs(4436)) and not (layer0_outputs(421));
    layer1_outputs(2930) <= not(layer0_outputs(2311)) or (layer0_outputs(422));
    layer1_outputs(2931) <= not(layer0_outputs(3254));
    layer1_outputs(2932) <= (layer0_outputs(439)) and (layer0_outputs(696));
    layer1_outputs(2933) <= not(layer0_outputs(1500));
    layer1_outputs(2934) <= (layer0_outputs(3252)) and not (layer0_outputs(4535));
    layer1_outputs(2935) <= '0';
    layer1_outputs(2936) <= layer0_outputs(1857);
    layer1_outputs(2937) <= (layer0_outputs(324)) and (layer0_outputs(948));
    layer1_outputs(2938) <= not(layer0_outputs(2368));
    layer1_outputs(2939) <= not((layer0_outputs(3538)) or (layer0_outputs(1656)));
    layer1_outputs(2940) <= (layer0_outputs(2322)) xor (layer0_outputs(4875));
    layer1_outputs(2941) <= not(layer0_outputs(1190)) or (layer0_outputs(1055));
    layer1_outputs(2942) <= (layer0_outputs(3355)) and not (layer0_outputs(4913));
    layer1_outputs(2943) <= layer0_outputs(2979);
    layer1_outputs(2944) <= not((layer0_outputs(1551)) and (layer0_outputs(1191)));
    layer1_outputs(2945) <= (layer0_outputs(2143)) xor (layer0_outputs(2117));
    layer1_outputs(2946) <= '0';
    layer1_outputs(2947) <= not(layer0_outputs(4139)) or (layer0_outputs(5080));
    layer1_outputs(2948) <= not((layer0_outputs(2825)) xor (layer0_outputs(2141)));
    layer1_outputs(2949) <= not(layer0_outputs(1485)) or (layer0_outputs(3396));
    layer1_outputs(2950) <= (layer0_outputs(1440)) and (layer0_outputs(4855));
    layer1_outputs(2951) <= layer0_outputs(2034);
    layer1_outputs(2952) <= not((layer0_outputs(4261)) or (layer0_outputs(4068)));
    layer1_outputs(2953) <= not(layer0_outputs(3686));
    layer1_outputs(2954) <= (layer0_outputs(1909)) and not (layer0_outputs(3174));
    layer1_outputs(2955) <= not(layer0_outputs(1612)) or (layer0_outputs(983));
    layer1_outputs(2956) <= not((layer0_outputs(3008)) or (layer0_outputs(2275)));
    layer1_outputs(2957) <= layer0_outputs(1122);
    layer1_outputs(2958) <= (layer0_outputs(915)) or (layer0_outputs(3975));
    layer1_outputs(2959) <= (layer0_outputs(1935)) and not (layer0_outputs(4947));
    layer1_outputs(2960) <= (layer0_outputs(1460)) and not (layer0_outputs(817));
    layer1_outputs(2961) <= not((layer0_outputs(2882)) or (layer0_outputs(3994)));
    layer1_outputs(2962) <= not(layer0_outputs(1848));
    layer1_outputs(2963) <= not((layer0_outputs(4047)) or (layer0_outputs(2086)));
    layer1_outputs(2964) <= not(layer0_outputs(260));
    layer1_outputs(2965) <= layer0_outputs(3027);
    layer1_outputs(2966) <= not((layer0_outputs(2922)) and (layer0_outputs(371)));
    layer1_outputs(2967) <= not(layer0_outputs(4092));
    layer1_outputs(2968) <= layer0_outputs(951);
    layer1_outputs(2969) <= (layer0_outputs(4168)) and not (layer0_outputs(4725));
    layer1_outputs(2970) <= layer0_outputs(2816);
    layer1_outputs(2971) <= not(layer0_outputs(4173));
    layer1_outputs(2972) <= not((layer0_outputs(224)) or (layer0_outputs(2744)));
    layer1_outputs(2973) <= (layer0_outputs(2935)) and not (layer0_outputs(2212));
    layer1_outputs(2974) <= not(layer0_outputs(4673)) or (layer0_outputs(83));
    layer1_outputs(2975) <= not(layer0_outputs(1574));
    layer1_outputs(2976) <= (layer0_outputs(59)) or (layer0_outputs(4166));
    layer1_outputs(2977) <= not(layer0_outputs(1033)) or (layer0_outputs(3052));
    layer1_outputs(2978) <= not(layer0_outputs(4581));
    layer1_outputs(2979) <= not(layer0_outputs(1008)) or (layer0_outputs(936));
    layer1_outputs(2980) <= not(layer0_outputs(1749));
    layer1_outputs(2981) <= (layer0_outputs(1393)) and not (layer0_outputs(4985));
    layer1_outputs(2982) <= not(layer0_outputs(572)) or (layer0_outputs(3259));
    layer1_outputs(2983) <= layer0_outputs(5073);
    layer1_outputs(2984) <= (layer0_outputs(2423)) and (layer0_outputs(3982));
    layer1_outputs(2985) <= not(layer0_outputs(4447));
    layer1_outputs(2986) <= not(layer0_outputs(3249));
    layer1_outputs(2987) <= not(layer0_outputs(2555)) or (layer0_outputs(293));
    layer1_outputs(2988) <= '1';
    layer1_outputs(2989) <= not(layer0_outputs(796));
    layer1_outputs(2990) <= (layer0_outputs(4393)) and not (layer0_outputs(2306));
    layer1_outputs(2991) <= (layer0_outputs(1187)) and (layer0_outputs(4677));
    layer1_outputs(2992) <= (layer0_outputs(329)) and not (layer0_outputs(1108));
    layer1_outputs(2993) <= layer0_outputs(786);
    layer1_outputs(2994) <= layer0_outputs(4963);
    layer1_outputs(2995) <= layer0_outputs(1744);
    layer1_outputs(2996) <= layer0_outputs(2491);
    layer1_outputs(2997) <= (layer0_outputs(2940)) and (layer0_outputs(641));
    layer1_outputs(2998) <= '0';
    layer1_outputs(2999) <= (layer0_outputs(265)) and not (layer0_outputs(3421));
    layer1_outputs(3000) <= not(layer0_outputs(2550));
    layer1_outputs(3001) <= (layer0_outputs(3313)) and (layer0_outputs(561));
    layer1_outputs(3002) <= layer0_outputs(377);
    layer1_outputs(3003) <= not((layer0_outputs(2270)) or (layer0_outputs(2033)));
    layer1_outputs(3004) <= not((layer0_outputs(2838)) or (layer0_outputs(2912)));
    layer1_outputs(3005) <= layer0_outputs(4699);
    layer1_outputs(3006) <= not(layer0_outputs(2032));
    layer1_outputs(3007) <= (layer0_outputs(3103)) xor (layer0_outputs(829));
    layer1_outputs(3008) <= not(layer0_outputs(4190));
    layer1_outputs(3009) <= not(layer0_outputs(2156)) or (layer0_outputs(4288));
    layer1_outputs(3010) <= not(layer0_outputs(865)) or (layer0_outputs(3872));
    layer1_outputs(3011) <= (layer0_outputs(4589)) or (layer0_outputs(4375));
    layer1_outputs(3012) <= not(layer0_outputs(3108)) or (layer0_outputs(2378));
    layer1_outputs(3013) <= not((layer0_outputs(1884)) and (layer0_outputs(1835)));
    layer1_outputs(3014) <= layer0_outputs(4902);
    layer1_outputs(3015) <= layer0_outputs(2757);
    layer1_outputs(3016) <= not(layer0_outputs(1502));
    layer1_outputs(3017) <= (layer0_outputs(3151)) and not (layer0_outputs(2211));
    layer1_outputs(3018) <= layer0_outputs(3360);
    layer1_outputs(3019) <= not(layer0_outputs(434)) or (layer0_outputs(4779));
    layer1_outputs(3020) <= not(layer0_outputs(3294));
    layer1_outputs(3021) <= layer0_outputs(3270);
    layer1_outputs(3022) <= layer0_outputs(3867);
    layer1_outputs(3023) <= layer0_outputs(4066);
    layer1_outputs(3024) <= not((layer0_outputs(2334)) and (layer0_outputs(1633)));
    layer1_outputs(3025) <= (layer0_outputs(2168)) and (layer0_outputs(2590));
    layer1_outputs(3026) <= '1';
    layer1_outputs(3027) <= (layer0_outputs(2383)) and (layer0_outputs(4409));
    layer1_outputs(3028) <= (layer0_outputs(119)) or (layer0_outputs(4491));
    layer1_outputs(3029) <= (layer0_outputs(3049)) and (layer0_outputs(3733));
    layer1_outputs(3030) <= '1';
    layer1_outputs(3031) <= not((layer0_outputs(4810)) or (layer0_outputs(3082)));
    layer1_outputs(3032) <= (layer0_outputs(2054)) and not (layer0_outputs(98));
    layer1_outputs(3033) <= not(layer0_outputs(3651)) or (layer0_outputs(1068));
    layer1_outputs(3034) <= layer0_outputs(202);
    layer1_outputs(3035) <= not((layer0_outputs(4466)) or (layer0_outputs(1816)));
    layer1_outputs(3036) <= not((layer0_outputs(1743)) or (layer0_outputs(2797)));
    layer1_outputs(3037) <= not((layer0_outputs(2950)) xor (layer0_outputs(4645)));
    layer1_outputs(3038) <= not(layer0_outputs(3321)) or (layer0_outputs(611));
    layer1_outputs(3039) <= not(layer0_outputs(90)) or (layer0_outputs(4882));
    layer1_outputs(3040) <= not((layer0_outputs(242)) or (layer0_outputs(4546)));
    layer1_outputs(3041) <= layer0_outputs(1146);
    layer1_outputs(3042) <= not((layer0_outputs(4446)) or (layer0_outputs(3238)));
    layer1_outputs(3043) <= not(layer0_outputs(5065));
    layer1_outputs(3044) <= '0';
    layer1_outputs(3045) <= (layer0_outputs(4424)) or (layer0_outputs(3833));
    layer1_outputs(3046) <= layer0_outputs(3491);
    layer1_outputs(3047) <= (layer0_outputs(4367)) and (layer0_outputs(1672));
    layer1_outputs(3048) <= not(layer0_outputs(5055));
    layer1_outputs(3049) <= '1';
    layer1_outputs(3050) <= (layer0_outputs(3242)) or (layer0_outputs(3326));
    layer1_outputs(3051) <= not((layer0_outputs(1335)) xor (layer0_outputs(762)));
    layer1_outputs(3052) <= not(layer0_outputs(4869));
    layer1_outputs(3053) <= not(layer0_outputs(4326));
    layer1_outputs(3054) <= (layer0_outputs(5009)) and not (layer0_outputs(2884));
    layer1_outputs(3055) <= '1';
    layer1_outputs(3056) <= not(layer0_outputs(4682));
    layer1_outputs(3057) <= (layer0_outputs(233)) and (layer0_outputs(4347));
    layer1_outputs(3058) <= (layer0_outputs(1563)) and not (layer0_outputs(4341));
    layer1_outputs(3059) <= (layer0_outputs(498)) and not (layer0_outputs(4100));
    layer1_outputs(3060) <= (layer0_outputs(1707)) xor (layer0_outputs(1556));
    layer1_outputs(3061) <= not((layer0_outputs(3380)) or (layer0_outputs(496)));
    layer1_outputs(3062) <= (layer0_outputs(956)) or (layer0_outputs(4250));
    layer1_outputs(3063) <= (layer0_outputs(3328)) and not (layer0_outputs(3060));
    layer1_outputs(3064) <= '1';
    layer1_outputs(3065) <= (layer0_outputs(295)) and not (layer0_outputs(4260));
    layer1_outputs(3066) <= not(layer0_outputs(994)) or (layer0_outputs(4298));
    layer1_outputs(3067) <= not(layer0_outputs(1260));
    layer1_outputs(3068) <= not((layer0_outputs(2330)) or (layer0_outputs(2217)));
    layer1_outputs(3069) <= (layer0_outputs(2474)) or (layer0_outputs(1154));
    layer1_outputs(3070) <= (layer0_outputs(4742)) and not (layer0_outputs(4668));
    layer1_outputs(3071) <= layer0_outputs(4468);
    layer1_outputs(3072) <= '1';
    layer1_outputs(3073) <= not(layer0_outputs(3557));
    layer1_outputs(3074) <= layer0_outputs(2793);
    layer1_outputs(3075) <= (layer0_outputs(3281)) and (layer0_outputs(1041));
    layer1_outputs(3076) <= (layer0_outputs(2954)) and not (layer0_outputs(2868));
    layer1_outputs(3077) <= not((layer0_outputs(3601)) or (layer0_outputs(4842)));
    layer1_outputs(3078) <= (layer0_outputs(2796)) and not (layer0_outputs(4424));
    layer1_outputs(3079) <= not(layer0_outputs(297)) or (layer0_outputs(1572));
    layer1_outputs(3080) <= layer0_outputs(3178);
    layer1_outputs(3081) <= layer0_outputs(800);
    layer1_outputs(3082) <= not(layer0_outputs(1667));
    layer1_outputs(3083) <= layer0_outputs(1753);
    layer1_outputs(3084) <= not(layer0_outputs(569)) or (layer0_outputs(3893));
    layer1_outputs(3085) <= layer0_outputs(4728);
    layer1_outputs(3086) <= layer0_outputs(1343);
    layer1_outputs(3087) <= not((layer0_outputs(2801)) or (layer0_outputs(4594)));
    layer1_outputs(3088) <= (layer0_outputs(1151)) and not (layer0_outputs(4425));
    layer1_outputs(3089) <= not(layer0_outputs(1950));
    layer1_outputs(3090) <= (layer0_outputs(3009)) and not (layer0_outputs(1407));
    layer1_outputs(3091) <= (layer0_outputs(1233)) and (layer0_outputs(1602));
    layer1_outputs(3092) <= layer0_outputs(1010);
    layer1_outputs(3093) <= not(layer0_outputs(4025)) or (layer0_outputs(392));
    layer1_outputs(3094) <= (layer0_outputs(4632)) and not (layer0_outputs(4282));
    layer1_outputs(3095) <= '0';
    layer1_outputs(3096) <= (layer0_outputs(650)) and (layer0_outputs(3282));
    layer1_outputs(3097) <= (layer0_outputs(3576)) xor (layer0_outputs(2745));
    layer1_outputs(3098) <= not(layer0_outputs(663)) or (layer0_outputs(2313));
    layer1_outputs(3099) <= not(layer0_outputs(1882));
    layer1_outputs(3100) <= not(layer0_outputs(3532));
    layer1_outputs(3101) <= layer0_outputs(1599);
    layer1_outputs(3102) <= layer0_outputs(4303);
    layer1_outputs(3103) <= (layer0_outputs(1974)) and (layer0_outputs(5));
    layer1_outputs(3104) <= layer0_outputs(1823);
    layer1_outputs(3105) <= (layer0_outputs(1585)) and (layer0_outputs(4642));
    layer1_outputs(3106) <= not(layer0_outputs(976)) or (layer0_outputs(342));
    layer1_outputs(3107) <= not(layer0_outputs(4277));
    layer1_outputs(3108) <= not(layer0_outputs(1493));
    layer1_outputs(3109) <= (layer0_outputs(2875)) and not (layer0_outputs(2704));
    layer1_outputs(3110) <= (layer0_outputs(4113)) and (layer0_outputs(3324));
    layer1_outputs(3111) <= not((layer0_outputs(1835)) xor (layer0_outputs(1467)));
    layer1_outputs(3112) <= (layer0_outputs(2696)) or (layer0_outputs(4255));
    layer1_outputs(3113) <= (layer0_outputs(967)) and not (layer0_outputs(1375));
    layer1_outputs(3114) <= (layer0_outputs(2616)) and not (layer0_outputs(1761));
    layer1_outputs(3115) <= not(layer0_outputs(1267));
    layer1_outputs(3116) <= layer0_outputs(418);
    layer1_outputs(3117) <= not((layer0_outputs(1274)) or (layer0_outputs(5058)));
    layer1_outputs(3118) <= not(layer0_outputs(1869));
    layer1_outputs(3119) <= not(layer0_outputs(1870)) or (layer0_outputs(4295));
    layer1_outputs(3120) <= not(layer0_outputs(543)) or (layer0_outputs(3462));
    layer1_outputs(3121) <= (layer0_outputs(5041)) xor (layer0_outputs(2061));
    layer1_outputs(3122) <= not((layer0_outputs(2021)) or (layer0_outputs(4611)));
    layer1_outputs(3123) <= not(layer0_outputs(592));
    layer1_outputs(3124) <= '0';
    layer1_outputs(3125) <= not(layer0_outputs(2812));
    layer1_outputs(3126) <= (layer0_outputs(4203)) and (layer0_outputs(3273));
    layer1_outputs(3127) <= not(layer0_outputs(1587));
    layer1_outputs(3128) <= not(layer0_outputs(130));
    layer1_outputs(3129) <= layer0_outputs(3127);
    layer1_outputs(3130) <= not((layer0_outputs(1783)) and (layer0_outputs(726)));
    layer1_outputs(3131) <= not(layer0_outputs(4563));
    layer1_outputs(3132) <= not(layer0_outputs(458));
    layer1_outputs(3133) <= (layer0_outputs(4707)) and not (layer0_outputs(3372));
    layer1_outputs(3134) <= layer0_outputs(2446);
    layer1_outputs(3135) <= (layer0_outputs(1578)) or (layer0_outputs(4265));
    layer1_outputs(3136) <= not(layer0_outputs(4782));
    layer1_outputs(3137) <= (layer0_outputs(1054)) and not (layer0_outputs(4187));
    layer1_outputs(3138) <= not(layer0_outputs(4475));
    layer1_outputs(3139) <= (layer0_outputs(1736)) and not (layer0_outputs(2908));
    layer1_outputs(3140) <= (layer0_outputs(1773)) or (layer0_outputs(1441));
    layer1_outputs(3141) <= '0';
    layer1_outputs(3142) <= not(layer0_outputs(900)) or (layer0_outputs(4864));
    layer1_outputs(3143) <= '0';
    layer1_outputs(3144) <= (layer0_outputs(4656)) and not (layer0_outputs(208));
    layer1_outputs(3145) <= not((layer0_outputs(284)) or (layer0_outputs(681)));
    layer1_outputs(3146) <= (layer0_outputs(4152)) or (layer0_outputs(2082));
    layer1_outputs(3147) <= not((layer0_outputs(2430)) or (layer0_outputs(1276)));
    layer1_outputs(3148) <= not(layer0_outputs(1977)) or (layer0_outputs(2989));
    layer1_outputs(3149) <= (layer0_outputs(3001)) or (layer0_outputs(4133));
    layer1_outputs(3150) <= (layer0_outputs(1469)) or (layer0_outputs(3652));
    layer1_outputs(3151) <= not((layer0_outputs(1065)) and (layer0_outputs(2798)));
    layer1_outputs(3152) <= not(layer0_outputs(1623));
    layer1_outputs(3153) <= not(layer0_outputs(778));
    layer1_outputs(3154) <= layer0_outputs(3057);
    layer1_outputs(3155) <= not(layer0_outputs(2375));
    layer1_outputs(3156) <= not(layer0_outputs(4065)) or (layer0_outputs(1577));
    layer1_outputs(3157) <= (layer0_outputs(1199)) and (layer0_outputs(1928));
    layer1_outputs(3158) <= not(layer0_outputs(41)) or (layer0_outputs(1998));
    layer1_outputs(3159) <= not(layer0_outputs(1604));
    layer1_outputs(3160) <= (layer0_outputs(496)) and not (layer0_outputs(5040));
    layer1_outputs(3161) <= (layer0_outputs(3639)) and not (layer0_outputs(1586));
    layer1_outputs(3162) <= not((layer0_outputs(3567)) and (layer0_outputs(571)));
    layer1_outputs(3163) <= (layer0_outputs(1389)) or (layer0_outputs(98));
    layer1_outputs(3164) <= not((layer0_outputs(2184)) and (layer0_outputs(2528)));
    layer1_outputs(3165) <= not((layer0_outputs(3109)) or (layer0_outputs(2114)));
    layer1_outputs(3166) <= not((layer0_outputs(2029)) or (layer0_outputs(1767)));
    layer1_outputs(3167) <= (layer0_outputs(408)) or (layer0_outputs(3677));
    layer1_outputs(3168) <= (layer0_outputs(4156)) or (layer0_outputs(2648));
    layer1_outputs(3169) <= not(layer0_outputs(3452)) or (layer0_outputs(4519));
    layer1_outputs(3170) <= (layer0_outputs(1504)) and not (layer0_outputs(690));
    layer1_outputs(3171) <= (layer0_outputs(481)) and not (layer0_outputs(1047));
    layer1_outputs(3172) <= (layer0_outputs(1145)) or (layer0_outputs(2116));
    layer1_outputs(3173) <= not(layer0_outputs(374));
    layer1_outputs(3174) <= (layer0_outputs(4402)) and not (layer0_outputs(3222));
    layer1_outputs(3175) <= not(layer0_outputs(2019));
    layer1_outputs(3176) <= not((layer0_outputs(4230)) or (layer0_outputs(558)));
    layer1_outputs(3177) <= not(layer0_outputs(2554));
    layer1_outputs(3178) <= not((layer0_outputs(4620)) and (layer0_outputs(18)));
    layer1_outputs(3179) <= not((layer0_outputs(2105)) or (layer0_outputs(378)));
    layer1_outputs(3180) <= (layer0_outputs(4942)) and (layer0_outputs(3108));
    layer1_outputs(3181) <= '0';
    layer1_outputs(3182) <= (layer0_outputs(3771)) and (layer0_outputs(1872));
    layer1_outputs(3183) <= not(layer0_outputs(4939)) or (layer0_outputs(3478));
    layer1_outputs(3184) <= layer0_outputs(233);
    layer1_outputs(3185) <= not(layer0_outputs(4682));
    layer1_outputs(3186) <= not(layer0_outputs(1876));
    layer1_outputs(3187) <= not((layer0_outputs(3548)) and (layer0_outputs(3012)));
    layer1_outputs(3188) <= (layer0_outputs(3091)) xor (layer0_outputs(3432));
    layer1_outputs(3189) <= (layer0_outputs(5094)) and (layer0_outputs(1247));
    layer1_outputs(3190) <= not(layer0_outputs(1406));
    layer1_outputs(3191) <= not(layer0_outputs(3911));
    layer1_outputs(3192) <= '0';
    layer1_outputs(3193) <= (layer0_outputs(2474)) and not (layer0_outputs(882));
    layer1_outputs(3194) <= layer0_outputs(3586);
    layer1_outputs(3195) <= (layer0_outputs(4658)) or (layer0_outputs(3711));
    layer1_outputs(3196) <= not((layer0_outputs(1285)) or (layer0_outputs(1370)));
    layer1_outputs(3197) <= (layer0_outputs(344)) and not (layer0_outputs(3359));
    layer1_outputs(3198) <= not(layer0_outputs(2440));
    layer1_outputs(3199) <= (layer0_outputs(2235)) and (layer0_outputs(3664));
    layer1_outputs(3200) <= (layer0_outputs(92)) xor (layer0_outputs(3548));
    layer1_outputs(3201) <= layer0_outputs(1832);
    layer1_outputs(3202) <= not(layer0_outputs(2199));
    layer1_outputs(3203) <= layer0_outputs(838);
    layer1_outputs(3204) <= not(layer0_outputs(2028));
    layer1_outputs(3205) <= layer0_outputs(750);
    layer1_outputs(3206) <= not((layer0_outputs(3430)) xor (layer0_outputs(1404)));
    layer1_outputs(3207) <= (layer0_outputs(3854)) and not (layer0_outputs(3209));
    layer1_outputs(3208) <= not(layer0_outputs(773));
    layer1_outputs(3209) <= (layer0_outputs(1648)) xor (layer0_outputs(4943));
    layer1_outputs(3210) <= not(layer0_outputs(5020));
    layer1_outputs(3211) <= layer0_outputs(4502);
    layer1_outputs(3212) <= layer0_outputs(4155);
    layer1_outputs(3213) <= (layer0_outputs(2431)) or (layer0_outputs(2261));
    layer1_outputs(3214) <= layer0_outputs(749);
    layer1_outputs(3215) <= '1';
    layer1_outputs(3216) <= not(layer0_outputs(966));
    layer1_outputs(3217) <= (layer0_outputs(4164)) and (layer0_outputs(2622));
    layer1_outputs(3218) <= (layer0_outputs(4803)) and not (layer0_outputs(4207));
    layer1_outputs(3219) <= layer0_outputs(600);
    layer1_outputs(3220) <= (layer0_outputs(2661)) and not (layer0_outputs(4513));
    layer1_outputs(3221) <= layer0_outputs(4845);
    layer1_outputs(3222) <= not((layer0_outputs(1286)) xor (layer0_outputs(3580)));
    layer1_outputs(3223) <= layer0_outputs(2090);
    layer1_outputs(3224) <= layer0_outputs(2898);
    layer1_outputs(3225) <= layer0_outputs(4898);
    layer1_outputs(3226) <= not(layer0_outputs(605)) or (layer0_outputs(2202));
    layer1_outputs(3227) <= not(layer0_outputs(3441));
    layer1_outputs(3228) <= layer0_outputs(3307);
    layer1_outputs(3229) <= (layer0_outputs(3162)) and (layer0_outputs(1299));
    layer1_outputs(3230) <= not(layer0_outputs(104)) or (layer0_outputs(2006));
    layer1_outputs(3231) <= not(layer0_outputs(2893));
    layer1_outputs(3232) <= not(layer0_outputs(2119));
    layer1_outputs(3233) <= '0';
    layer1_outputs(3234) <= not(layer0_outputs(1695));
    layer1_outputs(3235) <= not(layer0_outputs(1269)) or (layer0_outputs(206));
    layer1_outputs(3236) <= not(layer0_outputs(1350)) or (layer0_outputs(1606));
    layer1_outputs(3237) <= not((layer0_outputs(1144)) xor (layer0_outputs(207)));
    layer1_outputs(3238) <= not((layer0_outputs(1921)) or (layer0_outputs(754)));
    layer1_outputs(3239) <= (layer0_outputs(2292)) and (layer0_outputs(4368));
    layer1_outputs(3240) <= '1';
    layer1_outputs(3241) <= not(layer0_outputs(429));
    layer1_outputs(3242) <= '1';
    layer1_outputs(3243) <= (layer0_outputs(4882)) or (layer0_outputs(2423));
    layer1_outputs(3244) <= not(layer0_outputs(2098)) or (layer0_outputs(5061));
    layer1_outputs(3245) <= not(layer0_outputs(1259)) or (layer0_outputs(550));
    layer1_outputs(3246) <= not(layer0_outputs(4116));
    layer1_outputs(3247) <= (layer0_outputs(5083)) and not (layer0_outputs(811));
    layer1_outputs(3248) <= not(layer0_outputs(193));
    layer1_outputs(3249) <= (layer0_outputs(2226)) and not (layer0_outputs(4498));
    layer1_outputs(3250) <= (layer0_outputs(2918)) or (layer0_outputs(4556));
    layer1_outputs(3251) <= layer0_outputs(3045);
    layer1_outputs(3252) <= (layer0_outputs(2822)) and (layer0_outputs(3871));
    layer1_outputs(3253) <= (layer0_outputs(4618)) and not (layer0_outputs(3690));
    layer1_outputs(3254) <= layer0_outputs(351);
    layer1_outputs(3255) <= (layer0_outputs(1699)) and (layer0_outputs(1301));
    layer1_outputs(3256) <= not((layer0_outputs(4873)) and (layer0_outputs(675)));
    layer1_outputs(3257) <= layer0_outputs(3428);
    layer1_outputs(3258) <= (layer0_outputs(4404)) and not (layer0_outputs(857));
    layer1_outputs(3259) <= (layer0_outputs(2654)) and (layer0_outputs(1422));
    layer1_outputs(3260) <= not(layer0_outputs(586));
    layer1_outputs(3261) <= layer0_outputs(2341);
    layer1_outputs(3262) <= not(layer0_outputs(2370));
    layer1_outputs(3263) <= (layer0_outputs(502)) or (layer0_outputs(2264));
    layer1_outputs(3264) <= layer0_outputs(4703);
    layer1_outputs(3265) <= not(layer0_outputs(3830)) or (layer0_outputs(852));
    layer1_outputs(3266) <= not(layer0_outputs(2106));
    layer1_outputs(3267) <= (layer0_outputs(2452)) or (layer0_outputs(5005));
    layer1_outputs(3268) <= not(layer0_outputs(2820)) or (layer0_outputs(2103));
    layer1_outputs(3269) <= not(layer0_outputs(4304));
    layer1_outputs(3270) <= (layer0_outputs(3013)) and (layer0_outputs(3357));
    layer1_outputs(3271) <= (layer0_outputs(1457)) and (layer0_outputs(631));
    layer1_outputs(3272) <= (layer0_outputs(544)) or (layer0_outputs(2552));
    layer1_outputs(3273) <= (layer0_outputs(4380)) or (layer0_outputs(3536));
    layer1_outputs(3274) <= not(layer0_outputs(1189));
    layer1_outputs(3275) <= layer0_outputs(3176);
    layer1_outputs(3276) <= (layer0_outputs(5099)) and not (layer0_outputs(1265));
    layer1_outputs(3277) <= (layer0_outputs(3439)) or (layer0_outputs(3907));
    layer1_outputs(3278) <= layer0_outputs(1423);
    layer1_outputs(3279) <= layer0_outputs(4653);
    layer1_outputs(3280) <= (layer0_outputs(169)) and not (layer0_outputs(3359));
    layer1_outputs(3281) <= not(layer0_outputs(4192));
    layer1_outputs(3282) <= '0';
    layer1_outputs(3283) <= not(layer0_outputs(3482)) or (layer0_outputs(2923));
    layer1_outputs(3284) <= not((layer0_outputs(736)) and (layer0_outputs(3839)));
    layer1_outputs(3285) <= not(layer0_outputs(3584));
    layer1_outputs(3286) <= not(layer0_outputs(3063)) or (layer0_outputs(3969));
    layer1_outputs(3287) <= not(layer0_outputs(538));
    layer1_outputs(3288) <= not(layer0_outputs(1030));
    layer1_outputs(3289) <= not((layer0_outputs(5003)) or (layer0_outputs(3090)));
    layer1_outputs(3290) <= (layer0_outputs(4141)) and not (layer0_outputs(4849));
    layer1_outputs(3291) <= not((layer0_outputs(1960)) and (layer0_outputs(429)));
    layer1_outputs(3292) <= not((layer0_outputs(4151)) and (layer0_outputs(366)));
    layer1_outputs(3293) <= not(layer0_outputs(3271));
    layer1_outputs(3294) <= (layer0_outputs(5022)) or (layer0_outputs(4774));
    layer1_outputs(3295) <= (layer0_outputs(1048)) or (layer0_outputs(2295));
    layer1_outputs(3296) <= '1';
    layer1_outputs(3297) <= (layer0_outputs(254)) and not (layer0_outputs(2327));
    layer1_outputs(3298) <= (layer0_outputs(4517)) and not (layer0_outputs(2750));
    layer1_outputs(3299) <= layer0_outputs(3860);
    layer1_outputs(3300) <= (layer0_outputs(1440)) and not (layer0_outputs(1893));
    layer1_outputs(3301) <= '0';
    layer1_outputs(3302) <= not(layer0_outputs(1966));
    layer1_outputs(3303) <= not(layer0_outputs(2058));
    layer1_outputs(3304) <= not(layer0_outputs(4314)) or (layer0_outputs(975));
    layer1_outputs(3305) <= (layer0_outputs(148)) and not (layer0_outputs(4921));
    layer1_outputs(3306) <= not(layer0_outputs(3725)) or (layer0_outputs(4662));
    layer1_outputs(3307) <= (layer0_outputs(1988)) and not (layer0_outputs(4826));
    layer1_outputs(3308) <= not((layer0_outputs(1218)) xor (layer0_outputs(3101)));
    layer1_outputs(3309) <= not(layer0_outputs(1220));
    layer1_outputs(3310) <= (layer0_outputs(2699)) and (layer0_outputs(2183));
    layer1_outputs(3311) <= not((layer0_outputs(2266)) or (layer0_outputs(4943)));
    layer1_outputs(3312) <= not(layer0_outputs(2414));
    layer1_outputs(3313) <= not((layer0_outputs(1386)) and (layer0_outputs(2999)));
    layer1_outputs(3314) <= layer0_outputs(1050);
    layer1_outputs(3315) <= not(layer0_outputs(3873));
    layer1_outputs(3316) <= (layer0_outputs(4454)) and not (layer0_outputs(3788));
    layer1_outputs(3317) <= (layer0_outputs(2738)) and (layer0_outputs(3636));
    layer1_outputs(3318) <= not((layer0_outputs(1414)) or (layer0_outputs(3796)));
    layer1_outputs(3319) <= not(layer0_outputs(2176));
    layer1_outputs(3320) <= (layer0_outputs(2812)) and not (layer0_outputs(5006));
    layer1_outputs(3321) <= (layer0_outputs(2132)) and not (layer0_outputs(462));
    layer1_outputs(3322) <= layer0_outputs(3588);
    layer1_outputs(3323) <= not(layer0_outputs(1528));
    layer1_outputs(3324) <= not(layer0_outputs(2353)) or (layer0_outputs(2018));
    layer1_outputs(3325) <= (layer0_outputs(2282)) and not (layer0_outputs(2419));
    layer1_outputs(3326) <= layer0_outputs(3627);
    layer1_outputs(3327) <= not(layer0_outputs(321)) or (layer0_outputs(1537));
    layer1_outputs(3328) <= (layer0_outputs(3743)) and not (layer0_outputs(1028));
    layer1_outputs(3329) <= (layer0_outputs(1093)) and (layer0_outputs(4949));
    layer1_outputs(3330) <= layer0_outputs(2553);
    layer1_outputs(3331) <= (layer0_outputs(3891)) and not (layer0_outputs(1443));
    layer1_outputs(3332) <= not(layer0_outputs(482)) or (layer0_outputs(2174));
    layer1_outputs(3333) <= layer0_outputs(3210);
    layer1_outputs(3334) <= not((layer0_outputs(3167)) or (layer0_outputs(2523)));
    layer1_outputs(3335) <= layer0_outputs(2042);
    layer1_outputs(3336) <= (layer0_outputs(1419)) or (layer0_outputs(1699));
    layer1_outputs(3337) <= not(layer0_outputs(4316));
    layer1_outputs(3338) <= not(layer0_outputs(4696)) or (layer0_outputs(1663));
    layer1_outputs(3339) <= (layer0_outputs(3145)) xor (layer0_outputs(4990));
    layer1_outputs(3340) <= not((layer0_outputs(4807)) and (layer0_outputs(1904)));
    layer1_outputs(3341) <= not((layer0_outputs(4718)) xor (layer0_outputs(2151)));
    layer1_outputs(3342) <= not(layer0_outputs(1398));
    layer1_outputs(3343) <= layer0_outputs(2115);
    layer1_outputs(3344) <= (layer0_outputs(2325)) and not (layer0_outputs(149));
    layer1_outputs(3345) <= (layer0_outputs(174)) or (layer0_outputs(4845));
    layer1_outputs(3346) <= '0';
    layer1_outputs(3347) <= not((layer0_outputs(3244)) or (layer0_outputs(4846)));
    layer1_outputs(3348) <= (layer0_outputs(4873)) or (layer0_outputs(2591));
    layer1_outputs(3349) <= not(layer0_outputs(2783));
    layer1_outputs(3350) <= layer0_outputs(3602);
    layer1_outputs(3351) <= layer0_outputs(2267);
    layer1_outputs(3352) <= not(layer0_outputs(3244));
    layer1_outputs(3353) <= not(layer0_outputs(322)) or (layer0_outputs(2051));
    layer1_outputs(3354) <= not(layer0_outputs(2587));
    layer1_outputs(3355) <= not(layer0_outputs(17));
    layer1_outputs(3356) <= not(layer0_outputs(5050)) or (layer0_outputs(2470));
    layer1_outputs(3357) <= (layer0_outputs(547)) or (layer0_outputs(903));
    layer1_outputs(3358) <= (layer0_outputs(5050)) and not (layer0_outputs(500));
    layer1_outputs(3359) <= (layer0_outputs(2361)) or (layer0_outputs(3627));
    layer1_outputs(3360) <= layer0_outputs(441);
    layer1_outputs(3361) <= '1';
    layer1_outputs(3362) <= not(layer0_outputs(371)) or (layer0_outputs(2824));
    layer1_outputs(3363) <= layer0_outputs(3197);
    layer1_outputs(3364) <= layer0_outputs(1014);
    layer1_outputs(3365) <= layer0_outputs(3125);
    layer1_outputs(3366) <= not(layer0_outputs(3546));
    layer1_outputs(3367) <= layer0_outputs(2001);
    layer1_outputs(3368) <= (layer0_outputs(163)) xor (layer0_outputs(3942));
    layer1_outputs(3369) <= not(layer0_outputs(646)) or (layer0_outputs(3051));
    layer1_outputs(3370) <= not((layer0_outputs(4897)) or (layer0_outputs(2592)));
    layer1_outputs(3371) <= (layer0_outputs(1060)) and not (layer0_outputs(2588));
    layer1_outputs(3372) <= not(layer0_outputs(1965));
    layer1_outputs(3373) <= not(layer0_outputs(3013)) or (layer0_outputs(3979));
    layer1_outputs(3374) <= (layer0_outputs(2974)) or (layer0_outputs(4695));
    layer1_outputs(3375) <= (layer0_outputs(4890)) and (layer0_outputs(2319));
    layer1_outputs(3376) <= not(layer0_outputs(2444));
    layer1_outputs(3377) <= '0';
    layer1_outputs(3378) <= (layer0_outputs(3617)) and not (layer0_outputs(3499));
    layer1_outputs(3379) <= (layer0_outputs(1970)) and not (layer0_outputs(4234));
    layer1_outputs(3380) <= not(layer0_outputs(2062));
    layer1_outputs(3381) <= (layer0_outputs(3738)) and not (layer0_outputs(2359));
    layer1_outputs(3382) <= not((layer0_outputs(4406)) or (layer0_outputs(2786)));
    layer1_outputs(3383) <= not((layer0_outputs(824)) or (layer0_outputs(2562)));
    layer1_outputs(3384) <= not(layer0_outputs(1090)) or (layer0_outputs(2655));
    layer1_outputs(3385) <= (layer0_outputs(1655)) and not (layer0_outputs(2397));
    layer1_outputs(3386) <= (layer0_outputs(1640)) and (layer0_outputs(2673));
    layer1_outputs(3387) <= not(layer0_outputs(1730)) or (layer0_outputs(4995));
    layer1_outputs(3388) <= layer0_outputs(867);
    layer1_outputs(3389) <= not(layer0_outputs(4955)) or (layer0_outputs(3983));
    layer1_outputs(3390) <= layer0_outputs(40);
    layer1_outputs(3391) <= '0';
    layer1_outputs(3392) <= '0';
    layer1_outputs(3393) <= layer0_outputs(86);
    layer1_outputs(3394) <= not(layer0_outputs(1362));
    layer1_outputs(3395) <= (layer0_outputs(680)) and not (layer0_outputs(655));
    layer1_outputs(3396) <= not(layer0_outputs(2569)) or (layer0_outputs(2595));
    layer1_outputs(3397) <= layer0_outputs(1374);
    layer1_outputs(3398) <= not(layer0_outputs(2870));
    layer1_outputs(3399) <= not((layer0_outputs(3471)) or (layer0_outputs(904)));
    layer1_outputs(3400) <= layer0_outputs(1124);
    layer1_outputs(3401) <= not(layer0_outputs(703)) or (layer0_outputs(4669));
    layer1_outputs(3402) <= layer0_outputs(3395);
    layer1_outputs(3403) <= not(layer0_outputs(2907));
    layer1_outputs(3404) <= layer0_outputs(3672);
    layer1_outputs(3405) <= not((layer0_outputs(406)) and (layer0_outputs(4588)));
    layer1_outputs(3406) <= (layer0_outputs(1210)) and not (layer0_outputs(822));
    layer1_outputs(3407) <= (layer0_outputs(4956)) and not (layer0_outputs(4819));
    layer1_outputs(3408) <= not(layer0_outputs(590));
    layer1_outputs(3409) <= not((layer0_outputs(4359)) xor (layer0_outputs(1825)));
    layer1_outputs(3410) <= not(layer0_outputs(666));
    layer1_outputs(3411) <= not((layer0_outputs(4939)) and (layer0_outputs(2551)));
    layer1_outputs(3412) <= layer0_outputs(1710);
    layer1_outputs(3413) <= layer0_outputs(3601);
    layer1_outputs(3414) <= not((layer0_outputs(4458)) xor (layer0_outputs(2866)));
    layer1_outputs(3415) <= not(layer0_outputs(4220));
    layer1_outputs(3416) <= not(layer0_outputs(912));
    layer1_outputs(3417) <= not(layer0_outputs(4908));
    layer1_outputs(3418) <= not(layer0_outputs(4601));
    layer1_outputs(3419) <= not(layer0_outputs(3823)) or (layer0_outputs(122));
    layer1_outputs(3420) <= not((layer0_outputs(4020)) or (layer0_outputs(1916)));
    layer1_outputs(3421) <= layer0_outputs(133);
    layer1_outputs(3422) <= (layer0_outputs(1042)) xor (layer0_outputs(702));
    layer1_outputs(3423) <= not((layer0_outputs(1061)) and (layer0_outputs(3558)));
    layer1_outputs(3424) <= layer0_outputs(3272);
    layer1_outputs(3425) <= not((layer0_outputs(1830)) xor (layer0_outputs(3480)));
    layer1_outputs(3426) <= (layer0_outputs(2883)) and not (layer0_outputs(1546));
    layer1_outputs(3427) <= (layer0_outputs(4854)) xor (layer0_outputs(2189));
    layer1_outputs(3428) <= layer0_outputs(1683);
    layer1_outputs(3429) <= layer0_outputs(452);
    layer1_outputs(3430) <= (layer0_outputs(2443)) and not (layer0_outputs(101));
    layer1_outputs(3431) <= not(layer0_outputs(1652));
    layer1_outputs(3432) <= layer0_outputs(4583);
    layer1_outputs(3433) <= layer0_outputs(3384);
    layer1_outputs(3434) <= (layer0_outputs(3392)) and not (layer0_outputs(3340));
    layer1_outputs(3435) <= layer0_outputs(3445);
    layer1_outputs(3436) <= not(layer0_outputs(4754)) or (layer0_outputs(4890));
    layer1_outputs(3437) <= (layer0_outputs(4216)) and not (layer0_outputs(3935));
    layer1_outputs(3438) <= not(layer0_outputs(1462));
    layer1_outputs(3439) <= not(layer0_outputs(2162));
    layer1_outputs(3440) <= not((layer0_outputs(269)) xor (layer0_outputs(746)));
    layer1_outputs(3441) <= layer0_outputs(3618);
    layer1_outputs(3442) <= not(layer0_outputs(2849));
    layer1_outputs(3443) <= not(layer0_outputs(2044));
    layer1_outputs(3444) <= (layer0_outputs(2852)) xor (layer0_outputs(2900));
    layer1_outputs(3445) <= (layer0_outputs(2092)) and not (layer0_outputs(2973));
    layer1_outputs(3446) <= layer0_outputs(3987);
    layer1_outputs(3447) <= layer0_outputs(742);
    layer1_outputs(3448) <= not(layer0_outputs(3819)) or (layer0_outputs(956));
    layer1_outputs(3449) <= not((layer0_outputs(868)) xor (layer0_outputs(4536)));
    layer1_outputs(3450) <= not(layer0_outputs(701)) or (layer0_outputs(1106));
    layer1_outputs(3451) <= (layer0_outputs(2463)) and not (layer0_outputs(630));
    layer1_outputs(3452) <= (layer0_outputs(2863)) xor (layer0_outputs(2871));
    layer1_outputs(3453) <= layer0_outputs(1890);
    layer1_outputs(3454) <= not(layer0_outputs(4196)) or (layer0_outputs(4586));
    layer1_outputs(3455) <= layer0_outputs(4884);
    layer1_outputs(3456) <= not(layer0_outputs(4765)) or (layer0_outputs(1268));
    layer1_outputs(3457) <= not(layer0_outputs(4977));
    layer1_outputs(3458) <= (layer0_outputs(5032)) and (layer0_outputs(4525));
    layer1_outputs(3459) <= layer0_outputs(3259);
    layer1_outputs(3460) <= (layer0_outputs(191)) and (layer0_outputs(3467));
    layer1_outputs(3461) <= not((layer0_outputs(1420)) or (layer0_outputs(494)));
    layer1_outputs(3462) <= not(layer0_outputs(1734));
    layer1_outputs(3463) <= (layer0_outputs(2379)) xor (layer0_outputs(11));
    layer1_outputs(3464) <= (layer0_outputs(1625)) xor (layer0_outputs(4718));
    layer1_outputs(3465) <= not(layer0_outputs(4149)) or (layer0_outputs(3786));
    layer1_outputs(3466) <= not(layer0_outputs(2265));
    layer1_outputs(3467) <= not(layer0_outputs(1910));
    layer1_outputs(3468) <= layer0_outputs(3059);
    layer1_outputs(3469) <= not(layer0_outputs(2803)) or (layer0_outputs(4529));
    layer1_outputs(3470) <= not(layer0_outputs(2332));
    layer1_outputs(3471) <= not((layer0_outputs(3661)) and (layer0_outputs(780)));
    layer1_outputs(3472) <= not((layer0_outputs(1954)) or (layer0_outputs(4697)));
    layer1_outputs(3473) <= not(layer0_outputs(2827)) or (layer0_outputs(721));
    layer1_outputs(3474) <= (layer0_outputs(2019)) and not (layer0_outputs(4402));
    layer1_outputs(3475) <= (layer0_outputs(4992)) and not (layer0_outputs(2727));
    layer1_outputs(3476) <= (layer0_outputs(3785)) and (layer0_outputs(204));
    layer1_outputs(3477) <= not(layer0_outputs(4111));
    layer1_outputs(3478) <= not((layer0_outputs(71)) or (layer0_outputs(3376)));
    layer1_outputs(3479) <= not((layer0_outputs(182)) or (layer0_outputs(1328)));
    layer1_outputs(3480) <= (layer0_outputs(829)) and not (layer0_outputs(1134));
    layer1_outputs(3481) <= not(layer0_outputs(3248));
    layer1_outputs(3482) <= layer0_outputs(2716);
    layer1_outputs(3483) <= not(layer0_outputs(3689)) or (layer0_outputs(4911));
    layer1_outputs(3484) <= layer0_outputs(2834);
    layer1_outputs(3485) <= (layer0_outputs(4906)) and not (layer0_outputs(1579));
    layer1_outputs(3486) <= layer0_outputs(4062);
    layer1_outputs(3487) <= not(layer0_outputs(2779));
    layer1_outputs(3488) <= layer0_outputs(1116);
    layer1_outputs(3489) <= (layer0_outputs(357)) xor (layer0_outputs(458));
    layer1_outputs(3490) <= not((layer0_outputs(4683)) and (layer0_outputs(4944)));
    layer1_outputs(3491) <= layer0_outputs(1170);
    layer1_outputs(3492) <= layer0_outputs(1424);
    layer1_outputs(3493) <= layer0_outputs(1570);
    layer1_outputs(3494) <= '1';
    layer1_outputs(3495) <= not(layer0_outputs(3168));
    layer1_outputs(3496) <= not(layer0_outputs(3464)) or (layer0_outputs(2702));
    layer1_outputs(3497) <= layer0_outputs(4724);
    layer1_outputs(3498) <= not((layer0_outputs(4006)) xor (layer0_outputs(4356)));
    layer1_outputs(3499) <= layer0_outputs(2373);
    layer1_outputs(3500) <= not((layer0_outputs(4004)) or (layer0_outputs(123)));
    layer1_outputs(3501) <= layer0_outputs(2769);
    layer1_outputs(3502) <= not(layer0_outputs(1174));
    layer1_outputs(3503) <= not(layer0_outputs(2063)) or (layer0_outputs(3365));
    layer1_outputs(3504) <= layer0_outputs(3175);
    layer1_outputs(3505) <= not((layer0_outputs(4196)) or (layer0_outputs(2694)));
    layer1_outputs(3506) <= layer0_outputs(2340);
    layer1_outputs(3507) <= not(layer0_outputs(3310)) or (layer0_outputs(4671));
    layer1_outputs(3508) <= not((layer0_outputs(444)) and (layer0_outputs(4340)));
    layer1_outputs(3509) <= (layer0_outputs(68)) and not (layer0_outputs(5060));
    layer1_outputs(3510) <= (layer0_outputs(1883)) and not (layer0_outputs(3741));
    layer1_outputs(3511) <= not(layer0_outputs(1139));
    layer1_outputs(3512) <= (layer0_outputs(1344)) and (layer0_outputs(3822));
    layer1_outputs(3513) <= (layer0_outputs(1082)) and not (layer0_outputs(4554));
    layer1_outputs(3514) <= not((layer0_outputs(488)) or (layer0_outputs(2534)));
    layer1_outputs(3515) <= layer0_outputs(895);
    layer1_outputs(3516) <= not(layer0_outputs(1129)) or (layer0_outputs(317));
    layer1_outputs(3517) <= layer0_outputs(3279);
    layer1_outputs(3518) <= not((layer0_outputs(2676)) xor (layer0_outputs(4958)));
    layer1_outputs(3519) <= '0';
    layer1_outputs(3520) <= layer0_outputs(3992);
    layer1_outputs(3521) <= (layer0_outputs(1891)) xor (layer0_outputs(3083));
    layer1_outputs(3522) <= (layer0_outputs(384)) and not (layer0_outputs(971));
    layer1_outputs(3523) <= not(layer0_outputs(738));
    layer1_outputs(3524) <= not(layer0_outputs(1080));
    layer1_outputs(3525) <= not(layer0_outputs(2186));
    layer1_outputs(3526) <= layer0_outputs(3608);
    layer1_outputs(3527) <= not(layer0_outputs(1603));
    layer1_outputs(3528) <= not(layer0_outputs(1914));
    layer1_outputs(3529) <= layer0_outputs(4893);
    layer1_outputs(3530) <= not(layer0_outputs(54));
    layer1_outputs(3531) <= not((layer0_outputs(1359)) and (layer0_outputs(3133)));
    layer1_outputs(3532) <= not(layer0_outputs(235)) or (layer0_outputs(1251));
    layer1_outputs(3533) <= (layer0_outputs(2966)) xor (layer0_outputs(3418));
    layer1_outputs(3534) <= not((layer0_outputs(2206)) or (layer0_outputs(1790)));
    layer1_outputs(3535) <= (layer0_outputs(3390)) or (layer0_outputs(4320));
    layer1_outputs(3536) <= layer0_outputs(4372);
    layer1_outputs(3537) <= not((layer0_outputs(1996)) or (layer0_outputs(906)));
    layer1_outputs(3538) <= not(layer0_outputs(3748));
    layer1_outputs(3539) <= not(layer0_outputs(2605));
    layer1_outputs(3540) <= not(layer0_outputs(2007));
    layer1_outputs(3541) <= not(layer0_outputs(31)) or (layer0_outputs(1433));
    layer1_outputs(3542) <= '1';
    layer1_outputs(3543) <= not(layer0_outputs(4563)) or (layer0_outputs(2206));
    layer1_outputs(3544) <= (layer0_outputs(3299)) and (layer0_outputs(4877));
    layer1_outputs(3545) <= layer0_outputs(1877);
    layer1_outputs(3546) <= layer0_outputs(2420);
    layer1_outputs(3547) <= layer0_outputs(4700);
    layer1_outputs(3548) <= '1';
    layer1_outputs(3549) <= layer0_outputs(1580);
    layer1_outputs(3550) <= (layer0_outputs(3843)) or (layer0_outputs(1038));
    layer1_outputs(3551) <= not(layer0_outputs(2167));
    layer1_outputs(3552) <= (layer0_outputs(386)) and not (layer0_outputs(1979));
    layer1_outputs(3553) <= layer0_outputs(2546);
    layer1_outputs(3554) <= (layer0_outputs(1418)) or (layer0_outputs(1989));
    layer1_outputs(3555) <= layer0_outputs(447);
    layer1_outputs(3556) <= not(layer0_outputs(4602));
    layer1_outputs(3557) <= layer0_outputs(4924);
    layer1_outputs(3558) <= (layer0_outputs(3466)) and not (layer0_outputs(3718));
    layer1_outputs(3559) <= not(layer0_outputs(1565));
    layer1_outputs(3560) <= not(layer0_outputs(2396));
    layer1_outputs(3561) <= not((layer0_outputs(2599)) xor (layer0_outputs(4256)));
    layer1_outputs(3562) <= not(layer0_outputs(5076));
    layer1_outputs(3563) <= not(layer0_outputs(3524)) or (layer0_outputs(4991));
    layer1_outputs(3564) <= not(layer0_outputs(3073)) or (layer0_outputs(2905));
    layer1_outputs(3565) <= not(layer0_outputs(1412)) or (layer0_outputs(1781));
    layer1_outputs(3566) <= not(layer0_outputs(748));
    layer1_outputs(3567) <= layer0_outputs(2471);
    layer1_outputs(3568) <= layer0_outputs(4167);
    layer1_outputs(3569) <= layer0_outputs(4614);
    layer1_outputs(3570) <= layer0_outputs(530);
    layer1_outputs(3571) <= '1';
    layer1_outputs(3572) <= not(layer0_outputs(3241));
    layer1_outputs(3573) <= not(layer0_outputs(2481)) or (layer0_outputs(657));
    layer1_outputs(3574) <= layer0_outputs(3696);
    layer1_outputs(3575) <= layer0_outputs(5116);
    layer1_outputs(3576) <= not(layer0_outputs(1810));
    layer1_outputs(3577) <= not(layer0_outputs(3516));
    layer1_outputs(3578) <= not(layer0_outputs(4659));
    layer1_outputs(3579) <= '0';
    layer1_outputs(3580) <= (layer0_outputs(2369)) and not (layer0_outputs(4952));
    layer1_outputs(3581) <= not(layer0_outputs(3277));
    layer1_outputs(3582) <= not(layer0_outputs(3678)) or (layer0_outputs(3408));
    layer1_outputs(3583) <= not(layer0_outputs(2403));
    layer1_outputs(3584) <= (layer0_outputs(2371)) or (layer0_outputs(1211));
    layer1_outputs(3585) <= layer0_outputs(3390);
    layer1_outputs(3586) <= (layer0_outputs(4511)) and not (layer0_outputs(5053));
    layer1_outputs(3587) <= (layer0_outputs(3488)) and not (layer0_outputs(1653));
    layer1_outputs(3588) <= not(layer0_outputs(1843)) or (layer0_outputs(2683));
    layer1_outputs(3589) <= layer0_outputs(537);
    layer1_outputs(3590) <= layer0_outputs(241);
    layer1_outputs(3591) <= (layer0_outputs(1267)) and (layer0_outputs(3759));
    layer1_outputs(3592) <= not((layer0_outputs(2178)) or (layer0_outputs(2096)));
    layer1_outputs(3593) <= (layer0_outputs(1021)) and (layer0_outputs(3624));
    layer1_outputs(3594) <= not(layer0_outputs(646)) or (layer0_outputs(1773));
    layer1_outputs(3595) <= not(layer0_outputs(2823));
    layer1_outputs(3596) <= not(layer0_outputs(334));
    layer1_outputs(3597) <= (layer0_outputs(488)) and (layer0_outputs(2880));
    layer1_outputs(3598) <= (layer0_outputs(2961)) and not (layer0_outputs(3849));
    layer1_outputs(3599) <= (layer0_outputs(2675)) or (layer0_outputs(3311));
    layer1_outputs(3600) <= '1';
    layer1_outputs(3601) <= not((layer0_outputs(1073)) and (layer0_outputs(801)));
    layer1_outputs(3602) <= layer0_outputs(4502);
    layer1_outputs(3603) <= not(layer0_outputs(3930));
    layer1_outputs(3604) <= layer0_outputs(634);
    layer1_outputs(3605) <= layer0_outputs(37);
    layer1_outputs(3606) <= not((layer0_outputs(1814)) or (layer0_outputs(1261)));
    layer1_outputs(3607) <= (layer0_outputs(4362)) and (layer0_outputs(1892));
    layer1_outputs(3608) <= (layer0_outputs(42)) or (layer0_outputs(542));
    layer1_outputs(3609) <= not((layer0_outputs(1529)) or (layer0_outputs(5099)));
    layer1_outputs(3610) <= not(layer0_outputs(861));
    layer1_outputs(3611) <= not((layer0_outputs(1855)) and (layer0_outputs(665)));
    layer1_outputs(3612) <= not(layer0_outputs(1799)) or (layer0_outputs(2902));
    layer1_outputs(3613) <= '0';
    layer1_outputs(3614) <= not(layer0_outputs(2645));
    layer1_outputs(3615) <= layer0_outputs(4681);
    layer1_outputs(3616) <= layer0_outputs(2220);
    layer1_outputs(3617) <= not((layer0_outputs(1260)) or (layer0_outputs(898)));
    layer1_outputs(3618) <= (layer0_outputs(4712)) and not (layer0_outputs(4604));
    layer1_outputs(3619) <= (layer0_outputs(3656)) or (layer0_outputs(2030));
    layer1_outputs(3620) <= not(layer0_outputs(4809));
    layer1_outputs(3621) <= (layer0_outputs(1548)) and not (layer0_outputs(3610));
    layer1_outputs(3622) <= (layer0_outputs(2862)) and not (layer0_outputs(2755));
    layer1_outputs(3623) <= not(layer0_outputs(85));
    layer1_outputs(3624) <= (layer0_outputs(361)) or (layer0_outputs(777));
    layer1_outputs(3625) <= (layer0_outputs(3449)) or (layer0_outputs(3025));
    layer1_outputs(3626) <= layer0_outputs(1764);
    layer1_outputs(3627) <= not((layer0_outputs(4269)) or (layer0_outputs(3559)));
    layer1_outputs(3628) <= '0';
    layer1_outputs(3629) <= not(layer0_outputs(2600)) or (layer0_outputs(1943));
    layer1_outputs(3630) <= not(layer0_outputs(4315));
    layer1_outputs(3631) <= layer0_outputs(4031);
    layer1_outputs(3632) <= layer0_outputs(913);
    layer1_outputs(3633) <= not(layer0_outputs(1037));
    layer1_outputs(3634) <= '1';
    layer1_outputs(3635) <= not((layer0_outputs(3413)) and (layer0_outputs(3693)));
    layer1_outputs(3636) <= (layer0_outputs(2693)) or (layer0_outputs(3007));
    layer1_outputs(3637) <= not((layer0_outputs(4568)) or (layer0_outputs(908)));
    layer1_outputs(3638) <= not(layer0_outputs(661));
    layer1_outputs(3639) <= not(layer0_outputs(1204)) or (layer0_outputs(3534));
    layer1_outputs(3640) <= not(layer0_outputs(4111)) or (layer0_outputs(456));
    layer1_outputs(3641) <= not(layer0_outputs(2799));
    layer1_outputs(3642) <= layer0_outputs(1003);
    layer1_outputs(3643) <= not(layer0_outputs(4496));
    layer1_outputs(3644) <= not(layer0_outputs(1271));
    layer1_outputs(3645) <= layer0_outputs(1431);
    layer1_outputs(3646) <= not((layer0_outputs(2454)) or (layer0_outputs(710)));
    layer1_outputs(3647) <= not(layer0_outputs(1230));
    layer1_outputs(3648) <= (layer0_outputs(744)) and not (layer0_outputs(127));
    layer1_outputs(3649) <= layer0_outputs(667);
    layer1_outputs(3650) <= (layer0_outputs(4160)) and not (layer0_outputs(1538));
    layer1_outputs(3651) <= not(layer0_outputs(4138)) or (layer0_outputs(3186));
    layer1_outputs(3652) <= (layer0_outputs(1250)) and (layer0_outputs(582));
    layer1_outputs(3653) <= layer0_outputs(4723);
    layer1_outputs(3654) <= (layer0_outputs(3543)) and not (layer0_outputs(3410));
    layer1_outputs(3655) <= layer0_outputs(2118);
    layer1_outputs(3656) <= not((layer0_outputs(197)) or (layer0_outputs(3734)));
    layer1_outputs(3657) <= (layer0_outputs(128)) and (layer0_outputs(2011));
    layer1_outputs(3658) <= layer0_outputs(3722);
    layer1_outputs(3659) <= (layer0_outputs(1889)) and not (layer0_outputs(775));
    layer1_outputs(3660) <= layer0_outputs(4582);
    layer1_outputs(3661) <= not((layer0_outputs(810)) or (layer0_outputs(1660)));
    layer1_outputs(3662) <= layer0_outputs(3231);
    layer1_outputs(3663) <= '0';
    layer1_outputs(3664) <= not(layer0_outputs(538)) or (layer0_outputs(1966));
    layer1_outputs(3665) <= (layer0_outputs(356)) and not (layer0_outputs(4051));
    layer1_outputs(3666) <= (layer0_outputs(4599)) and (layer0_outputs(4396));
    layer1_outputs(3667) <= (layer0_outputs(5057)) and not (layer0_outputs(4338));
    layer1_outputs(3668) <= not((layer0_outputs(18)) and (layer0_outputs(2756)));
    layer1_outputs(3669) <= not(layer0_outputs(3853)) or (layer0_outputs(3205));
    layer1_outputs(3670) <= '1';
    layer1_outputs(3671) <= layer0_outputs(2343);
    layer1_outputs(3672) <= (layer0_outputs(397)) and not (layer0_outputs(3444));
    layer1_outputs(3673) <= (layer0_outputs(1125)) and not (layer0_outputs(2729));
    layer1_outputs(3674) <= not(layer0_outputs(209));
    layer1_outputs(3675) <= not((layer0_outputs(1303)) or (layer0_outputs(2415)));
    layer1_outputs(3676) <= (layer0_outputs(4354)) and not (layer0_outputs(4255));
    layer1_outputs(3677) <= not((layer0_outputs(3500)) or (layer0_outputs(1975)));
    layer1_outputs(3678) <= not(layer0_outputs(4028));
    layer1_outputs(3679) <= layer0_outputs(720);
    layer1_outputs(3680) <= not(layer0_outputs(1308));
    layer1_outputs(3681) <= layer0_outputs(4887);
    layer1_outputs(3682) <= not(layer0_outputs(843)) or (layer0_outputs(3046));
    layer1_outputs(3683) <= not(layer0_outputs(1609)) or (layer0_outputs(1544));
    layer1_outputs(3684) <= (layer0_outputs(3164)) or (layer0_outputs(2196));
    layer1_outputs(3685) <= not((layer0_outputs(4610)) xor (layer0_outputs(863)));
    layer1_outputs(3686) <= layer0_outputs(3692);
    layer1_outputs(3687) <= (layer0_outputs(2879)) and (layer0_outputs(4304));
    layer1_outputs(3688) <= not((layer0_outputs(1448)) and (layer0_outputs(970)));
    layer1_outputs(3689) <= not(layer0_outputs(4827));
    layer1_outputs(3690) <= layer0_outputs(3586);
    layer1_outputs(3691) <= not(layer0_outputs(1479)) or (layer0_outputs(1337));
    layer1_outputs(3692) <= not(layer0_outputs(3079));
    layer1_outputs(3693) <= layer0_outputs(3275);
    layer1_outputs(3694) <= not(layer0_outputs(271));
    layer1_outputs(3695) <= (layer0_outputs(1383)) and (layer0_outputs(1367));
    layer1_outputs(3696) <= layer0_outputs(3628);
    layer1_outputs(3697) <= not((layer0_outputs(712)) xor (layer0_outputs(2536)));
    layer1_outputs(3698) <= (layer0_outputs(2955)) or (layer0_outputs(3592));
    layer1_outputs(3699) <= layer0_outputs(1762);
    layer1_outputs(3700) <= (layer0_outputs(4648)) and (layer0_outputs(818));
    layer1_outputs(3701) <= '1';
    layer1_outputs(3702) <= not((layer0_outputs(55)) or (layer0_outputs(4373)));
    layer1_outputs(3703) <= not((layer0_outputs(1471)) or (layer0_outputs(1691)));
    layer1_outputs(3704) <= layer0_outputs(2134);
    layer1_outputs(3705) <= not(layer0_outputs(1520));
    layer1_outputs(3706) <= not((layer0_outputs(2618)) xor (layer0_outputs(3146)));
    layer1_outputs(3707) <= (layer0_outputs(3496)) and (layer0_outputs(1512));
    layer1_outputs(3708) <= (layer0_outputs(3258)) or (layer0_outputs(3426));
    layer1_outputs(3709) <= not(layer0_outputs(4660));
    layer1_outputs(3710) <= (layer0_outputs(1585)) and not (layer0_outputs(4879));
    layer1_outputs(3711) <= (layer0_outputs(1879)) or (layer0_outputs(3718));
    layer1_outputs(3712) <= layer0_outputs(3974);
    layer1_outputs(3713) <= not(layer0_outputs(625)) or (layer0_outputs(2015));
    layer1_outputs(3714) <= not(layer0_outputs(8));
    layer1_outputs(3715) <= not((layer0_outputs(1944)) or (layer0_outputs(4715)));
    layer1_outputs(3716) <= not(layer0_outputs(3106));
    layer1_outputs(3717) <= (layer0_outputs(4928)) or (layer0_outputs(788));
    layer1_outputs(3718) <= not(layer0_outputs(5093));
    layer1_outputs(3719) <= layer0_outputs(2998);
    layer1_outputs(3720) <= not(layer0_outputs(4883));
    layer1_outputs(3721) <= not(layer0_outputs(2303));
    layer1_outputs(3722) <= not(layer0_outputs(5010)) or (layer0_outputs(981));
    layer1_outputs(3723) <= not((layer0_outputs(3286)) and (layer0_outputs(4437)));
    layer1_outputs(3724) <= not((layer0_outputs(3315)) and (layer0_outputs(1555)));
    layer1_outputs(3725) <= '0';
    layer1_outputs(3726) <= not(layer0_outputs(4010)) or (layer0_outputs(3497));
    layer1_outputs(3727) <= not(layer0_outputs(4570));
    layer1_outputs(3728) <= layer0_outputs(2496);
    layer1_outputs(3729) <= layer0_outputs(4947);
    layer1_outputs(3730) <= (layer0_outputs(215)) and (layer0_outputs(438));
    layer1_outputs(3731) <= (layer0_outputs(3442)) and not (layer0_outputs(1513));
    layer1_outputs(3732) <= (layer0_outputs(3368)) xor (layer0_outputs(1836));
    layer1_outputs(3733) <= '0';
    layer1_outputs(3734) <= (layer0_outputs(4098)) and (layer0_outputs(3638));
    layer1_outputs(3735) <= layer0_outputs(797);
    layer1_outputs(3736) <= not((layer0_outputs(3011)) or (layer0_outputs(1083)));
    layer1_outputs(3737) <= (layer0_outputs(2174)) or (layer0_outputs(4321));
    layer1_outputs(3738) <= (layer0_outputs(1231)) and not (layer0_outputs(3195));
    layer1_outputs(3739) <= layer0_outputs(4061);
    layer1_outputs(3740) <= not((layer0_outputs(3304)) and (layer0_outputs(4252)));
    layer1_outputs(3741) <= not((layer0_outputs(3717)) and (layer0_outputs(639)));
    layer1_outputs(3742) <= not((layer0_outputs(2533)) and (layer0_outputs(645)));
    layer1_outputs(3743) <= not((layer0_outputs(4762)) or (layer0_outputs(2653)));
    layer1_outputs(3744) <= layer0_outputs(702);
    layer1_outputs(3745) <= (layer0_outputs(4980)) and not (layer0_outputs(4858));
    layer1_outputs(3746) <= (layer0_outputs(1923)) and (layer0_outputs(2209));
    layer1_outputs(3747) <= not(layer0_outputs(926));
    layer1_outputs(3748) <= not(layer0_outputs(2823));
    layer1_outputs(3749) <= layer0_outputs(2711);
    layer1_outputs(3750) <= not(layer0_outputs(5023)) or (layer0_outputs(2570));
    layer1_outputs(3751) <= not((layer0_outputs(2576)) and (layer0_outputs(1671)));
    layer1_outputs(3752) <= not((layer0_outputs(4941)) or (layer0_outputs(4456)));
    layer1_outputs(3753) <= (layer0_outputs(1091)) and not (layer0_outputs(3944));
    layer1_outputs(3754) <= (layer0_outputs(2494)) or (layer0_outputs(226));
    layer1_outputs(3755) <= not(layer0_outputs(3273)) or (layer0_outputs(3330));
    layer1_outputs(3756) <= not(layer0_outputs(3162));
    layer1_outputs(3757) <= (layer0_outputs(3793)) or (layer0_outputs(3824));
    layer1_outputs(3758) <= layer0_outputs(987);
    layer1_outputs(3759) <= (layer0_outputs(1407)) and not (layer0_outputs(5098));
    layer1_outputs(3760) <= not((layer0_outputs(4759)) or (layer0_outputs(2713)));
    layer1_outputs(3761) <= not(layer0_outputs(4750));
    layer1_outputs(3762) <= (layer0_outputs(2194)) and not (layer0_outputs(2242));
    layer1_outputs(3763) <= not(layer0_outputs(3750));
    layer1_outputs(3764) <= '1';
    layer1_outputs(3765) <= (layer0_outputs(4361)) and not (layer0_outputs(370));
    layer1_outputs(3766) <= (layer0_outputs(3988)) and not (layer0_outputs(2389));
    layer1_outputs(3767) <= not(layer0_outputs(1551));
    layer1_outputs(3768) <= (layer0_outputs(432)) or (layer0_outputs(2029));
    layer1_outputs(3769) <= (layer0_outputs(431)) and (layer0_outputs(881));
    layer1_outputs(3770) <= (layer0_outputs(4626)) and (layer0_outputs(2354));
    layer1_outputs(3771) <= (layer0_outputs(2766)) and not (layer0_outputs(3032));
    layer1_outputs(3772) <= (layer0_outputs(4210)) and not (layer0_outputs(4700));
    layer1_outputs(3773) <= not((layer0_outputs(4319)) or (layer0_outputs(887)));
    layer1_outputs(3774) <= not(layer0_outputs(1422)) or (layer0_outputs(3153));
    layer1_outputs(3775) <= layer0_outputs(826);
    layer1_outputs(3776) <= not(layer0_outputs(4417));
    layer1_outputs(3777) <= '0';
    layer1_outputs(3778) <= layer0_outputs(2308);
    layer1_outputs(3779) <= not(layer0_outputs(3583));
    layer1_outputs(3780) <= (layer0_outputs(982)) and not (layer0_outputs(1211));
    layer1_outputs(3781) <= (layer0_outputs(534)) and not (layer0_outputs(3066));
    layer1_outputs(3782) <= not(layer0_outputs(4541)) or (layer0_outputs(1557));
    layer1_outputs(3783) <= layer0_outputs(3256);
    layer1_outputs(3784) <= not((layer0_outputs(4467)) or (layer0_outputs(286)));
    layer1_outputs(3785) <= not(layer0_outputs(166)) or (layer0_outputs(4460));
    layer1_outputs(3786) <= not(layer0_outputs(2856));
    layer1_outputs(3787) <= layer0_outputs(1818);
    layer1_outputs(3788) <= not(layer0_outputs(1179)) or (layer0_outputs(1532));
    layer1_outputs(3789) <= (layer0_outputs(2948)) and not (layer0_outputs(89));
    layer1_outputs(3790) <= (layer0_outputs(479)) and not (layer0_outputs(2581));
    layer1_outputs(3791) <= not(layer0_outputs(1968)) or (layer0_outputs(15));
    layer1_outputs(3792) <= (layer0_outputs(2068)) and not (layer0_outputs(2083));
    layer1_outputs(3793) <= not(layer0_outputs(1736)) or (layer0_outputs(3069));
    layer1_outputs(3794) <= (layer0_outputs(5036)) and not (layer0_outputs(847));
    layer1_outputs(3795) <= (layer0_outputs(2228)) and not (layer0_outputs(4448));
    layer1_outputs(3796) <= not(layer0_outputs(4400)) or (layer0_outputs(2839));
    layer1_outputs(3797) <= not(layer0_outputs(474)) or (layer0_outputs(4137));
    layer1_outputs(3798) <= (layer0_outputs(2062)) or (layer0_outputs(2606));
    layer1_outputs(3799) <= (layer0_outputs(386)) or (layer0_outputs(721));
    layer1_outputs(3800) <= not(layer0_outputs(3202));
    layer1_outputs(3801) <= not(layer0_outputs(3515));
    layer1_outputs(3802) <= (layer0_outputs(354)) and not (layer0_outputs(1913));
    layer1_outputs(3803) <= not((layer0_outputs(2725)) or (layer0_outputs(389)));
    layer1_outputs(3804) <= '0';
    layer1_outputs(3805) <= '0';
    layer1_outputs(3806) <= (layer0_outputs(3334)) and not (layer0_outputs(3316));
    layer1_outputs(3807) <= (layer0_outputs(4084)) or (layer0_outputs(2081));
    layer1_outputs(3808) <= (layer0_outputs(3198)) and (layer0_outputs(2377));
    layer1_outputs(3809) <= (layer0_outputs(3071)) or (layer0_outputs(1840));
    layer1_outputs(3810) <= not(layer0_outputs(997)) or (layer0_outputs(339));
    layer1_outputs(3811) <= layer0_outputs(480);
    layer1_outputs(3812) <= layer0_outputs(4844);
    layer1_outputs(3813) <= (layer0_outputs(1472)) and not (layer0_outputs(253));
    layer1_outputs(3814) <= layer0_outputs(325);
    layer1_outputs(3815) <= not(layer0_outputs(2512));
    layer1_outputs(3816) <= not(layer0_outputs(1107));
    layer1_outputs(3817) <= not(layer0_outputs(355)) or (layer0_outputs(1033));
    layer1_outputs(3818) <= (layer0_outputs(3171)) and not (layer0_outputs(2072));
    layer1_outputs(3819) <= layer0_outputs(2545);
    layer1_outputs(3820) <= not(layer0_outputs(3056)) or (layer0_outputs(2082));
    layer1_outputs(3821) <= (layer0_outputs(875)) or (layer0_outputs(4911));
    layer1_outputs(3822) <= (layer0_outputs(4617)) and not (layer0_outputs(1484));
    layer1_outputs(3823) <= layer0_outputs(4017);
    layer1_outputs(3824) <= (layer0_outputs(4938)) and not (layer0_outputs(815));
    layer1_outputs(3825) <= layer0_outputs(2246);
    layer1_outputs(3826) <= not((layer0_outputs(1196)) and (layer0_outputs(2510)));
    layer1_outputs(3827) <= layer0_outputs(2888);
    layer1_outputs(3828) <= not((layer0_outputs(3506)) and (layer0_outputs(3655)));
    layer1_outputs(3829) <= not((layer0_outputs(1919)) xor (layer0_outputs(4656)));
    layer1_outputs(3830) <= (layer0_outputs(656)) and not (layer0_outputs(1223));
    layer1_outputs(3831) <= layer0_outputs(2338);
    layer1_outputs(3832) <= not(layer0_outputs(628));
    layer1_outputs(3833) <= not(layer0_outputs(725));
    layer1_outputs(3834) <= not(layer0_outputs(3409)) or (layer0_outputs(3475));
    layer1_outputs(3835) <= not(layer0_outputs(1214));
    layer1_outputs(3836) <= not(layer0_outputs(3848)) or (layer0_outputs(3976));
    layer1_outputs(3837) <= not((layer0_outputs(3878)) xor (layer0_outputs(1034)));
    layer1_outputs(3838) <= (layer0_outputs(4214)) and not (layer0_outputs(440));
    layer1_outputs(3839) <= not(layer0_outputs(376));
    layer1_outputs(3840) <= not(layer0_outputs(1500));
    layer1_outputs(3841) <= '0';
    layer1_outputs(3842) <= not((layer0_outputs(2397)) or (layer0_outputs(4153)));
    layer1_outputs(3843) <= (layer0_outputs(3381)) and (layer0_outputs(3121));
    layer1_outputs(3844) <= (layer0_outputs(3534)) and (layer0_outputs(2894));
    layer1_outputs(3845) <= layer0_outputs(4584);
    layer1_outputs(3846) <= not(layer0_outputs(1613));
    layer1_outputs(3847) <= not(layer0_outputs(3405)) or (layer0_outputs(4667));
    layer1_outputs(3848) <= not(layer0_outputs(2795));
    layer1_outputs(3849) <= not((layer0_outputs(1418)) or (layer0_outputs(3246)));
    layer1_outputs(3850) <= '1';
    layer1_outputs(3851) <= not((layer0_outputs(814)) or (layer0_outputs(2829)));
    layer1_outputs(3852) <= layer0_outputs(1599);
    layer1_outputs(3853) <= layer0_outputs(3163);
    layer1_outputs(3854) <= not(layer0_outputs(2345)) or (layer0_outputs(723));
    layer1_outputs(3855) <= layer0_outputs(2640);
    layer1_outputs(3856) <= not((layer0_outputs(2020)) or (layer0_outputs(2753)));
    layer1_outputs(3857) <= (layer0_outputs(4341)) or (layer0_outputs(3605));
    layer1_outputs(3858) <= (layer0_outputs(5068)) and not (layer0_outputs(2531));
    layer1_outputs(3859) <= layer0_outputs(3105);
    layer1_outputs(3860) <= not(layer0_outputs(4964));
    layer1_outputs(3861) <= layer0_outputs(4124);
    layer1_outputs(3862) <= (layer0_outputs(1099)) or (layer0_outputs(612));
    layer1_outputs(3863) <= not(layer0_outputs(2253)) or (layer0_outputs(75));
    layer1_outputs(3864) <= layer0_outputs(3031);
    layer1_outputs(3865) <= layer0_outputs(1463);
    layer1_outputs(3866) <= not((layer0_outputs(837)) or (layer0_outputs(2230)));
    layer1_outputs(3867) <= layer0_outputs(4597);
    layer1_outputs(3868) <= not(layer0_outputs(485));
    layer1_outputs(3869) <= not((layer0_outputs(2943)) or (layer0_outputs(4500)));
    layer1_outputs(3870) <= not(layer0_outputs(2833));
    layer1_outputs(3871) <= (layer0_outputs(2321)) or (layer0_outputs(3026));
    layer1_outputs(3872) <= not(layer0_outputs(3274));
    layer1_outputs(3873) <= (layer0_outputs(287)) and not (layer0_outputs(5094));
    layer1_outputs(3874) <= not(layer0_outputs(3268));
    layer1_outputs(3875) <= not(layer0_outputs(826));
    layer1_outputs(3876) <= not(layer0_outputs(21)) or (layer0_outputs(1229));
    layer1_outputs(3877) <= not(layer0_outputs(334));
    layer1_outputs(3878) <= not((layer0_outputs(1315)) or (layer0_outputs(984)));
    layer1_outputs(3879) <= (layer0_outputs(2502)) and (layer0_outputs(4476));
    layer1_outputs(3880) <= layer0_outputs(3212);
    layer1_outputs(3881) <= layer0_outputs(815);
    layer1_outputs(3882) <= not((layer0_outputs(2614)) and (layer0_outputs(1730)));
    layer1_outputs(3883) <= not((layer0_outputs(1779)) or (layer0_outputs(47)));
    layer1_outputs(3884) <= not(layer0_outputs(3460)) or (layer0_outputs(2992));
    layer1_outputs(3885) <= not(layer0_outputs(1745));
    layer1_outputs(3886) <= (layer0_outputs(4708)) and (layer0_outputs(2053));
    layer1_outputs(3887) <= not(layer0_outputs(3350)) or (layer0_outputs(4853));
    layer1_outputs(3888) <= not(layer0_outputs(1365)) or (layer0_outputs(4329));
    layer1_outputs(3889) <= layer0_outputs(4846);
    layer1_outputs(3890) <= layer0_outputs(1064);
    layer1_outputs(3891) <= layer0_outputs(1771);
    layer1_outputs(3892) <= (layer0_outputs(4755)) and not (layer0_outputs(1999));
    layer1_outputs(3893) <= (layer0_outputs(3072)) or (layer0_outputs(3419));
    layer1_outputs(3894) <= layer0_outputs(276);
    layer1_outputs(3895) <= layer0_outputs(589);
    layer1_outputs(3896) <= (layer0_outputs(2700)) and not (layer0_outputs(4757));
    layer1_outputs(3897) <= not(layer0_outputs(3553));
    layer1_outputs(3898) <= not(layer0_outputs(4734));
    layer1_outputs(3899) <= '1';
    layer1_outputs(3900) <= not(layer0_outputs(2514));
    layer1_outputs(3901) <= (layer0_outputs(4439)) and not (layer0_outputs(3078));
    layer1_outputs(3902) <= '1';
    layer1_outputs(3903) <= not(layer0_outputs(1894));
    layer1_outputs(3904) <= not(layer0_outputs(238));
    layer1_outputs(3905) <= not(layer0_outputs(314)) or (layer0_outputs(393));
    layer1_outputs(3906) <= layer0_outputs(4416);
    layer1_outputs(3907) <= (layer0_outputs(4592)) and (layer0_outputs(1600));
    layer1_outputs(3908) <= (layer0_outputs(1678)) and (layer0_outputs(3431));
    layer1_outputs(3909) <= not(layer0_outputs(3005));
    layer1_outputs(3910) <= not(layer0_outputs(4408));
    layer1_outputs(3911) <= layer0_outputs(876);
    layer1_outputs(3912) <= '0';
    layer1_outputs(3913) <= (layer0_outputs(1802)) xor (layer0_outputs(1643));
    layer1_outputs(3914) <= layer0_outputs(3599);
    layer1_outputs(3915) <= not(layer0_outputs(1503));
    layer1_outputs(3916) <= layer0_outputs(1669);
    layer1_outputs(3917) <= not(layer0_outputs(3545)) or (layer0_outputs(4655));
    layer1_outputs(3918) <= '0';
    layer1_outputs(3919) <= layer0_outputs(1171);
    layer1_outputs(3920) <= not(layer0_outputs(4809));
    layer1_outputs(3921) <= not((layer0_outputs(4126)) or (layer0_outputs(914)));
    layer1_outputs(3922) <= not((layer0_outputs(3803)) xor (layer0_outputs(2995)));
    layer1_outputs(3923) <= layer0_outputs(1549);
    layer1_outputs(3924) <= not(layer0_outputs(1492));
    layer1_outputs(3925) <= not(layer0_outputs(3871)) or (layer0_outputs(2166));
    layer1_outputs(3926) <= not(layer0_outputs(806)) or (layer0_outputs(4909));
    layer1_outputs(3927) <= (layer0_outputs(1356)) xor (layer0_outputs(1514));
    layer1_outputs(3928) <= (layer0_outputs(4669)) or (layer0_outputs(2749));
    layer1_outputs(3929) <= not(layer0_outputs(3882)) or (layer0_outputs(1917));
    layer1_outputs(3930) <= not((layer0_outputs(4773)) and (layer0_outputs(2489)));
    layer1_outputs(3931) <= layer0_outputs(4824);
    layer1_outputs(3932) <= not((layer0_outputs(100)) and (layer0_outputs(1246)));
    layer1_outputs(3933) <= layer0_outputs(4681);
    layer1_outputs(3934) <= '1';
    layer1_outputs(3935) <= not(layer0_outputs(3707));
    layer1_outputs(3936) <= not(layer0_outputs(859));
    layer1_outputs(3937) <= layer0_outputs(1203);
    layer1_outputs(3938) <= not(layer0_outputs(552)) or (layer0_outputs(1654));
    layer1_outputs(3939) <= not((layer0_outputs(3553)) xor (layer0_outputs(3986)));
    layer1_outputs(3940) <= (layer0_outputs(2603)) and not (layer0_outputs(3912));
    layer1_outputs(3941) <= not(layer0_outputs(3131));
    layer1_outputs(3942) <= not(layer0_outputs(2155));
    layer1_outputs(3943) <= layer0_outputs(1084);
    layer1_outputs(3944) <= layer0_outputs(4634);
    layer1_outputs(3945) <= not(layer0_outputs(1395)) or (layer0_outputs(4953));
    layer1_outputs(3946) <= (layer0_outputs(3889)) and (layer0_outputs(3772));
    layer1_outputs(3947) <= not(layer0_outputs(1566));
    layer1_outputs(3948) <= not((layer0_outputs(1137)) or (layer0_outputs(625)));
    layer1_outputs(3949) <= '0';
    layer1_outputs(3950) <= not(layer0_outputs(1502)) or (layer0_outputs(3088));
    layer1_outputs(3951) <= (layer0_outputs(4080)) and (layer0_outputs(1689));
    layer1_outputs(3952) <= not(layer0_outputs(172));
    layer1_outputs(3953) <= not(layer0_outputs(1044)) or (layer0_outputs(524));
    layer1_outputs(3954) <= not(layer0_outputs(4106));
    layer1_outputs(3955) <= not(layer0_outputs(2005));
    layer1_outputs(3956) <= not(layer0_outputs(864));
    layer1_outputs(3957) <= not((layer0_outputs(4934)) xor (layer0_outputs(336)));
    layer1_outputs(3958) <= not((layer0_outputs(2954)) or (layer0_outputs(3437)));
    layer1_outputs(3959) <= not((layer0_outputs(1831)) xor (layer0_outputs(1911)));
    layer1_outputs(3960) <= not((layer0_outputs(1245)) or (layer0_outputs(3965)));
    layer1_outputs(3961) <= not(layer0_outputs(3905));
    layer1_outputs(3962) <= not(layer0_outputs(4495)) or (layer0_outputs(3322));
    layer1_outputs(3963) <= not(layer0_outputs(3967)) or (layer0_outputs(3372));
    layer1_outputs(3964) <= layer0_outputs(3309);
    layer1_outputs(3965) <= not(layer0_outputs(4536));
    layer1_outputs(3966) <= not(layer0_outputs(3440)) or (layer0_outputs(2314));
    layer1_outputs(3967) <= (layer0_outputs(365)) xor (layer0_outputs(2803));
    layer1_outputs(3968) <= not(layer0_outputs(2743));
    layer1_outputs(3969) <= not(layer0_outputs(3780)) or (layer0_outputs(136));
    layer1_outputs(3970) <= layer0_outputs(4259);
    layer1_outputs(3971) <= (layer0_outputs(1470)) and not (layer0_outputs(1681));
    layer1_outputs(3972) <= not((layer0_outputs(999)) and (layer0_outputs(858)));
    layer1_outputs(3973) <= not(layer0_outputs(4828));
    layer1_outputs(3974) <= (layer0_outputs(1049)) and not (layer0_outputs(4257));
    layer1_outputs(3975) <= not(layer0_outputs(391)) or (layer0_outputs(4437));
    layer1_outputs(3976) <= '1';
    layer1_outputs(3977) <= layer0_outputs(3817);
    layer1_outputs(3978) <= (layer0_outputs(122)) xor (layer0_outputs(739));
    layer1_outputs(3979) <= layer0_outputs(4734);
    layer1_outputs(3980) <= not(layer0_outputs(4851));
    layer1_outputs(3981) <= not(layer0_outputs(1536)) or (layer0_outputs(5113));
    layer1_outputs(3982) <= not(layer0_outputs(220));
    layer1_outputs(3983) <= not(layer0_outputs(691));
    layer1_outputs(3984) <= (layer0_outputs(57)) xor (layer0_outputs(1620));
    layer1_outputs(3985) <= not(layer0_outputs(2690));
    layer1_outputs(3986) <= not((layer0_outputs(4915)) and (layer0_outputs(2628)));
    layer1_outputs(3987) <= layer0_outputs(4756);
    layer1_outputs(3988) <= not(layer0_outputs(4443)) or (layer0_outputs(1906));
    layer1_outputs(3989) <= layer0_outputs(4139);
    layer1_outputs(3990) <= not((layer0_outputs(2416)) xor (layer0_outputs(2929)));
    layer1_outputs(3991) <= (layer0_outputs(4560)) and not (layer0_outputs(1415));
    layer1_outputs(3992) <= (layer0_outputs(3027)) and not (layer0_outputs(1109));
    layer1_outputs(3993) <= layer0_outputs(4243);
    layer1_outputs(3994) <= (layer0_outputs(1259)) xor (layer0_outputs(4860));
    layer1_outputs(3995) <= layer0_outputs(773);
    layer1_outputs(3996) <= layer0_outputs(4120);
    layer1_outputs(3997) <= layer0_outputs(4821);
    layer1_outputs(3998) <= layer0_outputs(5063);
    layer1_outputs(3999) <= (layer0_outputs(1662)) and not (layer0_outputs(2261));
    layer1_outputs(4000) <= layer0_outputs(1826);
    layer1_outputs(4001) <= (layer0_outputs(4262)) and not (layer0_outputs(266));
    layer1_outputs(4002) <= layer0_outputs(1834);
    layer1_outputs(4003) <= layer0_outputs(2279);
    layer1_outputs(4004) <= (layer0_outputs(2662)) and (layer0_outputs(4215));
    layer1_outputs(4005) <= not(layer0_outputs(2669)) or (layer0_outputs(2320));
    layer1_outputs(4006) <= layer0_outputs(3494);
    layer1_outputs(4007) <= (layer0_outputs(4387)) and not (layer0_outputs(2291));
    layer1_outputs(4008) <= layer0_outputs(2925);
    layer1_outputs(4009) <= layer0_outputs(4055);
    layer1_outputs(4010) <= not((layer0_outputs(5077)) and (layer0_outputs(1115)));
    layer1_outputs(4011) <= '1';
    layer1_outputs(4012) <= '0';
    layer1_outputs(4013) <= (layer0_outputs(3339)) and not (layer0_outputs(991));
    layer1_outputs(4014) <= not(layer0_outputs(2629));
    layer1_outputs(4015) <= '0';
    layer1_outputs(4016) <= not((layer0_outputs(1091)) or (layer0_outputs(2027)));
    layer1_outputs(4017) <= layer0_outputs(1965);
    layer1_outputs(4018) <= '0';
    layer1_outputs(4019) <= '0';
    layer1_outputs(4020) <= layer0_outputs(3817);
    layer1_outputs(4021) <= not(layer0_outputs(3877));
    layer1_outputs(4022) <= '0';
    layer1_outputs(4023) <= not((layer0_outputs(4225)) and (layer0_outputs(321)));
    layer1_outputs(4024) <= not((layer0_outputs(4805)) and (layer0_outputs(1920)));
    layer1_outputs(4025) <= not(layer0_outputs(521)) or (layer0_outputs(3387));
    layer1_outputs(4026) <= '0';
    layer1_outputs(4027) <= not(layer0_outputs(3996)) or (layer0_outputs(5090));
    layer1_outputs(4028) <= layer0_outputs(3868);
    layer1_outputs(4029) <= (layer0_outputs(859)) xor (layer0_outputs(4493));
    layer1_outputs(4030) <= not((layer0_outputs(1733)) xor (layer0_outputs(4627)));
    layer1_outputs(4031) <= not(layer0_outputs(2475)) or (layer0_outputs(4144));
    layer1_outputs(4032) <= not(layer0_outputs(3936));
    layer1_outputs(4033) <= not((layer0_outputs(1595)) or (layer0_outputs(3388)));
    layer1_outputs(4034) <= not((layer0_outputs(4857)) xor (layer0_outputs(21)));
    layer1_outputs(4035) <= layer0_outputs(1078);
    layer1_outputs(4036) <= (layer0_outputs(1769)) and not (layer0_outputs(4431));
    layer1_outputs(4037) <= '0';
    layer1_outputs(4038) <= not(layer0_outputs(2630));
    layer1_outputs(4039) <= (layer0_outputs(2057)) and not (layer0_outputs(1813));
    layer1_outputs(4040) <= (layer0_outputs(5041)) and (layer0_outputs(1737));
    layer1_outputs(4041) <= (layer0_outputs(3134)) and (layer0_outputs(3870));
    layer1_outputs(4042) <= (layer0_outputs(3469)) or (layer0_outputs(3816));
    layer1_outputs(4043) <= not(layer0_outputs(3666)) or (layer0_outputs(1366));
    layer1_outputs(4044) <= not(layer0_outputs(674));
    layer1_outputs(4045) <= not(layer0_outputs(2400));
    layer1_outputs(4046) <= (layer0_outputs(1756)) or (layer0_outputs(2561));
    layer1_outputs(4047) <= (layer0_outputs(2659)) or (layer0_outputs(2677));
    layer1_outputs(4048) <= '0';
    layer1_outputs(4049) <= (layer0_outputs(3875)) and (layer0_outputs(3635));
    layer1_outputs(4050) <= layer0_outputs(1286);
    layer1_outputs(4051) <= layer0_outputs(3801);
    layer1_outputs(4052) <= (layer0_outputs(3211)) and not (layer0_outputs(1046));
    layer1_outputs(4053) <= (layer0_outputs(2712)) and (layer0_outputs(4524));
    layer1_outputs(4054) <= not(layer0_outputs(3479));
    layer1_outputs(4055) <= (layer0_outputs(2703)) and not (layer0_outputs(3364));
    layer1_outputs(4056) <= (layer0_outputs(3094)) and (layer0_outputs(3295));
    layer1_outputs(4057) <= not((layer0_outputs(1709)) and (layer0_outputs(1087)));
    layer1_outputs(4058) <= (layer0_outputs(457)) and not (layer0_outputs(3544));
    layer1_outputs(4059) <= not((layer0_outputs(1993)) and (layer0_outputs(2711)));
    layer1_outputs(4060) <= not(layer0_outputs(3270));
    layer1_outputs(4061) <= not((layer0_outputs(4446)) or (layer0_outputs(5021)));
    layer1_outputs(4062) <= '0';
    layer1_outputs(4063) <= not(layer0_outputs(2968)) or (layer0_outputs(2278));
    layer1_outputs(4064) <= (layer0_outputs(4230)) and not (layer0_outputs(2982));
    layer1_outputs(4065) <= (layer0_outputs(2587)) and not (layer0_outputs(2158));
    layer1_outputs(4066) <= (layer0_outputs(2489)) or (layer0_outputs(3147));
    layer1_outputs(4067) <= not(layer0_outputs(385)) or (layer0_outputs(2924));
    layer1_outputs(4068) <= not(layer0_outputs(559));
    layer1_outputs(4069) <= layer0_outputs(4137);
    layer1_outputs(4070) <= not(layer0_outputs(2152));
    layer1_outputs(4071) <= not(layer0_outputs(4271));
    layer1_outputs(4072) <= not(layer0_outputs(2367));
    layer1_outputs(4073) <= (layer0_outputs(2133)) and not (layer0_outputs(849));
    layer1_outputs(4074) <= (layer0_outputs(4614)) or (layer0_outputs(4463));
    layer1_outputs(4075) <= layer0_outputs(4422);
    layer1_outputs(4076) <= '0';
    layer1_outputs(4077) <= (layer0_outputs(364)) xor (layer0_outputs(1240));
    layer1_outputs(4078) <= not(layer0_outputs(4686));
    layer1_outputs(4079) <= not(layer0_outputs(4894)) or (layer0_outputs(4802));
    layer1_outputs(4080) <= (layer0_outputs(4993)) and not (layer0_outputs(4775));
    layer1_outputs(4081) <= not(layer0_outputs(1964));
    layer1_outputs(4082) <= not(layer0_outputs(1900)) or (layer0_outputs(390));
    layer1_outputs(4083) <= not(layer0_outputs(4114));
    layer1_outputs(4084) <= not(layer0_outputs(1307));
    layer1_outputs(4085) <= not(layer0_outputs(4241));
    layer1_outputs(4086) <= not((layer0_outputs(4836)) and (layer0_outputs(1131)));
    layer1_outputs(4087) <= not((layer0_outputs(2542)) and (layer0_outputs(4804)));
    layer1_outputs(4088) <= (layer0_outputs(4371)) or (layer0_outputs(3581));
    layer1_outputs(4089) <= not(layer0_outputs(1019));
    layer1_outputs(4090) <= not(layer0_outputs(3921));
    layer1_outputs(4091) <= (layer0_outputs(775)) or (layer0_outputs(1212));
    layer1_outputs(4092) <= not(layer0_outputs(3454));
    layer1_outputs(4093) <= not(layer0_outputs(1903));
    layer1_outputs(4094) <= layer0_outputs(3424);
    layer1_outputs(4095) <= not((layer0_outputs(3341)) or (layer0_outputs(5051)));
    layer1_outputs(4096) <= not((layer0_outputs(2517)) xor (layer0_outputs(1787)));
    layer1_outputs(4097) <= (layer0_outputs(1332)) and (layer0_outputs(3038));
    layer1_outputs(4098) <= layer0_outputs(4805);
    layer1_outputs(4099) <= not(layer0_outputs(4095)) or (layer0_outputs(3295));
    layer1_outputs(4100) <= not((layer0_outputs(3213)) and (layer0_outputs(4134)));
    layer1_outputs(4101) <= not(layer0_outputs(1102)) or (layer0_outputs(644));
    layer1_outputs(4102) <= (layer0_outputs(292)) and (layer0_outputs(5062));
    layer1_outputs(4103) <= not((layer0_outputs(730)) and (layer0_outputs(4147)));
    layer1_outputs(4104) <= layer0_outputs(1819);
    layer1_outputs(4105) <= (layer0_outputs(1570)) xor (layer0_outputs(350));
    layer1_outputs(4106) <= (layer0_outputs(597)) and not (layer0_outputs(4030));
    layer1_outputs(4107) <= layer0_outputs(2535);
    layer1_outputs(4108) <= layer0_outputs(3649);
    layer1_outputs(4109) <= (layer0_outputs(4108)) and not (layer0_outputs(235));
    layer1_outputs(4110) <= (layer0_outputs(528)) and (layer0_outputs(1138));
    layer1_outputs(4111) <= (layer0_outputs(2146)) or (layer0_outputs(880));
    layer1_outputs(4112) <= not((layer0_outputs(1582)) and (layer0_outputs(4838)));
    layer1_outputs(4113) <= (layer0_outputs(5027)) and not (layer0_outputs(1431));
    layer1_outputs(4114) <= layer0_outputs(1988);
    layer1_outputs(4115) <= (layer0_outputs(915)) and (layer0_outputs(3351));
    layer1_outputs(4116) <= not(layer0_outputs(2679)) or (layer0_outputs(1358));
    layer1_outputs(4117) <= (layer0_outputs(3849)) and not (layer0_outputs(146));
    layer1_outputs(4118) <= not(layer0_outputs(2790));
    layer1_outputs(4119) <= (layer0_outputs(4056)) or (layer0_outputs(16));
    layer1_outputs(4120) <= not((layer0_outputs(1112)) and (layer0_outputs(1401)));
    layer1_outputs(4121) <= layer0_outputs(3554);
    layer1_outputs(4122) <= layer0_outputs(3392);
    layer1_outputs(4123) <= layer0_outputs(1507);
    layer1_outputs(4124) <= (layer0_outputs(348)) or (layer0_outputs(3602));
    layer1_outputs(4125) <= not(layer0_outputs(3958));
    layer1_outputs(4126) <= not(layer0_outputs(3615));
    layer1_outputs(4127) <= not(layer0_outputs(4764));
    layer1_outputs(4128) <= not((layer0_outputs(4978)) or (layer0_outputs(1277)));
    layer1_outputs(4129) <= layer0_outputs(4832);
    layer1_outputs(4130) <= (layer0_outputs(2828)) xor (layer0_outputs(1488));
    layer1_outputs(4131) <= not(layer0_outputs(4885)) or (layer0_outputs(262));
    layer1_outputs(4132) <= layer0_outputs(1936);
    layer1_outputs(4133) <= not(layer0_outputs(3227)) or (layer0_outputs(2830));
    layer1_outputs(4134) <= (layer0_outputs(858)) and (layer0_outputs(2957));
    layer1_outputs(4135) <= not(layer0_outputs(2551)) or (layer0_outputs(5011));
    layer1_outputs(4136) <= not((layer0_outputs(4394)) and (layer0_outputs(1031)));
    layer1_outputs(4137) <= not(layer0_outputs(1580));
    layer1_outputs(4138) <= (layer0_outputs(4018)) or (layer0_outputs(1511));
    layer1_outputs(4139) <= not(layer0_outputs(229));
    layer1_outputs(4140) <= not(layer0_outputs(1205));
    layer1_outputs(4141) <= not(layer0_outputs(2885));
    layer1_outputs(4142) <= layer0_outputs(5118);
    layer1_outputs(4143) <= not(layer0_outputs(2806));
    layer1_outputs(4144) <= not(layer0_outputs(1510)) or (layer0_outputs(3786));
    layer1_outputs(4145) <= (layer0_outputs(175)) and not (layer0_outputs(1645));
    layer1_outputs(4146) <= layer0_outputs(4085);
    layer1_outputs(4147) <= layer0_outputs(1605);
    layer1_outputs(4148) <= not(layer0_outputs(4582));
    layer1_outputs(4149) <= not(layer0_outputs(3463));
    layer1_outputs(4150) <= layer0_outputs(4282);
    layer1_outputs(4151) <= '0';
    layer1_outputs(4152) <= layer0_outputs(251);
    layer1_outputs(4153) <= '1';
    layer1_outputs(4154) <= (layer0_outputs(785)) or (layer0_outputs(944));
    layer1_outputs(4155) <= not((layer0_outputs(3792)) and (layer0_outputs(2182)));
    layer1_outputs(4156) <= (layer0_outputs(2289)) and not (layer0_outputs(3959));
    layer1_outputs(4157) <= not(layer0_outputs(4804));
    layer1_outputs(4158) <= not(layer0_outputs(3746));
    layer1_outputs(4159) <= not(layer0_outputs(4889));
    layer1_outputs(4160) <= layer0_outputs(965);
    layer1_outputs(4161) <= not(layer0_outputs(440)) or (layer0_outputs(4916));
    layer1_outputs(4162) <= not(layer0_outputs(3115));
    layer1_outputs(4163) <= not((layer0_outputs(2113)) and (layer0_outputs(2109)));
    layer1_outputs(4164) <= layer0_outputs(1957);
    layer1_outputs(4165) <= layer0_outputs(2471);
    layer1_outputs(4166) <= (layer0_outputs(1083)) and (layer0_outputs(2207));
    layer1_outputs(4167) <= (layer0_outputs(1680)) and not (layer0_outputs(945));
    layer1_outputs(4168) <= (layer0_outputs(3452)) and not (layer0_outputs(1226));
    layer1_outputs(4169) <= (layer0_outputs(1774)) and not (layer0_outputs(2318));
    layer1_outputs(4170) <= not(layer0_outputs(410));
    layer1_outputs(4171) <= (layer0_outputs(1176)) and not (layer0_outputs(4043));
    layer1_outputs(4172) <= layer0_outputs(3149);
    layer1_outputs(4173) <= not((layer0_outputs(4598)) xor (layer0_outputs(3814)));
    layer1_outputs(4174) <= not(layer0_outputs(1143));
    layer1_outputs(4175) <= (layer0_outputs(3386)) or (layer0_outputs(3032));
    layer1_outputs(4176) <= (layer0_outputs(2394)) or (layer0_outputs(2296));
    layer1_outputs(4177) <= layer0_outputs(4777);
    layer1_outputs(4178) <= not(layer0_outputs(1162));
    layer1_outputs(4179) <= not(layer0_outputs(62));
    layer1_outputs(4180) <= '1';
    layer1_outputs(4181) <= not((layer0_outputs(2925)) and (layer0_outputs(2921)));
    layer1_outputs(4182) <= not((layer0_outputs(4826)) xor (layer0_outputs(2148)));
    layer1_outputs(4183) <= not(layer0_outputs(1808));
    layer1_outputs(4184) <= (layer0_outputs(2697)) xor (layer0_outputs(2077));
    layer1_outputs(4185) <= not(layer0_outputs(4187));
    layer1_outputs(4186) <= layer0_outputs(1006);
    layer1_outputs(4187) <= not(layer0_outputs(2666));
    layer1_outputs(4188) <= not(layer0_outputs(4477));
    layer1_outputs(4189) <= not(layer0_outputs(953));
    layer1_outputs(4190) <= not((layer0_outputs(765)) or (layer0_outputs(3528)));
    layer1_outputs(4191) <= not(layer0_outputs(2140));
    layer1_outputs(4192) <= not(layer0_outputs(2245));
    layer1_outputs(4193) <= not(layer0_outputs(3345));
    layer1_outputs(4194) <= layer0_outputs(4649);
    layer1_outputs(4195) <= layer0_outputs(987);
    layer1_outputs(4196) <= '1';
    layer1_outputs(4197) <= layer0_outputs(516);
    layer1_outputs(4198) <= (layer0_outputs(3805)) or (layer0_outputs(3842));
    layer1_outputs(4199) <= layer0_outputs(4224);
    layer1_outputs(4200) <= (layer0_outputs(1493)) and (layer0_outputs(2782));
    layer1_outputs(4201) <= not(layer0_outputs(4221)) or (layer0_outputs(443));
    layer1_outputs(4202) <= (layer0_outputs(4652)) and (layer0_outputs(3293));
    layer1_outputs(4203) <= not(layer0_outputs(2996));
    layer1_outputs(4204) <= layer0_outputs(4539);
    layer1_outputs(4205) <= not((layer0_outputs(1588)) and (layer0_outputs(2827)));
    layer1_outputs(4206) <= layer0_outputs(4202);
    layer1_outputs(4207) <= (layer0_outputs(1066)) and not (layer0_outputs(3275));
    layer1_outputs(4208) <= (layer0_outputs(3335)) and (layer0_outputs(1036));
    layer1_outputs(4209) <= not((layer0_outputs(5083)) and (layer0_outputs(1168)));
    layer1_outputs(4210) <= (layer0_outputs(4639)) or (layer0_outputs(153));
    layer1_outputs(4211) <= not(layer0_outputs(1434));
    layer1_outputs(4212) <= layer0_outputs(4726);
    layer1_outputs(4213) <= layer0_outputs(4540);
    layer1_outputs(4214) <= not((layer0_outputs(3407)) or (layer0_outputs(2389)));
    layer1_outputs(4215) <= layer0_outputs(707);
    layer1_outputs(4216) <= (layer0_outputs(924)) and (layer0_outputs(3385));
    layer1_outputs(4217) <= not(layer0_outputs(4535));
    layer1_outputs(4218) <= not(layer0_outputs(3246)) or (layer0_outputs(2061));
    layer1_outputs(4219) <= not((layer0_outputs(1368)) or (layer0_outputs(4988)));
    layer1_outputs(4220) <= layer0_outputs(504);
    layer1_outputs(4221) <= not(layer0_outputs(256));
    layer1_outputs(4222) <= layer0_outputs(2708);
    layer1_outputs(4223) <= layer0_outputs(2015);
    layer1_outputs(4224) <= (layer0_outputs(2243)) xor (layer0_outputs(3659));
    layer1_outputs(4225) <= not(layer0_outputs(1614)) or (layer0_outputs(4881));
    layer1_outputs(4226) <= layer0_outputs(430);
    layer1_outputs(4227) <= (layer0_outputs(1844)) or (layer0_outputs(2012));
    layer1_outputs(4228) <= layer0_outputs(4520);
    layer1_outputs(4229) <= layer0_outputs(2849);
    layer1_outputs(4230) <= layer0_outputs(3551);
    layer1_outputs(4231) <= (layer0_outputs(4074)) and not (layer0_outputs(1785));
    layer1_outputs(4232) <= (layer0_outputs(2730)) and not (layer0_outputs(4399));
    layer1_outputs(4233) <= not(layer0_outputs(1040));
    layer1_outputs(4234) <= not((layer0_outputs(1899)) and (layer0_outputs(682)));
    layer1_outputs(4235) <= (layer0_outputs(624)) and not (layer0_outputs(408));
    layer1_outputs(4236) <= not((layer0_outputs(3331)) or (layer0_outputs(3987)));
    layer1_outputs(4237) <= layer0_outputs(3128);
    layer1_outputs(4238) <= (layer0_outputs(781)) or (layer0_outputs(1465));
    layer1_outputs(4239) <= layer0_outputs(4105);
    layer1_outputs(4240) <= layer0_outputs(106);
    layer1_outputs(4241) <= (layer0_outputs(4670)) xor (layer0_outputs(3628));
    layer1_outputs(4242) <= not(layer0_outputs(3972)) or (layer0_outputs(70));
    layer1_outputs(4243) <= (layer0_outputs(2546)) or (layer0_outputs(3317));
    layer1_outputs(4244) <= not((layer0_outputs(471)) xor (layer0_outputs(3978)));
    layer1_outputs(4245) <= '1';
    layer1_outputs(4246) <= not(layer0_outputs(2191));
    layer1_outputs(4247) <= layer0_outputs(1967);
    layer1_outputs(4248) <= not(layer0_outputs(2763));
    layer1_outputs(4249) <= not(layer0_outputs(525));
    layer1_outputs(4250) <= not(layer0_outputs(2930));
    layer1_outputs(4251) <= not((layer0_outputs(3148)) and (layer0_outputs(369)));
    layer1_outputs(4252) <= layer0_outputs(3479);
    layer1_outputs(4253) <= layer0_outputs(1606);
    layer1_outputs(4254) <= not(layer0_outputs(3485));
    layer1_outputs(4255) <= not(layer0_outputs(459)) or (layer0_outputs(282));
    layer1_outputs(4256) <= layer0_outputs(541);
    layer1_outputs(4257) <= not(layer0_outputs(2472));
    layer1_outputs(4258) <= layer0_outputs(2653);
    layer1_outputs(4259) <= not(layer0_outputs(2944));
    layer1_outputs(4260) <= not((layer0_outputs(5045)) or (layer0_outputs(3962)));
    layer1_outputs(4261) <= layer0_outputs(4847);
    layer1_outputs(4262) <= not((layer0_outputs(3727)) and (layer0_outputs(2416)));
    layer1_outputs(4263) <= not((layer0_outputs(4971)) and (layer0_outputs(4251)));
    layer1_outputs(4264) <= layer0_outputs(2215);
    layer1_outputs(4265) <= (layer0_outputs(2701)) and not (layer0_outputs(3393));
    layer1_outputs(4266) <= (layer0_outputs(2904)) and not (layer0_outputs(3610));
    layer1_outputs(4267) <= (layer0_outputs(2589)) and not (layer0_outputs(3790));
    layer1_outputs(4268) <= not(layer0_outputs(736));
    layer1_outputs(4269) <= not(layer0_outputs(2234)) or (layer0_outputs(4862));
    layer1_outputs(4270) <= (layer0_outputs(1850)) and not (layer0_outputs(4955));
    layer1_outputs(4271) <= not(layer0_outputs(761));
    layer1_outputs(4272) <= (layer0_outputs(49)) and not (layer0_outputs(2643));
    layer1_outputs(4273) <= not((layer0_outputs(1625)) or (layer0_outputs(2232)));
    layer1_outputs(4274) <= not((layer0_outputs(4146)) and (layer0_outputs(2060)));
    layer1_outputs(4275) <= (layer0_outputs(993)) and (layer0_outputs(4180));
    layer1_outputs(4276) <= (layer0_outputs(3378)) and not (layer0_outputs(3112));
    layer1_outputs(4277) <= (layer0_outputs(3421)) or (layer0_outputs(2459));
    layer1_outputs(4278) <= not(layer0_outputs(3261)) or (layer0_outputs(1433));
    layer1_outputs(4279) <= layer0_outputs(288);
    layer1_outputs(4280) <= layer0_outputs(2715);
    layer1_outputs(4281) <= not((layer0_outputs(1073)) and (layer0_outputs(1416)));
    layer1_outputs(4282) <= not(layer0_outputs(3933));
    layer1_outputs(4283) <= not((layer0_outputs(1708)) and (layer0_outputs(695)));
    layer1_outputs(4284) <= not(layer0_outputs(2055)) or (layer0_outputs(1948));
    layer1_outputs(4285) <= not(layer0_outputs(3366));
    layer1_outputs(4286) <= not(layer0_outputs(5014)) or (layer0_outputs(3519));
    layer1_outputs(4287) <= not(layer0_outputs(3967)) or (layer0_outputs(4910));
    layer1_outputs(4288) <= not(layer0_outputs(575));
    layer1_outputs(4289) <= '1';
    layer1_outputs(4290) <= (layer0_outputs(4292)) and (layer0_outputs(2107));
    layer1_outputs(4291) <= not(layer0_outputs(939));
    layer1_outputs(4292) <= not(layer0_outputs(4054));
    layer1_outputs(4293) <= (layer0_outputs(1482)) and not (layer0_outputs(2326));
    layer1_outputs(4294) <= (layer0_outputs(763)) and (layer0_outputs(1680));
    layer1_outputs(4295) <= (layer0_outputs(2441)) and not (layer0_outputs(1059));
    layer1_outputs(4296) <= (layer0_outputs(1154)) and (layer0_outputs(2249));
    layer1_outputs(4297) <= layer0_outputs(3404);
    layer1_outputs(4298) <= (layer0_outputs(2198)) and not (layer0_outputs(2229));
    layer1_outputs(4299) <= not(layer0_outputs(4497)) or (layer0_outputs(2593));
    layer1_outputs(4300) <= not((layer0_outputs(4896)) or (layer0_outputs(4389)));
    layer1_outputs(4301) <= not(layer0_outputs(4570)) or (layer0_outputs(1918));
    layer1_outputs(4302) <= not(layer0_outputs(1264));
    layer1_outputs(4303) <= not((layer0_outputs(1652)) and (layer0_outputs(4238)));
    layer1_outputs(4304) <= not(layer0_outputs(477)) or (layer0_outputs(3198));
    layer1_outputs(4305) <= (layer0_outputs(695)) and (layer0_outputs(774));
    layer1_outputs(4306) <= (layer0_outputs(4951)) and (layer0_outputs(3040));
    layer1_outputs(4307) <= not(layer0_outputs(4770)) or (layer0_outputs(768));
    layer1_outputs(4308) <= (layer0_outputs(5097)) and (layer0_outputs(1426));
    layer1_outputs(4309) <= (layer0_outputs(5107)) and not (layer0_outputs(3941));
    layer1_outputs(4310) <= (layer0_outputs(2559)) and not (layer0_outputs(637));
    layer1_outputs(4311) <= not(layer0_outputs(1217));
    layer1_outputs(4312) <= not(layer0_outputs(1397));
    layer1_outputs(4313) <= not(layer0_outputs(3424)) or (layer0_outputs(36));
    layer1_outputs(4314) <= not(layer0_outputs(3044)) or (layer0_outputs(171));
    layer1_outputs(4315) <= '0';
    layer1_outputs(4316) <= not(layer0_outputs(4778));
    layer1_outputs(4317) <= not((layer0_outputs(969)) or (layer0_outputs(53)));
    layer1_outputs(4318) <= (layer0_outputs(4007)) and (layer0_outputs(314));
    layer1_outputs(4319) <= '1';
    layer1_outputs(4320) <= not(layer0_outputs(4923)) or (layer0_outputs(1042));
    layer1_outputs(4321) <= (layer0_outputs(4666)) and (layer0_outputs(3648));
    layer1_outputs(4322) <= layer0_outputs(2607);
    layer1_outputs(4323) <= (layer0_outputs(1343)) or (layer0_outputs(1581));
    layer1_outputs(4324) <= (layer0_outputs(1797)) or (layer0_outputs(2941));
    layer1_outputs(4325) <= not(layer0_outputs(3462)) or (layer0_outputs(1714));
    layer1_outputs(4326) <= not(layer0_outputs(971)) or (layer0_outputs(4842));
    layer1_outputs(4327) <= layer0_outputs(2287);
    layer1_outputs(4328) <= not(layer0_outputs(1781)) or (layer0_outputs(1518));
    layer1_outputs(4329) <= (layer0_outputs(219)) xor (layer0_outputs(4264));
    layer1_outputs(4330) <= not(layer0_outputs(688));
    layer1_outputs(4331) <= not((layer0_outputs(2053)) and (layer0_outputs(3074)));
    layer1_outputs(4332) <= not(layer0_outputs(1402));
    layer1_outputs(4333) <= (layer0_outputs(1589)) and (layer0_outputs(1392));
    layer1_outputs(4334) <= (layer0_outputs(1486)) and not (layer0_outputs(107));
    layer1_outputs(4335) <= (layer0_outputs(3190)) and not (layer0_outputs(3144));
    layer1_outputs(4336) <= not(layer0_outputs(1379)) or (layer0_outputs(2004));
    layer1_outputs(4337) <= layer0_outputs(856);
    layer1_outputs(4338) <= not(layer0_outputs(2644));
    layer1_outputs(4339) <= not(layer0_outputs(3926));
    layer1_outputs(4340) <= not((layer0_outputs(3815)) and (layer0_outputs(515)));
    layer1_outputs(4341) <= not(layer0_outputs(195));
    layer1_outputs(4342) <= not((layer0_outputs(2404)) or (layer0_outputs(3418)));
    layer1_outputs(4343) <= not((layer0_outputs(3980)) or (layer0_outputs(4657)));
    layer1_outputs(4344) <= layer0_outputs(1716);
    layer1_outputs(4345) <= layer0_outputs(4823);
    layer1_outputs(4346) <= not(layer0_outputs(2505)) or (layer0_outputs(4994));
    layer1_outputs(4347) <= layer0_outputs(2724);
    layer1_outputs(4348) <= (layer0_outputs(285)) and not (layer0_outputs(2131));
    layer1_outputs(4349) <= (layer0_outputs(3241)) xor (layer0_outputs(802));
    layer1_outputs(4350) <= (layer0_outputs(2014)) and (layer0_outputs(4218));
    layer1_outputs(4351) <= (layer0_outputs(2460)) and not (layer0_outputs(922));
    layer1_outputs(4352) <= (layer0_outputs(571)) and not (layer0_outputs(203));
    layer1_outputs(4353) <= (layer0_outputs(3229)) and not (layer0_outputs(1615));
    layer1_outputs(4354) <= (layer0_outputs(3643)) and (layer0_outputs(2122));
    layer1_outputs(4355) <= layer0_outputs(1684);
    layer1_outputs(4356) <= not((layer0_outputs(4330)) and (layer0_outputs(542)));
    layer1_outputs(4357) <= (layer0_outputs(4931)) and not (layer0_outputs(4746));
    layer1_outputs(4358) <= layer0_outputs(1127);
    layer1_outputs(4359) <= not(layer0_outputs(1810));
    layer1_outputs(4360) <= layer0_outputs(1692);
    layer1_outputs(4361) <= (layer0_outputs(2674)) or (layer0_outputs(1285));
    layer1_outputs(4362) <= not(layer0_outputs(1354));
    layer1_outputs(4363) <= not(layer0_outputs(2549));
    layer1_outputs(4364) <= not(layer0_outputs(2791));
    layer1_outputs(4365) <= not((layer0_outputs(1681)) and (layer0_outputs(1734)));
    layer1_outputs(4366) <= not((layer0_outputs(2760)) and (layer0_outputs(1086)));
    layer1_outputs(4367) <= not((layer0_outputs(3582)) and (layer0_outputs(4770)));
    layer1_outputs(4368) <= (layer0_outputs(3555)) and not (layer0_outputs(4760));
    layer1_outputs(4369) <= layer0_outputs(4749);
    layer1_outputs(4370) <= not(layer0_outputs(1215));
    layer1_outputs(4371) <= (layer0_outputs(2634)) or (layer0_outputs(4476));
    layer1_outputs(4372) <= layer0_outputs(3014);
    layer1_outputs(4373) <= layer0_outputs(460);
    layer1_outputs(4374) <= not(layer0_outputs(3928));
    layer1_outputs(4375) <= layer0_outputs(4643);
    layer1_outputs(4376) <= (layer0_outputs(4060)) or (layer0_outputs(4299));
    layer1_outputs(4377) <= not(layer0_outputs(1508)) or (layer0_outputs(1127));
    layer1_outputs(4378) <= not(layer0_outputs(4228));
    layer1_outputs(4379) <= not(layer0_outputs(2657));
    layer1_outputs(4380) <= not(layer0_outputs(3028));
    layer1_outputs(4381) <= layer0_outputs(552);
    layer1_outputs(4382) <= '0';
    layer1_outputs(4383) <= '1';
    layer1_outputs(4384) <= '1';
    layer1_outputs(4385) <= not((layer0_outputs(3337)) xor (layer0_outputs(3420)));
    layer1_outputs(4386) <= not(layer0_outputs(3363));
    layer1_outputs(4387) <= (layer0_outputs(5072)) and not (layer0_outputs(822));
    layer1_outputs(4388) <= not(layer0_outputs(1535)) or (layer0_outputs(1351));
    layer1_outputs(4389) <= (layer0_outputs(3155)) or (layer0_outputs(3360));
    layer1_outputs(4390) <= not((layer0_outputs(2233)) and (layer0_outputs(1616)));
    layer1_outputs(4391) <= (layer0_outputs(1536)) xor (layer0_outputs(1601));
    layer1_outputs(4392) <= not(layer0_outputs(2290)) or (layer0_outputs(893));
    layer1_outputs(4393) <= '0';
    layer1_outputs(4394) <= not((layer0_outputs(3130)) and (layer0_outputs(4229)));
    layer1_outputs(4395) <= '0';
    layer1_outputs(4396) <= (layer0_outputs(2040)) and not (layer0_outputs(3083));
    layer1_outputs(4397) <= not(layer0_outputs(1669));
    layer1_outputs(4398) <= layer0_outputs(3209);
    layer1_outputs(4399) <= layer0_outputs(629);
    layer1_outputs(4400) <= (layer0_outputs(2589)) and not (layer0_outputs(3207));
    layer1_outputs(4401) <= not(layer0_outputs(595));
    layer1_outputs(4402) <= (layer0_outputs(1631)) or (layer0_outputs(4439));
    layer1_outputs(4403) <= (layer0_outputs(1925)) and not (layer0_outputs(1634));
    layer1_outputs(4404) <= not(layer0_outputs(1788));
    layer1_outputs(4405) <= not((layer0_outputs(1702)) or (layer0_outputs(3075)));
    layer1_outputs(4406) <= (layer0_outputs(258)) or (layer0_outputs(4534));
    layer1_outputs(4407) <= not(layer0_outputs(4564));
    layer1_outputs(4408) <= (layer0_outputs(1366)) and not (layer0_outputs(3495));
    layer1_outputs(4409) <= not(layer0_outputs(165));
    layer1_outputs(4410) <= '0';
    layer1_outputs(4411) <= not((layer0_outputs(851)) or (layer0_outputs(1545)));
    layer1_outputs(4412) <= (layer0_outputs(1455)) and not (layer0_outputs(489));
    layer1_outputs(4413) <= not(layer0_outputs(2060)) or (layer0_outputs(659));
    layer1_outputs(4414) <= (layer0_outputs(5071)) and not (layer0_outputs(1443));
    layer1_outputs(4415) <= not(layer0_outputs(1704));
    layer1_outputs(4416) <= (layer0_outputs(905)) and (layer0_outputs(2079));
    layer1_outputs(4417) <= layer0_outputs(3455);
    layer1_outputs(4418) <= not(layer0_outputs(3455)) or (layer0_outputs(3716));
    layer1_outputs(4419) <= not(layer0_outputs(442));
    layer1_outputs(4420) <= not(layer0_outputs(2930)) or (layer0_outputs(2524));
    layer1_outputs(4421) <= not(layer0_outputs(156));
    layer1_outputs(4422) <= not(layer0_outputs(2170));
    layer1_outputs(4423) <= not(layer0_outputs(2350)) or (layer0_outputs(1558));
    layer1_outputs(4424) <= not(layer0_outputs(1940)) or (layer0_outputs(4177));
    layer1_outputs(4425) <= (layer0_outputs(4751)) or (layer0_outputs(1323));
    layer1_outputs(4426) <= layer0_outputs(1452);
    layer1_outputs(4427) <= not((layer0_outputs(1758)) or (layer0_outputs(1997)));
    layer1_outputs(4428) <= (layer0_outputs(164)) and not (layer0_outputs(279));
    layer1_outputs(4429) <= (layer0_outputs(2374)) or (layer0_outputs(3918));
    layer1_outputs(4430) <= not(layer0_outputs(336));
    layer1_outputs(4431) <= (layer0_outputs(2722)) or (layer0_outputs(4720));
    layer1_outputs(4432) <= layer0_outputs(1232);
    layer1_outputs(4433) <= layer0_outputs(4474);
    layer1_outputs(4434) <= not((layer0_outputs(108)) and (layer0_outputs(2567)));
    layer1_outputs(4435) <= (layer0_outputs(4457)) xor (layer0_outputs(1149));
    layer1_outputs(4436) <= '1';
    layer1_outputs(4437) <= (layer0_outputs(5073)) or (layer0_outputs(584));
    layer1_outputs(4438) <= layer0_outputs(1071);
    layer1_outputs(4439) <= layer0_outputs(4317);
    layer1_outputs(4440) <= layer0_outputs(2612);
    layer1_outputs(4441) <= not(layer0_outputs(678));
    layer1_outputs(4442) <= (layer0_outputs(3119)) and (layer0_outputs(2650));
    layer1_outputs(4443) <= layer0_outputs(4561);
    layer1_outputs(4444) <= not(layer0_outputs(3630));
    layer1_outputs(4445) <= not(layer0_outputs(165));
    layer1_outputs(4446) <= (layer0_outputs(1895)) and not (layer0_outputs(3675));
    layer1_outputs(4447) <= not(layer0_outputs(4600)) or (layer0_outputs(1087));
    layer1_outputs(4448) <= not(layer0_outputs(2853));
    layer1_outputs(4449) <= '0';
    layer1_outputs(4450) <= (layer0_outputs(4717)) and (layer0_outputs(2171));
    layer1_outputs(4451) <= (layer0_outputs(1241)) and (layer0_outputs(3181));
    layer1_outputs(4452) <= (layer0_outputs(2063)) xor (layer0_outputs(2380));
    layer1_outputs(4453) <= not((layer0_outputs(4291)) or (layer0_outputs(4934)));
    layer1_outputs(4454) <= not(layer0_outputs(1611));
    layer1_outputs(4455) <= not(layer0_outputs(2025)) or (layer0_outputs(1332));
    layer1_outputs(4456) <= not(layer0_outputs(1459)) or (layer0_outputs(405));
    layer1_outputs(4457) <= (layer0_outputs(1328)) and not (layer0_outputs(4865));
    layer1_outputs(4458) <= (layer0_outputs(616)) and (layer0_outputs(4824));
    layer1_outputs(4459) <= layer0_outputs(2927);
    layer1_outputs(4460) <= not(layer0_outputs(4997)) or (layer0_outputs(1482));
    layer1_outputs(4461) <= not((layer0_outputs(3505)) and (layer0_outputs(1814)));
    layer1_outputs(4462) <= not(layer0_outputs(4182));
    layer1_outputs(4463) <= not(layer0_outputs(1608));
    layer1_outputs(4464) <= (layer0_outputs(4987)) xor (layer0_outputs(3119));
    layer1_outputs(4465) <= not(layer0_outputs(3525));
    layer1_outputs(4466) <= '1';
    layer1_outputs(4467) <= not((layer0_outputs(197)) xor (layer0_outputs(3887)));
    layer1_outputs(4468) <= layer0_outputs(2254);
    layer1_outputs(4469) <= not(layer0_outputs(159));
    layer1_outputs(4470) <= not(layer0_outputs(2390));
    layer1_outputs(4471) <= (layer0_outputs(668)) and not (layer0_outputs(1262));
    layer1_outputs(4472) <= layer0_outputs(3135);
    layer1_outputs(4473) <= '1';
    layer1_outputs(4474) <= not((layer0_outputs(770)) or (layer0_outputs(699)));
    layer1_outputs(4475) <= (layer0_outputs(2012)) and not (layer0_outputs(743));
    layer1_outputs(4476) <= layer0_outputs(1819);
    layer1_outputs(4477) <= not(layer0_outputs(1905));
    layer1_outputs(4478) <= '0';
    layer1_outputs(4479) <= not((layer0_outputs(2398)) and (layer0_outputs(2013)));
    layer1_outputs(4480) <= (layer0_outputs(4858)) or (layer0_outputs(2046));
    layer1_outputs(4481) <= layer0_outputs(4857);
    layer1_outputs(4482) <= not(layer0_outputs(2942));
    layer1_outputs(4483) <= not(layer0_outputs(4885));
    layer1_outputs(4484) <= not((layer0_outputs(3006)) or (layer0_outputs(4962)));
    layer1_outputs(4485) <= (layer0_outputs(4249)) or (layer0_outputs(4636));
    layer1_outputs(4486) <= (layer0_outputs(4162)) and (layer0_outputs(2401));
    layer1_outputs(4487) <= not(layer0_outputs(3169));
    layer1_outputs(4488) <= not(layer0_outputs(4010));
    layer1_outputs(4489) <= layer0_outputs(2291);
    layer1_outputs(4490) <= not((layer0_outputs(1449)) or (layer0_outputs(3056)));
    layer1_outputs(4491) <= (layer0_outputs(212)) and not (layer0_outputs(248));
    layer1_outputs(4492) <= not(layer0_outputs(3301));
    layer1_outputs(4493) <= not(layer0_outputs(1723)) or (layer0_outputs(1862));
    layer1_outputs(4494) <= not(layer0_outputs(2480));
    layer1_outputs(4495) <= '0';
    layer1_outputs(4496) <= layer0_outputs(2905);
    layer1_outputs(4497) <= layer0_outputs(4335);
    layer1_outputs(4498) <= layer0_outputs(1524);
    layer1_outputs(4499) <= '0';
    layer1_outputs(4500) <= not((layer0_outputs(1305)) xor (layer0_outputs(3268)));
    layer1_outputs(4501) <= not(layer0_outputs(914)) or (layer0_outputs(2090));
    layer1_outputs(4502) <= (layer0_outputs(4309)) or (layer0_outputs(3047));
    layer1_outputs(4503) <= layer0_outputs(1474);
    layer1_outputs(4504) <= layer0_outputs(4687);
    layer1_outputs(4505) <= (layer0_outputs(2741)) or (layer0_outputs(2376));
    layer1_outputs(4506) <= not(layer0_outputs(1311));
    layer1_outputs(4507) <= layer0_outputs(3759);
    layer1_outputs(4508) <= not(layer0_outputs(1792));
    layer1_outputs(4509) <= (layer0_outputs(3644)) and not (layer0_outputs(1978));
    layer1_outputs(4510) <= not(layer0_outputs(3931)) or (layer0_outputs(1367));
    layer1_outputs(4511) <= not((layer0_outputs(3537)) and (layer0_outputs(3637)));
    layer1_outputs(4512) <= (layer0_outputs(4441)) xor (layer0_outputs(1961));
    layer1_outputs(4513) <= not(layer0_outputs(2898));
    layer1_outputs(4514) <= not((layer0_outputs(3124)) or (layer0_outputs(3297)));
    layer1_outputs(4515) <= not(layer0_outputs(4732));
    layer1_outputs(4516) <= (layer0_outputs(4637)) and not (layer0_outputs(3280));
    layer1_outputs(4517) <= (layer0_outputs(4052)) and (layer0_outputs(1161));
    layer1_outputs(4518) <= not((layer0_outputs(3011)) or (layer0_outputs(4543)));
    layer1_outputs(4519) <= not(layer0_outputs(3000));
    layer1_outputs(4520) <= not(layer0_outputs(3773));
    layer1_outputs(4521) <= (layer0_outputs(4917)) and not (layer0_outputs(2165));
    layer1_outputs(4522) <= not(layer0_outputs(2097));
    layer1_outputs(4523) <= '1';
    layer1_outputs(4524) <= '0';
    layer1_outputs(4525) <= not((layer0_outputs(1791)) xor (layer0_outputs(1491)));
    layer1_outputs(4526) <= not(layer0_outputs(5092));
    layer1_outputs(4527) <= not(layer0_outputs(897)) or (layer0_outputs(4096));
    layer1_outputs(4528) <= layer0_outputs(885);
    layer1_outputs(4529) <= (layer0_outputs(2247)) or (layer0_outputs(905));
    layer1_outputs(4530) <= (layer0_outputs(4555)) xor (layer0_outputs(1284));
    layer1_outputs(4531) <= not(layer0_outputs(439));
    layer1_outputs(4532) <= '1';
    layer1_outputs(4533) <= (layer0_outputs(3539)) and not (layer0_outputs(960));
    layer1_outputs(4534) <= '1';
    layer1_outputs(4535) <= layer0_outputs(1240);
    layer1_outputs(4536) <= not(layer0_outputs(5085));
    layer1_outputs(4537) <= not(layer0_outputs(1297));
    layer1_outputs(4538) <= not(layer0_outputs(1764)) or (layer0_outputs(1257));
    layer1_outputs(4539) <= not((layer0_outputs(849)) xor (layer0_outputs(4976)));
    layer1_outputs(4540) <= (layer0_outputs(493)) and not (layer0_outputs(3188));
    layer1_outputs(4541) <= (layer0_outputs(4253)) or (layer0_outputs(297));
    layer1_outputs(4542) <= layer0_outputs(3676);
    layer1_outputs(4543) <= not(layer0_outputs(3915));
    layer1_outputs(4544) <= layer0_outputs(323);
    layer1_outputs(4545) <= (layer0_outputs(5096)) or (layer0_outputs(1647));
    layer1_outputs(4546) <= (layer0_outputs(4900)) and not (layer0_outputs(728));
    layer1_outputs(4547) <= (layer0_outputs(4929)) and not (layer0_outputs(3293));
    layer1_outputs(4548) <= not((layer0_outputs(4829)) and (layer0_outputs(4705)));
    layer1_outputs(4549) <= not(layer0_outputs(4000)) or (layer0_outputs(1933));
    layer1_outputs(4550) <= layer0_outputs(4867);
    layer1_outputs(4551) <= layer0_outputs(273);
    layer1_outputs(4552) <= '1';
    layer1_outputs(4553) <= layer0_outputs(927);
    layer1_outputs(4554) <= layer0_outputs(265);
    layer1_outputs(4555) <= not(layer0_outputs(4736)) or (layer0_outputs(1860));
    layer1_outputs(4556) <= (layer0_outputs(2563)) and not (layer0_outputs(5060));
    layer1_outputs(4557) <= (layer0_outputs(3925)) and not (layer0_outputs(2244));
    layer1_outputs(4558) <= layer0_outputs(1824);
    layer1_outputs(4559) <= not((layer0_outputs(4379)) or (layer0_outputs(145)));
    layer1_outputs(4560) <= layer0_outputs(1013);
    layer1_outputs(4561) <= not(layer0_outputs(4290)) or (layer0_outputs(1908));
    layer1_outputs(4562) <= not(layer0_outputs(4473));
    layer1_outputs(4563) <= (layer0_outputs(3597)) and (layer0_outputs(1537));
    layer1_outputs(4564) <= (layer0_outputs(186)) and not (layer0_outputs(3526));
    layer1_outputs(4565) <= not(layer0_outputs(163));
    layer1_outputs(4566) <= not((layer0_outputs(1243)) and (layer0_outputs(2672)));
    layer1_outputs(4567) <= not((layer0_outputs(4219)) or (layer0_outputs(1782)));
    layer1_outputs(4568) <= not((layer0_outputs(540)) or (layer0_outputs(4215)));
    layer1_outputs(4569) <= not(layer0_outputs(149)) or (layer0_outputs(3305));
    layer1_outputs(4570) <= '1';
    layer1_outputs(4571) <= not(layer0_outputs(2439));
    layer1_outputs(4572) <= layer0_outputs(3188);
    layer1_outputs(4573) <= not(layer0_outputs(1980));
    layer1_outputs(4574) <= not(layer0_outputs(3256)) or (layer0_outputs(1719));
    layer1_outputs(4575) <= not(layer0_outputs(4515));
    layer1_outputs(4576) <= (layer0_outputs(3903)) and (layer0_outputs(3766));
    layer1_outputs(4577) <= layer0_outputs(587);
    layer1_outputs(4578) <= (layer0_outputs(175)) or (layer0_outputs(4811));
    layer1_outputs(4579) <= not((layer0_outputs(3022)) and (layer0_outputs(2099)));
    layer1_outputs(4580) <= not(layer0_outputs(4843));
    layer1_outputs(4581) <= layer0_outputs(1962);
    layer1_outputs(4582) <= not(layer0_outputs(3747)) or (layer0_outputs(3036));
    layer1_outputs(4583) <= layer0_outputs(735);
    layer1_outputs(4584) <= (layer0_outputs(4428)) and not (layer0_outputs(2158));
    layer1_outputs(4585) <= '1';
    layer1_outputs(4586) <= not((layer0_outputs(1696)) or (layer0_outputs(3329)));
    layer1_outputs(4587) <= not((layer0_outputs(982)) or (layer0_outputs(2728)));
    layer1_outputs(4588) <= not((layer0_outputs(1731)) or (layer0_outputs(2084)));
    layer1_outputs(4589) <= layer0_outputs(3500);
    layer1_outputs(4590) <= not(layer0_outputs(3033)) or (layer0_outputs(462));
    layer1_outputs(4591) <= (layer0_outputs(2529)) or (layer0_outputs(1972));
    layer1_outputs(4592) <= (layer0_outputs(1194)) and not (layer0_outputs(2163));
    layer1_outputs(4593) <= not(layer0_outputs(1610)) or (layer0_outputs(652));
    layer1_outputs(4594) <= not(layer0_outputs(4641));
    layer1_outputs(4595) <= (layer0_outputs(4432)) or (layer0_outputs(400));
    layer1_outputs(4596) <= not(layer0_outputs(1796));
    layer1_outputs(4597) <= not(layer0_outputs(1576)) or (layer0_outputs(1654));
    layer1_outputs(4598) <= layer0_outputs(1926);
    layer1_outputs(4599) <= (layer0_outputs(3689)) and not (layer0_outputs(3990));
    layer1_outputs(4600) <= layer0_outputs(2732);
    layer1_outputs(4601) <= (layer0_outputs(3755)) xor (layer0_outputs(559));
    layer1_outputs(4602) <= (layer0_outputs(3907)) and not (layer0_outputs(3089));
    layer1_outputs(4603) <= '1';
    layer1_outputs(4604) <= layer0_outputs(2920);
    layer1_outputs(4605) <= not(layer0_outputs(4641));
    layer1_outputs(4606) <= not((layer0_outputs(1051)) or (layer0_outputs(3142)));
    layer1_outputs(4607) <= layer0_outputs(72);
    layer1_outputs(4608) <= layer0_outputs(1886);
    layer1_outputs(4609) <= not(layer0_outputs(3004)) or (layer0_outputs(699));
    layer1_outputs(4610) <= (layer0_outputs(2733)) and not (layer0_outputs(347));
    layer1_outputs(4611) <= not((layer0_outputs(1193)) or (layer0_outputs(3740)));
    layer1_outputs(4612) <= layer0_outputs(1882);
    layer1_outputs(4613) <= not(layer0_outputs(1577));
    layer1_outputs(4614) <= not((layer0_outputs(1432)) or (layer0_outputs(1726)));
    layer1_outputs(4615) <= '1';
    layer1_outputs(4616) <= (layer0_outputs(2259)) xor (layer0_outputs(2686));
    layer1_outputs(4617) <= not(layer0_outputs(4569));
    layer1_outputs(4618) <= '1';
    layer1_outputs(4619) <= '1';
    layer1_outputs(4620) <= not(layer0_outputs(791));
    layer1_outputs(4621) <= not(layer0_outputs(2687));
    layer1_outputs(4622) <= layer0_outputs(4946);
    layer1_outputs(4623) <= (layer0_outputs(340)) and not (layer0_outputs(4686));
    layer1_outputs(4624) <= not(layer0_outputs(865)) or (layer0_outputs(3302));
    layer1_outputs(4625) <= (layer0_outputs(4363)) and (layer0_outputs(2560));
    layer1_outputs(4626) <= layer0_outputs(3064);
    layer1_outputs(4627) <= (layer0_outputs(3250)) or (layer0_outputs(3159));
    layer1_outputs(4628) <= not(layer0_outputs(1906)) or (layer0_outputs(1828));
    layer1_outputs(4629) <= (layer0_outputs(988)) and (layer0_outputs(379));
    layer1_outputs(4630) <= layer0_outputs(535);
    layer1_outputs(4631) <= not(layer0_outputs(463));
    layer1_outputs(4632) <= not(layer0_outputs(2525));
    layer1_outputs(4633) <= not(layer0_outputs(4077));
    layer1_outputs(4634) <= (layer0_outputs(2373)) and not (layer0_outputs(5003));
    layer1_outputs(4635) <= not(layer0_outputs(862));
    layer1_outputs(4636) <= not(layer0_outputs(3364));
    layer1_outputs(4637) <= not((layer0_outputs(2705)) and (layer0_outputs(2472)));
    layer1_outputs(4638) <= not((layer0_outputs(1270)) or (layer0_outputs(2130)));
    layer1_outputs(4639) <= not(layer0_outputs(3255));
    layer1_outputs(4640) <= not((layer0_outputs(1844)) and (layer0_outputs(2656)));
    layer1_outputs(4641) <= (layer0_outputs(1994)) and (layer0_outputs(3850));
    layer1_outputs(4642) <= not(layer0_outputs(426));
    layer1_outputs(4643) <= layer0_outputs(1180);
    layer1_outputs(4644) <= not((layer0_outputs(221)) xor (layer0_outputs(4463)));
    layer1_outputs(4645) <= not(layer0_outputs(417));
    layer1_outputs(4646) <= layer0_outputs(1339);
    layer1_outputs(4647) <= not(layer0_outputs(4316));
    layer1_outputs(4648) <= not((layer0_outputs(4670)) and (layer0_outputs(1124)));
    layer1_outputs(4649) <= not(layer0_outputs(3879));
    layer1_outputs(4650) <= not(layer0_outputs(1410));
    layer1_outputs(4651) <= (layer0_outputs(1266)) or (layer0_outputs(511));
    layer1_outputs(4652) <= (layer0_outputs(3842)) or (layer0_outputs(3541));
    layer1_outputs(4653) <= '1';
    layer1_outputs(4654) <= (layer0_outputs(3533)) or (layer0_outputs(679));
    layer1_outputs(4655) <= (layer0_outputs(3960)) and (layer0_outputs(2280));
    layer1_outputs(4656) <= not(layer0_outputs(164)) or (layer0_outputs(2096));
    layer1_outputs(4657) <= not(layer0_outputs(294));
    layer1_outputs(4658) <= not(layer0_outputs(836));
    layer1_outputs(4659) <= not((layer0_outputs(2411)) or (layer0_outputs(3294)));
    layer1_outputs(4660) <= not(layer0_outputs(2239));
    layer1_outputs(4661) <= (layer0_outputs(3431)) and not (layer0_outputs(4257));
    layer1_outputs(4662) <= layer0_outputs(1724);
    layer1_outputs(4663) <= layer0_outputs(2260);
    layer1_outputs(4664) <= not(layer0_outputs(3914));
    layer1_outputs(4665) <= not(layer0_outputs(1830)) or (layer0_outputs(4870));
    layer1_outputs(4666) <= layer0_outputs(2488);
    layer1_outputs(4667) <= (layer0_outputs(4027)) and not (layer0_outputs(1081));
    layer1_outputs(4668) <= layer0_outputs(1451);
    layer1_outputs(4669) <= (layer0_outputs(1743)) or (layer0_outputs(2422));
    layer1_outputs(4670) <= not(layer0_outputs(1055));
    layer1_outputs(4671) <= not(layer0_outputs(823)) or (layer0_outputs(193));
    layer1_outputs(4672) <= not(layer0_outputs(4180));
    layer1_outputs(4673) <= not((layer0_outputs(4426)) or (layer0_outputs(4254)));
    layer1_outputs(4674) <= layer0_outputs(2683);
    layer1_outputs(4675) <= (layer0_outputs(4450)) and not (layer0_outputs(1414));
    layer1_outputs(4676) <= not((layer0_outputs(3297)) and (layer0_outputs(3200)));
    layer1_outputs(4677) <= not(layer0_outputs(3391)) or (layer0_outputs(2642));
    layer1_outputs(4678) <= not((layer0_outputs(4494)) or (layer0_outputs(1813)));
    layer1_outputs(4679) <= (layer0_outputs(1883)) and not (layer0_outputs(668));
    layer1_outputs(4680) <= not((layer0_outputs(2706)) or (layer0_outputs(4575)));
    layer1_outputs(4681) <= not((layer0_outputs(3694)) and (layer0_outputs(747)));
    layer1_outputs(4682) <= not(layer0_outputs(4322)) or (layer0_outputs(4840));
    layer1_outputs(4683) <= not((layer0_outputs(2347)) xor (layer0_outputs(901)));
    layer1_outputs(4684) <= not((layer0_outputs(3092)) and (layer0_outputs(3024)));
    layer1_outputs(4685) <= (layer0_outputs(3820)) and not (layer0_outputs(2109));
    layer1_outputs(4686) <= (layer0_outputs(3910)) and not (layer0_outputs(497));
    layer1_outputs(4687) <= not(layer0_outputs(320));
    layer1_outputs(4688) <= layer0_outputs(2218);
    layer1_outputs(4689) <= (layer0_outputs(255)) or (layer0_outputs(3018));
    layer1_outputs(4690) <= layer0_outputs(1234);
    layer1_outputs(4691) <= not(layer0_outputs(1130)) or (layer0_outputs(3949));
    layer1_outputs(4692) <= not(layer0_outputs(4284));
    layer1_outputs(4693) <= layer0_outputs(3177);
    layer1_outputs(4694) <= layer0_outputs(3858);
    layer1_outputs(4695) <= not((layer0_outputs(4342)) and (layer0_outputs(3232)));
    layer1_outputs(4696) <= not(layer0_outputs(2516));
    layer1_outputs(4697) <= not(layer0_outputs(63));
    layer1_outputs(4698) <= not((layer0_outputs(2443)) and (layer0_outputs(655)));
    layer1_outputs(4699) <= not(layer0_outputs(752)) or (layer0_outputs(1302));
    layer1_outputs(4700) <= layer0_outputs(4711);
    layer1_outputs(4701) <= not(layer0_outputs(1892));
    layer1_outputs(4702) <= not(layer0_outputs(997)) or (layer0_outputs(2986));
    layer1_outputs(4703) <= layer0_outputs(4191);
    layer1_outputs(4704) <= not(layer0_outputs(4273)) or (layer0_outputs(4399));
    layer1_outputs(4705) <= '0';
    layer1_outputs(4706) <= not(layer0_outputs(3618)) or (layer0_outputs(3741));
    layer1_outputs(4707) <= not(layer0_outputs(3880));
    layer1_outputs(4708) <= not(layer0_outputs(577)) or (layer0_outputs(3752));
    layer1_outputs(4709) <= not(layer0_outputs(3237));
    layer1_outputs(4710) <= not(layer0_outputs(4376));
    layer1_outputs(4711) <= (layer0_outputs(2120)) or (layer0_outputs(3437));
    layer1_outputs(4712) <= (layer0_outputs(2463)) and (layer0_outputs(2089));
    layer1_outputs(4713) <= not(layer0_outputs(2810));
    layer1_outputs(4714) <= layer0_outputs(1614);
    layer1_outputs(4715) <= not((layer0_outputs(3471)) and (layer0_outputs(4622)));
    layer1_outputs(4716) <= not(layer0_outputs(4243)) or (layer0_outputs(991));
    layer1_outputs(4717) <= (layer0_outputs(812)) xor (layer0_outputs(1487));
    layer1_outputs(4718) <= not(layer0_outputs(1172));
    layer1_outputs(4719) <= not(layer0_outputs(1888)) or (layer0_outputs(4990));
    layer1_outputs(4720) <= not(layer0_outputs(4392));
    layer1_outputs(4721) <= not((layer0_outputs(2022)) or (layer0_outputs(2550)));
    layer1_outputs(4722) <= not(layer0_outputs(589)) or (layer0_outputs(189));
    layer1_outputs(4723) <= not(layer0_outputs(676));
    layer1_outputs(4724) <= (layer0_outputs(3481)) and (layer0_outputs(3096));
    layer1_outputs(4725) <= '1';
    layer1_outputs(4726) <= not(layer0_outputs(506)) or (layer0_outputs(3899));
    layer1_outputs(4727) <= (layer0_outputs(2815)) or (layer0_outputs(3934));
    layer1_outputs(4728) <= not((layer0_outputs(2006)) xor (layer0_outputs(1003)));
    layer1_outputs(4729) <= layer0_outputs(607);
    layer1_outputs(4730) <= layer0_outputs(87);
    layer1_outputs(4731) <= (layer0_outputs(1437)) or (layer0_outputs(4572));
    layer1_outputs(4732) <= layer0_outputs(1476);
    layer1_outputs(4733) <= layer0_outputs(3131);
    layer1_outputs(4734) <= not(layer0_outputs(3514)) or (layer0_outputs(4948));
    layer1_outputs(4735) <= not((layer0_outputs(2603)) or (layer0_outputs(2722)));
    layer1_outputs(4736) <= (layer0_outputs(2979)) and not (layer0_outputs(3327));
    layer1_outputs(4737) <= not(layer0_outputs(536)) or (layer0_outputs(362));
    layer1_outputs(4738) <= layer0_outputs(247);
    layer1_outputs(4739) <= not(layer0_outputs(551));
    layer1_outputs(4740) <= (layer0_outputs(2903)) xor (layer0_outputs(2777));
    layer1_outputs(4741) <= not((layer0_outputs(2889)) or (layer0_outputs(1006)));
    layer1_outputs(4742) <= (layer0_outputs(3193)) and (layer0_outputs(3923));
    layer1_outputs(4743) <= layer0_outputs(4081);
    layer1_outputs(4744) <= layer0_outputs(4698);
    layer1_outputs(4745) <= not((layer0_outputs(2363)) or (layer0_outputs(593)));
    layer1_outputs(4746) <= not(layer0_outputs(4459));
    layer1_outputs(4747) <= layer0_outputs(2196);
    layer1_outputs(4748) <= not(layer0_outputs(4292)) or (layer0_outputs(224));
    layer1_outputs(4749) <= (layer0_outputs(1202)) or (layer0_outputs(2106));
    layer1_outputs(4750) <= (layer0_outputs(4044)) and not (layer0_outputs(526));
    layer1_outputs(4751) <= not(layer0_outputs(1400)) or (layer0_outputs(3660));
    layer1_outputs(4752) <= not(layer0_outputs(2424)) or (layer0_outputs(3621));
    layer1_outputs(4753) <= not((layer0_outputs(3568)) or (layer0_outputs(367)));
    layer1_outputs(4754) <= layer0_outputs(2971);
    layer1_outputs(4755) <= (layer0_outputs(394)) and (layer0_outputs(3569));
    layer1_outputs(4756) <= '1';
    layer1_outputs(4757) <= not(layer0_outputs(2636)) or (layer0_outputs(4905));
    layer1_outputs(4758) <= not(layer0_outputs(2059));
    layer1_outputs(4759) <= '0';
    layer1_outputs(4760) <= (layer0_outputs(2717)) and (layer0_outputs(980));
    layer1_outputs(4761) <= not(layer0_outputs(4769));
    layer1_outputs(4762) <= not((layer0_outputs(520)) or (layer0_outputs(890)));
    layer1_outputs(4763) <= not(layer0_outputs(425)) or (layer0_outputs(111));
    layer1_outputs(4764) <= not((layer0_outputs(2288)) or (layer0_outputs(1338)));
    layer1_outputs(4765) <= not(layer0_outputs(482)) or (layer0_outputs(4311));
    layer1_outputs(4766) <= not(layer0_outputs(3158)) or (layer0_outputs(1043));
    layer1_outputs(4767) <= not(layer0_outputs(2761));
    layer1_outputs(4768) <= not(layer0_outputs(406)) or (layer0_outputs(89));
    layer1_outputs(4769) <= not((layer0_outputs(3916)) xor (layer0_outputs(4861)));
    layer1_outputs(4770) <= not(layer0_outputs(5015));
    layer1_outputs(4771) <= layer0_outputs(4432);
    layer1_outputs(4772) <= layer0_outputs(3048);
    layer1_outputs(4773) <= not(layer0_outputs(1370)) or (layer0_outputs(1758));
    layer1_outputs(4774) <= not(layer0_outputs(3456)) or (layer0_outputs(2439));
    layer1_outputs(4775) <= layer0_outputs(4517);
    layer1_outputs(4776) <= not(layer0_outputs(5027));
    layer1_outputs(4777) <= not((layer0_outputs(4996)) or (layer0_outputs(2789)));
    layer1_outputs(4778) <= not(layer0_outputs(1780)) or (layer0_outputs(3539));
    layer1_outputs(4779) <= layer0_outputs(3622);
    layer1_outputs(4780) <= layer0_outputs(298);
    layer1_outputs(4781) <= not(layer0_outputs(3017));
    layer1_outputs(4782) <= layer0_outputs(3596);
    layer1_outputs(4783) <= not(layer0_outputs(565));
    layer1_outputs(4784) <= (layer0_outputs(992)) and (layer0_outputs(1952));
    layer1_outputs(4785) <= not(layer0_outputs(1038));
    layer1_outputs(4786) <= (layer0_outputs(1281)) and not (layer0_outputs(2730));
    layer1_outputs(4787) <= (layer0_outputs(3353)) and not (layer0_outputs(3105));
    layer1_outputs(4788) <= not(layer0_outputs(465)) or (layer0_outputs(874));
    layer1_outputs(4789) <= not(layer0_outputs(886));
    layer1_outputs(4790) <= (layer0_outputs(2077)) and not (layer0_outputs(719));
    layer1_outputs(4791) <= (layer0_outputs(3435)) and (layer0_outputs(4260));
    layer1_outputs(4792) <= (layer0_outputs(537)) and not (layer0_outputs(4970));
    layer1_outputs(4793) <= (layer0_outputs(1553)) and not (layer0_outputs(4927));
    layer1_outputs(4794) <= (layer0_outputs(1772)) and (layer0_outputs(4241));
    layer1_outputs(4795) <= not(layer0_outputs(2216));
    layer1_outputs(4796) <= '1';
    layer1_outputs(4797) <= not(layer0_outputs(553));
    layer1_outputs(4798) <= (layer0_outputs(134)) and (layer0_outputs(3757));
    layer1_outputs(4799) <= not((layer0_outputs(153)) xor (layer0_outputs(1254)));
    layer1_outputs(4800) <= not(layer0_outputs(3631)) or (layer0_outputs(4574));
    layer1_outputs(4801) <= not(layer0_outputs(275));
    layer1_outputs(4802) <= not(layer0_outputs(5056));
    layer1_outputs(4803) <= (layer0_outputs(1938)) and (layer0_outputs(4876));
    layer1_outputs(4804) <= layer0_outputs(3203);
    layer1_outputs(4805) <= layer0_outputs(3474);
    layer1_outputs(4806) <= (layer0_outputs(1177)) or (layer0_outputs(4113));
    layer1_outputs(4807) <= not((layer0_outputs(669)) and (layer0_outputs(850)));
    layer1_outputs(4808) <= not(layer0_outputs(3525)) or (layer0_outputs(799));
    layer1_outputs(4809) <= not(layer0_outputs(1081)) or (layer0_outputs(2391));
    layer1_outputs(4810) <= (layer0_outputs(4806)) and (layer0_outputs(3153));
    layer1_outputs(4811) <= layer0_outputs(4175);
    layer1_outputs(4812) <= layer0_outputs(409);
    layer1_outputs(4813) <= not(layer0_outputs(2469));
    layer1_outputs(4814) <= not(layer0_outputs(4183));
    layer1_outputs(4815) <= layer0_outputs(4593);
    layer1_outputs(4816) <= layer0_outputs(644);
    layer1_outputs(4817) <= layer0_outputs(484);
    layer1_outputs(4818) <= not((layer0_outputs(4566)) or (layer0_outputs(4831)));
    layer1_outputs(4819) <= not(layer0_outputs(1629)) or (layer0_outputs(1071));
    layer1_outputs(4820) <= (layer0_outputs(2681)) and not (layer0_outputs(896));
    layer1_outputs(4821) <= (layer0_outputs(241)) and (layer0_outputs(554));
    layer1_outputs(4822) <= not(layer0_outputs(888));
    layer1_outputs(4823) <= (layer0_outputs(1527)) and not (layer0_outputs(71));
    layer1_outputs(4824) <= not(layer0_outputs(3578)) or (layer0_outputs(857));
    layer1_outputs(4825) <= not((layer0_outputs(3095)) xor (layer0_outputs(2529)));
    layer1_outputs(4826) <= not(layer0_outputs(4415));
    layer1_outputs(4827) <= (layer0_outputs(3547)) or (layer0_outputs(3248));
    layer1_outputs(4828) <= not(layer0_outputs(4138));
    layer1_outputs(4829) <= (layer0_outputs(2030)) or (layer0_outputs(4585));
    layer1_outputs(4830) <= '0';
    layer1_outputs(4831) <= layer0_outputs(1317);
    layer1_outputs(4832) <= not(layer0_outputs(2002)) or (layer0_outputs(1133));
    layer1_outputs(4833) <= (layer0_outputs(83)) and (layer0_outputs(2485));
    layer1_outputs(4834) <= not(layer0_outputs(472));
    layer1_outputs(4835) <= not(layer0_outputs(24)) or (layer0_outputs(1691));
    layer1_outputs(4836) <= not(layer0_outputs(129)) or (layer0_outputs(4217));
    layer1_outputs(4837) <= layer0_outputs(3848);
    layer1_outputs(4838) <= layer0_outputs(842);
    layer1_outputs(4839) <= not((layer0_outputs(5068)) xor (layer0_outputs(5007)));
    layer1_outputs(4840) <= (layer0_outputs(2021)) or (layer0_outputs(4313));
    layer1_outputs(4841) <= (layer0_outputs(1494)) and (layer0_outputs(2769));
    layer1_outputs(4842) <= (layer0_outputs(2434)) xor (layer0_outputs(4494));
    layer1_outputs(4843) <= (layer0_outputs(560)) and not (layer0_outputs(992));
    layer1_outputs(4844) <= layer0_outputs(4090);
    layer1_outputs(4845) <= not(layer0_outputs(3678));
    layer1_outputs(4846) <= '1';
    layer1_outputs(4847) <= layer0_outputs(3977);
    layer1_outputs(4848) <= (layer0_outputs(1123)) and (layer0_outputs(3287));
    layer1_outputs(4849) <= layer0_outputs(5119);
    layer1_outputs(4850) <= not((layer0_outputs(405)) xor (layer0_outputs(1884)));
    layer1_outputs(4851) <= (layer0_outputs(363)) and not (layer0_outputs(2259));
    layer1_outputs(4852) <= '0';
    layer1_outputs(4853) <= (layer0_outputs(1659)) and not (layer0_outputs(1363));
    layer1_outputs(4854) <= (layer0_outputs(2054)) and not (layer0_outputs(3604));
    layer1_outputs(4855) <= not((layer0_outputs(3117)) and (layer0_outputs(3000)));
    layer1_outputs(4856) <= layer0_outputs(3735);
    layer1_outputs(4857) <= (layer0_outputs(1628)) and not (layer0_outputs(2819));
    layer1_outputs(4858) <= not(layer0_outputs(2372)) or (layer0_outputs(1032));
    layer1_outputs(4859) <= not((layer0_outputs(4352)) and (layer0_outputs(2449)));
    layer1_outputs(4860) <= not((layer0_outputs(2665)) or (layer0_outputs(2426)));
    layer1_outputs(4861) <= '0';
    layer1_outputs(4862) <= (layer0_outputs(1893)) and (layer0_outputs(2441));
    layer1_outputs(4863) <= not(layer0_outputs(2235)) or (layer0_outputs(1917));
    layer1_outputs(4864) <= (layer0_outputs(3296)) and (layer0_outputs(115));
    layer1_outputs(4865) <= layer0_outputs(3084);
    layer1_outputs(4866) <= '0';
    layer1_outputs(4867) <= (layer0_outputs(4336)) and (layer0_outputs(3031));
    layer1_outputs(4868) <= (layer0_outputs(4976)) and not (layer0_outputs(114));
    layer1_outputs(4869) <= not(layer0_outputs(5030)) or (layer0_outputs(3429));
    layer1_outputs(4870) <= (layer0_outputs(2110)) or (layer0_outputs(29));
    layer1_outputs(4871) <= not((layer0_outputs(3859)) and (layer0_outputs(3620)));
    layer1_outputs(4872) <= layer0_outputs(3186);
    layer1_outputs(4873) <= not(layer0_outputs(2157)) or (layer0_outputs(4946));
    layer1_outputs(4874) <= layer0_outputs(4312);
    layer1_outputs(4875) <= '0';
    layer1_outputs(4876) <= (layer0_outputs(835)) and (layer0_outputs(3184));
    layer1_outputs(4877) <= layer0_outputs(25);
    layer1_outputs(4878) <= layer0_outputs(2124);
    layer1_outputs(4879) <= (layer0_outputs(1698)) or (layer0_outputs(4328));
    layer1_outputs(4880) <= not((layer0_outputs(2786)) or (layer0_outputs(2236)));
    layer1_outputs(4881) <= not(layer0_outputs(3394)) or (layer0_outputs(512));
    layer1_outputs(4882) <= not(layer0_outputs(5081));
    layer1_outputs(4883) <= not((layer0_outputs(1483)) or (layer0_outputs(3312)));
    layer1_outputs(4884) <= not(layer0_outputs(3702));
    layer1_outputs(4885) <= not(layer0_outputs(1800)) or (layer0_outputs(4285));
    layer1_outputs(4886) <= '1';
    layer1_outputs(4887) <= '0';
    layer1_outputs(4888) <= not(layer0_outputs(4962));
    layer1_outputs(4889) <= '1';
    layer1_outputs(4890) <= (layer0_outputs(1963)) and not (layer0_outputs(2187));
    layer1_outputs(4891) <= not(layer0_outputs(2317));
    layer1_outputs(4892) <= not(layer0_outputs(4129)) or (layer0_outputs(929));
    layer1_outputs(4893) <= not((layer0_outputs(3180)) or (layer0_outputs(4381)));
    layer1_outputs(4894) <= layer0_outputs(4898);
    layer1_outputs(4895) <= not(layer0_outputs(554)) or (layer0_outputs(3642));
    layer1_outputs(4896) <= (layer0_outputs(1940)) and not (layer0_outputs(1963));
    layer1_outputs(4897) <= (layer0_outputs(4083)) and not (layer0_outputs(4248));
    layer1_outputs(4898) <= not(layer0_outputs(4901));
    layer1_outputs(4899) <= not(layer0_outputs(46));
    layer1_outputs(4900) <= (layer0_outputs(4727)) and not (layer0_outputs(3403));
    layer1_outputs(4901) <= layer0_outputs(4674);
    layer1_outputs(4902) <= '0';
    layer1_outputs(4903) <= not((layer0_outputs(541)) and (layer0_outputs(2781)));
    layer1_outputs(4904) <= not(layer0_outputs(4083));
    layer1_outputs(4905) <= layer0_outputs(988);
    layer1_outputs(4906) <= not(layer0_outputs(2549)) or (layer0_outputs(130));
    layer1_outputs(4907) <= not(layer0_outputs(4878));
    layer1_outputs(4908) <= not(layer0_outputs(751));
    layer1_outputs(4909) <= not((layer0_outputs(2360)) or (layer0_outputs(4249)));
    layer1_outputs(4910) <= not(layer0_outputs(5111)) or (layer0_outputs(4375));
    layer1_outputs(4911) <= (layer0_outputs(1930)) and not (layer0_outputs(2633));
    layer1_outputs(4912) <= not((layer0_outputs(2706)) and (layer0_outputs(1092)));
    layer1_outputs(4913) <= not(layer0_outputs(3050)) or (layer0_outputs(5051));
    layer1_outputs(4914) <= not(layer0_outputs(2442));
    layer1_outputs(4915) <= (layer0_outputs(3519)) and not (layer0_outputs(238));
    layer1_outputs(4916) <= not((layer0_outputs(781)) or (layer0_outputs(1642)));
    layer1_outputs(4917) <= '0';
    layer1_outputs(4918) <= not((layer0_outputs(619)) and (layer0_outputs(1032)));
    layer1_outputs(4919) <= (layer0_outputs(2265)) and (layer0_outputs(2514));
    layer1_outputs(4920) <= not(layer0_outputs(4810));
    layer1_outputs(4921) <= not((layer0_outputs(4800)) and (layer0_outputs(517)));
    layer1_outputs(4922) <= not(layer0_outputs(3177)) or (layer0_outputs(5015));
    layer1_outputs(4923) <= not(layer0_outputs(2179)) or (layer0_outputs(612));
    layer1_outputs(4924) <= layer0_outputs(3835);
    layer1_outputs(4925) <= (layer0_outputs(1621)) and (layer0_outputs(1357));
    layer1_outputs(4926) <= not(layer0_outputs(382));
    layer1_outputs(4927) <= layer0_outputs(4294);
    layer1_outputs(4928) <= (layer0_outputs(1881)) and not (layer0_outputs(549));
    layer1_outputs(4929) <= layer0_outputs(1657);
    layer1_outputs(4930) <= '1';
    layer1_outputs(4931) <= layer0_outputs(2944);
    layer1_outputs(4932) <= layer0_outputs(690);
    layer1_outputs(4933) <= not(layer0_outputs(1863));
    layer1_outputs(4934) <= not(layer0_outputs(2457)) or (layer0_outputs(3771));
    layer1_outputs(4935) <= not(layer0_outputs(3712));
    layer1_outputs(4936) <= (layer0_outputs(1389)) and not (layer0_outputs(3884));
    layer1_outputs(4937) <= layer0_outputs(179);
    layer1_outputs(4938) <= not(layer0_outputs(2934));
    layer1_outputs(4939) <= not(layer0_outputs(1880));
    layer1_outputs(4940) <= (layer0_outputs(3939)) and (layer0_outputs(3937));
    layer1_outputs(4941) <= (layer0_outputs(2507)) and not (layer0_outputs(4041));
    layer1_outputs(4942) <= '0';
    layer1_outputs(4943) <= not(layer0_outputs(3968)) or (layer0_outputs(2121));
    layer1_outputs(4944) <= not(layer0_outputs(4226));
    layer1_outputs(4945) <= not((layer0_outputs(4925)) or (layer0_outputs(5033)));
    layer1_outputs(4946) <= not(layer0_outputs(2475));
    layer1_outputs(4947) <= layer0_outputs(1160);
    layer1_outputs(4948) <= (layer0_outputs(4741)) and not (layer0_outputs(3815));
    layer1_outputs(4949) <= layer0_outputs(4608);
    layer1_outputs(4950) <= layer0_outputs(1253);
    layer1_outputs(4951) <= (layer0_outputs(1902)) and (layer0_outputs(3423));
    layer1_outputs(4952) <= (layer0_outputs(3531)) and (layer0_outputs(1834));
    layer1_outputs(4953) <= not(layer0_outputs(3739)) or (layer0_outputs(1229));
    layer1_outputs(4954) <= not(layer0_outputs(2476)) or (layer0_outputs(383));
    layer1_outputs(4955) <= not(layer0_outputs(268)) or (layer0_outputs(316));
    layer1_outputs(4956) <= layer0_outputs(4690);
    layer1_outputs(4957) <= layer0_outputs(798);
    layer1_outputs(4958) <= (layer0_outputs(2342)) and not (layer0_outputs(42));
    layer1_outputs(4959) <= (layer0_outputs(1473)) and not (layer0_outputs(2842));
    layer1_outputs(4960) <= '1';
    layer1_outputs(4961) <= not(layer0_outputs(995)) or (layer0_outputs(2670));
    layer1_outputs(4962) <= not(layer0_outputs(2257));
    layer1_outputs(4963) <= layer0_outputs(3423);
    layer1_outputs(4964) <= not(layer0_outputs(3609));
    layer1_outputs(4965) <= layer0_outputs(677);
    layer1_outputs(4966) <= layer0_outputs(2352);
    layer1_outputs(4967) <= not(layer0_outputs(2996)) or (layer0_outputs(4195));
    layer1_outputs(4968) <= layer0_outputs(3366);
    layer1_outputs(4969) <= not((layer0_outputs(375)) and (layer0_outputs(4984)));
    layer1_outputs(4970) <= (layer0_outputs(3767)) or (layer0_outputs(1406));
    layer1_outputs(4971) <= not(layer0_outputs(855)) or (layer0_outputs(3956));
    layer1_outputs(4972) <= not((layer0_outputs(797)) and (layer0_outputs(1880)));
    layer1_outputs(4973) <= not((layer0_outputs(907)) and (layer0_outputs(4398)));
    layer1_outputs(4974) <= (layer0_outputs(2680)) or (layer0_outputs(3144));
    layer1_outputs(4975) <= not((layer0_outputs(3616)) and (layer0_outputs(4121)));
    layer1_outputs(4976) <= layer0_outputs(2771);
    layer1_outputs(4977) <= (layer0_outputs(4348)) and not (layer0_outputs(26));
    layer1_outputs(4978) <= not((layer0_outputs(2307)) or (layer0_outputs(4591)));
    layer1_outputs(4979) <= layer0_outputs(45);
    layer1_outputs(4980) <= (layer0_outputs(3199)) and not (layer0_outputs(2227));
    layer1_outputs(4981) <= not((layer0_outputs(4719)) or (layer0_outputs(4938)));
    layer1_outputs(4982) <= not(layer0_outputs(3807)) or (layer0_outputs(3457));
    layer1_outputs(4983) <= not((layer0_outputs(3304)) and (layer0_outputs(932)));
    layer1_outputs(4984) <= not(layer0_outputs(276));
    layer1_outputs(4985) <= layer0_outputs(957);
    layer1_outputs(4986) <= not(layer0_outputs(4580));
    layer1_outputs(4987) <= not(layer0_outputs(1860));
    layer1_outputs(4988) <= not(layer0_outputs(1263));
    layer1_outputs(4989) <= not(layer0_outputs(3042)) or (layer0_outputs(1336));
    layer1_outputs(4990) <= not((layer0_outputs(919)) and (layer0_outputs(2777)));
    layer1_outputs(4991) <= '1';
    layer1_outputs(4992) <= not((layer0_outputs(181)) or (layer0_outputs(2333)));
    layer1_outputs(4993) <= not(layer0_outputs(3508));
    layer1_outputs(4994) <= layer0_outputs(3888);
    layer1_outputs(4995) <= layer0_outputs(3138);
    layer1_outputs(4996) <= layer0_outputs(582);
    layer1_outputs(4997) <= not(layer0_outputs(4343));
    layer1_outputs(4998) <= not(layer0_outputs(1246));
    layer1_outputs(4999) <= (layer0_outputs(2597)) or (layer0_outputs(693));
    layer1_outputs(5000) <= '1';
    layer1_outputs(5001) <= (layer0_outputs(667)) and not (layer0_outputs(343));
    layer1_outputs(5002) <= (layer0_outputs(1301)) or (layer0_outputs(225));
    layer1_outputs(5003) <= layer0_outputs(1522);
    layer1_outputs(5004) <= (layer0_outputs(4510)) and not (layer0_outputs(4561));
    layer1_outputs(5005) <= layer0_outputs(1105);
    layer1_outputs(5006) <= layer0_outputs(3159);
    layer1_outputs(5007) <= (layer0_outputs(549)) and not (layer0_outputs(1480));
    layer1_outputs(5008) <= (layer0_outputs(3632)) or (layer0_outputs(168));
    layer1_outputs(5009) <= layer0_outputs(4827);
    layer1_outputs(5010) <= (layer0_outputs(3154)) and not (layer0_outputs(4871));
    layer1_outputs(5011) <= layer0_outputs(4335);
    layer1_outputs(5012) <= not(layer0_outputs(2807));
    layer1_outputs(5013) <= layer0_outputs(2532);
    layer1_outputs(5014) <= (layer0_outputs(3517)) and not (layer0_outputs(3343));
    layer1_outputs(5015) <= not(layer0_outputs(1735)) or (layer0_outputs(4722));
    layer1_outputs(5016) <= not(layer0_outputs(2792));
    layer1_outputs(5017) <= not((layer0_outputs(1201)) xor (layer0_outputs(2178)));
    layer1_outputs(5018) <= not(layer0_outputs(364));
    layer1_outputs(5019) <= (layer0_outputs(4880)) and not (layer0_outputs(4638));
    layer1_outputs(5020) <= not(layer0_outputs(4096));
    layer1_outputs(5021) <= layer0_outputs(136);
    layer1_outputs(5022) <= not(layer0_outputs(22));
    layer1_outputs(5023) <= (layer0_outputs(2757)) and not (layer0_outputs(574));
    layer1_outputs(5024) <= layer0_outputs(1018);
    layer1_outputs(5025) <= (layer0_outputs(553)) and (layer0_outputs(3381));
    layer1_outputs(5026) <= not((layer0_outputs(1045)) or (layer0_outputs(4357)));
    layer1_outputs(5027) <= (layer0_outputs(161)) and not (layer0_outputs(316));
    layer1_outputs(5028) <= not((layer0_outputs(3600)) and (layer0_outputs(2495)));
    layer1_outputs(5029) <= not((layer0_outputs(2024)) or (layer0_outputs(3934)));
    layer1_outputs(5030) <= (layer0_outputs(1941)) xor (layer0_outputs(3076));
    layer1_outputs(5031) <= (layer0_outputs(1815)) and (layer0_outputs(3102));
    layer1_outputs(5032) <= not(layer0_outputs(3595));
    layer1_outputs(5033) <= (layer0_outputs(2782)) or (layer0_outputs(4008));
    layer1_outputs(5034) <= layer0_outputs(4231);
    layer1_outputs(5035) <= not(layer0_outputs(1365));
    layer1_outputs(5036) <= (layer0_outputs(4680)) and not (layer0_outputs(2339));
    layer1_outputs(5037) <= not(layer0_outputs(5064));
    layer1_outputs(5038) <= layer0_outputs(1598);
    layer1_outputs(5039) <= (layer0_outputs(4721)) and not (layer0_outputs(847));
    layer1_outputs(5040) <= not(layer0_outputs(4959));
    layer1_outputs(5041) <= not(layer0_outputs(613));
    layer1_outputs(5042) <= (layer0_outputs(622)) and not (layer0_outputs(841));
    layer1_outputs(5043) <= '0';
    layer1_outputs(5044) <= (layer0_outputs(4210)) or (layer0_outputs(990));
    layer1_outputs(5045) <= '1';
    layer1_outputs(5046) <= (layer0_outputs(2572)) and not (layer0_outputs(2787));
    layer1_outputs(5047) <= layer0_outputs(1954);
    layer1_outputs(5048) <= layer0_outputs(2864);
    layer1_outputs(5049) <= not(layer0_outputs(477));
    layer1_outputs(5050) <= layer0_outputs(2746);
    layer1_outputs(5051) <= layer0_outputs(4613);
    layer1_outputs(5052) <= not(layer0_outputs(2026)) or (layer0_outputs(2157));
    layer1_outputs(5053) <= not((layer0_outputs(4049)) or (layer0_outputs(2059)));
    layer1_outputs(5054) <= not((layer0_outputs(3041)) or (layer0_outputs(4067)));
    layer1_outputs(5055) <= not(layer0_outputs(4063)) or (layer0_outputs(1761));
    layer1_outputs(5056) <= not(layer0_outputs(2176));
    layer1_outputs(5057) <= (layer0_outputs(4834)) and not (layer0_outputs(1846));
    layer1_outputs(5058) <= layer0_outputs(4122);
    layer1_outputs(5059) <= not(layer0_outputs(1520));
    layer1_outputs(5060) <= '0';
    layer1_outputs(5061) <= not(layer0_outputs(86));
    layer1_outputs(5062) <= layer0_outputs(1849);
    layer1_outputs(5063) <= layer0_outputs(4933);
    layer1_outputs(5064) <= layer0_outputs(2762);
    layer1_outputs(5065) <= (layer0_outputs(1924)) and not (layer0_outputs(3795));
    layer1_outputs(5066) <= layer0_outputs(1929);
    layer1_outputs(5067) <= not(layer0_outputs(4654));
    layer1_outputs(5068) <= not((layer0_outputs(2461)) or (layer0_outputs(1468)));
    layer1_outputs(5069) <= (layer0_outputs(909)) or (layer0_outputs(4568));
    layer1_outputs(5070) <= not(layer0_outputs(2351));
    layer1_outputs(5071) <= (layer0_outputs(3026)) or (layer0_outputs(403));
    layer1_outputs(5072) <= not(layer0_outputs(4957));
    layer1_outputs(5073) <= layer0_outputs(4565);
    layer1_outputs(5074) <= (layer0_outputs(1636)) and not (layer0_outputs(2086));
    layer1_outputs(5075) <= '1';
    layer1_outputs(5076) <= (layer0_outputs(1501)) and (layer0_outputs(295));
    layer1_outputs(5077) <= not((layer0_outputs(2480)) xor (layer0_outputs(3491)));
    layer1_outputs(5078) <= not(layer0_outputs(1755));
    layer1_outputs(5079) <= not(layer0_outputs(2445)) or (layer0_outputs(4242));
    layer1_outputs(5080) <= not(layer0_outputs(303));
    layer1_outputs(5081) <= layer0_outputs(4359);
    layer1_outputs(5082) <= (layer0_outputs(4817)) xor (layer0_outputs(3063));
    layer1_outputs(5083) <= not(layer0_outputs(381)) or (layer0_outputs(4350));
    layer1_outputs(5084) <= not(layer0_outputs(1566));
    layer1_outputs(5085) <= not(layer0_outputs(3991)) or (layer0_outputs(1530));
    layer1_outputs(5086) <= (layer0_outputs(2916)) and (layer0_outputs(1626));
    layer1_outputs(5087) <= not(layer0_outputs(1959));
    layer1_outputs(5088) <= (layer0_outputs(2177)) and not (layer0_outputs(1228));
    layer1_outputs(5089) <= layer0_outputs(10);
    layer1_outputs(5090) <= (layer0_outputs(5103)) or (layer0_outputs(88));
    layer1_outputs(5091) <= (layer0_outputs(4954)) and not (layer0_outputs(4204));
    layer1_outputs(5092) <= '1';
    layer1_outputs(5093) <= layer0_outputs(1134);
    layer1_outputs(5094) <= not(layer0_outputs(2959)) or (layer0_outputs(1207));
    layer1_outputs(5095) <= not(layer0_outputs(2044));
    layer1_outputs(5096) <= layer0_outputs(1869);
    layer1_outputs(5097) <= not(layer0_outputs(4102));
    layer1_outputs(5098) <= layer0_outputs(410);
    layer1_outputs(5099) <= not(layer0_outputs(2328));
    layer1_outputs(5100) <= layer0_outputs(3224);
    layer1_outputs(5101) <= layer0_outputs(701);
    layer1_outputs(5102) <= not((layer0_outputs(1368)) and (layer0_outputs(3504)));
    layer1_outputs(5103) <= not((layer0_outputs(4109)) xor (layer0_outputs(1983)));
    layer1_outputs(5104) <= not(layer0_outputs(2805)) or (layer0_outputs(2821));
    layer1_outputs(5105) <= not(layer0_outputs(2531)) or (layer0_outputs(832));
    layer1_outputs(5106) <= not((layer0_outputs(2874)) or (layer0_outputs(5109)));
    layer1_outputs(5107) <= not(layer0_outputs(3391)) or (layer0_outputs(3118));
    layer1_outputs(5108) <= not(layer0_outputs(2254));
    layer1_outputs(5109) <= (layer0_outputs(416)) and not (layer0_outputs(2468));
    layer1_outputs(5110) <= (layer0_outputs(3865)) or (layer0_outputs(935));
    layer1_outputs(5111) <= not(layer0_outputs(1063));
    layer1_outputs(5112) <= not(layer0_outputs(1986));
    layer1_outputs(5113) <= not((layer0_outputs(1558)) and (layer0_outputs(19)));
    layer1_outputs(5114) <= (layer0_outputs(313)) and not (layer0_outputs(1611));
    layer1_outputs(5115) <= (layer0_outputs(501)) and not (layer0_outputs(4492));
    layer1_outputs(5116) <= (layer0_outputs(2784)) xor (layer0_outputs(995));
    layer1_outputs(5117) <= not(layer0_outputs(1484));
    layer1_outputs(5118) <= layer0_outputs(1870);
    layer1_outputs(5119) <= (layer0_outputs(1853)) and not (layer0_outputs(3147));
    layer2_outputs(0) <= (layer1_outputs(1812)) or (layer1_outputs(109));
    layer2_outputs(1) <= layer1_outputs(4927);
    layer2_outputs(2) <= (layer1_outputs(166)) and not (layer1_outputs(3865));
    layer2_outputs(3) <= (layer1_outputs(3210)) xor (layer1_outputs(335));
    layer2_outputs(4) <= not(layer1_outputs(2434));
    layer2_outputs(5) <= (layer1_outputs(4796)) xor (layer1_outputs(4732));
    layer2_outputs(6) <= (layer1_outputs(3513)) and (layer1_outputs(1076));
    layer2_outputs(7) <= (layer1_outputs(3110)) and not (layer1_outputs(2184));
    layer2_outputs(8) <= not(layer1_outputs(3746)) or (layer1_outputs(2245));
    layer2_outputs(9) <= layer1_outputs(4231);
    layer2_outputs(10) <= layer1_outputs(839);
    layer2_outputs(11) <= '0';
    layer2_outputs(12) <= '0';
    layer2_outputs(13) <= not(layer1_outputs(5029));
    layer2_outputs(14) <= not(layer1_outputs(1275)) or (layer1_outputs(4553));
    layer2_outputs(15) <= not(layer1_outputs(4239)) or (layer1_outputs(21));
    layer2_outputs(16) <= (layer1_outputs(3015)) or (layer1_outputs(2651));
    layer2_outputs(17) <= not((layer1_outputs(4142)) or (layer1_outputs(2279)));
    layer2_outputs(18) <= not(layer1_outputs(1585));
    layer2_outputs(19) <= not(layer1_outputs(902));
    layer2_outputs(20) <= layer1_outputs(1129);
    layer2_outputs(21) <= (layer1_outputs(263)) and (layer1_outputs(1965));
    layer2_outputs(22) <= not(layer1_outputs(3796)) or (layer1_outputs(1868));
    layer2_outputs(23) <= not(layer1_outputs(2484)) or (layer1_outputs(948));
    layer2_outputs(24) <= not((layer1_outputs(1735)) xor (layer1_outputs(2195)));
    layer2_outputs(25) <= not(layer1_outputs(3380)) or (layer1_outputs(2740));
    layer2_outputs(26) <= (layer1_outputs(1432)) or (layer1_outputs(5031));
    layer2_outputs(27) <= '1';
    layer2_outputs(28) <= not(layer1_outputs(2270));
    layer2_outputs(29) <= (layer1_outputs(1950)) and (layer1_outputs(1163));
    layer2_outputs(30) <= (layer1_outputs(4407)) or (layer1_outputs(3118));
    layer2_outputs(31) <= layer1_outputs(4298);
    layer2_outputs(32) <= not(layer1_outputs(4306));
    layer2_outputs(33) <= (layer1_outputs(3712)) or (layer1_outputs(2549));
    layer2_outputs(34) <= (layer1_outputs(3662)) and not (layer1_outputs(4882));
    layer2_outputs(35) <= not(layer1_outputs(134)) or (layer1_outputs(1886));
    layer2_outputs(36) <= not(layer1_outputs(685));
    layer2_outputs(37) <= layer1_outputs(2596);
    layer2_outputs(38) <= (layer1_outputs(2916)) and not (layer1_outputs(1632));
    layer2_outputs(39) <= layer1_outputs(3562);
    layer2_outputs(40) <= not(layer1_outputs(2638));
    layer2_outputs(41) <= not((layer1_outputs(3039)) and (layer1_outputs(1930)));
    layer2_outputs(42) <= layer1_outputs(3384);
    layer2_outputs(43) <= not((layer1_outputs(3042)) xor (layer1_outputs(4487)));
    layer2_outputs(44) <= not(layer1_outputs(3190)) or (layer1_outputs(3650));
    layer2_outputs(45) <= layer1_outputs(347);
    layer2_outputs(46) <= not(layer1_outputs(4973));
    layer2_outputs(47) <= (layer1_outputs(2618)) and not (layer1_outputs(492));
    layer2_outputs(48) <= not((layer1_outputs(2903)) or (layer1_outputs(833)));
    layer2_outputs(49) <= not(layer1_outputs(3553));
    layer2_outputs(50) <= (layer1_outputs(2697)) and not (layer1_outputs(1405));
    layer2_outputs(51) <= layer1_outputs(3057);
    layer2_outputs(52) <= layer1_outputs(1396);
    layer2_outputs(53) <= not(layer1_outputs(1064));
    layer2_outputs(54) <= not((layer1_outputs(1319)) or (layer1_outputs(384)));
    layer2_outputs(55) <= not(layer1_outputs(1126));
    layer2_outputs(56) <= (layer1_outputs(2969)) or (layer1_outputs(2347));
    layer2_outputs(57) <= layer1_outputs(2771);
    layer2_outputs(58) <= not(layer1_outputs(1648));
    layer2_outputs(59) <= not((layer1_outputs(139)) and (layer1_outputs(2025)));
    layer2_outputs(60) <= not((layer1_outputs(4730)) and (layer1_outputs(502)));
    layer2_outputs(61) <= not((layer1_outputs(4532)) and (layer1_outputs(1862)));
    layer2_outputs(62) <= not(layer1_outputs(2215));
    layer2_outputs(63) <= not((layer1_outputs(1594)) xor (layer1_outputs(1409)));
    layer2_outputs(64) <= not(layer1_outputs(3737));
    layer2_outputs(65) <= not(layer1_outputs(4817));
    layer2_outputs(66) <= (layer1_outputs(4237)) or (layer1_outputs(362));
    layer2_outputs(67) <= not(layer1_outputs(4819));
    layer2_outputs(68) <= layer1_outputs(2200);
    layer2_outputs(69) <= layer1_outputs(2608);
    layer2_outputs(70) <= not(layer1_outputs(4955));
    layer2_outputs(71) <= layer1_outputs(2837);
    layer2_outputs(72) <= not(layer1_outputs(5004));
    layer2_outputs(73) <= layer1_outputs(2216);
    layer2_outputs(74) <= layer1_outputs(1875);
    layer2_outputs(75) <= not(layer1_outputs(194));
    layer2_outputs(76) <= not(layer1_outputs(1499));
    layer2_outputs(77) <= not((layer1_outputs(1374)) and (layer1_outputs(2569)));
    layer2_outputs(78) <= not(layer1_outputs(20));
    layer2_outputs(79) <= layer1_outputs(1591);
    layer2_outputs(80) <= not(layer1_outputs(2306)) or (layer1_outputs(1954));
    layer2_outputs(81) <= not((layer1_outputs(1417)) xor (layer1_outputs(2422)));
    layer2_outputs(82) <= layer1_outputs(2304);
    layer2_outputs(83) <= '1';
    layer2_outputs(84) <= not(layer1_outputs(4661));
    layer2_outputs(85) <= layer1_outputs(2060);
    layer2_outputs(86) <= not(layer1_outputs(1200)) or (layer1_outputs(4753));
    layer2_outputs(87) <= layer1_outputs(2837);
    layer2_outputs(88) <= (layer1_outputs(439)) and not (layer1_outputs(3873));
    layer2_outputs(89) <= layer1_outputs(925);
    layer2_outputs(90) <= layer1_outputs(2096);
    layer2_outputs(91) <= layer1_outputs(303);
    layer2_outputs(92) <= not(layer1_outputs(2906)) or (layer1_outputs(4369));
    layer2_outputs(93) <= (layer1_outputs(5041)) or (layer1_outputs(4796));
    layer2_outputs(94) <= '1';
    layer2_outputs(95) <= (layer1_outputs(509)) and not (layer1_outputs(3614));
    layer2_outputs(96) <= not(layer1_outputs(2721));
    layer2_outputs(97) <= not((layer1_outputs(2937)) and (layer1_outputs(3626)));
    layer2_outputs(98) <= not(layer1_outputs(1838));
    layer2_outputs(99) <= not(layer1_outputs(3853));
    layer2_outputs(100) <= layer1_outputs(4474);
    layer2_outputs(101) <= not(layer1_outputs(253));
    layer2_outputs(102) <= layer1_outputs(1778);
    layer2_outputs(103) <= layer1_outputs(1741);
    layer2_outputs(104) <= layer1_outputs(790);
    layer2_outputs(105) <= not(layer1_outputs(2577));
    layer2_outputs(106) <= layer1_outputs(89);
    layer2_outputs(107) <= layer1_outputs(1819);
    layer2_outputs(108) <= not(layer1_outputs(1505));
    layer2_outputs(109) <= not(layer1_outputs(1470));
    layer2_outputs(110) <= not((layer1_outputs(3112)) and (layer1_outputs(4184)));
    layer2_outputs(111) <= not(layer1_outputs(4631));
    layer2_outputs(112) <= not(layer1_outputs(1324));
    layer2_outputs(113) <= layer1_outputs(1142);
    layer2_outputs(114) <= layer1_outputs(363);
    layer2_outputs(115) <= '0';
    layer2_outputs(116) <= not(layer1_outputs(2462));
    layer2_outputs(117) <= not(layer1_outputs(120));
    layer2_outputs(118) <= layer1_outputs(4629);
    layer2_outputs(119) <= layer1_outputs(4897);
    layer2_outputs(120) <= (layer1_outputs(2912)) and not (layer1_outputs(4147));
    layer2_outputs(121) <= not((layer1_outputs(2953)) xor (layer1_outputs(4348)));
    layer2_outputs(122) <= not((layer1_outputs(3800)) xor (layer1_outputs(3923)));
    layer2_outputs(123) <= layer1_outputs(2487);
    layer2_outputs(124) <= not(layer1_outputs(2365)) or (layer1_outputs(1898));
    layer2_outputs(125) <= (layer1_outputs(2643)) and not (layer1_outputs(533));
    layer2_outputs(126) <= not(layer1_outputs(412));
    layer2_outputs(127) <= not(layer1_outputs(1284)) or (layer1_outputs(762));
    layer2_outputs(128) <= layer1_outputs(503);
    layer2_outputs(129) <= not((layer1_outputs(1343)) and (layer1_outputs(1652)));
    layer2_outputs(130) <= not(layer1_outputs(2090));
    layer2_outputs(131) <= (layer1_outputs(115)) and not (layer1_outputs(2188));
    layer2_outputs(132) <= (layer1_outputs(3883)) and not (layer1_outputs(1402));
    layer2_outputs(133) <= (layer1_outputs(261)) and (layer1_outputs(2201));
    layer2_outputs(134) <= layer1_outputs(826);
    layer2_outputs(135) <= layer1_outputs(4719);
    layer2_outputs(136) <= not(layer1_outputs(2174));
    layer2_outputs(137) <= not(layer1_outputs(727));
    layer2_outputs(138) <= not(layer1_outputs(125));
    layer2_outputs(139) <= not(layer1_outputs(3540));
    layer2_outputs(140) <= layer1_outputs(837);
    layer2_outputs(141) <= (layer1_outputs(3843)) and (layer1_outputs(2486));
    layer2_outputs(142) <= '1';
    layer2_outputs(143) <= not(layer1_outputs(3837));
    layer2_outputs(144) <= layer1_outputs(4885);
    layer2_outputs(145) <= (layer1_outputs(2717)) and (layer1_outputs(3474));
    layer2_outputs(146) <= '0';
    layer2_outputs(147) <= not(layer1_outputs(787)) or (layer1_outputs(3694));
    layer2_outputs(148) <= (layer1_outputs(1067)) and not (layer1_outputs(2198));
    layer2_outputs(149) <= not(layer1_outputs(1110)) or (layer1_outputs(2066));
    layer2_outputs(150) <= layer1_outputs(2539);
    layer2_outputs(151) <= (layer1_outputs(2680)) and not (layer1_outputs(1127));
    layer2_outputs(152) <= not(layer1_outputs(3079));
    layer2_outputs(153) <= not(layer1_outputs(2228));
    layer2_outputs(154) <= not(layer1_outputs(3315));
    layer2_outputs(155) <= layer1_outputs(1697);
    layer2_outputs(156) <= layer1_outputs(4672);
    layer2_outputs(157) <= layer1_outputs(2969);
    layer2_outputs(158) <= not((layer1_outputs(817)) xor (layer1_outputs(4768)));
    layer2_outputs(159) <= layer1_outputs(1465);
    layer2_outputs(160) <= not((layer1_outputs(1228)) or (layer1_outputs(2971)));
    layer2_outputs(161) <= not(layer1_outputs(4430));
    layer2_outputs(162) <= not((layer1_outputs(3947)) and (layer1_outputs(4673)));
    layer2_outputs(163) <= not(layer1_outputs(2748));
    layer2_outputs(164) <= not((layer1_outputs(3844)) or (layer1_outputs(945)));
    layer2_outputs(165) <= (layer1_outputs(4933)) or (layer1_outputs(94));
    layer2_outputs(166) <= layer1_outputs(3301);
    layer2_outputs(167) <= layer1_outputs(534);
    layer2_outputs(168) <= not(layer1_outputs(686));
    layer2_outputs(169) <= not(layer1_outputs(273));
    layer2_outputs(170) <= not(layer1_outputs(2836));
    layer2_outputs(171) <= not(layer1_outputs(4596));
    layer2_outputs(172) <= layer1_outputs(1015);
    layer2_outputs(173) <= not(layer1_outputs(3920));
    layer2_outputs(174) <= layer1_outputs(1961);
    layer2_outputs(175) <= not(layer1_outputs(3103)) or (layer1_outputs(1686));
    layer2_outputs(176) <= '0';
    layer2_outputs(177) <= layer1_outputs(1288);
    layer2_outputs(178) <= not(layer1_outputs(3569)) or (layer1_outputs(1776));
    layer2_outputs(179) <= layer1_outputs(458);
    layer2_outputs(180) <= layer1_outputs(4894);
    layer2_outputs(181) <= not(layer1_outputs(4887));
    layer2_outputs(182) <= not(layer1_outputs(3324));
    layer2_outputs(183) <= not(layer1_outputs(1439));
    layer2_outputs(184) <= not(layer1_outputs(3759)) or (layer1_outputs(1588));
    layer2_outputs(185) <= (layer1_outputs(1182)) and (layer1_outputs(3060));
    layer2_outputs(186) <= not(layer1_outputs(1499)) or (layer1_outputs(3871));
    layer2_outputs(187) <= not((layer1_outputs(3425)) or (layer1_outputs(1599)));
    layer2_outputs(188) <= not((layer1_outputs(3276)) or (layer1_outputs(1069)));
    layer2_outputs(189) <= not(layer1_outputs(1186));
    layer2_outputs(190) <= (layer1_outputs(3129)) or (layer1_outputs(3197));
    layer2_outputs(191) <= (layer1_outputs(4384)) and not (layer1_outputs(2978));
    layer2_outputs(192) <= not(layer1_outputs(4309));
    layer2_outputs(193) <= (layer1_outputs(49)) and (layer1_outputs(412));
    layer2_outputs(194) <= layer1_outputs(3256);
    layer2_outputs(195) <= layer1_outputs(423);
    layer2_outputs(196) <= layer1_outputs(1658);
    layer2_outputs(197) <= (layer1_outputs(1639)) and (layer1_outputs(4104));
    layer2_outputs(198) <= not(layer1_outputs(2079));
    layer2_outputs(199) <= (layer1_outputs(4566)) and not (layer1_outputs(2945));
    layer2_outputs(200) <= layer1_outputs(4513);
    layer2_outputs(201) <= not(layer1_outputs(1895));
    layer2_outputs(202) <= not(layer1_outputs(2742)) or (layer1_outputs(4462));
    layer2_outputs(203) <= not(layer1_outputs(4173));
    layer2_outputs(204) <= not(layer1_outputs(954));
    layer2_outputs(205) <= not(layer1_outputs(631));
    layer2_outputs(206) <= (layer1_outputs(2878)) and (layer1_outputs(753));
    layer2_outputs(207) <= not(layer1_outputs(2370));
    layer2_outputs(208) <= '1';
    layer2_outputs(209) <= not(layer1_outputs(1062));
    layer2_outputs(210) <= (layer1_outputs(1530)) or (layer1_outputs(718));
    layer2_outputs(211) <= not((layer1_outputs(1311)) xor (layer1_outputs(151)));
    layer2_outputs(212) <= layer1_outputs(22);
    layer2_outputs(213) <= not(layer1_outputs(2891));
    layer2_outputs(214) <= not(layer1_outputs(1381));
    layer2_outputs(215) <= layer1_outputs(4554);
    layer2_outputs(216) <= not(layer1_outputs(3382));
    layer2_outputs(217) <= (layer1_outputs(1298)) and (layer1_outputs(2439));
    layer2_outputs(218) <= layer1_outputs(991);
    layer2_outputs(219) <= (layer1_outputs(3112)) xor (layer1_outputs(1885));
    layer2_outputs(220) <= not(layer1_outputs(3801)) or (layer1_outputs(1003));
    layer2_outputs(221) <= layer1_outputs(2065);
    layer2_outputs(222) <= layer1_outputs(3778);
    layer2_outputs(223) <= layer1_outputs(1195);
    layer2_outputs(224) <= (layer1_outputs(3407)) xor (layer1_outputs(2641));
    layer2_outputs(225) <= not(layer1_outputs(819));
    layer2_outputs(226) <= layer1_outputs(2447);
    layer2_outputs(227) <= layer1_outputs(4677);
    layer2_outputs(228) <= not(layer1_outputs(1573)) or (layer1_outputs(307));
    layer2_outputs(229) <= not(layer1_outputs(454)) or (layer1_outputs(67));
    layer2_outputs(230) <= not(layer1_outputs(799)) or (layer1_outputs(1357));
    layer2_outputs(231) <= (layer1_outputs(1571)) and not (layer1_outputs(3566));
    layer2_outputs(232) <= (layer1_outputs(3251)) or (layer1_outputs(3853));
    layer2_outputs(233) <= not(layer1_outputs(2746));
    layer2_outputs(234) <= not(layer1_outputs(2802));
    layer2_outputs(235) <= (layer1_outputs(99)) or (layer1_outputs(2912));
    layer2_outputs(236) <= not(layer1_outputs(2498));
    layer2_outputs(237) <= not(layer1_outputs(1763));
    layer2_outputs(238) <= not(layer1_outputs(4381));
    layer2_outputs(239) <= not(layer1_outputs(4396)) or (layer1_outputs(526));
    layer2_outputs(240) <= layer1_outputs(538);
    layer2_outputs(241) <= (layer1_outputs(113)) or (layer1_outputs(2063));
    layer2_outputs(242) <= (layer1_outputs(5058)) or (layer1_outputs(1572));
    layer2_outputs(243) <= layer1_outputs(3714);
    layer2_outputs(244) <= layer1_outputs(950);
    layer2_outputs(245) <= not(layer1_outputs(2687));
    layer2_outputs(246) <= not(layer1_outputs(1912));
    layer2_outputs(247) <= '1';
    layer2_outputs(248) <= layer1_outputs(4905);
    layer2_outputs(249) <= layer1_outputs(678);
    layer2_outputs(250) <= not(layer1_outputs(3710));
    layer2_outputs(251) <= not(layer1_outputs(3044));
    layer2_outputs(252) <= not(layer1_outputs(1773));
    layer2_outputs(253) <= '0';
    layer2_outputs(254) <= not(layer1_outputs(4474)) or (layer1_outputs(3482));
    layer2_outputs(255) <= layer1_outputs(2892);
    layer2_outputs(256) <= layer1_outputs(3055);
    layer2_outputs(257) <= layer1_outputs(3050);
    layer2_outputs(258) <= (layer1_outputs(2888)) and (layer1_outputs(114));
    layer2_outputs(259) <= (layer1_outputs(2420)) xor (layer1_outputs(3296));
    layer2_outputs(260) <= not(layer1_outputs(4028));
    layer2_outputs(261) <= (layer1_outputs(2290)) and not (layer1_outputs(320));
    layer2_outputs(262) <= not(layer1_outputs(4133));
    layer2_outputs(263) <= not(layer1_outputs(2040)) or (layer1_outputs(4169));
    layer2_outputs(264) <= not(layer1_outputs(534));
    layer2_outputs(265) <= layer1_outputs(453);
    layer2_outputs(266) <= not(layer1_outputs(3067));
    layer2_outputs(267) <= layer1_outputs(3205);
    layer2_outputs(268) <= layer1_outputs(3176);
    layer2_outputs(269) <= layer1_outputs(3515);
    layer2_outputs(270) <= layer1_outputs(4116);
    layer2_outputs(271) <= layer1_outputs(2993);
    layer2_outputs(272) <= layer1_outputs(2726);
    layer2_outputs(273) <= not(layer1_outputs(741));
    layer2_outputs(274) <= not((layer1_outputs(3624)) or (layer1_outputs(3911)));
    layer2_outputs(275) <= layer1_outputs(497);
    layer2_outputs(276) <= not(layer1_outputs(3036));
    layer2_outputs(277) <= not(layer1_outputs(4192)) or (layer1_outputs(3487));
    layer2_outputs(278) <= (layer1_outputs(508)) and not (layer1_outputs(613));
    layer2_outputs(279) <= not(layer1_outputs(1281));
    layer2_outputs(280) <= not(layer1_outputs(2132));
    layer2_outputs(281) <= (layer1_outputs(3635)) and not (layer1_outputs(1257));
    layer2_outputs(282) <= layer1_outputs(4029);
    layer2_outputs(283) <= not(layer1_outputs(971));
    layer2_outputs(284) <= not((layer1_outputs(1006)) and (layer1_outputs(2571)));
    layer2_outputs(285) <= not(layer1_outputs(3383));
    layer2_outputs(286) <= layer1_outputs(1846);
    layer2_outputs(287) <= not(layer1_outputs(5068));
    layer2_outputs(288) <= not(layer1_outputs(4567));
    layer2_outputs(289) <= not((layer1_outputs(769)) or (layer1_outputs(322)));
    layer2_outputs(290) <= (layer1_outputs(864)) or (layer1_outputs(3827));
    layer2_outputs(291) <= layer1_outputs(4454);
    layer2_outputs(292) <= not((layer1_outputs(1326)) or (layer1_outputs(16)));
    layer2_outputs(293) <= not(layer1_outputs(4086));
    layer2_outputs(294) <= not((layer1_outputs(3930)) and (layer1_outputs(177)));
    layer2_outputs(295) <= (layer1_outputs(329)) and not (layer1_outputs(4439));
    layer2_outputs(296) <= layer1_outputs(2110);
    layer2_outputs(297) <= not(layer1_outputs(2767));
    layer2_outputs(298) <= not(layer1_outputs(1971)) or (layer1_outputs(3288));
    layer2_outputs(299) <= layer1_outputs(2190);
    layer2_outputs(300) <= not(layer1_outputs(1213));
    layer2_outputs(301) <= (layer1_outputs(3201)) and not (layer1_outputs(2694));
    layer2_outputs(302) <= (layer1_outputs(1219)) and (layer1_outputs(1938));
    layer2_outputs(303) <= (layer1_outputs(2792)) or (layer1_outputs(4203));
    layer2_outputs(304) <= not(layer1_outputs(1065));
    layer2_outputs(305) <= layer1_outputs(906);
    layer2_outputs(306) <= layer1_outputs(4379);
    layer2_outputs(307) <= not(layer1_outputs(466));
    layer2_outputs(308) <= not((layer1_outputs(1678)) or (layer1_outputs(117)));
    layer2_outputs(309) <= (layer1_outputs(2350)) or (layer1_outputs(311));
    layer2_outputs(310) <= (layer1_outputs(4315)) and not (layer1_outputs(1239));
    layer2_outputs(311) <= not(layer1_outputs(35));
    layer2_outputs(312) <= not((layer1_outputs(2195)) or (layer1_outputs(1662)));
    layer2_outputs(313) <= not(layer1_outputs(931));
    layer2_outputs(314) <= not(layer1_outputs(4299)) or (layer1_outputs(3752));
    layer2_outputs(315) <= not((layer1_outputs(1454)) or (layer1_outputs(2286)));
    layer2_outputs(316) <= not((layer1_outputs(885)) xor (layer1_outputs(2964)));
    layer2_outputs(317) <= not(layer1_outputs(3536));
    layer2_outputs(318) <= layer1_outputs(80);
    layer2_outputs(319) <= not((layer1_outputs(4113)) and (layer1_outputs(638)));
    layer2_outputs(320) <= not(layer1_outputs(1594)) or (layer1_outputs(4594));
    layer2_outputs(321) <= '1';
    layer2_outputs(322) <= layer1_outputs(245);
    layer2_outputs(323) <= not(layer1_outputs(2627));
    layer2_outputs(324) <= (layer1_outputs(1124)) and not (layer1_outputs(3818));
    layer2_outputs(325) <= (layer1_outputs(963)) and not (layer1_outputs(3453));
    layer2_outputs(326) <= (layer1_outputs(1961)) and (layer1_outputs(185));
    layer2_outputs(327) <= not(layer1_outputs(4929));
    layer2_outputs(328) <= not(layer1_outputs(1045));
    layer2_outputs(329) <= not((layer1_outputs(1916)) or (layer1_outputs(2375)));
    layer2_outputs(330) <= (layer1_outputs(1041)) and not (layer1_outputs(1974));
    layer2_outputs(331) <= not((layer1_outputs(4131)) xor (layer1_outputs(3062)));
    layer2_outputs(332) <= not(layer1_outputs(4459));
    layer2_outputs(333) <= not((layer1_outputs(3027)) and (layer1_outputs(3343)));
    layer2_outputs(334) <= layer1_outputs(3520);
    layer2_outputs(335) <= (layer1_outputs(1094)) and not (layer1_outputs(4690));
    layer2_outputs(336) <= layer1_outputs(4212);
    layer2_outputs(337) <= not(layer1_outputs(93));
    layer2_outputs(338) <= not((layer1_outputs(972)) and (layer1_outputs(1473)));
    layer2_outputs(339) <= (layer1_outputs(3665)) or (layer1_outputs(729));
    layer2_outputs(340) <= layer1_outputs(4828);
    layer2_outputs(341) <= not(layer1_outputs(2444));
    layer2_outputs(342) <= not(layer1_outputs(4865));
    layer2_outputs(343) <= not((layer1_outputs(4820)) and (layer1_outputs(2666)));
    layer2_outputs(344) <= not(layer1_outputs(2283));
    layer2_outputs(345) <= layer1_outputs(4918);
    layer2_outputs(346) <= layer1_outputs(1285);
    layer2_outputs(347) <= layer1_outputs(768);
    layer2_outputs(348) <= not((layer1_outputs(695)) xor (layer1_outputs(4529)));
    layer2_outputs(349) <= not(layer1_outputs(1270));
    layer2_outputs(350) <= layer1_outputs(1915);
    layer2_outputs(351) <= layer1_outputs(756);
    layer2_outputs(352) <= layer1_outputs(3554);
    layer2_outputs(353) <= not(layer1_outputs(2763));
    layer2_outputs(354) <= (layer1_outputs(353)) and not (layer1_outputs(2221));
    layer2_outputs(355) <= not((layer1_outputs(3974)) and (layer1_outputs(1230)));
    layer2_outputs(356) <= layer1_outputs(3455);
    layer2_outputs(357) <= not(layer1_outputs(1887));
    layer2_outputs(358) <= layer1_outputs(4431);
    layer2_outputs(359) <= not(layer1_outputs(3146));
    layer2_outputs(360) <= not((layer1_outputs(2316)) or (layer1_outputs(1869)));
    layer2_outputs(361) <= not(layer1_outputs(65));
    layer2_outputs(362) <= layer1_outputs(1739);
    layer2_outputs(363) <= not(layer1_outputs(1577)) or (layer1_outputs(1444));
    layer2_outputs(364) <= (layer1_outputs(1838)) or (layer1_outputs(4849));
    layer2_outputs(365) <= (layer1_outputs(4555)) and not (layer1_outputs(3570));
    layer2_outputs(366) <= not(layer1_outputs(3095));
    layer2_outputs(367) <= not(layer1_outputs(4559));
    layer2_outputs(368) <= (layer1_outputs(466)) and not (layer1_outputs(3848));
    layer2_outputs(369) <= (layer1_outputs(650)) and (layer1_outputs(5014));
    layer2_outputs(370) <= not(layer1_outputs(830)) or (layer1_outputs(1939));
    layer2_outputs(371) <= layer1_outputs(1750);
    layer2_outputs(372) <= not((layer1_outputs(4276)) or (layer1_outputs(521)));
    layer2_outputs(373) <= layer1_outputs(147);
    layer2_outputs(374) <= layer1_outputs(4602);
    layer2_outputs(375) <= (layer1_outputs(3242)) xor (layer1_outputs(4152));
    layer2_outputs(376) <= not(layer1_outputs(749)) or (layer1_outputs(4117));
    layer2_outputs(377) <= not(layer1_outputs(4420)) or (layer1_outputs(1453));
    layer2_outputs(378) <= (layer1_outputs(4616)) and not (layer1_outputs(2715));
    layer2_outputs(379) <= layer1_outputs(4061);
    layer2_outputs(380) <= layer1_outputs(3352);
    layer2_outputs(381) <= layer1_outputs(1205);
    layer2_outputs(382) <= not(layer1_outputs(5004)) or (layer1_outputs(1188));
    layer2_outputs(383) <= (layer1_outputs(132)) and not (layer1_outputs(148));
    layer2_outputs(384) <= layer1_outputs(2115);
    layer2_outputs(385) <= layer1_outputs(2155);
    layer2_outputs(386) <= not(layer1_outputs(2743)) or (layer1_outputs(3085));
    layer2_outputs(387) <= layer1_outputs(4813);
    layer2_outputs(388) <= not(layer1_outputs(429)) or (layer1_outputs(4922));
    layer2_outputs(389) <= not(layer1_outputs(4322));
    layer2_outputs(390) <= not(layer1_outputs(355));
    layer2_outputs(391) <= layer1_outputs(3177);
    layer2_outputs(392) <= (layer1_outputs(5074)) and not (layer1_outputs(846));
    layer2_outputs(393) <= not(layer1_outputs(4634)) or (layer1_outputs(1496));
    layer2_outputs(394) <= layer1_outputs(5057);
    layer2_outputs(395) <= not((layer1_outputs(2326)) or (layer1_outputs(2730)));
    layer2_outputs(396) <= layer1_outputs(2185);
    layer2_outputs(397) <= not(layer1_outputs(211)) or (layer1_outputs(228));
    layer2_outputs(398) <= layer1_outputs(3134);
    layer2_outputs(399) <= not(layer1_outputs(2111)) or (layer1_outputs(1925));
    layer2_outputs(400) <= layer1_outputs(969);
    layer2_outputs(401) <= (layer1_outputs(4974)) and (layer1_outputs(3526));
    layer2_outputs(402) <= (layer1_outputs(1705)) and not (layer1_outputs(4534));
    layer2_outputs(403) <= not(layer1_outputs(668));
    layer2_outputs(404) <= not(layer1_outputs(1696)) or (layer1_outputs(3617));
    layer2_outputs(405) <= (layer1_outputs(465)) or (layer1_outputs(1129));
    layer2_outputs(406) <= not(layer1_outputs(4617));
    layer2_outputs(407) <= not(layer1_outputs(3961)) or (layer1_outputs(4132));
    layer2_outputs(408) <= not(layer1_outputs(1244));
    layer2_outputs(409) <= (layer1_outputs(3128)) and (layer1_outputs(3018));
    layer2_outputs(410) <= layer1_outputs(2949);
    layer2_outputs(411) <= not(layer1_outputs(2368));
    layer2_outputs(412) <= not(layer1_outputs(385)) or (layer1_outputs(3577));
    layer2_outputs(413) <= layer1_outputs(1984);
    layer2_outputs(414) <= (layer1_outputs(474)) and (layer1_outputs(2441));
    layer2_outputs(415) <= not(layer1_outputs(2695)) or (layer1_outputs(101));
    layer2_outputs(416) <= layer1_outputs(2387);
    layer2_outputs(417) <= layer1_outputs(2539);
    layer2_outputs(418) <= layer1_outputs(2898);
    layer2_outputs(419) <= (layer1_outputs(2605)) or (layer1_outputs(3264));
    layer2_outputs(420) <= layer1_outputs(1374);
    layer2_outputs(421) <= not((layer1_outputs(115)) and (layer1_outputs(2312)));
    layer2_outputs(422) <= not(layer1_outputs(1134)) or (layer1_outputs(2007));
    layer2_outputs(423) <= not(layer1_outputs(4857)) or (layer1_outputs(3645));
    layer2_outputs(424) <= not(layer1_outputs(2110));
    layer2_outputs(425) <= not(layer1_outputs(1853));
    layer2_outputs(426) <= not((layer1_outputs(1800)) and (layer1_outputs(2246)));
    layer2_outputs(427) <= not((layer1_outputs(4020)) or (layer1_outputs(1968)));
    layer2_outputs(428) <= (layer1_outputs(3140)) and not (layer1_outputs(1260));
    layer2_outputs(429) <= not(layer1_outputs(2793));
    layer2_outputs(430) <= (layer1_outputs(5001)) or (layer1_outputs(4192));
    layer2_outputs(431) <= (layer1_outputs(874)) and not (layer1_outputs(3615));
    layer2_outputs(432) <= layer1_outputs(2761);
    layer2_outputs(433) <= not(layer1_outputs(696));
    layer2_outputs(434) <= layer1_outputs(2208);
    layer2_outputs(435) <= not((layer1_outputs(2672)) xor (layer1_outputs(197)));
    layer2_outputs(436) <= layer1_outputs(2033);
    layer2_outputs(437) <= not(layer1_outputs(2441)) or (layer1_outputs(4181));
    layer2_outputs(438) <= '0';
    layer2_outputs(439) <= not(layer1_outputs(759)) or (layer1_outputs(13));
    layer2_outputs(440) <= not(layer1_outputs(194));
    layer2_outputs(441) <= layer1_outputs(4909);
    layer2_outputs(442) <= (layer1_outputs(4026)) xor (layer1_outputs(395));
    layer2_outputs(443) <= (layer1_outputs(2839)) and not (layer1_outputs(95));
    layer2_outputs(444) <= not(layer1_outputs(1447));
    layer2_outputs(445) <= layer1_outputs(3495);
    layer2_outputs(446) <= layer1_outputs(2301);
    layer2_outputs(447) <= (layer1_outputs(164)) or (layer1_outputs(1128));
    layer2_outputs(448) <= (layer1_outputs(2193)) or (layer1_outputs(2489));
    layer2_outputs(449) <= not((layer1_outputs(1635)) or (layer1_outputs(2432)));
    layer2_outputs(450) <= not(layer1_outputs(4388)) or (layer1_outputs(2477));
    layer2_outputs(451) <= (layer1_outputs(3240)) or (layer1_outputs(3649));
    layer2_outputs(452) <= not(layer1_outputs(853));
    layer2_outputs(453) <= not((layer1_outputs(1626)) or (layer1_outputs(2654)));
    layer2_outputs(454) <= not(layer1_outputs(1652));
    layer2_outputs(455) <= (layer1_outputs(3544)) and (layer1_outputs(4134));
    layer2_outputs(456) <= layer1_outputs(3954);
    layer2_outputs(457) <= not(layer1_outputs(4671)) or (layer1_outputs(1642));
    layer2_outputs(458) <= (layer1_outputs(2549)) and (layer1_outputs(349));
    layer2_outputs(459) <= not(layer1_outputs(4645));
    layer2_outputs(460) <= not(layer1_outputs(1481));
    layer2_outputs(461) <= layer1_outputs(5072);
    layer2_outputs(462) <= (layer1_outputs(138)) and not (layer1_outputs(3527));
    layer2_outputs(463) <= not(layer1_outputs(4327));
    layer2_outputs(464) <= not((layer1_outputs(4692)) xor (layer1_outputs(3633)));
    layer2_outputs(465) <= not(layer1_outputs(3097));
    layer2_outputs(466) <= '0';
    layer2_outputs(467) <= (layer1_outputs(2756)) and not (layer1_outputs(730));
    layer2_outputs(468) <= not(layer1_outputs(2289)) or (layer1_outputs(542));
    layer2_outputs(469) <= layer1_outputs(3081);
    layer2_outputs(470) <= not(layer1_outputs(3449));
    layer2_outputs(471) <= not((layer1_outputs(1937)) and (layer1_outputs(719)));
    layer2_outputs(472) <= not(layer1_outputs(2327)) or (layer1_outputs(3259));
    layer2_outputs(473) <= not((layer1_outputs(1848)) and (layer1_outputs(1452)));
    layer2_outputs(474) <= not(layer1_outputs(866));
    layer2_outputs(475) <= layer1_outputs(1824);
    layer2_outputs(476) <= not(layer1_outputs(1958)) or (layer1_outputs(3697));
    layer2_outputs(477) <= not(layer1_outputs(4032));
    layer2_outputs(478) <= (layer1_outputs(1723)) and not (layer1_outputs(4168));
    layer2_outputs(479) <= not(layer1_outputs(2570)) or (layer1_outputs(2973));
    layer2_outputs(480) <= layer1_outputs(3811);
    layer2_outputs(481) <= layer1_outputs(964);
    layer2_outputs(482) <= '0';
    layer2_outputs(483) <= not((layer1_outputs(2360)) or (layer1_outputs(3427)));
    layer2_outputs(484) <= not((layer1_outputs(3688)) and (layer1_outputs(3513)));
    layer2_outputs(485) <= not(layer1_outputs(3946));
    layer2_outputs(486) <= layer1_outputs(4581);
    layer2_outputs(487) <= not((layer1_outputs(75)) and (layer1_outputs(505)));
    layer2_outputs(488) <= (layer1_outputs(577)) and (layer1_outputs(5005));
    layer2_outputs(489) <= not(layer1_outputs(3799)) or (layer1_outputs(3838));
    layer2_outputs(490) <= not((layer1_outputs(3982)) xor (layer1_outputs(1243)));
    layer2_outputs(491) <= not(layer1_outputs(520)) or (layer1_outputs(3960));
    layer2_outputs(492) <= not((layer1_outputs(242)) and (layer1_outputs(404)));
    layer2_outputs(493) <= layer1_outputs(4003);
    layer2_outputs(494) <= (layer1_outputs(2826)) and (layer1_outputs(3058));
    layer2_outputs(495) <= not(layer1_outputs(5021)) or (layer1_outputs(1412));
    layer2_outputs(496) <= not((layer1_outputs(3159)) or (layer1_outputs(1610)));
    layer2_outputs(497) <= (layer1_outputs(416)) and not (layer1_outputs(2471));
    layer2_outputs(498) <= not((layer1_outputs(1036)) and (layer1_outputs(3545)));
    layer2_outputs(499) <= layer1_outputs(2800);
    layer2_outputs(500) <= layer1_outputs(1879);
    layer2_outputs(501) <= layer1_outputs(1934);
    layer2_outputs(502) <= (layer1_outputs(676)) and not (layer1_outputs(4625));
    layer2_outputs(503) <= (layer1_outputs(489)) and (layer1_outputs(1721));
    layer2_outputs(504) <= not((layer1_outputs(3953)) or (layer1_outputs(370)));
    layer2_outputs(505) <= not(layer1_outputs(2461));
    layer2_outputs(506) <= not((layer1_outputs(1411)) xor (layer1_outputs(4197)));
    layer2_outputs(507) <= (layer1_outputs(3530)) and not (layer1_outputs(1783));
    layer2_outputs(508) <= layer1_outputs(2092);
    layer2_outputs(509) <= layer1_outputs(319);
    layer2_outputs(510) <= not(layer1_outputs(2815)) or (layer1_outputs(3815));
    layer2_outputs(511) <= (layer1_outputs(3689)) or (layer1_outputs(1339));
    layer2_outputs(512) <= (layer1_outputs(3936)) and not (layer1_outputs(3100));
    layer2_outputs(513) <= not((layer1_outputs(1158)) xor (layer1_outputs(4881)));
    layer2_outputs(514) <= (layer1_outputs(3565)) and not (layer1_outputs(2171));
    layer2_outputs(515) <= not(layer1_outputs(3678)) or (layer1_outputs(1195));
    layer2_outputs(516) <= (layer1_outputs(2500)) and not (layer1_outputs(1816));
    layer2_outputs(517) <= not(layer1_outputs(2609));
    layer2_outputs(518) <= (layer1_outputs(3664)) and not (layer1_outputs(1106));
    layer2_outputs(519) <= (layer1_outputs(1474)) and (layer1_outputs(18));
    layer2_outputs(520) <= (layer1_outputs(3054)) and not (layer1_outputs(3505));
    layer2_outputs(521) <= not((layer1_outputs(5038)) or (layer1_outputs(816)));
    layer2_outputs(522) <= layer1_outputs(3246);
    layer2_outputs(523) <= '1';
    layer2_outputs(524) <= (layer1_outputs(2175)) or (layer1_outputs(3660));
    layer2_outputs(525) <= (layer1_outputs(2962)) and not (layer1_outputs(3479));
    layer2_outputs(526) <= (layer1_outputs(1163)) and not (layer1_outputs(3225));
    layer2_outputs(527) <= (layer1_outputs(2014)) and not (layer1_outputs(2693));
    layer2_outputs(528) <= (layer1_outputs(4698)) and not (layer1_outputs(1462));
    layer2_outputs(529) <= (layer1_outputs(217)) and (layer1_outputs(2861));
    layer2_outputs(530) <= not(layer1_outputs(3374));
    layer2_outputs(531) <= layer1_outputs(951);
    layer2_outputs(532) <= not(layer1_outputs(1178));
    layer2_outputs(533) <= layer1_outputs(1157);
    layer2_outputs(534) <= not((layer1_outputs(5095)) xor (layer1_outputs(2954)));
    layer2_outputs(535) <= (layer1_outputs(2606)) and not (layer1_outputs(3736));
    layer2_outputs(536) <= not(layer1_outputs(2153));
    layer2_outputs(537) <= not(layer1_outputs(4392));
    layer2_outputs(538) <= not((layer1_outputs(3971)) or (layer1_outputs(2509)));
    layer2_outputs(539) <= layer1_outputs(112);
    layer2_outputs(540) <= layer1_outputs(544);
    layer2_outputs(541) <= not(layer1_outputs(1898));
    layer2_outputs(542) <= not((layer1_outputs(1638)) xor (layer1_outputs(3717)));
    layer2_outputs(543) <= (layer1_outputs(19)) and (layer1_outputs(4402));
    layer2_outputs(544) <= not(layer1_outputs(4958));
    layer2_outputs(545) <= not(layer1_outputs(3276));
    layer2_outputs(546) <= not((layer1_outputs(4626)) and (layer1_outputs(828)));
    layer2_outputs(547) <= layer1_outputs(2702);
    layer2_outputs(548) <= (layer1_outputs(2006)) and not (layer1_outputs(271));
    layer2_outputs(549) <= not(layer1_outputs(1121));
    layer2_outputs(550) <= not((layer1_outputs(133)) and (layer1_outputs(623)));
    layer2_outputs(551) <= not(layer1_outputs(3556)) or (layer1_outputs(2760));
    layer2_outputs(552) <= not((layer1_outputs(174)) and (layer1_outputs(3136)));
    layer2_outputs(553) <= (layer1_outputs(2528)) xor (layer1_outputs(20));
    layer2_outputs(554) <= not(layer1_outputs(2795));
    layer2_outputs(555) <= not(layer1_outputs(1524));
    layer2_outputs(556) <= layer1_outputs(5085);
    layer2_outputs(557) <= (layer1_outputs(5056)) or (layer1_outputs(2046));
    layer2_outputs(558) <= not(layer1_outputs(1166)) or (layer1_outputs(5022));
    layer2_outputs(559) <= layer1_outputs(1117);
    layer2_outputs(560) <= layer1_outputs(2986);
    layer2_outputs(561) <= layer1_outputs(1742);
    layer2_outputs(562) <= layer1_outputs(1649);
    layer2_outputs(563) <= layer1_outputs(4950);
    layer2_outputs(564) <= (layer1_outputs(4023)) and not (layer1_outputs(469));
    layer2_outputs(565) <= not(layer1_outputs(4979));
    layer2_outputs(566) <= not((layer1_outputs(448)) xor (layer1_outputs(3792)));
    layer2_outputs(567) <= not(layer1_outputs(671));
    layer2_outputs(568) <= not((layer1_outputs(4866)) xor (layer1_outputs(1864)));
    layer2_outputs(569) <= layer1_outputs(3908);
    layer2_outputs(570) <= (layer1_outputs(3629)) and not (layer1_outputs(2975));
    layer2_outputs(571) <= not((layer1_outputs(2963)) xor (layer1_outputs(846)));
    layer2_outputs(572) <= layer1_outputs(2877);
    layer2_outputs(573) <= layer1_outputs(2132);
    layer2_outputs(574) <= not(layer1_outputs(2738));
    layer2_outputs(575) <= layer1_outputs(2956);
    layer2_outputs(576) <= layer1_outputs(3779);
    layer2_outputs(577) <= not(layer1_outputs(2318));
    layer2_outputs(578) <= layer1_outputs(3129);
    layer2_outputs(579) <= (layer1_outputs(4069)) and not (layer1_outputs(3470));
    layer2_outputs(580) <= not(layer1_outputs(3534));
    layer2_outputs(581) <= layer1_outputs(1338);
    layer2_outputs(582) <= not(layer1_outputs(4573));
    layer2_outputs(583) <= not(layer1_outputs(429));
    layer2_outputs(584) <= not(layer1_outputs(1973));
    layer2_outputs(585) <= not(layer1_outputs(1362));
    layer2_outputs(586) <= not((layer1_outputs(1074)) and (layer1_outputs(728)));
    layer2_outputs(587) <= layer1_outputs(2395);
    layer2_outputs(588) <= not(layer1_outputs(4824));
    layer2_outputs(589) <= layer1_outputs(3423);
    layer2_outputs(590) <= layer1_outputs(167);
    layer2_outputs(591) <= not(layer1_outputs(1038));
    layer2_outputs(592) <= not(layer1_outputs(2644)) or (layer1_outputs(813));
    layer2_outputs(593) <= (layer1_outputs(1282)) or (layer1_outputs(1391));
    layer2_outputs(594) <= not(layer1_outputs(758)) or (layer1_outputs(229));
    layer2_outputs(595) <= not((layer1_outputs(2658)) or (layer1_outputs(2919)));
    layer2_outputs(596) <= layer1_outputs(3202);
    layer2_outputs(597) <= not(layer1_outputs(104));
    layer2_outputs(598) <= not(layer1_outputs(557));
    layer2_outputs(599) <= not(layer1_outputs(4008));
    layer2_outputs(600) <= not(layer1_outputs(1631));
    layer2_outputs(601) <= not(layer1_outputs(1955));
    layer2_outputs(602) <= not(layer1_outputs(1889));
    layer2_outputs(603) <= layer1_outputs(7);
    layer2_outputs(604) <= not(layer1_outputs(4189));
    layer2_outputs(605) <= layer1_outputs(1492);
    layer2_outputs(606) <= layer1_outputs(2514);
    layer2_outputs(607) <= not(layer1_outputs(1689));
    layer2_outputs(608) <= (layer1_outputs(1301)) and not (layer1_outputs(2240));
    layer2_outputs(609) <= layer1_outputs(2146);
    layer2_outputs(610) <= not((layer1_outputs(3669)) or (layer1_outputs(4185)));
    layer2_outputs(611) <= layer1_outputs(1822);
    layer2_outputs(612) <= not(layer1_outputs(4670));
    layer2_outputs(613) <= not((layer1_outputs(3932)) and (layer1_outputs(3924)));
    layer2_outputs(614) <= not((layer1_outputs(12)) or (layer1_outputs(2624)));
    layer2_outputs(615) <= not((layer1_outputs(777)) xor (layer1_outputs(3969)));
    layer2_outputs(616) <= not(layer1_outputs(3431)) or (layer1_outputs(545));
    layer2_outputs(617) <= not(layer1_outputs(50));
    layer2_outputs(618) <= layer1_outputs(2761);
    layer2_outputs(619) <= (layer1_outputs(1827)) xor (layer1_outputs(608));
    layer2_outputs(620) <= not(layer1_outputs(856));
    layer2_outputs(621) <= (layer1_outputs(1422)) and (layer1_outputs(3417));
    layer2_outputs(622) <= not(layer1_outputs(1428));
    layer2_outputs(623) <= layer1_outputs(1651);
    layer2_outputs(624) <= layer1_outputs(2592);
    layer2_outputs(625) <= (layer1_outputs(3433)) and not (layer1_outputs(4267));
    layer2_outputs(626) <= not(layer1_outputs(2664)) or (layer1_outputs(352));
    layer2_outputs(627) <= not(layer1_outputs(638));
    layer2_outputs(628) <= (layer1_outputs(3181)) or (layer1_outputs(2414));
    layer2_outputs(629) <= not(layer1_outputs(2382));
    layer2_outputs(630) <= layer1_outputs(2364);
    layer2_outputs(631) <= not((layer1_outputs(1861)) xor (layer1_outputs(1415)));
    layer2_outputs(632) <= (layer1_outputs(4054)) or (layer1_outputs(759));
    layer2_outputs(633) <= not(layer1_outputs(3302));
    layer2_outputs(634) <= (layer1_outputs(1269)) and not (layer1_outputs(2880));
    layer2_outputs(635) <= (layer1_outputs(1302)) or (layer1_outputs(1778));
    layer2_outputs(636) <= layer1_outputs(1459);
    layer2_outputs(637) <= not(layer1_outputs(2133)) or (layer1_outputs(4386));
    layer2_outputs(638) <= not(layer1_outputs(11));
    layer2_outputs(639) <= (layer1_outputs(299)) and (layer1_outputs(4381));
    layer2_outputs(640) <= not(layer1_outputs(2463));
    layer2_outputs(641) <= layer1_outputs(24);
    layer2_outputs(642) <= layer1_outputs(1032);
    layer2_outputs(643) <= not((layer1_outputs(1268)) or (layer1_outputs(482)));
    layer2_outputs(644) <= (layer1_outputs(1839)) and not (layer1_outputs(2292));
    layer2_outputs(645) <= not(layer1_outputs(3521)) or (layer1_outputs(402));
    layer2_outputs(646) <= (layer1_outputs(946)) and not (layer1_outputs(406));
    layer2_outputs(647) <= (layer1_outputs(1714)) or (layer1_outputs(1799));
    layer2_outputs(648) <= not((layer1_outputs(2330)) xor (layer1_outputs(3014)));
    layer2_outputs(649) <= not(layer1_outputs(334));
    layer2_outputs(650) <= (layer1_outputs(2189)) xor (layer1_outputs(3411));
    layer2_outputs(651) <= not(layer1_outputs(2209)) or (layer1_outputs(1192));
    layer2_outputs(652) <= (layer1_outputs(5019)) and not (layer1_outputs(1866));
    layer2_outputs(653) <= not((layer1_outputs(2900)) and (layer1_outputs(3747)));
    layer2_outputs(654) <= not(layer1_outputs(3000));
    layer2_outputs(655) <= not(layer1_outputs(1944)) or (layer1_outputs(323));
    layer2_outputs(656) <= layer1_outputs(4786);
    layer2_outputs(657) <= not(layer1_outputs(3180));
    layer2_outputs(658) <= not(layer1_outputs(622));
    layer2_outputs(659) <= not(layer1_outputs(560)) or (layer1_outputs(1786));
    layer2_outputs(660) <= layer1_outputs(4596);
    layer2_outputs(661) <= not(layer1_outputs(2973));
    layer2_outputs(662) <= not((layer1_outputs(4639)) and (layer1_outputs(4205)));
    layer2_outputs(663) <= layer1_outputs(2596);
    layer2_outputs(664) <= not(layer1_outputs(3388)) or (layer1_outputs(1953));
    layer2_outputs(665) <= not(layer1_outputs(3200)) or (layer1_outputs(1641));
    layer2_outputs(666) <= not((layer1_outputs(287)) and (layer1_outputs(3953)));
    layer2_outputs(667) <= not(layer1_outputs(1384));
    layer2_outputs(668) <= not((layer1_outputs(3757)) xor (layer1_outputs(2165)));
    layer2_outputs(669) <= (layer1_outputs(751)) and not (layer1_outputs(4668));
    layer2_outputs(670) <= not(layer1_outputs(106));
    layer2_outputs(671) <= not(layer1_outputs(1782));
    layer2_outputs(672) <= layer1_outputs(4272);
    layer2_outputs(673) <= layer1_outputs(1079);
    layer2_outputs(674) <= layer1_outputs(592);
    layer2_outputs(675) <= not(layer1_outputs(259));
    layer2_outputs(676) <= (layer1_outputs(2257)) xor (layer1_outputs(3182));
    layer2_outputs(677) <= not(layer1_outputs(1681));
    layer2_outputs(678) <= layer1_outputs(1921);
    layer2_outputs(679) <= not(layer1_outputs(4091)) or (layer1_outputs(3990));
    layer2_outputs(680) <= layer1_outputs(3489);
    layer2_outputs(681) <= not((layer1_outputs(5072)) and (layer1_outputs(4215)));
    layer2_outputs(682) <= (layer1_outputs(1874)) and (layer1_outputs(328));
    layer2_outputs(683) <= (layer1_outputs(1947)) or (layer1_outputs(4476));
    layer2_outputs(684) <= not(layer1_outputs(2378)) or (layer1_outputs(1061));
    layer2_outputs(685) <= not((layer1_outputs(1606)) and (layer1_outputs(3368)));
    layer2_outputs(686) <= (layer1_outputs(4177)) and not (layer1_outputs(2945));
    layer2_outputs(687) <= layer1_outputs(2928);
    layer2_outputs(688) <= not(layer1_outputs(3243));
    layer2_outputs(689) <= not(layer1_outputs(1772)) or (layer1_outputs(882));
    layer2_outputs(690) <= not((layer1_outputs(4365)) or (layer1_outputs(3636)));
    layer2_outputs(691) <= layer1_outputs(3366);
    layer2_outputs(692) <= not((layer1_outputs(1097)) xor (layer1_outputs(686)));
    layer2_outputs(693) <= layer1_outputs(1420);
    layer2_outputs(694) <= not(layer1_outputs(3487));
    layer2_outputs(695) <= (layer1_outputs(1976)) or (layer1_outputs(313));
    layer2_outputs(696) <= '1';
    layer2_outputs(697) <= (layer1_outputs(4222)) or (layer1_outputs(178));
    layer2_outputs(698) <= not((layer1_outputs(2707)) and (layer1_outputs(4435)));
    layer2_outputs(699) <= not(layer1_outputs(3563));
    layer2_outputs(700) <= not(layer1_outputs(1556));
    layer2_outputs(701) <= (layer1_outputs(4458)) and (layer1_outputs(2752));
    layer2_outputs(702) <= layer1_outputs(1791);
    layer2_outputs(703) <= (layer1_outputs(2310)) and not (layer1_outputs(4794));
    layer2_outputs(704) <= not(layer1_outputs(845)) or (layer1_outputs(2210));
    layer2_outputs(705) <= not(layer1_outputs(4257));
    layer2_outputs(706) <= layer1_outputs(3818);
    layer2_outputs(707) <= layer1_outputs(2833);
    layer2_outputs(708) <= not((layer1_outputs(2247)) or (layer1_outputs(527)));
    layer2_outputs(709) <= layer1_outputs(3052);
    layer2_outputs(710) <= layer1_outputs(657);
    layer2_outputs(711) <= not((layer1_outputs(1925)) or (layer1_outputs(4128)));
    layer2_outputs(712) <= (layer1_outputs(1634)) and not (layer1_outputs(1484));
    layer2_outputs(713) <= not(layer1_outputs(4870)) or (layer1_outputs(2481));
    layer2_outputs(714) <= (layer1_outputs(2858)) and (layer1_outputs(4227));
    layer2_outputs(715) <= layer1_outputs(253);
    layer2_outputs(716) <= not(layer1_outputs(557)) or (layer1_outputs(4748));
    layer2_outputs(717) <= not(layer1_outputs(356));
    layer2_outputs(718) <= not((layer1_outputs(3660)) or (layer1_outputs(2169)));
    layer2_outputs(719) <= not((layer1_outputs(46)) or (layer1_outputs(99)));
    layer2_outputs(720) <= layer1_outputs(2831);
    layer2_outputs(721) <= not((layer1_outputs(831)) and (layer1_outputs(2801)));
    layer2_outputs(722) <= layer1_outputs(4634);
    layer2_outputs(723) <= (layer1_outputs(146)) xor (layer1_outputs(1517));
    layer2_outputs(724) <= not(layer1_outputs(4405));
    layer2_outputs(725) <= not(layer1_outputs(360));
    layer2_outputs(726) <= not(layer1_outputs(4792));
    layer2_outputs(727) <= not((layer1_outputs(149)) xor (layer1_outputs(4123)));
    layer2_outputs(728) <= not(layer1_outputs(2561));
    layer2_outputs(729) <= (layer1_outputs(3779)) or (layer1_outputs(562));
    layer2_outputs(730) <= not((layer1_outputs(4476)) and (layer1_outputs(4427)));
    layer2_outputs(731) <= layer1_outputs(1506);
    layer2_outputs(732) <= not(layer1_outputs(313));
    layer2_outputs(733) <= not(layer1_outputs(1310));
    layer2_outputs(734) <= not(layer1_outputs(4913));
    layer2_outputs(735) <= layer1_outputs(2896);
    layer2_outputs(736) <= layer1_outputs(4987);
    layer2_outputs(737) <= layer1_outputs(3456);
    layer2_outputs(738) <= not((layer1_outputs(3415)) or (layer1_outputs(4304)));
    layer2_outputs(739) <= (layer1_outputs(3001)) and not (layer1_outputs(3842));
    layer2_outputs(740) <= (layer1_outputs(2076)) and (layer1_outputs(2740));
    layer2_outputs(741) <= '0';
    layer2_outputs(742) <= not(layer1_outputs(4607));
    layer2_outputs(743) <= not(layer1_outputs(4094));
    layer2_outputs(744) <= not((layer1_outputs(996)) and (layer1_outputs(4167)));
    layer2_outputs(745) <= layer1_outputs(2238);
    layer2_outputs(746) <= layer1_outputs(4398);
    layer2_outputs(747) <= layer1_outputs(4842);
    layer2_outputs(748) <= (layer1_outputs(4810)) or (layer1_outputs(3459));
    layer2_outputs(749) <= not((layer1_outputs(2206)) xor (layer1_outputs(1455)));
    layer2_outputs(750) <= not((layer1_outputs(1621)) or (layer1_outputs(620)));
    layer2_outputs(751) <= layer1_outputs(4105);
    layer2_outputs(752) <= (layer1_outputs(2894)) and (layer1_outputs(4210));
    layer2_outputs(753) <= (layer1_outputs(2674)) or (layer1_outputs(3727));
    layer2_outputs(754) <= '1';
    layer2_outputs(755) <= not((layer1_outputs(2871)) and (layer1_outputs(1710)));
    layer2_outputs(756) <= not(layer1_outputs(3207));
    layer2_outputs(757) <= not(layer1_outputs(2060)) or (layer1_outputs(2583));
    layer2_outputs(758) <= layer1_outputs(3640);
    layer2_outputs(759) <= not((layer1_outputs(4832)) or (layer1_outputs(3702)));
    layer2_outputs(760) <= not(layer1_outputs(2348));
    layer2_outputs(761) <= not(layer1_outputs(5037));
    layer2_outputs(762) <= not(layer1_outputs(4973));
    layer2_outputs(763) <= (layer1_outputs(1472)) and not (layer1_outputs(4626));
    layer2_outputs(764) <= layer1_outputs(3697);
    layer2_outputs(765) <= layer1_outputs(4720);
    layer2_outputs(766) <= layer1_outputs(3699);
    layer2_outputs(767) <= (layer1_outputs(3939)) and not (layer1_outputs(3651));
    layer2_outputs(768) <= not(layer1_outputs(4660));
    layer2_outputs(769) <= layer1_outputs(4556);
    layer2_outputs(770) <= layer1_outputs(1493);
    layer2_outputs(771) <= not(layer1_outputs(5104)) or (layer1_outputs(4145));
    layer2_outputs(772) <= not(layer1_outputs(809)) or (layer1_outputs(4028));
    layer2_outputs(773) <= layer1_outputs(791);
    layer2_outputs(774) <= layer1_outputs(4923);
    layer2_outputs(775) <= (layer1_outputs(621)) and (layer1_outputs(4014));
    layer2_outputs(776) <= layer1_outputs(4090);
    layer2_outputs(777) <= layer1_outputs(2315);
    layer2_outputs(778) <= not(layer1_outputs(294));
    layer2_outputs(779) <= layer1_outputs(5027);
    layer2_outputs(780) <= not(layer1_outputs(1981));
    layer2_outputs(781) <= layer1_outputs(1815);
    layer2_outputs(782) <= (layer1_outputs(4910)) and not (layer1_outputs(3354));
    layer2_outputs(783) <= not((layer1_outputs(4629)) or (layer1_outputs(4044)));
    layer2_outputs(784) <= (layer1_outputs(3857)) and not (layer1_outputs(3530));
    layer2_outputs(785) <= layer1_outputs(3532);
    layer2_outputs(786) <= not(layer1_outputs(4082));
    layer2_outputs(787) <= layer1_outputs(1000);
    layer2_outputs(788) <= not((layer1_outputs(2595)) and (layer1_outputs(164)));
    layer2_outputs(789) <= not(layer1_outputs(438));
    layer2_outputs(790) <= layer1_outputs(4311);
    layer2_outputs(791) <= not(layer1_outputs(962)) or (layer1_outputs(3253));
    layer2_outputs(792) <= not(layer1_outputs(4972)) or (layer1_outputs(3750));
    layer2_outputs(793) <= (layer1_outputs(4051)) and not (layer1_outputs(2210));
    layer2_outputs(794) <= not(layer1_outputs(1346)) or (layer1_outputs(1732));
    layer2_outputs(795) <= not((layer1_outputs(251)) xor (layer1_outputs(5105)));
    layer2_outputs(796) <= layer1_outputs(2861);
    layer2_outputs(797) <= not((layer1_outputs(2039)) and (layer1_outputs(5106)));
    layer2_outputs(798) <= not(layer1_outputs(1347)) or (layer1_outputs(199));
    layer2_outputs(799) <= not(layer1_outputs(2112));
    layer2_outputs(800) <= not(layer1_outputs(3260)) or (layer1_outputs(3167));
    layer2_outputs(801) <= layer1_outputs(2863);
    layer2_outputs(802) <= not(layer1_outputs(1574));
    layer2_outputs(803) <= layer1_outputs(4536);
    layer2_outputs(804) <= (layer1_outputs(2246)) and (layer1_outputs(2821));
    layer2_outputs(805) <= not(layer1_outputs(1196));
    layer2_outputs(806) <= not(layer1_outputs(3734));
    layer2_outputs(807) <= (layer1_outputs(2447)) and not (layer1_outputs(3133));
    layer2_outputs(808) <= not(layer1_outputs(4005)) or (layer1_outputs(123));
    layer2_outputs(809) <= layer1_outputs(4639);
    layer2_outputs(810) <= not((layer1_outputs(829)) and (layer1_outputs(3330)));
    layer2_outputs(811) <= not(layer1_outputs(1717));
    layer2_outputs(812) <= layer1_outputs(3965);
    layer2_outputs(813) <= not(layer1_outputs(4123));
    layer2_outputs(814) <= not(layer1_outputs(2890));
    layer2_outputs(815) <= layer1_outputs(4341);
    layer2_outputs(816) <= (layer1_outputs(4293)) and not (layer1_outputs(1901));
    layer2_outputs(817) <= not(layer1_outputs(1823)) or (layer1_outputs(3466));
    layer2_outputs(818) <= not((layer1_outputs(3673)) and (layer1_outputs(2884)));
    layer2_outputs(819) <= layer1_outputs(4689);
    layer2_outputs(820) <= (layer1_outputs(41)) and (layer1_outputs(1854));
    layer2_outputs(821) <= not(layer1_outputs(3725)) or (layer1_outputs(2499));
    layer2_outputs(822) <= not(layer1_outputs(3099)) or (layer1_outputs(2131));
    layer2_outputs(823) <= not((layer1_outputs(116)) xor (layer1_outputs(3648)));
    layer2_outputs(824) <= (layer1_outputs(628)) and (layer1_outputs(257));
    layer2_outputs(825) <= not(layer1_outputs(2562));
    layer2_outputs(826) <= not((layer1_outputs(1834)) and (layer1_outputs(4604)));
    layer2_outputs(827) <= (layer1_outputs(1344)) and not (layer1_outputs(4238));
    layer2_outputs(828) <= not((layer1_outputs(2121)) or (layer1_outputs(4176)));
    layer2_outputs(829) <= (layer1_outputs(2529)) or (layer1_outputs(2895));
    layer2_outputs(830) <= not(layer1_outputs(2183));
    layer2_outputs(831) <= not(layer1_outputs(3709));
    layer2_outputs(832) <= layer1_outputs(4439);
    layer2_outputs(833) <= (layer1_outputs(1256)) and (layer1_outputs(304));
    layer2_outputs(834) <= (layer1_outputs(985)) and (layer1_outputs(4108));
    layer2_outputs(835) <= not(layer1_outputs(3600)) or (layer1_outputs(4912));
    layer2_outputs(836) <= not(layer1_outputs(2984)) or (layer1_outputs(3460));
    layer2_outputs(837) <= (layer1_outputs(1554)) and not (layer1_outputs(2053));
    layer2_outputs(838) <= not(layer1_outputs(4854)) or (layer1_outputs(3160));
    layer2_outputs(839) <= layer1_outputs(4999);
    layer2_outputs(840) <= not(layer1_outputs(1104));
    layer2_outputs(841) <= not(layer1_outputs(2419));
    layer2_outputs(842) <= layer1_outputs(1865);
    layer2_outputs(843) <= not(layer1_outputs(1180));
    layer2_outputs(844) <= not(layer1_outputs(4720)) or (layer1_outputs(1286));
    layer2_outputs(845) <= '0';
    layer2_outputs(846) <= not(layer1_outputs(4767));
    layer2_outputs(847) <= not(layer1_outputs(2278));
    layer2_outputs(848) <= not(layer1_outputs(805));
    layer2_outputs(849) <= (layer1_outputs(1288)) and (layer1_outputs(1665));
    layer2_outputs(850) <= not(layer1_outputs(2008)) or (layer1_outputs(135));
    layer2_outputs(851) <= not(layer1_outputs(990)) or (layer1_outputs(2388));
    layer2_outputs(852) <= layer1_outputs(3026);
    layer2_outputs(853) <= not(layer1_outputs(2516));
    layer2_outputs(854) <= layer1_outputs(5081);
    layer2_outputs(855) <= layer1_outputs(1341);
    layer2_outputs(856) <= not(layer1_outputs(4083)) or (layer1_outputs(5025));
    layer2_outputs(857) <= (layer1_outputs(4265)) or (layer1_outputs(1502));
    layer2_outputs(858) <= not((layer1_outputs(4619)) or (layer1_outputs(642)));
    layer2_outputs(859) <= (layer1_outputs(4850)) and (layer1_outputs(2056));
    layer2_outputs(860) <= (layer1_outputs(2463)) and (layer1_outputs(2736));
    layer2_outputs(861) <= layer1_outputs(1553);
    layer2_outputs(862) <= (layer1_outputs(1267)) and not (layer1_outputs(2254));
    layer2_outputs(863) <= not(layer1_outputs(2234)) or (layer1_outputs(1476));
    layer2_outputs(864) <= not(layer1_outputs(4780));
    layer2_outputs(865) <= not(layer1_outputs(1451)) or (layer1_outputs(13));
    layer2_outputs(866) <= not((layer1_outputs(1172)) and (layer1_outputs(293)));
    layer2_outputs(867) <= not(layer1_outputs(2859)) or (layer1_outputs(3364));
    layer2_outputs(868) <= not(layer1_outputs(4545)) or (layer1_outputs(1464));
    layer2_outputs(869) <= (layer1_outputs(628)) and (layer1_outputs(2840));
    layer2_outputs(870) <= not((layer1_outputs(4869)) and (layer1_outputs(2010)));
    layer2_outputs(871) <= not((layer1_outputs(3428)) and (layer1_outputs(209)));
    layer2_outputs(872) <= not(layer1_outputs(1419));
    layer2_outputs(873) <= (layer1_outputs(890)) and not (layer1_outputs(332));
    layer2_outputs(874) <= not(layer1_outputs(316));
    layer2_outputs(875) <= not((layer1_outputs(2051)) and (layer1_outputs(4835)));
    layer2_outputs(876) <= layer1_outputs(2013);
    layer2_outputs(877) <= not(layer1_outputs(4177));
    layer2_outputs(878) <= not(layer1_outputs(671));
    layer2_outputs(879) <= layer1_outputs(1024);
    layer2_outputs(880) <= not(layer1_outputs(4859));
    layer2_outputs(881) <= not(layer1_outputs(1716));
    layer2_outputs(882) <= layer1_outputs(1212);
    layer2_outputs(883) <= not(layer1_outputs(583));
    layer2_outputs(884) <= not(layer1_outputs(4655));
    layer2_outputs(885) <= layer1_outputs(4119);
    layer2_outputs(886) <= '0';
    layer2_outputs(887) <= (layer1_outputs(2157)) and (layer1_outputs(4960));
    layer2_outputs(888) <= layer1_outputs(3215);
    layer2_outputs(889) <= (layer1_outputs(1770)) and (layer1_outputs(5025));
    layer2_outputs(890) <= not(layer1_outputs(1133));
    layer2_outputs(891) <= (layer1_outputs(4522)) xor (layer1_outputs(4675));
    layer2_outputs(892) <= layer1_outputs(4714);
    layer2_outputs(893) <= (layer1_outputs(1724)) xor (layer1_outputs(2834));
    layer2_outputs(894) <= layer1_outputs(3359);
    layer2_outputs(895) <= not((layer1_outputs(1334)) or (layer1_outputs(92)));
    layer2_outputs(896) <= layer1_outputs(4752);
    layer2_outputs(897) <= '0';
    layer2_outputs(898) <= not(layer1_outputs(4191)) or (layer1_outputs(5049));
    layer2_outputs(899) <= '1';
    layer2_outputs(900) <= layer1_outputs(1148);
    layer2_outputs(901) <= not(layer1_outputs(2972));
    layer2_outputs(902) <= (layer1_outputs(1303)) xor (layer1_outputs(4358));
    layer2_outputs(903) <= layer1_outputs(3237);
    layer2_outputs(904) <= (layer1_outputs(3247)) or (layer1_outputs(2444));
    layer2_outputs(905) <= layer1_outputs(2035);
    layer2_outputs(906) <= not(layer1_outputs(3220));
    layer2_outputs(907) <= (layer1_outputs(2338)) or (layer1_outputs(1795));
    layer2_outputs(908) <= not(layer1_outputs(4862)) or (layer1_outputs(361));
    layer2_outputs(909) <= layer1_outputs(64);
    layer2_outputs(910) <= (layer1_outputs(281)) or (layer1_outputs(1423));
    layer2_outputs(911) <= layer1_outputs(4993);
    layer2_outputs(912) <= (layer1_outputs(1537)) and (layer1_outputs(3290));
    layer2_outputs(913) <= not(layer1_outputs(4115)) or (layer1_outputs(5010));
    layer2_outputs(914) <= not(layer1_outputs(1028));
    layer2_outputs(915) <= (layer1_outputs(4574)) and not (layer1_outputs(757));
    layer2_outputs(916) <= (layer1_outputs(3477)) and (layer1_outputs(1072));
    layer2_outputs(917) <= layer1_outputs(2344);
    layer2_outputs(918) <= (layer1_outputs(2509)) and not (layer1_outputs(4368));
    layer2_outputs(919) <= not(layer1_outputs(2383)) or (layer1_outputs(2081));
    layer2_outputs(920) <= not(layer1_outputs(4723)) or (layer1_outputs(3210));
    layer2_outputs(921) <= not(layer1_outputs(2487));
    layer2_outputs(922) <= not(layer1_outputs(1941)) or (layer1_outputs(4146));
    layer2_outputs(923) <= not(layer1_outputs(1053));
    layer2_outputs(924) <= not(layer1_outputs(3084));
    layer2_outputs(925) <= layer1_outputs(3284);
    layer2_outputs(926) <= (layer1_outputs(3348)) and not (layer1_outputs(707));
    layer2_outputs(927) <= (layer1_outputs(4302)) xor (layer1_outputs(4140));
    layer2_outputs(928) <= (layer1_outputs(84)) and not (layer1_outputs(1382));
    layer2_outputs(929) <= layer1_outputs(2982);
    layer2_outputs(930) <= layer1_outputs(1300);
    layer2_outputs(931) <= layer1_outputs(2359);
    layer2_outputs(932) <= not((layer1_outputs(2518)) and (layer1_outputs(2231)));
    layer2_outputs(933) <= (layer1_outputs(2925)) xor (layer1_outputs(3283));
    layer2_outputs(934) <= not(layer1_outputs(2169));
    layer2_outputs(935) <= layer1_outputs(2433);
    layer2_outputs(936) <= '1';
    layer2_outputs(937) <= not((layer1_outputs(4677)) or (layer1_outputs(4302)));
    layer2_outputs(938) <= '0';
    layer2_outputs(939) <= layer1_outputs(3649);
    layer2_outputs(940) <= not(layer1_outputs(4024)) or (layer1_outputs(4265));
    layer2_outputs(941) <= not((layer1_outputs(1023)) or (layer1_outputs(130)));
    layer2_outputs(942) <= layer1_outputs(4298);
    layer2_outputs(943) <= not(layer1_outputs(380)) or (layer1_outputs(3286));
    layer2_outputs(944) <= not((layer1_outputs(1837)) and (layer1_outputs(3754)));
    layer2_outputs(945) <= layer1_outputs(1014);
    layer2_outputs(946) <= not((layer1_outputs(174)) and (layer1_outputs(2808)));
    layer2_outputs(947) <= (layer1_outputs(378)) and not (layer1_outputs(877));
    layer2_outputs(948) <= (layer1_outputs(1236)) xor (layer1_outputs(3667));
    layer2_outputs(949) <= layer1_outputs(4235);
    layer2_outputs(950) <= (layer1_outputs(679)) or (layer1_outputs(4086));
    layer2_outputs(951) <= (layer1_outputs(3653)) or (layer1_outputs(4121));
    layer2_outputs(952) <= not((layer1_outputs(4212)) xor (layer1_outputs(445)));
    layer2_outputs(953) <= layer1_outputs(4016);
    layer2_outputs(954) <= (layer1_outputs(4623)) and (layer1_outputs(4899));
    layer2_outputs(955) <= not(layer1_outputs(3556));
    layer2_outputs(956) <= layer1_outputs(4674);
    layer2_outputs(957) <= not(layer1_outputs(1311));
    layer2_outputs(958) <= layer1_outputs(2367);
    layer2_outputs(959) <= not(layer1_outputs(4500));
    layer2_outputs(960) <= not(layer1_outputs(2704)) or (layer1_outputs(3087));
    layer2_outputs(961) <= not(layer1_outputs(4900));
    layer2_outputs(962) <= not(layer1_outputs(5074));
    layer2_outputs(963) <= not(layer1_outputs(3144));
    layer2_outputs(964) <= layer1_outputs(506);
    layer2_outputs(965) <= (layer1_outputs(889)) or (layer1_outputs(555));
    layer2_outputs(966) <= (layer1_outputs(2956)) and (layer1_outputs(3820));
    layer2_outputs(967) <= not((layer1_outputs(2102)) and (layer1_outputs(3496)));
    layer2_outputs(968) <= not(layer1_outputs(922));
    layer2_outputs(969) <= not(layer1_outputs(4424));
    layer2_outputs(970) <= not((layer1_outputs(949)) and (layer1_outputs(3245)));
    layer2_outputs(971) <= (layer1_outputs(2316)) and not (layer1_outputs(4080));
    layer2_outputs(972) <= not(layer1_outputs(697));
    layer2_outputs(973) <= layer1_outputs(2725);
    layer2_outputs(974) <= layer1_outputs(3502);
    layer2_outputs(975) <= layer1_outputs(1873);
    layer2_outputs(976) <= not(layer1_outputs(4621));
    layer2_outputs(977) <= not(layer1_outputs(4549));
    layer2_outputs(978) <= not(layer1_outputs(3862));
    layer2_outputs(979) <= not((layer1_outputs(3989)) or (layer1_outputs(414)));
    layer2_outputs(980) <= layer1_outputs(2996);
    layer2_outputs(981) <= (layer1_outputs(1878)) and not (layer1_outputs(2309));
    layer2_outputs(982) <= (layer1_outputs(1176)) or (layer1_outputs(874));
    layer2_outputs(983) <= layer1_outputs(3538);
    layer2_outputs(984) <= not((layer1_outputs(2737)) and (layer1_outputs(2183)));
    layer2_outputs(985) <= (layer1_outputs(4485)) and not (layer1_outputs(1869));
    layer2_outputs(986) <= not(layer1_outputs(660));
    layer2_outputs(987) <= (layer1_outputs(2802)) or (layer1_outputs(4828));
    layer2_outputs(988) <= (layer1_outputs(125)) or (layer1_outputs(2319));
    layer2_outputs(989) <= (layer1_outputs(1879)) and not (layer1_outputs(1558));
    layer2_outputs(990) <= not(layer1_outputs(4323)) or (layer1_outputs(937));
    layer2_outputs(991) <= (layer1_outputs(3804)) xor (layer1_outputs(4681));
    layer2_outputs(992) <= layer1_outputs(2944);
    layer2_outputs(993) <= not(layer1_outputs(659));
    layer2_outputs(994) <= not(layer1_outputs(1460));
    layer2_outputs(995) <= '1';
    layer2_outputs(996) <= not(layer1_outputs(5002));
    layer2_outputs(997) <= (layer1_outputs(1031)) xor (layer1_outputs(687));
    layer2_outputs(998) <= not(layer1_outputs(658));
    layer2_outputs(999) <= not(layer1_outputs(3033));
    layer2_outputs(1000) <= not(layer1_outputs(221)) or (layer1_outputs(4997));
    layer2_outputs(1001) <= layer1_outputs(76);
    layer2_outputs(1002) <= not(layer1_outputs(2437));
    layer2_outputs(1003) <= layer1_outputs(1776);
    layer2_outputs(1004) <= not(layer1_outputs(2553)) or (layer1_outputs(3839));
    layer2_outputs(1005) <= not(layer1_outputs(3109));
    layer2_outputs(1006) <= not(layer1_outputs(4856));
    layer2_outputs(1007) <= layer1_outputs(2142);
    layer2_outputs(1008) <= (layer1_outputs(4030)) or (layer1_outputs(4527));
    layer2_outputs(1009) <= (layer1_outputs(4255)) and not (layer1_outputs(233));
    layer2_outputs(1010) <= not(layer1_outputs(180));
    layer2_outputs(1011) <= (layer1_outputs(3457)) xor (layer1_outputs(2608));
    layer2_outputs(1012) <= not(layer1_outputs(5075)) or (layer1_outputs(45));
    layer2_outputs(1013) <= not(layer1_outputs(2313));
    layer2_outputs(1014) <= not((layer1_outputs(1068)) and (layer1_outputs(4791)));
    layer2_outputs(1015) <= not(layer1_outputs(4842));
    layer2_outputs(1016) <= layer1_outputs(3686);
    layer2_outputs(1017) <= (layer1_outputs(4547)) xor (layer1_outputs(876));
    layer2_outputs(1018) <= layer1_outputs(5008);
    layer2_outputs(1019) <= not(layer1_outputs(1159));
    layer2_outputs(1020) <= not((layer1_outputs(141)) and (layer1_outputs(3473)));
    layer2_outputs(1021) <= not(layer1_outputs(4609));
    layer2_outputs(1022) <= (layer1_outputs(3341)) and not (layer1_outputs(4696));
    layer2_outputs(1023) <= not(layer1_outputs(3142));
    layer2_outputs(1024) <= not(layer1_outputs(2482)) or (layer1_outputs(3463));
    layer2_outputs(1025) <= (layer1_outputs(4295)) and not (layer1_outputs(2380));
    layer2_outputs(1026) <= (layer1_outputs(680)) or (layer1_outputs(4248));
    layer2_outputs(1027) <= not(layer1_outputs(1756));
    layer2_outputs(1028) <= layer1_outputs(230);
    layer2_outputs(1029) <= (layer1_outputs(4242)) or (layer1_outputs(2735));
    layer2_outputs(1030) <= not((layer1_outputs(2378)) or (layer1_outputs(1145)));
    layer2_outputs(1031) <= (layer1_outputs(4645)) or (layer1_outputs(647));
    layer2_outputs(1032) <= layer1_outputs(2429);
    layer2_outputs(1033) <= not((layer1_outputs(3579)) and (layer1_outputs(2064)));
    layer2_outputs(1034) <= not(layer1_outputs(1788));
    layer2_outputs(1035) <= (layer1_outputs(5009)) and not (layer1_outputs(5086));
    layer2_outputs(1036) <= not((layer1_outputs(2122)) and (layer1_outputs(4942)));
    layer2_outputs(1037) <= not(layer1_outputs(2827)) or (layer1_outputs(30));
    layer2_outputs(1038) <= layer1_outputs(1754);
    layer2_outputs(1039) <= (layer1_outputs(923)) and not (layer1_outputs(2917));
    layer2_outputs(1040) <= not(layer1_outputs(2374));
    layer2_outputs(1041) <= not((layer1_outputs(918)) and (layer1_outputs(3834)));
    layer2_outputs(1042) <= not(layer1_outputs(699));
    layer2_outputs(1043) <= not(layer1_outputs(1842)) or (layer1_outputs(2894));
    layer2_outputs(1044) <= not(layer1_outputs(263));
    layer2_outputs(1045) <= not(layer1_outputs(2534)) or (layer1_outputs(1397));
    layer2_outputs(1046) <= (layer1_outputs(512)) and (layer1_outputs(1533));
    layer2_outputs(1047) <= not(layer1_outputs(649));
    layer2_outputs(1048) <= not(layer1_outputs(4964));
    layer2_outputs(1049) <= not((layer1_outputs(457)) xor (layer1_outputs(1468)));
    layer2_outputs(1050) <= not(layer1_outputs(4098));
    layer2_outputs(1051) <= not(layer1_outputs(2506)) or (layer1_outputs(4566));
    layer2_outputs(1052) <= layer1_outputs(2580);
    layer2_outputs(1053) <= not(layer1_outputs(808));
    layer2_outputs(1054) <= layer1_outputs(625);
    layer2_outputs(1055) <= not(layer1_outputs(1534)) or (layer1_outputs(2630));
    layer2_outputs(1056) <= not(layer1_outputs(1253)) or (layer1_outputs(3602));
    layer2_outputs(1057) <= (layer1_outputs(4146)) and not (layer1_outputs(1214));
    layer2_outputs(1058) <= (layer1_outputs(2914)) and not (layer1_outputs(2901));
    layer2_outputs(1059) <= (layer1_outputs(3983)) and not (layer1_outputs(3475));
    layer2_outputs(1060) <= layer1_outputs(4819);
    layer2_outputs(1061) <= not((layer1_outputs(1233)) and (layer1_outputs(184)));
    layer2_outputs(1062) <= not(layer1_outputs(3057));
    layer2_outputs(1063) <= layer1_outputs(18);
    layer2_outputs(1064) <= not((layer1_outputs(5036)) and (layer1_outputs(994)));
    layer2_outputs(1065) <= not((layer1_outputs(1309)) and (layer1_outputs(481)));
    layer2_outputs(1066) <= layer1_outputs(2265);
    layer2_outputs(1067) <= (layer1_outputs(1055)) or (layer1_outputs(1277));
    layer2_outputs(1068) <= not(layer1_outputs(2697));
    layer2_outputs(1069) <= layer1_outputs(2669);
    layer2_outputs(1070) <= not(layer1_outputs(1033));
    layer2_outputs(1071) <= layer1_outputs(304);
    layer2_outputs(1072) <= (layer1_outputs(1099)) and not (layer1_outputs(1451));
    layer2_outputs(1073) <= layer1_outputs(3252);
    layer2_outputs(1074) <= (layer1_outputs(4633)) or (layer1_outputs(275));
    layer2_outputs(1075) <= not(layer1_outputs(3674));
    layer2_outputs(1076) <= (layer1_outputs(3406)) and not (layer1_outputs(523));
    layer2_outputs(1077) <= not(layer1_outputs(2752));
    layer2_outputs(1078) <= not(layer1_outputs(3119));
    layer2_outputs(1079) <= (layer1_outputs(2468)) and (layer1_outputs(3564));
    layer2_outputs(1080) <= not(layer1_outputs(1239)) or (layer1_outputs(1429));
    layer2_outputs(1081) <= (layer1_outputs(4768)) xor (layer1_outputs(3283));
    layer2_outputs(1082) <= not(layer1_outputs(1001)) or (layer1_outputs(4777));
    layer2_outputs(1083) <= not(layer1_outputs(3713)) or (layer1_outputs(2399));
    layer2_outputs(1084) <= (layer1_outputs(4100)) or (layer1_outputs(4078));
    layer2_outputs(1085) <= layer1_outputs(4150);
    layer2_outputs(1086) <= not((layer1_outputs(4013)) and (layer1_outputs(1986)));
    layer2_outputs(1087) <= (layer1_outputs(4851)) and (layer1_outputs(3858));
    layer2_outputs(1088) <= not(layer1_outputs(2308)) or (layer1_outputs(1386));
    layer2_outputs(1089) <= (layer1_outputs(610)) or (layer1_outputs(2242));
    layer2_outputs(1090) <= layer1_outputs(1991);
    layer2_outputs(1091) <= (layer1_outputs(2910)) and not (layer1_outputs(4283));
    layer2_outputs(1092) <= not(layer1_outputs(3079));
    layer2_outputs(1093) <= not(layer1_outputs(3294));
    layer2_outputs(1094) <= not(layer1_outputs(1189));
    layer2_outputs(1095) <= (layer1_outputs(1165)) and not (layer1_outputs(1520));
    layer2_outputs(1096) <= not((layer1_outputs(3490)) and (layer1_outputs(1782)));
    layer2_outputs(1097) <= (layer1_outputs(3320)) or (layer1_outputs(2391));
    layer2_outputs(1098) <= layer1_outputs(1077);
    layer2_outputs(1099) <= not(layer1_outputs(1119));
    layer2_outputs(1100) <= (layer1_outputs(3580)) and (layer1_outputs(554));
    layer2_outputs(1101) <= layer1_outputs(2868);
    layer2_outputs(1102) <= not((layer1_outputs(3955)) or (layer1_outputs(2028)));
    layer2_outputs(1103) <= not(layer1_outputs(141));
    layer2_outputs(1104) <= layer1_outputs(4575);
    layer2_outputs(1105) <= not(layer1_outputs(3404));
    layer2_outputs(1106) <= not(layer1_outputs(2225));
    layer2_outputs(1107) <= layer1_outputs(4924);
    layer2_outputs(1108) <= layer1_outputs(3399);
    layer2_outputs(1109) <= not((layer1_outputs(3999)) or (layer1_outputs(4400)));
    layer2_outputs(1110) <= layer1_outputs(2225);
    layer2_outputs(1111) <= not(layer1_outputs(1602));
    layer2_outputs(1112) <= layer1_outputs(4120);
    layer2_outputs(1113) <= layer1_outputs(812);
    layer2_outputs(1114) <= not((layer1_outputs(4892)) and (layer1_outputs(4853)));
    layer2_outputs(1115) <= layer1_outputs(2043);
    layer2_outputs(1116) <= layer1_outputs(2253);
    layer2_outputs(1117) <= (layer1_outputs(4273)) and not (layer1_outputs(742));
    layer2_outputs(1118) <= (layer1_outputs(2665)) or (layer1_outputs(3026));
    layer2_outputs(1119) <= not(layer1_outputs(1997)) or (layer1_outputs(1169));
    layer2_outputs(1120) <= not((layer1_outputs(5033)) or (layer1_outputs(3274)));
    layer2_outputs(1121) <= not(layer1_outputs(2028));
    layer2_outputs(1122) <= not(layer1_outputs(4380));
    layer2_outputs(1123) <= (layer1_outputs(2915)) or (layer1_outputs(351));
    layer2_outputs(1124) <= (layer1_outputs(515)) and not (layer1_outputs(3913));
    layer2_outputs(1125) <= layer1_outputs(2921);
    layer2_outputs(1126) <= (layer1_outputs(849)) or (layer1_outputs(3656));
    layer2_outputs(1127) <= not(layer1_outputs(3333));
    layer2_outputs(1128) <= layer1_outputs(1812);
    layer2_outputs(1129) <= layer1_outputs(4429);
    layer2_outputs(1130) <= not(layer1_outputs(4598));
    layer2_outputs(1131) <= not((layer1_outputs(5070)) xor (layer1_outputs(3076)));
    layer2_outputs(1132) <= not((layer1_outputs(4747)) or (layer1_outputs(2798)));
    layer2_outputs(1133) <= layer1_outputs(3491);
    layer2_outputs(1134) <= not(layer1_outputs(2452)) or (layer1_outputs(2293));
    layer2_outputs(1135) <= not(layer1_outputs(4246));
    layer2_outputs(1136) <= not(layer1_outputs(3350)) or (layer1_outputs(3208));
    layer2_outputs(1137) <= layer1_outputs(2265);
    layer2_outputs(1138) <= not(layer1_outputs(397)) or (layer1_outputs(2691));
    layer2_outputs(1139) <= not(layer1_outputs(4435));
    layer2_outputs(1140) <= (layer1_outputs(858)) and not (layer1_outputs(711));
    layer2_outputs(1141) <= not(layer1_outputs(1658)) or (layer1_outputs(4694));
    layer2_outputs(1142) <= layer1_outputs(1113);
    layer2_outputs(1143) <= layer1_outputs(283);
    layer2_outputs(1144) <= (layer1_outputs(5089)) or (layer1_outputs(1624));
    layer2_outputs(1145) <= layer1_outputs(3434);
    layer2_outputs(1146) <= (layer1_outputs(1222)) or (layer1_outputs(1371));
    layer2_outputs(1147) <= not((layer1_outputs(1687)) xor (layer1_outputs(1391)));
    layer2_outputs(1148) <= layer1_outputs(2749);
    layer2_outputs(1149) <= (layer1_outputs(3250)) xor (layer1_outputs(643));
    layer2_outputs(1150) <= not(layer1_outputs(211));
    layer2_outputs(1151) <= not(layer1_outputs(51));
    layer2_outputs(1152) <= (layer1_outputs(792)) and not (layer1_outputs(1349));
    layer2_outputs(1153) <= (layer1_outputs(1437)) and not (layer1_outputs(44));
    layer2_outputs(1154) <= not((layer1_outputs(4697)) or (layer1_outputs(937)));
    layer2_outputs(1155) <= layer1_outputs(1755);
    layer2_outputs(1156) <= not(layer1_outputs(5081)) or (layer1_outputs(367));
    layer2_outputs(1157) <= (layer1_outputs(19)) and not (layer1_outputs(519));
    layer2_outputs(1158) <= not((layer1_outputs(1306)) xor (layer1_outputs(3003)));
    layer2_outputs(1159) <= not(layer1_outputs(3729)) or (layer1_outputs(705));
    layer2_outputs(1160) <= not(layer1_outputs(873));
    layer2_outputs(1161) <= not((layer1_outputs(4815)) and (layer1_outputs(517)));
    layer2_outputs(1162) <= not(layer1_outputs(237)) or (layer1_outputs(1809));
    layer2_outputs(1163) <= not((layer1_outputs(4096)) or (layer1_outputs(2263)));
    layer2_outputs(1164) <= not((layer1_outputs(6)) xor (layer1_outputs(2926)));
    layer2_outputs(1165) <= layer1_outputs(4623);
    layer2_outputs(1166) <= layer1_outputs(4632);
    layer2_outputs(1167) <= not((layer1_outputs(2326)) and (layer1_outputs(1913)));
    layer2_outputs(1168) <= not((layer1_outputs(1992)) and (layer1_outputs(3641)));
    layer2_outputs(1169) <= (layer1_outputs(3925)) and not (layer1_outputs(2839));
    layer2_outputs(1170) <= not(layer1_outputs(4988));
    layer2_outputs(1171) <= (layer1_outputs(635)) and (layer1_outputs(4148));
    layer2_outputs(1172) <= not(layer1_outputs(4818));
    layer2_outputs(1173) <= not((layer1_outputs(4877)) xor (layer1_outputs(4647)));
    layer2_outputs(1174) <= not(layer1_outputs(38)) or (layer1_outputs(476));
    layer2_outputs(1175) <= (layer1_outputs(2578)) and not (layer1_outputs(1608));
    layer2_outputs(1176) <= not(layer1_outputs(4885));
    layer2_outputs(1177) <= not((layer1_outputs(2349)) and (layer1_outputs(683)));
    layer2_outputs(1178) <= not((layer1_outputs(651)) xor (layer1_outputs(3870)));
    layer2_outputs(1179) <= not(layer1_outputs(311));
    layer2_outputs(1180) <= not(layer1_outputs(1215));
    layer2_outputs(1181) <= not(layer1_outputs(4610));
    layer2_outputs(1182) <= not(layer1_outputs(1854));
    layer2_outputs(1183) <= not(layer1_outputs(1863));
    layer2_outputs(1184) <= (layer1_outputs(366)) and not (layer1_outputs(4360));
    layer2_outputs(1185) <= not((layer1_outputs(123)) or (layer1_outputs(5070)));
    layer2_outputs(1186) <= (layer1_outputs(1008)) and not (layer1_outputs(2148));
    layer2_outputs(1187) <= layer1_outputs(3099);
    layer2_outputs(1188) <= layer1_outputs(378);
    layer2_outputs(1189) <= (layer1_outputs(1631)) or (layer1_outputs(4945));
    layer2_outputs(1190) <= (layer1_outputs(2097)) xor (layer1_outputs(1779));
    layer2_outputs(1191) <= not(layer1_outputs(1212));
    layer2_outputs(1192) <= (layer1_outputs(3825)) or (layer1_outputs(4170));
    layer2_outputs(1193) <= (layer1_outputs(1575)) or (layer1_outputs(1963));
    layer2_outputs(1194) <= layer1_outputs(1137);
    layer2_outputs(1195) <= not(layer1_outputs(4376)) or (layer1_outputs(84));
    layer2_outputs(1196) <= not(layer1_outputs(1674));
    layer2_outputs(1197) <= (layer1_outputs(1897)) and not (layer1_outputs(2576));
    layer2_outputs(1198) <= layer1_outputs(1808);
    layer2_outputs(1199) <= (layer1_outputs(1357)) and not (layer1_outputs(4052));
    layer2_outputs(1200) <= not(layer1_outputs(5036)) or (layer1_outputs(4656));
    layer2_outputs(1201) <= layer1_outputs(3983);
    layer2_outputs(1202) <= layer1_outputs(1565);
    layer2_outputs(1203) <= layer1_outputs(1146);
    layer2_outputs(1204) <= not((layer1_outputs(961)) xor (layer1_outputs(2705)));
    layer2_outputs(1205) <= not(layer1_outputs(2902));
    layer2_outputs(1206) <= '0';
    layer2_outputs(1207) <= not(layer1_outputs(3131));
    layer2_outputs(1208) <= (layer1_outputs(238)) and (layer1_outputs(1583));
    layer2_outputs(1209) <= (layer1_outputs(4556)) or (layer1_outputs(3068));
    layer2_outputs(1210) <= not(layer1_outputs(3492));
    layer2_outputs(1211) <= not(layer1_outputs(420));
    layer2_outputs(1212) <= not(layer1_outputs(2163));
    layer2_outputs(1213) <= not(layer1_outputs(4207));
    layer2_outputs(1214) <= (layer1_outputs(3436)) xor (layer1_outputs(2488));
    layer2_outputs(1215) <= (layer1_outputs(3241)) or (layer1_outputs(924));
    layer2_outputs(1216) <= not(layer1_outputs(1203)) or (layer1_outputs(2777));
    layer2_outputs(1217) <= not(layer1_outputs(4805)) or (layer1_outputs(1749));
    layer2_outputs(1218) <= not(layer1_outputs(1090));
    layer2_outputs(1219) <= not(layer1_outputs(4074)) or (layer1_outputs(2890));
    layer2_outputs(1220) <= layer1_outputs(3373);
    layer2_outputs(1221) <= layer1_outputs(2574);
    layer2_outputs(1222) <= (layer1_outputs(2143)) or (layer1_outputs(3637));
    layer2_outputs(1223) <= (layer1_outputs(3861)) and not (layer1_outputs(1970));
    layer2_outputs(1224) <= (layer1_outputs(3595)) or (layer1_outputs(1548));
    layer2_outputs(1225) <= layer1_outputs(2021);
    layer2_outputs(1226) <= (layer1_outputs(2974)) and (layer1_outputs(2583));
    layer2_outputs(1227) <= not(layer1_outputs(2754));
    layer2_outputs(1228) <= not(layer1_outputs(692)) or (layer1_outputs(4183));
    layer2_outputs(1229) <= layer1_outputs(122);
    layer2_outputs(1230) <= (layer1_outputs(3287)) or (layer1_outputs(3245));
    layer2_outputs(1231) <= not(layer1_outputs(4443));
    layer2_outputs(1232) <= not(layer1_outputs(543));
    layer2_outputs(1233) <= not((layer1_outputs(109)) or (layer1_outputs(267)));
    layer2_outputs(1234) <= (layer1_outputs(4205)) and not (layer1_outputs(801));
    layer2_outputs(1235) <= layer1_outputs(2860);
    layer2_outputs(1236) <= layer1_outputs(2957);
    layer2_outputs(1237) <= not(layer1_outputs(4227));
    layer2_outputs(1238) <= '1';
    layer2_outputs(1239) <= not((layer1_outputs(250)) xor (layer1_outputs(1340)));
    layer2_outputs(1240) <= not((layer1_outputs(701)) or (layer1_outputs(4880)));
    layer2_outputs(1241) <= (layer1_outputs(3315)) or (layer1_outputs(589));
    layer2_outputs(1242) <= (layer1_outputs(2940)) or (layer1_outputs(3387));
    layer2_outputs(1243) <= '0';
    layer2_outputs(1244) <= not(layer1_outputs(2730));
    layer2_outputs(1245) <= layer1_outputs(339);
    layer2_outputs(1246) <= (layer1_outputs(4666)) and (layer1_outputs(540));
    layer2_outputs(1247) <= layer1_outputs(2999);
    layer2_outputs(1248) <= not(layer1_outputs(3782));
    layer2_outputs(1249) <= not(layer1_outputs(2586)) or (layer1_outputs(3860));
    layer2_outputs(1250) <= layer1_outputs(3271);
    layer2_outputs(1251) <= not(layer1_outputs(2590));
    layer2_outputs(1252) <= layer1_outputs(2318);
    layer2_outputs(1253) <= layer1_outputs(3947);
    layer2_outputs(1254) <= not(layer1_outputs(1769)) or (layer1_outputs(421));
    layer2_outputs(1255) <= (layer1_outputs(3910)) and not (layer1_outputs(2747));
    layer2_outputs(1256) <= not(layer1_outputs(1111)) or (layer1_outputs(3867));
    layer2_outputs(1257) <= layer1_outputs(1259);
    layer2_outputs(1258) <= not(layer1_outputs(1725));
    layer2_outputs(1259) <= not((layer1_outputs(4936)) xor (layer1_outputs(2676)));
    layer2_outputs(1260) <= '0';
    layer2_outputs(1261) <= not(layer1_outputs(4210));
    layer2_outputs(1262) <= not(layer1_outputs(2994)) or (layer1_outputs(5077));
    layer2_outputs(1263) <= not(layer1_outputs(3998));
    layer2_outputs(1264) <= (layer1_outputs(2806)) xor (layer1_outputs(3823));
    layer2_outputs(1265) <= not(layer1_outputs(398));
    layer2_outputs(1266) <= (layer1_outputs(3302)) xor (layer1_outputs(2328));
    layer2_outputs(1267) <= not(layer1_outputs(3341));
    layer2_outputs(1268) <= layer1_outputs(3887);
    layer2_outputs(1269) <= not(layer1_outputs(4266));
    layer2_outputs(1270) <= (layer1_outputs(4437)) and not (layer1_outputs(666));
    layer2_outputs(1271) <= not(layer1_outputs(746));
    layer2_outputs(1272) <= not(layer1_outputs(4126));
    layer2_outputs(1273) <= (layer1_outputs(1191)) and (layer1_outputs(946));
    layer2_outputs(1274) <= not(layer1_outputs(1483));
    layer2_outputs(1275) <= not(layer1_outputs(2630));
    layer2_outputs(1276) <= (layer1_outputs(1177)) and (layer1_outputs(2879));
    layer2_outputs(1277) <= not(layer1_outputs(1906));
    layer2_outputs(1278) <= layer1_outputs(880);
    layer2_outputs(1279) <= layer1_outputs(798);
    layer2_outputs(1280) <= (layer1_outputs(3226)) or (layer1_outputs(4878));
    layer2_outputs(1281) <= layer1_outputs(454);
    layer2_outputs(1282) <= not(layer1_outputs(2980));
    layer2_outputs(1283) <= not((layer1_outputs(4077)) or (layer1_outputs(871)));
    layer2_outputs(1284) <= layer1_outputs(2568);
    layer2_outputs(1285) <= (layer1_outputs(3514)) or (layer1_outputs(4217));
    layer2_outputs(1286) <= (layer1_outputs(949)) and (layer1_outputs(4595));
    layer2_outputs(1287) <= not(layer1_outputs(629));
    layer2_outputs(1288) <= not(layer1_outputs(4970));
    layer2_outputs(1289) <= layer1_outputs(3847);
    layer2_outputs(1290) <= not(layer1_outputs(252));
    layer2_outputs(1291) <= not((layer1_outputs(2636)) or (layer1_outputs(2836)));
    layer2_outputs(1292) <= not((layer1_outputs(3666)) or (layer1_outputs(201)));
    layer2_outputs(1293) <= not(layer1_outputs(4662)) or (layer1_outputs(4477));
    layer2_outputs(1294) <= not((layer1_outputs(3575)) and (layer1_outputs(4466)));
    layer2_outputs(1295) <= not(layer1_outputs(1633)) or (layer1_outputs(1229));
    layer2_outputs(1296) <= not((layer1_outputs(4659)) or (layer1_outputs(991)));
    layer2_outputs(1297) <= layer1_outputs(1408);
    layer2_outputs(1298) <= not(layer1_outputs(4727)) or (layer1_outputs(936));
    layer2_outputs(1299) <= (layer1_outputs(4863)) or (layer1_outputs(3574));
    layer2_outputs(1300) <= (layer1_outputs(1605)) xor (layer1_outputs(2490));
    layer2_outputs(1301) <= not(layer1_outputs(4209));
    layer2_outputs(1302) <= (layer1_outputs(2418)) or (layer1_outputs(1098));
    layer2_outputs(1303) <= layer1_outputs(2480);
    layer2_outputs(1304) <= layer1_outputs(4513);
    layer2_outputs(1305) <= not(layer1_outputs(4288));
    layer2_outputs(1306) <= layer1_outputs(2434);
    layer2_outputs(1307) <= not(layer1_outputs(3756)) or (layer1_outputs(4673));
    layer2_outputs(1308) <= not(layer1_outputs(1445)) or (layer1_outputs(1857));
    layer2_outputs(1309) <= (layer1_outputs(5088)) and not (layer1_outputs(2113));
    layer2_outputs(1310) <= layer1_outputs(867);
    layer2_outputs(1311) <= layer1_outputs(1026);
    layer2_outputs(1312) <= not(layer1_outputs(1535));
    layer2_outputs(1313) <= not(layer1_outputs(1589));
    layer2_outputs(1314) <= not(layer1_outputs(1807));
    layer2_outputs(1315) <= not(layer1_outputs(3345)) or (layer1_outputs(550));
    layer2_outputs(1316) <= (layer1_outputs(2059)) or (layer1_outputs(4552));
    layer2_outputs(1317) <= not(layer1_outputs(3885)) or (layer1_outputs(960));
    layer2_outputs(1318) <= not(layer1_outputs(2656));
    layer2_outputs(1319) <= layer1_outputs(1520);
    layer2_outputs(1320) <= not(layer1_outputs(3138));
    layer2_outputs(1321) <= not(layer1_outputs(3476)) or (layer1_outputs(4644));
    layer2_outputs(1322) <= (layer1_outputs(4116)) and not (layer1_outputs(2475));
    layer2_outputs(1323) <= not(layer1_outputs(2338));
    layer2_outputs(1324) <= (layer1_outputs(3400)) xor (layer1_outputs(2144));
    layer2_outputs(1325) <= (layer1_outputs(3817)) and (layer1_outputs(4800));
    layer2_outputs(1326) <= (layer1_outputs(2662)) or (layer1_outputs(1412));
    layer2_outputs(1327) <= layer1_outputs(4459);
    layer2_outputs(1328) <= (layer1_outputs(3407)) and not (layer1_outputs(4147));
    layer2_outputs(1329) <= '0';
    layer2_outputs(1330) <= layer1_outputs(1535);
    layer2_outputs(1331) <= not(layer1_outputs(45));
    layer2_outputs(1332) <= layer1_outputs(3658);
    layer2_outputs(1333) <= layer1_outputs(2461);
    layer2_outputs(1334) <= (layer1_outputs(3017)) or (layer1_outputs(4748));
    layer2_outputs(1335) <= layer1_outputs(3906);
    layer2_outputs(1336) <= (layer1_outputs(1549)) or (layer1_outputs(3608));
    layer2_outputs(1337) <= layer1_outputs(2769);
    layer2_outputs(1338) <= (layer1_outputs(3884)) and (layer1_outputs(3574));
    layer2_outputs(1339) <= (layer1_outputs(2030)) and (layer1_outputs(4635));
    layer2_outputs(1340) <= (layer1_outputs(3317)) and not (layer1_outputs(3397));
    layer2_outputs(1341) <= (layer1_outputs(269)) and not (layer1_outputs(3695));
    layer2_outputs(1342) <= (layer1_outputs(634)) and not (layer1_outputs(3393));
    layer2_outputs(1343) <= not(layer1_outputs(487));
    layer2_outputs(1344) <= not(layer1_outputs(4224));
    layer2_outputs(1345) <= not(layer1_outputs(3662)) or (layer1_outputs(1410));
    layer2_outputs(1346) <= not(layer1_outputs(3219));
    layer2_outputs(1347) <= not(layer1_outputs(4035)) or (layer1_outputs(1909));
    layer2_outputs(1348) <= layer1_outputs(4219);
    layer2_outputs(1349) <= not((layer1_outputs(1222)) xor (layer1_outputs(3029)));
    layer2_outputs(1350) <= not(layer1_outputs(3771));
    layer2_outputs(1351) <= layer1_outputs(945);
    layer2_outputs(1352) <= not(layer1_outputs(3424));
    layer2_outputs(1353) <= not(layer1_outputs(1784));
    layer2_outputs(1354) <= (layer1_outputs(1518)) or (layer1_outputs(1963));
    layer2_outputs(1355) <= layer1_outputs(5095);
    layer2_outputs(1356) <= (layer1_outputs(3731)) and not (layer1_outputs(1820));
    layer2_outputs(1357) <= (layer1_outputs(1004)) and not (layer1_outputs(794));
    layer2_outputs(1358) <= not(layer1_outputs(491));
    layer2_outputs(1359) <= layer1_outputs(5096);
    layer2_outputs(1360) <= not(layer1_outputs(54));
    layer2_outputs(1361) <= not(layer1_outputs(339));
    layer2_outputs(1362) <= layer1_outputs(2294);
    layer2_outputs(1363) <= layer1_outputs(3034);
    layer2_outputs(1364) <= (layer1_outputs(1368)) and not (layer1_outputs(2130));
    layer2_outputs(1365) <= layer1_outputs(1069);
    layer2_outputs(1366) <= not(layer1_outputs(1985));
    layer2_outputs(1367) <= layer1_outputs(2714);
    layer2_outputs(1368) <= not(layer1_outputs(1530));
    layer2_outputs(1369) <= not(layer1_outputs(2087));
    layer2_outputs(1370) <= not((layer1_outputs(4793)) or (layer1_outputs(2930)));
    layer2_outputs(1371) <= layer1_outputs(3178);
    layer2_outputs(1372) <= layer1_outputs(4422);
    layer2_outputs(1373) <= not(layer1_outputs(774));
    layer2_outputs(1374) <= not((layer1_outputs(4576)) or (layer1_outputs(572)));
    layer2_outputs(1375) <= (layer1_outputs(3854)) and not (layer1_outputs(1639));
    layer2_outputs(1376) <= not(layer1_outputs(4413));
    layer2_outputs(1377) <= layer1_outputs(2046);
    layer2_outputs(1378) <= (layer1_outputs(1353)) and (layer1_outputs(2803));
    layer2_outputs(1379) <= not(layer1_outputs(4168));
    layer2_outputs(1380) <= (layer1_outputs(2071)) and (layer1_outputs(2341));
    layer2_outputs(1381) <= not(layer1_outputs(886)) or (layer1_outputs(1078));
    layer2_outputs(1382) <= layer1_outputs(5094);
    layer2_outputs(1383) <= not((layer1_outputs(2664)) xor (layer1_outputs(2285)));
    layer2_outputs(1384) <= layer1_outputs(2877);
    layer2_outputs(1385) <= not(layer1_outputs(1551));
    layer2_outputs(1386) <= not(layer1_outputs(2699)) or (layer1_outputs(715));
    layer2_outputs(1387) <= not(layer1_outputs(2988));
    layer2_outputs(1388) <= layer1_outputs(923);
    layer2_outputs(1389) <= not(layer1_outputs(450)) or (layer1_outputs(4006));
    layer2_outputs(1390) <= not(layer1_outputs(1401));
    layer2_outputs(1391) <= not(layer1_outputs(2251));
    layer2_outputs(1392) <= (layer1_outputs(782)) and (layer1_outputs(4059));
    layer2_outputs(1393) <= not(layer1_outputs(1888)) or (layer1_outputs(3705));
    layer2_outputs(1394) <= '0';
    layer2_outputs(1395) <= (layer1_outputs(4313)) or (layer1_outputs(3115));
    layer2_outputs(1396) <= (layer1_outputs(4343)) and not (layer1_outputs(1071));
    layer2_outputs(1397) <= (layer1_outputs(31)) or (layer1_outputs(1081));
    layer2_outputs(1398) <= not(layer1_outputs(578));
    layer2_outputs(1399) <= (layer1_outputs(694)) or (layer1_outputs(4583));
    layer2_outputs(1400) <= not((layer1_outputs(163)) and (layer1_outputs(3384)));
    layer2_outputs(1401) <= not(layer1_outputs(2085));
    layer2_outputs(1402) <= layer1_outputs(2714);
    layer2_outputs(1403) <= not(layer1_outputs(1188));
    layer2_outputs(1404) <= not((layer1_outputs(56)) xor (layer1_outputs(3900)));
    layer2_outputs(1405) <= not((layer1_outputs(2416)) and (layer1_outputs(1299)));
    layer2_outputs(1406) <= '0';
    layer2_outputs(1407) <= layer1_outputs(4947);
    layer2_outputs(1408) <= not(layer1_outputs(82));
    layer2_outputs(1409) <= (layer1_outputs(3421)) and (layer1_outputs(1904));
    layer2_outputs(1410) <= (layer1_outputs(1567)) or (layer1_outputs(3164));
    layer2_outputs(1411) <= layer1_outputs(117);
    layer2_outputs(1412) <= not(layer1_outputs(2708)) or (layer1_outputs(5100));
    layer2_outputs(1413) <= not(layer1_outputs(2499)) or (layer1_outputs(3588));
    layer2_outputs(1414) <= layer1_outputs(1052);
    layer2_outputs(1415) <= (layer1_outputs(4576)) or (layer1_outputs(4614));
    layer2_outputs(1416) <= not(layer1_outputs(4847)) or (layer1_outputs(4251));
    layer2_outputs(1417) <= (layer1_outputs(2745)) or (layer1_outputs(4546));
    layer2_outputs(1418) <= not(layer1_outputs(3744)) or (layer1_outputs(2959));
    layer2_outputs(1419) <= (layer1_outputs(4605)) or (layer1_outputs(2152));
    layer2_outputs(1420) <= layer1_outputs(446);
    layer2_outputs(1421) <= not(layer1_outputs(3989));
    layer2_outputs(1422) <= not(layer1_outputs(409)) or (layer1_outputs(1100));
    layer2_outputs(1423) <= (layer1_outputs(2271)) xor (layer1_outputs(2481));
    layer2_outputs(1424) <= layer1_outputs(2972);
    layer2_outputs(1425) <= not((layer1_outputs(2152)) or (layer1_outputs(1135)));
    layer2_outputs(1426) <= layer1_outputs(486);
    layer2_outputs(1427) <= not(layer1_outputs(973)) or (layer1_outputs(1331));
    layer2_outputs(1428) <= layer1_outputs(4962);
    layer2_outputs(1429) <= not(layer1_outputs(3497));
    layer2_outputs(1430) <= (layer1_outputs(3101)) xor (layer1_outputs(3255));
    layer2_outputs(1431) <= layer1_outputs(1785);
    layer2_outputs(1432) <= layer1_outputs(4551);
    layer2_outputs(1433) <= layer1_outputs(3891);
    layer2_outputs(1434) <= (layer1_outputs(3165)) and not (layer1_outputs(4915));
    layer2_outputs(1435) <= (layer1_outputs(2402)) and (layer1_outputs(2188));
    layer2_outputs(1436) <= not((layer1_outputs(3548)) xor (layer1_outputs(2665)));
    layer2_outputs(1437) <= layer1_outputs(92);
    layer2_outputs(1438) <= not((layer1_outputs(3713)) and (layer1_outputs(1774)));
    layer2_outputs(1439) <= not((layer1_outputs(59)) or (layer1_outputs(1630)));
    layer2_outputs(1440) <= not(layer1_outputs(1051));
    layer2_outputs(1441) <= not(layer1_outputs(3874));
    layer2_outputs(1442) <= layer1_outputs(2071);
    layer2_outputs(1443) <= layer1_outputs(1418);
    layer2_outputs(1444) <= layer1_outputs(4593);
    layer2_outputs(1445) <= (layer1_outputs(602)) xor (layer1_outputs(4092));
    layer2_outputs(1446) <= (layer1_outputs(1382)) and not (layer1_outputs(4220));
    layer2_outputs(1447) <= not(layer1_outputs(855));
    layer2_outputs(1448) <= layer1_outputs(1153);
    layer2_outputs(1449) <= (layer1_outputs(3485)) and not (layer1_outputs(2948));
    layer2_outputs(1450) <= layer1_outputs(3258);
    layer2_outputs(1451) <= not(layer1_outputs(3682));
    layer2_outputs(1452) <= not(layer1_outputs(4765));
    layer2_outputs(1453) <= not(layer1_outputs(2611)) or (layer1_outputs(3647));
    layer2_outputs(1454) <= '1';
    layer2_outputs(1455) <= not(layer1_outputs(3850));
    layer2_outputs(1456) <= (layer1_outputs(1456)) and (layer1_outputs(4010));
    layer2_outputs(1457) <= not(layer1_outputs(2625));
    layer2_outputs(1458) <= layer1_outputs(4068);
    layer2_outputs(1459) <= not(layer1_outputs(3108)) or (layer1_outputs(102));
    layer2_outputs(1460) <= not(layer1_outputs(2106));
    layer2_outputs(1461) <= layer1_outputs(4465);
    layer2_outputs(1462) <= layer1_outputs(3541);
    layer2_outputs(1463) <= not(layer1_outputs(4294)) or (layer1_outputs(2392));
    layer2_outputs(1464) <= not(layer1_outputs(5065));
    layer2_outputs(1465) <= (layer1_outputs(3127)) or (layer1_outputs(4943));
    layer2_outputs(1466) <= not(layer1_outputs(967));
    layer2_outputs(1467) <= not(layer1_outputs(1247)) or (layer1_outputs(914));
    layer2_outputs(1468) <= layer1_outputs(2426);
    layer2_outputs(1469) <= layer1_outputs(4282);
    layer2_outputs(1470) <= not((layer1_outputs(2009)) and (layer1_outputs(3751)));
    layer2_outputs(1471) <= layer1_outputs(1787);
    layer2_outputs(1472) <= not(layer1_outputs(4019)) or (layer1_outputs(2331));
    layer2_outputs(1473) <= layer1_outputs(2983);
    layer2_outputs(1474) <= not((layer1_outputs(3716)) xor (layer1_outputs(4788)));
    layer2_outputs(1475) <= not(layer1_outputs(3467));
    layer2_outputs(1476) <= not((layer1_outputs(5064)) and (layer1_outputs(4671)));
    layer2_outputs(1477) <= (layer1_outputs(1197)) and not (layer1_outputs(415));
    layer2_outputs(1478) <= layer1_outputs(3795);
    layer2_outputs(1479) <= (layer1_outputs(3655)) or (layer1_outputs(4271));
    layer2_outputs(1480) <= (layer1_outputs(2340)) and (layer1_outputs(841));
    layer2_outputs(1481) <= (layer1_outputs(2849)) and not (layer1_outputs(3694));
    layer2_outputs(1482) <= not(layer1_outputs(4499)) or (layer1_outputs(533));
    layer2_outputs(1483) <= layer1_outputs(4158);
    layer2_outputs(1484) <= not(layer1_outputs(3016));
    layer2_outputs(1485) <= not(layer1_outputs(413)) or (layer1_outputs(3000));
    layer2_outputs(1486) <= (layer1_outputs(4984)) or (layer1_outputs(2870));
    layer2_outputs(1487) <= not(layer1_outputs(2604));
    layer2_outputs(1488) <= layer1_outputs(4923);
    layer2_outputs(1489) <= not(layer1_outputs(2227));
    layer2_outputs(1490) <= (layer1_outputs(3670)) or (layer1_outputs(390));
    layer2_outputs(1491) <= not(layer1_outputs(2626)) or (layer1_outputs(315));
    layer2_outputs(1492) <= layer1_outputs(4942);
    layer2_outputs(1493) <= not(layer1_outputs(3375));
    layer2_outputs(1494) <= not((layer1_outputs(4802)) and (layer1_outputs(2135)));
    layer2_outputs(1495) <= not(layer1_outputs(3347));
    layer2_outputs(1496) <= not(layer1_outputs(1644));
    layer2_outputs(1497) <= not(layer1_outputs(3826));
    layer2_outputs(1498) <= layer1_outputs(3611);
    layer2_outputs(1499) <= not(layer1_outputs(2846));
    layer2_outputs(1500) <= layer1_outputs(820);
    layer2_outputs(1501) <= (layer1_outputs(4347)) or (layer1_outputs(4353));
    layer2_outputs(1502) <= (layer1_outputs(3253)) and not (layer1_outputs(565));
    layer2_outputs(1503) <= not(layer1_outputs(2521));
    layer2_outputs(1504) <= layer1_outputs(2663);
    layer2_outputs(1505) <= not(layer1_outputs(4675));
    layer2_outputs(1506) <= not(layer1_outputs(4007)) or (layer1_outputs(1355));
    layer2_outputs(1507) <= layer1_outputs(2427);
    layer2_outputs(1508) <= not(layer1_outputs(3068));
    layer2_outputs(1509) <= layer1_outputs(5028);
    layer2_outputs(1510) <= not(layer1_outputs(100));
    layer2_outputs(1511) <= layer1_outputs(4102);
    layer2_outputs(1512) <= '1';
    layer2_outputs(1513) <= (layer1_outputs(2029)) and not (layer1_outputs(1755));
    layer2_outputs(1514) <= (layer1_outputs(2804)) and not (layer1_outputs(4110));
    layer2_outputs(1515) <= not(layer1_outputs(3632));
    layer2_outputs(1516) <= not((layer1_outputs(2625)) and (layer1_outputs(887)));
    layer2_outputs(1517) <= layer1_outputs(3218);
    layer2_outputs(1518) <= not(layer1_outputs(3623));
    layer2_outputs(1519) <= (layer1_outputs(3578)) or (layer1_outputs(1418));
    layer2_outputs(1520) <= (layer1_outputs(2397)) xor (layer1_outputs(1101));
    layer2_outputs(1521) <= not(layer1_outputs(4897));
    layer2_outputs(1522) <= not(layer1_outputs(2910)) or (layer1_outputs(1568));
    layer2_outputs(1523) <= not(layer1_outputs(546));
    layer2_outputs(1524) <= not(layer1_outputs(203));
    layer2_outputs(1525) <= not((layer1_outputs(4344)) or (layer1_outputs(4009)));
    layer2_outputs(1526) <= not((layer1_outputs(432)) and (layer1_outputs(2200)));
    layer2_outputs(1527) <= (layer1_outputs(710)) and not (layer1_outputs(3730));
    layer2_outputs(1528) <= (layer1_outputs(2516)) and not (layer1_outputs(3533));
    layer2_outputs(1529) <= not((layer1_outputs(1211)) and (layer1_outputs(2612)));
    layer2_outputs(1530) <= not((layer1_outputs(4313)) and (layer1_outputs(1915)));
    layer2_outputs(1531) <= not(layer1_outputs(4281));
    layer2_outputs(1532) <= (layer1_outputs(4652)) xor (layer1_outputs(5092));
    layer2_outputs(1533) <= not(layer1_outputs(1193));
    layer2_outputs(1534) <= not(layer1_outputs(3749));
    layer2_outputs(1535) <= layer1_outputs(299);
    layer2_outputs(1536) <= not(layer1_outputs(249));
    layer2_outputs(1537) <= layer1_outputs(673);
    layer2_outputs(1538) <= not(layer1_outputs(797));
    layer2_outputs(1539) <= not((layer1_outputs(667)) and (layer1_outputs(1073)));
    layer2_outputs(1540) <= layer1_outputs(4557);
    layer2_outputs(1541) <= (layer1_outputs(1804)) and (layer1_outputs(408));
    layer2_outputs(1542) <= (layer1_outputs(3668)) and not (layer1_outputs(4739));
    layer2_outputs(1543) <= not((layer1_outputs(4112)) and (layer1_outputs(3927)));
    layer2_outputs(1544) <= not(layer1_outputs(4551));
    layer2_outputs(1545) <= (layer1_outputs(1486)) or (layer1_outputs(4368));
    layer2_outputs(1546) <= layer1_outputs(4833);
    layer2_outputs(1547) <= layer1_outputs(4004);
    layer2_outputs(1548) <= (layer1_outputs(649)) and not (layer1_outputs(655));
    layer2_outputs(1549) <= layer1_outputs(2307);
    layer2_outputs(1550) <= layer1_outputs(3943);
    layer2_outputs(1551) <= not(layer1_outputs(3591));
    layer2_outputs(1552) <= layer1_outputs(2337);
    layer2_outputs(1553) <= (layer1_outputs(3888)) or (layer1_outputs(5));
    layer2_outputs(1554) <= layer1_outputs(3015);
    layer2_outputs(1555) <= (layer1_outputs(3735)) and not (layer1_outputs(4481));
    layer2_outputs(1556) <= layer1_outputs(3097);
    layer2_outputs(1557) <= not(layer1_outputs(2160));
    layer2_outputs(1558) <= layer1_outputs(3454);
    layer2_outputs(1559) <= not((layer1_outputs(4806)) and (layer1_outputs(4434)));
    layer2_outputs(1560) <= (layer1_outputs(358)) or (layer1_outputs(669));
    layer2_outputs(1561) <= (layer1_outputs(1935)) or (layer1_outputs(2967));
    layer2_outputs(1562) <= (layer1_outputs(507)) or (layer1_outputs(1852));
    layer2_outputs(1563) <= not((layer1_outputs(904)) and (layer1_outputs(3261)));
    layer2_outputs(1564) <= not(layer1_outputs(1634));
    layer2_outputs(1565) <= layer1_outputs(491);
    layer2_outputs(1566) <= not(layer1_outputs(4284));
    layer2_outputs(1567) <= not(layer1_outputs(1991)) or (layer1_outputs(4773));
    layer2_outputs(1568) <= layer1_outputs(1911);
    layer2_outputs(1569) <= layer1_outputs(4224);
    layer2_outputs(1570) <= (layer1_outputs(3447)) and not (layer1_outputs(2334));
    layer2_outputs(1571) <= '1';
    layer2_outputs(1572) <= not(layer1_outputs(3249)) or (layer1_outputs(36));
    layer2_outputs(1573) <= not((layer1_outputs(2975)) or (layer1_outputs(3544)));
    layer2_outputs(1574) <= layer1_outputs(1323);
    layer2_outputs(1575) <= not(layer1_outputs(1066));
    layer2_outputs(1576) <= not(layer1_outputs(316));
    layer2_outputs(1577) <= layer1_outputs(5098);
    layer2_outputs(1578) <= layer1_outputs(1089);
    layer2_outputs(1579) <= not(layer1_outputs(4364)) or (layer1_outputs(1007));
    layer2_outputs(1580) <= layer1_outputs(4903);
    layer2_outputs(1581) <= layer1_outputs(2537);
    layer2_outputs(1582) <= not(layer1_outputs(1378)) or (layer1_outputs(998));
    layer2_outputs(1583) <= (layer1_outputs(3360)) or (layer1_outputs(3736));
    layer2_outputs(1584) <= not(layer1_outputs(4574));
    layer2_outputs(1585) <= not(layer1_outputs(4081)) or (layer1_outputs(1122));
    layer2_outputs(1586) <= not(layer1_outputs(4731));
    layer2_outputs(1587) <= not(layer1_outputs(2290));
    layer2_outputs(1588) <= not(layer1_outputs(1498));
    layer2_outputs(1589) <= not(layer1_outputs(2919)) or (layer1_outputs(2872));
    layer2_outputs(1590) <= not(layer1_outputs(3004)) or (layer1_outputs(3893));
    layer2_outputs(1591) <= (layer1_outputs(2406)) xor (layer1_outputs(1942));
    layer2_outputs(1592) <= layer1_outputs(4358);
    layer2_outputs(1593) <= (layer1_outputs(4935)) and not (layer1_outputs(4401));
    layer2_outputs(1594) <= not(layer1_outputs(870));
    layer2_outputs(1595) <= not((layer1_outputs(3430)) or (layer1_outputs(1401)));
    layer2_outputs(1596) <= not((layer1_outputs(411)) and (layer1_outputs(5103)));
    layer2_outputs(1597) <= (layer1_outputs(2647)) or (layer1_outputs(2935));
    layer2_outputs(1598) <= layer1_outputs(3936);
    layer2_outputs(1599) <= layer1_outputs(2628);
    layer2_outputs(1600) <= '0';
    layer2_outputs(1601) <= (layer1_outputs(2830)) and not (layer1_outputs(1427));
    layer2_outputs(1602) <= not(layer1_outputs(1147)) or (layer1_outputs(1555));
    layer2_outputs(1603) <= not((layer1_outputs(1232)) or (layer1_outputs(1109)));
    layer2_outputs(1604) <= not(layer1_outputs(2947));
    layer2_outputs(1605) <= not(layer1_outputs(1708));
    layer2_outputs(1606) <= layer1_outputs(780);
    layer2_outputs(1607) <= layer1_outputs(2347);
    layer2_outputs(1608) <= layer1_outputs(1373);
    layer2_outputs(1609) <= not(layer1_outputs(4127)) or (layer1_outputs(4494));
    layer2_outputs(1610) <= not(layer1_outputs(2105));
    layer2_outputs(1611) <= layer1_outputs(584);
    layer2_outputs(1612) <= layer1_outputs(4269);
    layer2_outputs(1613) <= (layer1_outputs(3342)) and (layer1_outputs(2363));
    layer2_outputs(1614) <= not(layer1_outputs(2384)) or (layer1_outputs(2768));
    layer2_outputs(1615) <= not(layer1_outputs(3107)) or (layer1_outputs(297));
    layer2_outputs(1616) <= (layer1_outputs(4065)) and not (layer1_outputs(1680));
    layer2_outputs(1617) <= not((layer1_outputs(1640)) or (layer1_outputs(1232)));
    layer2_outputs(1618) <= (layer1_outputs(1937)) and not (layer1_outputs(4442));
    layer2_outputs(1619) <= (layer1_outputs(895)) and not (layer1_outputs(4314));
    layer2_outputs(1620) <= not(layer1_outputs(619));
    layer2_outputs(1621) <= '0';
    layer2_outputs(1622) <= layer1_outputs(3077);
    layer2_outputs(1623) <= layer1_outputs(1645);
    layer2_outputs(1624) <= not((layer1_outputs(738)) xor (layer1_outputs(1233)));
    layer2_outputs(1625) <= not(layer1_outputs(5059));
    layer2_outputs(1626) <= not(layer1_outputs(2779));
    layer2_outputs(1627) <= not(layer1_outputs(5018));
    layer2_outputs(1628) <= not(layer1_outputs(1067));
    layer2_outputs(1629) <= not(layer1_outputs(3553));
    layer2_outputs(1630) <= layer1_outputs(4586);
    layer2_outputs(1631) <= layer1_outputs(2476);
    layer2_outputs(1632) <= not(layer1_outputs(1153));
    layer2_outputs(1633) <= not(layer1_outputs(824));
    layer2_outputs(1634) <= (layer1_outputs(1561)) or (layer1_outputs(2709));
    layer2_outputs(1635) <= (layer1_outputs(4654)) or (layer1_outputs(1675));
    layer2_outputs(1636) <= layer1_outputs(325);
    layer2_outputs(1637) <= (layer1_outputs(3996)) and (layer1_outputs(2700));
    layer2_outputs(1638) <= (layer1_outputs(64)) or (layer1_outputs(39));
    layer2_outputs(1639) <= '0';
    layer2_outputs(1640) <= not(layer1_outputs(1911));
    layer2_outputs(1641) <= (layer1_outputs(1678)) and (layer1_outputs(2264));
    layer2_outputs(1642) <= not(layer1_outputs(3783));
    layer2_outputs(1643) <= not(layer1_outputs(57)) or (layer1_outputs(1445));
    layer2_outputs(1644) <= (layer1_outputs(2068)) or (layer1_outputs(5017));
    layer2_outputs(1645) <= not((layer1_outputs(55)) and (layer1_outputs(107)));
    layer2_outputs(1646) <= (layer1_outputs(714)) and (layer1_outputs(1760));
    layer2_outputs(1647) <= layer1_outputs(4867);
    layer2_outputs(1648) <= layer1_outputs(547);
    layer2_outputs(1649) <= not(layer1_outputs(2785));
    layer2_outputs(1650) <= not(layer1_outputs(1536));
    layer2_outputs(1651) <= not(layer1_outputs(1109));
    layer2_outputs(1652) <= layer1_outputs(2926);
    layer2_outputs(1653) <= not((layer1_outputs(1977)) or (layer1_outputs(3451)));
    layer2_outputs(1654) <= not(layer1_outputs(3813)) or (layer1_outputs(2819));
    layer2_outputs(1655) <= layer1_outputs(2342);
    layer2_outputs(1656) <= layer1_outputs(4320);
    layer2_outputs(1657) <= not((layer1_outputs(3260)) and (layer1_outputs(5003)));
    layer2_outputs(1658) <= layer1_outputs(3693);
    layer2_outputs(1659) <= (layer1_outputs(4686)) and not (layer1_outputs(3603));
    layer2_outputs(1660) <= layer1_outputs(3410);
    layer2_outputs(1661) <= not(layer1_outputs(2887));
    layer2_outputs(1662) <= layer1_outputs(4737);
    layer2_outputs(1663) <= layer1_outputs(1681);
    layer2_outputs(1664) <= (layer1_outputs(1964)) or (layer1_outputs(1882));
    layer2_outputs(1665) <= layer1_outputs(4254);
    layer2_outputs(1666) <= (layer1_outputs(5016)) xor (layer1_outputs(4755));
    layer2_outputs(1667) <= not(layer1_outputs(970)) or (layer1_outputs(1201));
    layer2_outputs(1668) <= not((layer1_outputs(2510)) or (layer1_outputs(4775)));
    layer2_outputs(1669) <= layer1_outputs(3935);
    layer2_outputs(1670) <= layer1_outputs(2140);
    layer2_outputs(1671) <= not(layer1_outputs(521)) or (layer1_outputs(1803));
    layer2_outputs(1672) <= (layer1_outputs(4478)) and not (layer1_outputs(4628));
    layer2_outputs(1673) <= layer1_outputs(2866);
    layer2_outputs(1674) <= layer1_outputs(2832);
    layer2_outputs(1675) <= layer1_outputs(3379);
    layer2_outputs(1676) <= (layer1_outputs(4404)) and not (layer1_outputs(3053));
    layer2_outputs(1677) <= layer1_outputs(382);
    layer2_outputs(1678) <= (layer1_outputs(4102)) or (layer1_outputs(4907));
    layer2_outputs(1679) <= not(layer1_outputs(1576));
    layer2_outputs(1680) <= (layer1_outputs(3027)) xor (layer1_outputs(4362));
    layer2_outputs(1681) <= not((layer1_outputs(3774)) and (layer1_outputs(2557)));
    layer2_outputs(1682) <= not(layer1_outputs(2298));
    layer2_outputs(1683) <= (layer1_outputs(2932)) and (layer1_outputs(1749));
    layer2_outputs(1684) <= not(layer1_outputs(1379));
    layer2_outputs(1685) <= not(layer1_outputs(1450));
    layer2_outputs(1686) <= (layer1_outputs(3348)) and not (layer1_outputs(204));
    layer2_outputs(1687) <= not(layer1_outputs(1112));
    layer2_outputs(1688) <= not(layer1_outputs(305)) or (layer1_outputs(4511));
    layer2_outputs(1689) <= (layer1_outputs(322)) or (layer1_outputs(1402));
    layer2_outputs(1690) <= layer1_outputs(2698);
    layer2_outputs(1691) <= (layer1_outputs(4223)) and not (layer1_outputs(1733));
    layer2_outputs(1692) <= not(layer1_outputs(831));
    layer2_outputs(1693) <= layer1_outputs(3543);
    layer2_outputs(1694) <= layer1_outputs(1492);
    layer2_outputs(1695) <= not(layer1_outputs(2868)) or (layer1_outputs(2465));
    layer2_outputs(1696) <= not(layer1_outputs(2237));
    layer2_outputs(1697) <= layer1_outputs(4950);
    layer2_outputs(1698) <= layer1_outputs(1643);
    layer2_outputs(1699) <= layer1_outputs(415);
    layer2_outputs(1700) <= layer1_outputs(1648);
    layer2_outputs(1701) <= not(layer1_outputs(5006)) or (layer1_outputs(90));
    layer2_outputs(1702) <= layer1_outputs(1224);
    layer2_outputs(1703) <= (layer1_outputs(4784)) or (layer1_outputs(830));
    layer2_outputs(1704) <= not(layer1_outputs(241));
    layer2_outputs(1705) <= not(layer1_outputs(1065));
    layer2_outputs(1706) <= layer1_outputs(5054);
    layer2_outputs(1707) <= (layer1_outputs(3838)) and (layer1_outputs(2605));
    layer2_outputs(1708) <= layer1_outputs(269);
    layer2_outputs(1709) <= (layer1_outputs(1940)) or (layer1_outputs(2122));
    layer2_outputs(1710) <= not(layer1_outputs(647));
    layer2_outputs(1711) <= not(layer1_outputs(4065));
    layer2_outputs(1712) <= not(layer1_outputs(4782)) or (layer1_outputs(2803));
    layer2_outputs(1713) <= not(layer1_outputs(4408));
    layer2_outputs(1714) <= not((layer1_outputs(2979)) and (layer1_outputs(2437)));
    layer2_outputs(1715) <= (layer1_outputs(2963)) xor (layer1_outputs(2034));
    layer2_outputs(1716) <= not(layer1_outputs(2352));
    layer2_outputs(1717) <= layer1_outputs(2182);
    layer2_outputs(1718) <= not(layer1_outputs(2818));
    layer2_outputs(1719) <= layer1_outputs(2124);
    layer2_outputs(1720) <= not(layer1_outputs(4528)) or (layer1_outputs(3206));
    layer2_outputs(1721) <= (layer1_outputs(4422)) and not (layer1_outputs(4510));
    layer2_outputs(1722) <= not(layer1_outputs(1383)) or (layer1_outputs(4061));
    layer2_outputs(1723) <= layer1_outputs(4284);
    layer2_outputs(1724) <= not(layer1_outputs(959));
    layer2_outputs(1725) <= layer1_outputs(1623);
    layer2_outputs(1726) <= (layer1_outputs(4470)) xor (layer1_outputs(1252));
    layer2_outputs(1727) <= (layer1_outputs(3894)) and not (layer1_outputs(4428));
    layer2_outputs(1728) <= not(layer1_outputs(1260));
    layer2_outputs(1729) <= not(layer1_outputs(2675));
    layer2_outputs(1730) <= (layer1_outputs(2090)) and not (layer1_outputs(1967));
    layer2_outputs(1731) <= not(layer1_outputs(4525)) or (layer1_outputs(483));
    layer2_outputs(1732) <= layer1_outputs(4247);
    layer2_outputs(1733) <= not(layer1_outputs(2672));
    layer2_outputs(1734) <= layer1_outputs(3184);
    layer2_outputs(1735) <= (layer1_outputs(4758)) xor (layer1_outputs(3160));
    layer2_outputs(1736) <= not(layer1_outputs(4179)) or (layer1_outputs(902));
    layer2_outputs(1737) <= not((layer1_outputs(2971)) and (layer1_outputs(2927)));
    layer2_outputs(1738) <= not(layer1_outputs(200));
    layer2_outputs(1739) <= (layer1_outputs(5022)) and not (layer1_outputs(5037));
    layer2_outputs(1740) <= layer1_outputs(256);
    layer2_outputs(1741) <= not((layer1_outputs(239)) or (layer1_outputs(2379)));
    layer2_outputs(1742) <= layer1_outputs(1836);
    layer2_outputs(1743) <= not(layer1_outputs(4637));
    layer2_outputs(1744) <= (layer1_outputs(4321)) and (layer1_outputs(2787));
    layer2_outputs(1745) <= not(layer1_outputs(60));
    layer2_outputs(1746) <= not(layer1_outputs(2857));
    layer2_outputs(1747) <= layer1_outputs(772);
    layer2_outputs(1748) <= layer1_outputs(3979);
    layer2_outputs(1749) <= not(layer1_outputs(3405)) or (layer1_outputs(3203));
    layer2_outputs(1750) <= not(layer1_outputs(2091));
    layer2_outputs(1751) <= (layer1_outputs(1716)) and (layer1_outputs(4717));
    layer2_outputs(1752) <= not(layer1_outputs(1181));
    layer2_outputs(1753) <= layer1_outputs(2572);
    layer2_outputs(1754) <= layer1_outputs(3464);
    layer2_outputs(1755) <= not(layer1_outputs(2336)) or (layer1_outputs(198));
    layer2_outputs(1756) <= not(layer1_outputs(3769)) or (layer1_outputs(441));
    layer2_outputs(1757) <= '0';
    layer2_outputs(1758) <= not(layer1_outputs(3190));
    layer2_outputs(1759) <= not((layer1_outputs(698)) or (layer1_outputs(2513)));
    layer2_outputs(1760) <= not(layer1_outputs(1978));
    layer2_outputs(1761) <= not((layer1_outputs(4310)) or (layer1_outputs(135)));
    layer2_outputs(1762) <= (layer1_outputs(2449)) and not (layer1_outputs(1011));
    layer2_outputs(1763) <= not(layer1_outputs(4832)) or (layer1_outputs(1448));
    layer2_outputs(1764) <= not(layer1_outputs(3501));
    layer2_outputs(1765) <= layer1_outputs(282);
    layer2_outputs(1766) <= '1';
    layer2_outputs(1767) <= not((layer1_outputs(388)) or (layer1_outputs(680)));
    layer2_outputs(1768) <= (layer1_outputs(2451)) and not (layer1_outputs(3472));
    layer2_outputs(1769) <= layer1_outputs(3314);
    layer2_outputs(1770) <= (layer1_outputs(4362)) and not (layer1_outputs(1811));
    layer2_outputs(1771) <= not(layer1_outputs(3467));
    layer2_outputs(1772) <= (layer1_outputs(3495)) or (layer1_outputs(1706));
    layer2_outputs(1773) <= not((layer1_outputs(1626)) and (layer1_outputs(1291)));
    layer2_outputs(1774) <= not(layer1_outputs(2401)) or (layer1_outputs(931));
    layer2_outputs(1775) <= layer1_outputs(4138);
    layer2_outputs(1776) <= layer1_outputs(1516);
    layer2_outputs(1777) <= layer1_outputs(2541);
    layer2_outputs(1778) <= layer1_outputs(2423);
    layer2_outputs(1779) <= not(layer1_outputs(4258));
    layer2_outputs(1780) <= not(layer1_outputs(3431));
    layer2_outputs(1781) <= not(layer1_outputs(1184)) or (layer1_outputs(4237));
    layer2_outputs(1782) <= (layer1_outputs(1273)) xor (layer1_outputs(3972));
    layer2_outputs(1783) <= not(layer1_outputs(1619));
    layer2_outputs(1784) <= not(layer1_outputs(3929));
    layer2_outputs(1785) <= not((layer1_outputs(496)) and (layer1_outputs(1817)));
    layer2_outputs(1786) <= (layer1_outputs(614)) xor (layer1_outputs(1729));
    layer2_outputs(1787) <= not(layer1_outputs(529)) or (layer1_outputs(2957));
    layer2_outputs(1788) <= (layer1_outputs(2898)) xor (layer1_outputs(2496));
    layer2_outputs(1789) <= (layer1_outputs(3622)) and not (layer1_outputs(696));
    layer2_outputs(1790) <= not(layer1_outputs(3090));
    layer2_outputs(1791) <= layer1_outputs(4385);
    layer2_outputs(1792) <= (layer1_outputs(4932)) or (layer1_outputs(1315));
    layer2_outputs(1793) <= not((layer1_outputs(3524)) or (layer1_outputs(1393)));
    layer2_outputs(1794) <= not(layer1_outputs(3879));
    layer2_outputs(1795) <= not((layer1_outputs(1432)) xor (layer1_outputs(1313)));
    layer2_outputs(1796) <= not((layer1_outputs(1333)) or (layer1_outputs(879)));
    layer2_outputs(1797) <= not(layer1_outputs(364));
    layer2_outputs(1798) <= (layer1_outputs(215)) and not (layer1_outputs(2339));
    layer2_outputs(1799) <= not(layer1_outputs(3237));
    layer2_outputs(1800) <= layer1_outputs(2377);
    layer2_outputs(1801) <= layer1_outputs(4734);
    layer2_outputs(1802) <= not(layer1_outputs(3334)) or (layer1_outputs(2741));
    layer2_outputs(1803) <= not(layer1_outputs(185));
    layer2_outputs(1804) <= layer1_outputs(4512);
    layer2_outputs(1805) <= not(layer1_outputs(3719));
    layer2_outputs(1806) <= not((layer1_outputs(350)) or (layer1_outputs(4866)));
    layer2_outputs(1807) <= not(layer1_outputs(5067));
    layer2_outputs(1808) <= layer1_outputs(3435);
    layer2_outputs(1809) <= layer1_outputs(2017);
    layer2_outputs(1810) <= not(layer1_outputs(1956));
    layer2_outputs(1811) <= not(layer1_outputs(2681)) or (layer1_outputs(4803));
    layer2_outputs(1812) <= (layer1_outputs(12)) xor (layer1_outputs(1638));
    layer2_outputs(1813) <= not((layer1_outputs(5046)) or (layer1_outputs(4907)));
    layer2_outputs(1814) <= not(layer1_outputs(110));
    layer2_outputs(1815) <= (layer1_outputs(5075)) xor (layer1_outputs(4421));
    layer2_outputs(1816) <= (layer1_outputs(5111)) xor (layer1_outputs(1702));
    layer2_outputs(1817) <= not(layer1_outputs(941));
    layer2_outputs(1818) <= not((layer1_outputs(4643)) and (layer1_outputs(83)));
    layer2_outputs(1819) <= layer1_outputs(1202);
    layer2_outputs(1820) <= not(layer1_outputs(4908));
    layer2_outputs(1821) <= not(layer1_outputs(1831)) or (layer1_outputs(4215));
    layer2_outputs(1822) <= (layer1_outputs(769)) and (layer1_outputs(3535));
    layer2_outputs(1823) <= '1';
    layer2_outputs(1824) <= (layer1_outputs(4047)) and not (layer1_outputs(4867));
    layer2_outputs(1825) <= not(layer1_outputs(4131));
    layer2_outputs(1826) <= not(layer1_outputs(1274));
    layer2_outputs(1827) <= layer1_outputs(2064);
    layer2_outputs(1828) <= not((layer1_outputs(2258)) and (layer1_outputs(3343)));
    layer2_outputs(1829) <= not(layer1_outputs(2369));
    layer2_outputs(1830) <= not(layer1_outputs(4956));
    layer2_outputs(1831) <= (layer1_outputs(987)) and not (layer1_outputs(5014));
    layer2_outputs(1832) <= not(layer1_outputs(4871));
    layer2_outputs(1833) <= (layer1_outputs(425)) and (layer1_outputs(2362));
    layer2_outputs(1834) <= not(layer1_outputs(4246)) or (layer1_outputs(1676));
    layer2_outputs(1835) <= (layer1_outputs(1226)) and (layer1_outputs(2763));
    layer2_outputs(1836) <= layer1_outputs(2833);
    layer2_outputs(1837) <= (layer1_outputs(3153)) and not (layer1_outputs(2077));
    layer2_outputs(1838) <= not((layer1_outputs(4745)) or (layer1_outputs(3617)));
    layer2_outputs(1839) <= layer1_outputs(4248);
    layer2_outputs(1840) <= not(layer1_outputs(2216));
    layer2_outputs(1841) <= layer1_outputs(1017);
    layer2_outputs(1842) <= (layer1_outputs(2938)) or (layer1_outputs(301));
    layer2_outputs(1843) <= layer1_outputs(3680);
    layer2_outputs(1844) <= not((layer1_outputs(3759)) or (layer1_outputs(4651)));
    layer2_outputs(1845) <= not((layer1_outputs(4060)) and (layer1_outputs(2831)));
    layer2_outputs(1846) <= not(layer1_outputs(1157));
    layer2_outputs(1847) <= not(layer1_outputs(2690));
    layer2_outputs(1848) <= not(layer1_outputs(2790)) or (layer1_outputs(1141));
    layer2_outputs(1849) <= not(layer1_outputs(929)) or (layer1_outputs(3794));
    layer2_outputs(1850) <= not((layer1_outputs(1016)) or (layer1_outputs(1604)));
    layer2_outputs(1851) <= (layer1_outputs(804)) or (layer1_outputs(3025));
    layer2_outputs(1852) <= not((layer1_outputs(2189)) or (layer1_outputs(908)));
    layer2_outputs(1853) <= not(layer1_outputs(3954));
    layer2_outputs(1854) <= (layer1_outputs(2020)) xor (layer1_outputs(2119));
    layer2_outputs(1855) <= not(layer1_outputs(2178));
    layer2_outputs(1856) <= '1';
    layer2_outputs(1857) <= (layer1_outputs(1994)) and (layer1_outputs(2501));
    layer2_outputs(1858) <= not((layer1_outputs(975)) or (layer1_outputs(1656)));
    layer2_outputs(1859) <= not((layer1_outputs(2747)) or (layer1_outputs(144)));
    layer2_outputs(1860) <= layer1_outputs(486);
    layer2_outputs(1861) <= (layer1_outputs(2944)) or (layer1_outputs(2591));
    layer2_outputs(1862) <= not(layer1_outputs(3968)) or (layer1_outputs(3696));
    layer2_outputs(1863) <= not((layer1_outputs(4414)) xor (layer1_outputs(2417)));
    layer2_outputs(1864) <= layer1_outputs(2330);
    layer2_outputs(1865) <= layer1_outputs(3919);
    layer2_outputs(1866) <= '1';
    layer2_outputs(1867) <= (layer1_outputs(2116)) or (layer1_outputs(3985));
    layer2_outputs(1868) <= not(layer1_outputs(1578)) or (layer1_outputs(3765));
    layer2_outputs(1869) <= '1';
    layer2_outputs(1870) <= (layer1_outputs(1354)) and (layer1_outputs(2637));
    layer2_outputs(1871) <= (layer1_outputs(2099)) or (layer1_outputs(4943));
    layer2_outputs(1872) <= layer1_outputs(1210);
    layer2_outputs(1873) <= not(layer1_outputs(4125));
    layer2_outputs(1874) <= layer1_outputs(1539);
    layer2_outputs(1875) <= not(layer1_outputs(2597));
    layer2_outputs(1876) <= not(layer1_outputs(2388));
    layer2_outputs(1877) <= not(layer1_outputs(4959));
    layer2_outputs(1878) <= (layer1_outputs(417)) and not (layer1_outputs(4444));
    layer2_outputs(1879) <= not((layer1_outputs(1813)) and (layer1_outputs(2095)));
    layer2_outputs(1880) <= layer1_outputs(3896);
    layer2_outputs(1881) <= not(layer1_outputs(4567));
    layer2_outputs(1882) <= not((layer1_outputs(3187)) or (layer1_outputs(189)));
    layer2_outputs(1883) <= layer1_outputs(4725);
    layer2_outputs(1884) <= not((layer1_outputs(1669)) or (layer1_outputs(3839)));
    layer2_outputs(1885) <= not(layer1_outputs(226)) or (layer1_outputs(5102));
    layer2_outputs(1886) <= not(layer1_outputs(151)) or (layer1_outputs(2936));
    layer2_outputs(1887) <= (layer1_outputs(433)) and not (layer1_outputs(1966));
    layer2_outputs(1888) <= (layer1_outputs(143)) xor (layer1_outputs(5101));
    layer2_outputs(1889) <= layer1_outputs(2232);
    layer2_outputs(1890) <= not((layer1_outputs(4113)) or (layer1_outputs(1712)));
    layer2_outputs(1891) <= not(layer1_outputs(187));
    layer2_outputs(1892) <= not(layer1_outputs(1345));
    layer2_outputs(1893) <= not((layer1_outputs(3515)) and (layer1_outputs(3232)));
    layer2_outputs(1894) <= (layer1_outputs(1392)) xor (layer1_outputs(2303));
    layer2_outputs(1895) <= not(layer1_outputs(1395));
    layer2_outputs(1896) <= (layer1_outputs(2901)) or (layer1_outputs(580));
    layer2_outputs(1897) <= not((layer1_outputs(1978)) and (layer1_outputs(4420)));
    layer2_outputs(1898) <= not(layer1_outputs(225)) or (layer1_outputs(4944));
    layer2_outputs(1899) <= not(layer1_outputs(3272));
    layer2_outputs(1900) <= '1';
    layer2_outputs(1901) <= not(layer1_outputs(2655)) or (layer1_outputs(4911));
    layer2_outputs(1902) <= not(layer1_outputs(2118)) or (layer1_outputs(4926));
    layer2_outputs(1903) <= (layer1_outputs(2578)) and (layer1_outputs(2180));
    layer2_outputs(1904) <= (layer1_outputs(2311)) and not (layer1_outputs(3646));
    layer2_outputs(1905) <= (layer1_outputs(4143)) and (layer1_outputs(3832));
    layer2_outputs(1906) <= not(layer1_outputs(440));
    layer2_outputs(1907) <= not(layer1_outputs(3901)) or (layer1_outputs(1328));
    layer2_outputs(1908) <= not(layer1_outputs(2379)) or (layer1_outputs(4912));
    layer2_outputs(1909) <= layer1_outputs(4515);
    layer2_outputs(1910) <= not(layer1_outputs(1140));
    layer2_outputs(1911) <= layer1_outputs(1939);
    layer2_outputs(1912) <= not(layer1_outputs(3812));
    layer2_outputs(1913) <= not(layer1_outputs(1510));
    layer2_outputs(1914) <= layer1_outputs(2864);
    layer2_outputs(1915) <= not(layer1_outputs(2702)) or (layer1_outputs(665));
    layer2_outputs(1916) <= layer1_outputs(3496);
    layer2_outputs(1917) <= not((layer1_outputs(591)) or (layer1_outputs(4665)));
    layer2_outputs(1918) <= not(layer1_outputs(805));
    layer2_outputs(1919) <= (layer1_outputs(1612)) and (layer1_outputs(3362));
    layer2_outputs(1920) <= layer1_outputs(1352);
    layer2_outputs(1921) <= not((layer1_outputs(5010)) or (layer1_outputs(4009)));
    layer2_outputs(1922) <= layer1_outputs(4649);
    layer2_outputs(1923) <= not((layer1_outputs(3949)) and (layer1_outputs(4917)));
    layer2_outputs(1924) <= layer1_outputs(1294);
    layer2_outputs(1925) <= not(layer1_outputs(2835));
    layer2_outputs(1926) <= not(layer1_outputs(2816));
    layer2_outputs(1927) <= not(layer1_outputs(2488));
    layer2_outputs(1928) <= (layer1_outputs(4430)) and (layer1_outputs(3851));
    layer2_outputs(1929) <= not(layer1_outputs(663));
    layer2_outputs(1930) <= not(layer1_outputs(4165));
    layer2_outputs(1931) <= layer1_outputs(985);
    layer2_outputs(1932) <= (layer1_outputs(4300)) and not (layer1_outputs(1282));
    layer2_outputs(1933) <= layer1_outputs(4164);
    layer2_outputs(1934) <= (layer1_outputs(453)) and not (layer1_outputs(4366));
    layer2_outputs(1935) <= layer1_outputs(2078);
    layer2_outputs(1936) <= layer1_outputs(2829);
    layer2_outputs(1937) <= not(layer1_outputs(4769));
    layer2_outputs(1938) <= layer1_outputs(2374);
    layer2_outputs(1939) <= not(layer1_outputs(2074));
    layer2_outputs(1940) <= not(layer1_outputs(4204));
    layer2_outputs(1941) <= not((layer1_outputs(761)) xor (layer1_outputs(495)));
    layer2_outputs(1942) <= not(layer1_outputs(2854));
    layer2_outputs(1943) <= not(layer1_outputs(1155)) or (layer1_outputs(1787));
    layer2_outputs(1944) <= layer1_outputs(400);
    layer2_outputs(1945) <= layer1_outputs(3778);
    layer2_outputs(1946) <= (layer1_outputs(2977)) and (layer1_outputs(1877));
    layer2_outputs(1947) <= layer1_outputs(155);
    layer2_outputs(1948) <= not(layer1_outputs(1995));
    layer2_outputs(1949) <= not(layer1_outputs(3885));
    layer2_outputs(1950) <= not((layer1_outputs(4679)) or (layer1_outputs(726)));
    layer2_outputs(1951) <= not(layer1_outputs(903)) or (layer1_outputs(1091));
    layer2_outputs(1952) <= (layer1_outputs(2642)) and not (layer1_outputs(3086));
    layer2_outputs(1953) <= not((layer1_outputs(2899)) and (layer1_outputs(3772)));
    layer2_outputs(1954) <= layer1_outputs(1570);
    layer2_outputs(1955) <= layer1_outputs(4760);
    layer2_outputs(1956) <= not((layer1_outputs(4228)) and (layer1_outputs(2862)));
    layer2_outputs(1957) <= (layer1_outputs(2779)) or (layer1_outputs(368));
    layer2_outputs(1958) <= layer1_outputs(2000);
    layer2_outputs(1959) <= not(layer1_outputs(3744)) or (layer1_outputs(2297));
    layer2_outputs(1960) <= not(layer1_outputs(2365));
    layer2_outputs(1961) <= not((layer1_outputs(3925)) xor (layer1_outputs(42)));
    layer2_outputs(1962) <= (layer1_outputs(653)) or (layer1_outputs(721));
    layer2_outputs(1963) <= not(layer1_outputs(430)) or (layer1_outputs(3471));
    layer2_outputs(1964) <= not(layer1_outputs(351));
    layer2_outputs(1965) <= not(layer1_outputs(745));
    layer2_outputs(1966) <= (layer1_outputs(3576)) or (layer1_outputs(2734));
    layer2_outputs(1967) <= not((layer1_outputs(3389)) and (layer1_outputs(4940)));
    layer2_outputs(1968) <= layer1_outputs(4868);
    layer2_outputs(1969) <= not(layer1_outputs(364));
    layer2_outputs(1970) <= not((layer1_outputs(3151)) xor (layer1_outputs(2531)));
    layer2_outputs(1971) <= layer1_outputs(2557);
    layer2_outputs(1972) <= not(layer1_outputs(1892));
    layer2_outputs(1973) <= '1';
    layer2_outputs(1974) <= not((layer1_outputs(2311)) xor (layer1_outputs(3020)));
    layer2_outputs(1975) <= not(layer1_outputs(948)) or (layer1_outputs(3639));
    layer2_outputs(1976) <= not(layer1_outputs(748));
    layer2_outputs(1977) <= not(layer1_outputs(3774));
    layer2_outputs(1978) <= layer1_outputs(4043);
    layer2_outputs(1979) <= not((layer1_outputs(4814)) or (layer1_outputs(1537)));
    layer2_outputs(1980) <= not(layer1_outputs(2082));
    layer2_outputs(1981) <= (layer1_outputs(3950)) and not (layer1_outputs(3801));
    layer2_outputs(1982) <= layer1_outputs(4042);
    layer2_outputs(1983) <= layer1_outputs(3939);
    layer2_outputs(1984) <= layer1_outputs(3154);
    layer2_outputs(1985) <= (layer1_outputs(2727)) and not (layer1_outputs(4145));
    layer2_outputs(1986) <= '1';
    layer2_outputs(1987) <= (layer1_outputs(61)) and (layer1_outputs(1431));
    layer2_outputs(1988) <= not(layer1_outputs(4005)) or (layer1_outputs(4821));
    layer2_outputs(1989) <= not(layer1_outputs(2999));
    layer2_outputs(1990) <= not((layer1_outputs(511)) or (layer1_outputs(3577)));
    layer2_outputs(1991) <= not(layer1_outputs(3716)) or (layer1_outputs(1540));
    layer2_outputs(1992) <= layer1_outputs(1026);
    layer2_outputs(1993) <= layer1_outputs(2683);
    layer2_outputs(1994) <= not(layer1_outputs(2981)) or (layer1_outputs(1563));
    layer2_outputs(1995) <= (layer1_outputs(1810)) and not (layer1_outputs(3761));
    layer2_outputs(1996) <= not(layer1_outputs(4635));
    layer2_outputs(1997) <= (layer1_outputs(152)) xor (layer1_outputs(566));
    layer2_outputs(1998) <= (layer1_outputs(5035)) and not (layer1_outputs(1230));
    layer2_outputs(1999) <= (layer1_outputs(2346)) and not (layer1_outputs(834));
    layer2_outputs(2000) <= not((layer1_outputs(2873)) or (layer1_outputs(4715)));
    layer2_outputs(2001) <= not((layer1_outputs(3956)) or (layer1_outputs(2217)));
    layer2_outputs(2002) <= not(layer1_outputs(4454));
    layer2_outputs(2003) <= not(layer1_outputs(493));
    layer2_outputs(2004) <= not(layer1_outputs(900));
    layer2_outputs(2005) <= not(layer1_outputs(4961)) or (layer1_outputs(128));
    layer2_outputs(2006) <= layer1_outputs(3216);
    layer2_outputs(2007) <= (layer1_outputs(3715)) and not (layer1_outputs(4499));
    layer2_outputs(2008) <= (layer1_outputs(2494)) and (layer1_outputs(2135));
    layer2_outputs(2009) <= (layer1_outputs(5035)) and not (layer1_outputs(1122));
    layer2_outputs(2010) <= not((layer1_outputs(2772)) xor (layer1_outputs(863)));
    layer2_outputs(2011) <= (layer1_outputs(4199)) or (layer1_outputs(4199));
    layer2_outputs(2012) <= (layer1_outputs(137)) or (layer1_outputs(617));
    layer2_outputs(2013) <= (layer1_outputs(335)) and not (layer1_outputs(2396));
    layer2_outputs(2014) <= layer1_outputs(218);
    layer2_outputs(2015) <= layer1_outputs(586);
    layer2_outputs(2016) <= (layer1_outputs(3506)) and (layer1_outputs(883));
    layer2_outputs(2017) <= (layer1_outputs(2321)) and not (layer1_outputs(97));
    layer2_outputs(2018) <= not(layer1_outputs(2554));
    layer2_outputs(2019) <= (layer1_outputs(1446)) and not (layer1_outputs(2032));
    layer2_outputs(2020) <= not(layer1_outputs(1713)) or (layer1_outputs(567));
    layer2_outputs(2021) <= not(layer1_outputs(4592)) or (layer1_outputs(2976));
    layer2_outputs(2022) <= not(layer1_outputs(1923));
    layer2_outputs(2023) <= (layer1_outputs(2227)) and (layer1_outputs(2652));
    layer2_outputs(2024) <= (layer1_outputs(5011)) xor (layer1_outputs(3712));
    layer2_outputs(2025) <= (layer1_outputs(1358)) and (layer1_outputs(1830));
    layer2_outputs(2026) <= (layer1_outputs(2305)) and not (layer1_outputs(1194));
    layer2_outputs(2027) <= not(layer1_outputs(2651)) or (layer1_outputs(1318));
    layer2_outputs(2028) <= layer1_outputs(2047);
    layer2_outputs(2029) <= layer1_outputs(529);
    layer2_outputs(2030) <= layer1_outputs(1169);
    layer2_outputs(2031) <= layer1_outputs(69);
    layer2_outputs(2032) <= layer1_outputs(37);
    layer2_outputs(2033) <= not(layer1_outputs(3525));
    layer2_outputs(2034) <= not(layer1_outputs(1987));
    layer2_outputs(2035) <= not((layer1_outputs(548)) or (layer1_outputs(3807)));
    layer2_outputs(2036) <= not((layer1_outputs(1123)) or (layer1_outputs(4085)));
    layer2_outputs(2037) <= (layer1_outputs(1366)) or (layer1_outputs(1020));
    layer2_outputs(2038) <= not((layer1_outputs(309)) xor (layer1_outputs(254)));
    layer2_outputs(2039) <= not((layer1_outputs(4759)) and (layer1_outputs(939)));
    layer2_outputs(2040) <= not(layer1_outputs(1258)) or (layer1_outputs(3254));
    layer2_outputs(2041) <= not(layer1_outputs(800)) or (layer1_outputs(3162));
    layer2_outputs(2042) <= not(layer1_outputs(2424)) or (layer1_outputs(3014));
    layer2_outputs(2043) <= layer1_outputs(4158);
    layer2_outputs(2044) <= layer1_outputs(659);
    layer2_outputs(2045) <= layer1_outputs(3189);
    layer2_outputs(2046) <= not(layer1_outputs(2788));
    layer2_outputs(2047) <= layer1_outputs(74);
    layer2_outputs(2048) <= not(layer1_outputs(2239));
    layer2_outputs(2049) <= layer1_outputs(1389);
    layer2_outputs(2050) <= not(layer1_outputs(1409)) or (layer1_outputs(2932));
    layer2_outputs(2051) <= not(layer1_outputs(2075));
    layer2_outputs(2052) <= not(layer1_outputs(80));
    layer2_outputs(2053) <= (layer1_outputs(582)) and not (layer1_outputs(3755));
    layer2_outputs(2054) <= layer1_outputs(1180);
    layer2_outputs(2055) <= layer1_outputs(3546);
    layer2_outputs(2056) <= not((layer1_outputs(3122)) or (layer1_outputs(706)));
    layer2_outputs(2057) <= (layer1_outputs(1162)) xor (layer1_outputs(130));
    layer2_outputs(2058) <= not((layer1_outputs(645)) and (layer1_outputs(4664)));
    layer2_outputs(2059) <= layer1_outputs(4956);
    layer2_outputs(2060) <= not(layer1_outputs(3427));
    layer2_outputs(2061) <= not(layer1_outputs(3365));
    layer2_outputs(2062) <= layer1_outputs(1149);
    layer2_outputs(2063) <= not(layer1_outputs(881));
    layer2_outputs(2064) <= layer1_outputs(3940);
    layer2_outputs(2065) <= layer1_outputs(3447);
    layer2_outputs(2066) <= not(layer1_outputs(4738));
    layer2_outputs(2067) <= layer1_outputs(3602);
    layer2_outputs(2068) <= not(layer1_outputs(4191));
    layer2_outputs(2069) <= not(layer1_outputs(1497));
    layer2_outputs(2070) <= (layer1_outputs(1857)) xor (layer1_outputs(1745));
    layer2_outputs(2071) <= not(layer1_outputs(2266));
    layer2_outputs(2072) <= not(layer1_outputs(1355)) or (layer1_outputs(3468));
    layer2_outputs(2073) <= (layer1_outputs(3625)) and (layer1_outputs(1952));
    layer2_outputs(2074) <= not(layer1_outputs(4614));
    layer2_outputs(2075) <= not(layer1_outputs(3708)) or (layer1_outputs(4962));
    layer2_outputs(2076) <= not(layer1_outputs(1698));
    layer2_outputs(2077) <= not(layer1_outputs(4448));
    layer2_outputs(2078) <= layer1_outputs(832);
    layer2_outputs(2079) <= (layer1_outputs(726)) or (layer1_outputs(2856));
    layer2_outputs(2080) <= not((layer1_outputs(3878)) or (layer1_outputs(4872)));
    layer2_outputs(2081) <= not(layer1_outputs(4058)) or (layer1_outputs(1312));
    layer2_outputs(2082) <= layer1_outputs(3196);
    layer2_outputs(2083) <= layer1_outputs(3390);
    layer2_outputs(2084) <= not(layer1_outputs(3426));
    layer2_outputs(2085) <= layer1_outputs(1995);
    layer2_outputs(2086) <= not(layer1_outputs(3040)) or (layer1_outputs(1801));
    layer2_outputs(2087) <= layer1_outputs(4492);
    layer2_outputs(2088) <= layer1_outputs(3727);
    layer2_outputs(2089) <= not(layer1_outputs(3008));
    layer2_outputs(2090) <= (layer1_outputs(697)) and not (layer1_outputs(3652));
    layer2_outputs(2091) <= not(layer1_outputs(3529));
    layer2_outputs(2092) <= layer1_outputs(4934);
    layer2_outputs(2093) <= not(layer1_outputs(3367));
    layer2_outputs(2094) <= layer1_outputs(1115);
    layer2_outputs(2095) <= layer1_outputs(4531);
    layer2_outputs(2096) <= not(layer1_outputs(3107));
    layer2_outputs(2097) <= not(layer1_outputs(662));
    layer2_outputs(2098) <= not(layer1_outputs(4095));
    layer2_outputs(2099) <= not(layer1_outputs(739)) or (layer1_outputs(522));
    layer2_outputs(2100) <= layer1_outputs(4357);
    layer2_outputs(2101) <= not(layer1_outputs(1821));
    layer2_outputs(2102) <= (layer1_outputs(1835)) and (layer1_outputs(572));
    layer2_outputs(2103) <= not((layer1_outputs(3828)) and (layer1_outputs(862)));
    layer2_outputs(2104) <= (layer1_outputs(4243)) or (layer1_outputs(3635));
    layer2_outputs(2105) <= not(layer1_outputs(598));
    layer2_outputs(2106) <= (layer1_outputs(1509)) and not (layer1_outputs(3963));
    layer2_outputs(2107) <= not(layer1_outputs(1934));
    layer2_outputs(2108) <= (layer1_outputs(1425)) xor (layer1_outputs(2989));
    layer2_outputs(2109) <= not(layer1_outputs(349));
    layer2_outputs(2110) <= not(layer1_outputs(3156));
    layer2_outputs(2111) <= not(layer1_outputs(1406));
    layer2_outputs(2112) <= (layer1_outputs(4807)) and not (layer1_outputs(3036));
    layer2_outputs(2113) <= not(layer1_outputs(3233));
    layer2_outputs(2114) <= (layer1_outputs(326)) or (layer1_outputs(1829));
    layer2_outputs(2115) <= not(layer1_outputs(1575));
    layer2_outputs(2116) <= not(layer1_outputs(1790));
    layer2_outputs(2117) <= (layer1_outputs(3295)) and (layer1_outputs(1025));
    layer2_outputs(2118) <= layer1_outputs(477);
    layer2_outputs(2119) <= not((layer1_outputs(3310)) xor (layer1_outputs(4928)));
    layer2_outputs(2120) <= layer1_outputs(5116);
    layer2_outputs(2121) <= layer1_outputs(4968);
    layer2_outputs(2122) <= not(layer1_outputs(1849));
    layer2_outputs(2123) <= not(layer1_outputs(3323));
    layer2_outputs(2124) <= (layer1_outputs(514)) and not (layer1_outputs(3959));
    layer2_outputs(2125) <= not(layer1_outputs(2590));
    layer2_outputs(2126) <= (layer1_outputs(4092)) xor (layer1_outputs(4830));
    layer2_outputs(2127) <= not(layer1_outputs(2970)) or (layer1_outputs(3006));
    layer2_outputs(2128) <= layer1_outputs(1372);
    layer2_outputs(2129) <= not((layer1_outputs(3182)) or (layer1_outputs(645)));
    layer2_outputs(2130) <= layer1_outputs(3935);
    layer2_outputs(2131) <= (layer1_outputs(2258)) and (layer1_outputs(234));
    layer2_outputs(2132) <= not((layer1_outputs(173)) and (layer1_outputs(2062)));
    layer2_outputs(2133) <= not(layer1_outputs(2641));
    layer2_outputs(2134) <= not(layer1_outputs(3528)) or (layer1_outputs(97));
    layer2_outputs(2135) <= (layer1_outputs(2328)) or (layer1_outputs(3105));
    layer2_outputs(2136) <= (layer1_outputs(827)) and not (layer1_outputs(1203));
    layer2_outputs(2137) <= not(layer1_outputs(4569));
    layer2_outputs(2138) <= not(layer1_outputs(4765));
    layer2_outputs(2139) <= layer1_outputs(1560);
    layer2_outputs(2140) <= (layer1_outputs(1351)) and (layer1_outputs(3193));
    layer2_outputs(2141) <= not(layer1_outputs(4291)) or (layer1_outputs(4638));
    layer2_outputs(2142) <= not(layer1_outputs(2442));
    layer2_outputs(2143) <= layer1_outputs(1272);
    layer2_outputs(2144) <= not(layer1_outputs(3921)) or (layer1_outputs(913));
    layer2_outputs(2145) <= layer1_outputs(2211);
    layer2_outputs(2146) <= layer1_outputs(4727);
    layer2_outputs(2147) <= not((layer1_outputs(1610)) or (layer1_outputs(4965)));
    layer2_outputs(2148) <= not(layer1_outputs(808)) or (layer1_outputs(732));
    layer2_outputs(2149) <= not(layer1_outputs(3272));
    layer2_outputs(2150) <= layer1_outputs(2147);
    layer2_outputs(2151) <= layer1_outputs(3789);
    layer2_outputs(2152) <= not(layer1_outputs(2164)) or (layer1_outputs(3603));
    layer2_outputs(2153) <= not(layer1_outputs(4283));
    layer2_outputs(2154) <= (layer1_outputs(2632)) and not (layer1_outputs(3760));
    layer2_outputs(2155) <= layer1_outputs(2438);
    layer2_outputs(2156) <= layer1_outputs(1824);
    layer2_outputs(2157) <= not(layer1_outputs(2256)) or (layer1_outputs(1390));
    layer2_outputs(2158) <= '0';
    layer2_outputs(2159) <= not(layer1_outputs(4780)) or (layer1_outputs(4854));
    layer2_outputs(2160) <= not((layer1_outputs(744)) or (layer1_outputs(1765)));
    layer2_outputs(2161) <= not(layer1_outputs(4827));
    layer2_outputs(2162) <= layer1_outputs(385);
    layer2_outputs(2163) <= (layer1_outputs(3583)) xor (layer1_outputs(3228));
    layer2_outputs(2164) <= (layer1_outputs(4627)) and not (layer1_outputs(3445));
    layer2_outputs(2165) <= not(layer1_outputs(289));
    layer2_outputs(2166) <= not(layer1_outputs(3673));
    layer2_outputs(2167) <= not(layer1_outputs(4250));
    layer2_outputs(2168) <= not((layer1_outputs(392)) and (layer1_outputs(4419)));
    layer2_outputs(2169) <= not((layer1_outputs(1485)) or (layer1_outputs(2673)));
    layer2_outputs(2170) <= (layer1_outputs(2479)) and not (layer1_outputs(3444));
    layer2_outputs(2171) <= layer1_outputs(1750);
    layer2_outputs(2172) <= (layer1_outputs(5048)) and (layer1_outputs(1161));
    layer2_outputs(2173) <= (layer1_outputs(4602)) and (layer1_outputs(4879));
    layer2_outputs(2174) <= not(layer1_outputs(2398));
    layer2_outputs(2175) <= not((layer1_outputs(4377)) or (layer1_outputs(3758)));
    layer2_outputs(2176) <= not(layer1_outputs(2419));
    layer2_outputs(2177) <= layer1_outputs(4805);
    layer2_outputs(2178) <= (layer1_outputs(3593)) and (layer1_outputs(2824));
    layer2_outputs(2179) <= (layer1_outputs(3010)) and not (layer1_outputs(1603));
    layer2_outputs(2180) <= (layer1_outputs(3882)) and not (layer1_outputs(1060));
    layer2_outputs(2181) <= not(layer1_outputs(395));
    layer2_outputs(2182) <= not(layer1_outputs(3299));
    layer2_outputs(2183) <= not(layer1_outputs(4287));
    layer2_outputs(2184) <= not(layer1_outputs(4101));
    layer2_outputs(2185) <= not((layer1_outputs(3517)) or (layer1_outputs(2312)));
    layer2_outputs(2186) <= (layer1_outputs(2340)) and (layer1_outputs(2016));
    layer2_outputs(2187) <= '1';
    layer2_outputs(2188) <= not(layer1_outputs(2037));
    layer2_outputs(2189) <= not(layer1_outputs(1429));
    layer2_outputs(2190) <= not((layer1_outputs(1508)) and (layer1_outputs(827)));
    layer2_outputs(2191) <= not(layer1_outputs(432));
    layer2_outputs(2192) <= (layer1_outputs(1361)) or (layer1_outputs(2492));
    layer2_outputs(2193) <= not(layer1_outputs(4097));
    layer2_outputs(2194) <= (layer1_outputs(1979)) and not (layer1_outputs(2653));
    layer2_outputs(2195) <= (layer1_outputs(3439)) and not (layer1_outputs(3665));
    layer2_outputs(2196) <= layer1_outputs(500);
    layer2_outputs(2197) <= not(layer1_outputs(812));
    layer2_outputs(2198) <= (layer1_outputs(3964)) and (layer1_outputs(4988));
    layer2_outputs(2199) <= not(layer1_outputs(3509));
    layer2_outputs(2200) <= not(layer1_outputs(3731));
    layer2_outputs(2201) <= not((layer1_outputs(441)) and (layer1_outputs(2517)));
    layer2_outputs(2202) <= (layer1_outputs(4483)) and not (layer1_outputs(2268));
    layer2_outputs(2203) <= not(layer1_outputs(271));
    layer2_outputs(2204) <= not(layer1_outputs(4873));
    layer2_outputs(2205) <= layer1_outputs(4599);
    layer2_outputs(2206) <= layer1_outputs(2235);
    layer2_outputs(2207) <= (layer1_outputs(1785)) xor (layer1_outputs(4687));
    layer2_outputs(2208) <= layer1_outputs(4372);
    layer2_outputs(2209) <= not((layer1_outputs(1722)) or (layer1_outputs(2774)));
    layer2_outputs(2210) <= not(layer1_outputs(68)) or (layer1_outputs(1276));
    layer2_outputs(2211) <= not(layer1_outputs(1523));
    layer2_outputs(2212) <= not(layer1_outputs(1346)) or (layer1_outputs(242));
    layer2_outputs(2213) <= not(layer1_outputs(438)) or (layer1_outputs(3845));
    layer2_outputs(2214) <= (layer1_outputs(1294)) and (layer1_outputs(1784));
    layer2_outputs(2215) <= (layer1_outputs(1120)) or (layer1_outputs(1752));
    layer2_outputs(2216) <= not(layer1_outputs(3248));
    layer2_outputs(2217) <= not(layer1_outputs(1531));
    layer2_outputs(2218) <= not((layer1_outputs(5110)) or (layer1_outputs(765)));
    layer2_outputs(2219) <= (layer1_outputs(4529)) and not (layer1_outputs(1581));
    layer2_outputs(2220) <= not(layer1_outputs(3521)) or (layer1_outputs(815));
    layer2_outputs(2221) <= layer1_outputs(2556);
    layer2_outputs(2222) <= layer1_outputs(3357);
    layer2_outputs(2223) <= layer1_outputs(1343);
    layer2_outputs(2224) <= not(layer1_outputs(712)) or (layer1_outputs(1728));
    layer2_outputs(2225) <= '0';
    layer2_outputs(2226) <= layer1_outputs(4848);
    layer2_outputs(2227) <= layer1_outputs(624);
    layer2_outputs(2228) <= not((layer1_outputs(4022)) xor (layer1_outputs(1166)));
    layer2_outputs(2229) <= layer1_outputs(4530);
    layer2_outputs(2230) <= (layer1_outputs(1532)) xor (layer1_outputs(3436));
    layer2_outputs(2231) <= not(layer1_outputs(4990));
    layer2_outputs(2232) <= not((layer1_outputs(1956)) and (layer1_outputs(1375)));
    layer2_outputs(2233) <= not(layer1_outputs(4668));
    layer2_outputs(2234) <= not(layer1_outputs(1054));
    layer2_outputs(2235) <= not(layer1_outputs(4658));
    layer2_outputs(2236) <= layer1_outputs(4751);
    layer2_outputs(2237) <= (layer1_outputs(2478)) and (layer1_outputs(4996));
    layer2_outputs(2238) <= not((layer1_outputs(1094)) or (layer1_outputs(4941)));
    layer2_outputs(2239) <= not((layer1_outputs(2436)) and (layer1_outputs(1016)));
    layer2_outputs(2240) <= (layer1_outputs(4403)) and not (layer1_outputs(2507));
    layer2_outputs(2241) <= not((layer1_outputs(3970)) or (layer1_outputs(3679)));
    layer2_outputs(2242) <= not((layer1_outputs(3724)) or (layer1_outputs(1448)));
    layer2_outputs(2243) <= not(layer1_outputs(3969)) or (layer1_outputs(3164));
    layer2_outputs(2244) <= (layer1_outputs(3573)) and not (layer1_outputs(492));
    layer2_outputs(2245) <= (layer1_outputs(692)) and not (layer1_outputs(4939));
    layer2_outputs(2246) <= layer1_outputs(1883);
    layer2_outputs(2247) <= not(layer1_outputs(1974)) or (layer1_outputs(3628));
    layer2_outputs(2248) <= layer1_outputs(1474);
    layer2_outputs(2249) <= layer1_outputs(3378);
    layer2_outputs(2250) <= layer1_outputs(1736);
    layer2_outputs(2251) <= not((layer1_outputs(4733)) and (layer1_outputs(2655)));
    layer2_outputs(2252) <= not(layer1_outputs(3266));
    layer2_outputs(2253) <= layer1_outputs(1076);
    layer2_outputs(2254) <= (layer1_outputs(1164)) and not (layer1_outputs(3106));
    layer2_outputs(2255) <= not(layer1_outputs(4839));
    layer2_outputs(2256) <= not(layer1_outputs(1560)) or (layer1_outputs(2670));
    layer2_outputs(2257) <= (layer1_outputs(3350)) and not (layer1_outputs(1751));
    layer2_outputs(2258) <= '1';
    layer2_outputs(2259) <= layer1_outputs(2192);
    layer2_outputs(2260) <= not(layer1_outputs(3690));
    layer2_outputs(2261) <= not(layer1_outputs(3310)) or (layer1_outputs(702));
    layer2_outputs(2262) <= not(layer1_outputs(2649));
    layer2_outputs(2263) <= layer1_outputs(2118);
    layer2_outputs(2264) <= not(layer1_outputs(3964));
    layer2_outputs(2265) <= layer1_outputs(995);
    layer2_outputs(2266) <= (layer1_outputs(3222)) xor (layer1_outputs(1193));
    layer2_outputs(2267) <= not(layer1_outputs(1840)) or (layer1_outputs(4949));
    layer2_outputs(2268) <= (layer1_outputs(4249)) and not (layer1_outputs(3633));
    layer2_outputs(2269) <= layer1_outputs(3040);
    layer2_outputs(2270) <= not(layer1_outputs(4544));
    layer2_outputs(2271) <= not((layer1_outputs(2562)) xor (layer1_outputs(1148)));
    layer2_outputs(2272) <= layer1_outputs(1833);
    layer2_outputs(2273) <= (layer1_outputs(2629)) and (layer1_outputs(4978));
    layer2_outputs(2274) <= not(layer1_outputs(2575));
    layer2_outputs(2275) <= layer1_outputs(832);
    layer2_outputs(2276) <= not((layer1_outputs(3917)) and (layer1_outputs(4710)));
    layer2_outputs(2277) <= not(layer1_outputs(2164));
    layer2_outputs(2278) <= (layer1_outputs(1564)) xor (layer1_outputs(4254));
    layer2_outputs(2279) <= not((layer1_outputs(1579)) and (layer1_outputs(3952)));
    layer2_outputs(2280) <= not(layer1_outputs(4363)) or (layer1_outputs(760));
    layer2_outputs(2281) <= not(layer1_outputs(1837));
    layer2_outputs(2282) <= (layer1_outputs(3822)) and not (layer1_outputs(4296));
    layer2_outputs(2283) <= layer1_outputs(82);
    layer2_outputs(2284) <= not(layer1_outputs(4404)) or (layer1_outputs(4876));
    layer2_outputs(2285) <= layer1_outputs(2279);
    layer2_outputs(2286) <= layer1_outputs(1362);
    layer2_outputs(2287) <= not((layer1_outputs(4011)) or (layer1_outputs(1388)));
    layer2_outputs(2288) <= (layer1_outputs(192)) or (layer1_outputs(2355));
    layer2_outputs(2289) <= not((layer1_outputs(1007)) and (layer1_outputs(1249)));
    layer2_outputs(2290) <= (layer1_outputs(1029)) xor (layer1_outputs(3524));
    layer2_outputs(2291) <= not(layer1_outputs(4031));
    layer2_outputs(2292) <= not((layer1_outputs(3331)) or (layer1_outputs(4543)));
    layer2_outputs(2293) <= layer1_outputs(3268);
    layer2_outputs(2294) <= (layer1_outputs(1134)) xor (layer1_outputs(4416));
    layer2_outputs(2295) <= '1';
    layer2_outputs(2296) <= (layer1_outputs(2917)) or (layer1_outputs(4751));
    layer2_outputs(2297) <= not(layer1_outputs(4572));
    layer2_outputs(2298) <= not(layer1_outputs(2828));
    layer2_outputs(2299) <= (layer1_outputs(528)) xor (layer1_outputs(773));
    layer2_outputs(2300) <= not(layer1_outputs(3637)) or (layer1_outputs(2946));
    layer2_outputs(2301) <= (layer1_outputs(4789)) or (layer1_outputs(3591));
    layer2_outputs(2302) <= (layer1_outputs(4021)) and not (layer1_outputs(3335));
    layer2_outputs(2303) <= (layer1_outputs(2632)) and not (layer1_outputs(4636));
    layer2_outputs(2304) <= '1';
    layer2_outputs(2305) <= layer1_outputs(4925);
    layer2_outputs(2306) <= (layer1_outputs(1539)) or (layer1_outputs(2351));
    layer2_outputs(2307) <= (layer1_outputs(2404)) or (layer1_outputs(4890));
    layer2_outputs(2308) <= (layer1_outputs(2140)) or (layer1_outputs(4393));
    layer2_outputs(2309) <= not(layer1_outputs(3604));
    layer2_outputs(2310) <= not((layer1_outputs(703)) or (layer1_outputs(3370)));
    layer2_outputs(2311) <= not(layer1_outputs(4047));
    layer2_outputs(2312) <= not((layer1_outputs(98)) and (layer1_outputs(1191)));
    layer2_outputs(2313) <= (layer1_outputs(3620)) and not (layer1_outputs(3351));
    layer2_outputs(2314) <= not(layer1_outputs(119));
    layer2_outputs(2315) <= not((layer1_outputs(2891)) and (layer1_outputs(3204)));
    layer2_outputs(2316) <= not(layer1_outputs(244));
    layer2_outputs(2317) <= not(layer1_outputs(2271));
    layer2_outputs(2318) <= not(layer1_outputs(4954));
    layer2_outputs(2319) <= layer1_outputs(1104);
    layer2_outputs(2320) <= (layer1_outputs(2010)) and not (layer1_outputs(3791));
    layer2_outputs(2321) <= layer1_outputs(1116);
    layer2_outputs(2322) <= not((layer1_outputs(1559)) and (layer1_outputs(407)));
    layer2_outputs(2323) <= not(layer1_outputs(3542)) or (layer1_outputs(2689));
    layer2_outputs(2324) <= layer1_outputs(3537);
    layer2_outputs(2325) <= not(layer1_outputs(2440));
    layer2_outputs(2326) <= layer1_outputs(1396);
    layer2_outputs(2327) <= not((layer1_outputs(3082)) and (layer1_outputs(1245)));
    layer2_outputs(2328) <= layer1_outputs(4172);
    layer2_outputs(2329) <= layer1_outputs(610);
    layer2_outputs(2330) <= layer1_outputs(2320);
    layer2_outputs(2331) <= layer1_outputs(3339);
    layer2_outputs(2332) <= (layer1_outputs(2403)) and not (layer1_outputs(2202));
    layer2_outputs(2333) <= layer1_outputs(2423);
    layer2_outputs(2334) <= not(layer1_outputs(4174)) or (layer1_outputs(1093));
    layer2_outputs(2335) <= not(layer1_outputs(2525));
    layer2_outputs(2336) <= (layer1_outputs(337)) or (layer1_outputs(4264));
    layer2_outputs(2337) <= (layer1_outputs(793)) and not (layer1_outputs(4109));
    layer2_outputs(2338) <= not((layer1_outputs(2840)) and (layer1_outputs(3976)));
    layer2_outputs(2339) <= layer1_outputs(2107);
    layer2_outputs(2340) <= not((layer1_outputs(2675)) and (layer1_outputs(4572)));
    layer2_outputs(2341) <= not((layer1_outputs(1528)) or (layer1_outputs(1496)));
    layer2_outputs(2342) <= not(layer1_outputs(4260)) or (layer1_outputs(3214));
    layer2_outputs(2343) <= layer1_outputs(4160);
    layer2_outputs(2344) <= not(layer1_outputs(4170));
    layer2_outputs(2345) <= not((layer1_outputs(4594)) xor (layer1_outputs(3093)));
    layer2_outputs(2346) <= not(layer1_outputs(1806)) or (layer1_outputs(3217));
    layer2_outputs(2347) <= (layer1_outputs(427)) or (layer1_outputs(4549));
    layer2_outputs(2348) <= not((layer1_outputs(420)) or (layer1_outputs(4505)));
    layer2_outputs(2349) <= (layer1_outputs(433)) and not (layer1_outputs(3259));
    layer2_outputs(2350) <= not(layer1_outputs(4178));
    layer2_outputs(2351) <= not(layer1_outputs(606));
    layer2_outputs(2352) <= not((layer1_outputs(1607)) and (layer1_outputs(1798)));
    layer2_outputs(2353) <= layer1_outputs(1884);
    layer2_outputs(2354) <= (layer1_outputs(2243)) or (layer1_outputs(4046));
    layer2_outputs(2355) <= not(layer1_outputs(3321)) or (layer1_outputs(3429));
    layer2_outputs(2356) <= (layer1_outputs(3830)) xor (layer1_outputs(3958));
    layer2_outputs(2357) <= (layer1_outputs(4710)) and not (layer1_outputs(1672));
    layer2_outputs(2358) <= not(layer1_outputs(1013));
    layer2_outputs(2359) <= layer1_outputs(1542);
    layer2_outputs(2360) <= not(layer1_outputs(795));
    layer2_outputs(2361) <= not(layer1_outputs(2493));
    layer2_outputs(2362) <= not(layer1_outputs(460));
    layer2_outputs(2363) <= layer1_outputs(3363);
    layer2_outputs(2364) <= not(layer1_outputs(3048));
    layer2_outputs(2365) <= layer1_outputs(3265);
    layer2_outputs(2366) <= not(layer1_outputs(2679)) or (layer1_outputs(4031));
    layer2_outputs(2367) <= not(layer1_outputs(3452));
    layer2_outputs(2368) <= not(layer1_outputs(3884)) or (layer1_outputs(2457));
    layer2_outputs(2369) <= (layer1_outputs(3401)) or (layer1_outputs(3620));
    layer2_outputs(2370) <= (layer1_outputs(4792)) or (layer1_outputs(4127));
    layer2_outputs(2371) <= layer1_outputs(4230);
    layer2_outputs(2372) <= layer1_outputs(3863);
    layer2_outputs(2373) <= (layer1_outputs(3836)) or (layer1_outputs(544));
    layer2_outputs(2374) <= (layer1_outputs(2523)) or (layer1_outputs(4578));
    layer2_outputs(2375) <= not(layer1_outputs(3498)) or (layer1_outputs(2257));
    layer2_outputs(2376) <= (layer1_outputs(2297)) or (layer1_outputs(1254));
    layer2_outputs(2377) <= not(layer1_outputs(4954));
    layer2_outputs(2378) <= not((layer1_outputs(2001)) or (layer1_outputs(321)));
    layer2_outputs(2379) <= not(layer1_outputs(4186));
    layer2_outputs(2380) <= (layer1_outputs(2109)) or (layer1_outputs(2150));
    layer2_outputs(2381) <= (layer1_outputs(716)) and not (layer1_outputs(4893));
    layer2_outputs(2382) <= not(layer1_outputs(2775));
    layer2_outputs(2383) <= layer1_outputs(5079);
    layer2_outputs(2384) <= not((layer1_outputs(2221)) or (layer1_outputs(2908)));
    layer2_outputs(2385) <= layer1_outputs(2145);
    layer2_outputs(2386) <= layer1_outputs(859);
    layer2_outputs(2387) <= not(layer1_outputs(3909));
    layer2_outputs(2388) <= not((layer1_outputs(2106)) and (layer1_outputs(4322)));
    layer2_outputs(2389) <= not(layer1_outputs(781)) or (layer1_outputs(2685));
    layer2_outputs(2390) <= '0';
    layer2_outputs(2391) <= not(layer1_outputs(452));
    layer2_outputs(2392) <= not((layer1_outputs(4438)) xor (layer1_outputs(2464)));
    layer2_outputs(2393) <= not(layer1_outputs(2838));
    layer2_outputs(2394) <= (layer1_outputs(2883)) and not (layer1_outputs(2636));
    layer2_outputs(2395) <= not(layer1_outputs(3747));
    layer2_outputs(2396) <= not(layer1_outputs(3481));
    layer2_outputs(2397) <= not(layer1_outputs(3846));
    layer2_outputs(2398) <= layer1_outputs(1855);
    layer2_outputs(2399) <= not(layer1_outputs(3604)) or (layer1_outputs(4565));
    layer2_outputs(2400) <= not(layer1_outputs(3880));
    layer2_outputs(2401) <= '0';
    layer2_outputs(2402) <= (layer1_outputs(3005)) or (layer1_outputs(3559));
    layer2_outputs(2403) <= layer1_outputs(1936);
    layer2_outputs(2404) <= layer1_outputs(86);
    layer2_outputs(2405) <= not(layer1_outputs(2393));
    layer2_outputs(2406) <= (layer1_outputs(2855)) and not (layer1_outputs(3549));
    layer2_outputs(2407) <= (layer1_outputs(2459)) or (layer1_outputs(2451));
    layer2_outputs(2408) <= layer1_outputs(1906);
    layer2_outputs(2409) <= not(layer1_outputs(338));
    layer2_outputs(2410) <= (layer1_outputs(4724)) or (layer1_outputs(4405));
    layer2_outputs(2411) <= not(layer1_outputs(1528)) or (layer1_outputs(1035));
    layer2_outputs(2412) <= layer1_outputs(3700);
    layer2_outputs(2413) <= not((layer1_outputs(545)) or (layer1_outputs(3292)));
    layer2_outputs(2414) <= layer1_outputs(1712);
    layer2_outputs(2415) <= not((layer1_outputs(1892)) and (layer1_outputs(2339)));
    layer2_outputs(2416) <= (layer1_outputs(1446)) xor (layer1_outputs(1822));
    layer2_outputs(2417) <= not(layer1_outputs(3738));
    layer2_outputs(2418) <= layer1_outputs(2666);
    layer2_outputs(2419) <= layer1_outputs(4338);
    layer2_outputs(2420) <= layer1_outputs(930);
    layer2_outputs(2421) <= not(layer1_outputs(2647)) or (layer1_outputs(953));
    layer2_outputs(2422) <= layer1_outputs(4783);
    layer2_outputs(2423) <= layer1_outputs(280);
    layer2_outputs(2424) <= layer1_outputs(103);
    layer2_outputs(2425) <= not(layer1_outputs(3372));
    layer2_outputs(2426) <= not((layer1_outputs(4925)) or (layer1_outputs(4099)));
    layer2_outputs(2427) <= layer1_outputs(3230);
    layer2_outputs(2428) <= not(layer1_outputs(4672));
    layer2_outputs(2429) <= not(layer1_outputs(1219));
    layer2_outputs(2430) <= (layer1_outputs(2012)) or (layer1_outputs(1663));
    layer2_outputs(2431) <= not(layer1_outputs(3150)) or (layer1_outputs(4321));
    layer2_outputs(2432) <= not(layer1_outputs(3119));
    layer2_outputs(2433) <= (layer1_outputs(2117)) and not (layer1_outputs(4017));
    layer2_outputs(2434) <= layer1_outputs(2817);
    layer2_outputs(2435) <= layer1_outputs(3559);
    layer2_outputs(2436) <= (layer1_outputs(4920)) or (layer1_outputs(2155));
    layer2_outputs(2437) <= not((layer1_outputs(5050)) or (layer1_outputs(4477)));
    layer2_outputs(2438) <= not(layer1_outputs(1666));
    layer2_outputs(2439) <= layer1_outputs(1434);
    layer2_outputs(2440) <= not((layer1_outputs(4338)) and (layer1_outputs(2392)));
    layer2_outputs(2441) <= (layer1_outputs(1549)) and not (layer1_outputs(891));
    layer2_outputs(2442) <= '0';
    layer2_outputs(2443) <= not(layer1_outputs(652));
    layer2_outputs(2444) <= '0';
    layer2_outputs(2445) <= (layer1_outputs(1211)) and not (layer1_outputs(1818));
    layer2_outputs(2446) <= (layer1_outputs(1259)) and not (layer1_outputs(3102));
    layer2_outputs(2447) <= (layer1_outputs(3103)) or (layer1_outputs(699));
    layer2_outputs(2448) <= not(layer1_outputs(3433)) or (layer1_outputs(2719));
    layer2_outputs(2449) <= (layer1_outputs(3725)) xor (layer1_outputs(2547));
    layer2_outputs(2450) <= not(layer1_outputs(4229)) or (layer1_outputs(146));
    layer2_outputs(2451) <= (layer1_outputs(1273)) or (layer1_outputs(2470));
    layer2_outputs(2452) <= not(layer1_outputs(2723));
    layer2_outputs(2453) <= layer1_outputs(2230);
    layer2_outputs(2454) <= layer1_outputs(693);
    layer2_outputs(2455) <= not(layer1_outputs(880));
    layer2_outputs(2456) <= (layer1_outputs(1933)) or (layer1_outputs(2513));
    layer2_outputs(2457) <= not(layer1_outputs(2958));
    layer2_outputs(2458) <= (layer1_outputs(4621)) and (layer1_outputs(1439));
    layer2_outputs(2459) <= not((layer1_outputs(2978)) or (layer1_outputs(1795)));
    layer2_outputs(2460) <= not(layer1_outputs(4296));
    layer2_outputs(2461) <= not((layer1_outputs(2528)) xor (layer1_outputs(1766)));
    layer2_outputs(2462) <= not(layer1_outputs(1644));
    layer2_outputs(2463) <= not(layer1_outputs(4862));
    layer2_outputs(2464) <= (layer1_outputs(4136)) or (layer1_outputs(2954));
    layer2_outputs(2465) <= not(layer1_outputs(1986));
    layer2_outputs(2466) <= layer1_outputs(3229);
    layer2_outputs(2467) <= not(layer1_outputs(4279));
    layer2_outputs(2468) <= layer1_outputs(3405);
    layer2_outputs(2469) <= not(layer1_outputs(2960));
    layer2_outputs(2470) <= not((layer1_outputs(2645)) xor (layer1_outputs(419)));
    layer2_outputs(2471) <= (layer1_outputs(4663)) and not (layer1_outputs(1672));
    layer2_outputs(2472) <= layer1_outputs(399);
    layer2_outputs(2473) <= not((layer1_outputs(3041)) and (layer1_outputs(4506)));
    layer2_outputs(2474) <= (layer1_outputs(2823)) and not (layer1_outputs(4735));
    layer2_outputs(2475) <= layer1_outputs(2800);
    layer2_outputs(2476) <= not(layer1_outputs(4038));
    layer2_outputs(2477) <= '0';
    layer2_outputs(2478) <= not(layer1_outputs(4661)) or (layer1_outputs(2540));
    layer2_outputs(2479) <= not(layer1_outputs(5032)) or (layer1_outputs(523));
    layer2_outputs(2480) <= not(layer1_outputs(4290)) or (layer1_outputs(2052));
    layer2_outputs(2481) <= not((layer1_outputs(1598)) or (layer1_outputs(2621)));
    layer2_outputs(2482) <= (layer1_outputs(961)) and (layer1_outputs(2411));
    layer2_outputs(2483) <= not(layer1_outputs(576));
    layer2_outputs(2484) <= '1';
    layer2_outputs(2485) <= not(layer1_outputs(980));
    layer2_outputs(2486) <= not(layer1_outputs(3578));
    layer2_outputs(2487) <= not(layer1_outputs(4787)) or (layer1_outputs(4803));
    layer2_outputs(2488) <= (layer1_outputs(4622)) and (layer1_outputs(4171));
    layer2_outputs(2489) <= not(layer1_outputs(2134));
    layer2_outputs(2490) <= not((layer1_outputs(156)) xor (layer1_outputs(1106)));
    layer2_outputs(2491) <= not((layer1_outputs(1217)) and (layer1_outputs(664)));
    layer2_outputs(2492) <= layer1_outputs(928);
    layer2_outputs(2493) <= not(layer1_outputs(2065));
    layer2_outputs(2494) <= (layer1_outputs(524)) and not (layer1_outputs(2567));
    layer2_outputs(2495) <= layer1_outputs(3831);
    layer2_outputs(2496) <= layer1_outputs(979);
    layer2_outputs(2497) <= not(layer1_outputs(2390)) or (layer1_outputs(5118));
    layer2_outputs(2498) <= (layer1_outputs(3104)) and not (layer1_outputs(4679));
    layer2_outputs(2499) <= (layer1_outputs(2428)) or (layer1_outputs(4716));
    layer2_outputs(2500) <= not(layer1_outputs(764));
    layer2_outputs(2501) <= not(layer1_outputs(3455));
    layer2_outputs(2502) <= layer1_outputs(2726);
    layer2_outputs(2503) <= not(layer1_outputs(3833));
    layer2_outputs(2504) <= not(layer1_outputs(63)) or (layer1_outputs(1569));
    layer2_outputs(2505) <= layer1_outputs(3748);
    layer2_outputs(2506) <= layer1_outputs(2547);
    layer2_outputs(2507) <= (layer1_outputs(33)) xor (layer1_outputs(3022));
    layer2_outputs(2508) <= not(layer1_outputs(1454));
    layer2_outputs(2509) <= not(layer1_outputs(1057));
    layer2_outputs(2510) <= (layer1_outputs(1628)) xor (layer1_outputs(2998));
    layer2_outputs(2511) <= not(layer1_outputs(1993));
    layer2_outputs(2512) <= (layer1_outputs(5026)) or (layer1_outputs(3292));
    layer2_outputs(2513) <= not((layer1_outputs(2256)) or (layer1_outputs(2077)));
    layer2_outputs(2514) <= (layer1_outputs(223)) or (layer1_outputs(3669));
    layer2_outputs(2515) <= not(layer1_outputs(4706));
    layer2_outputs(2516) <= not(layer1_outputs(4490));
    layer2_outputs(2517) <= layer1_outputs(3465);
    layer2_outputs(2518) <= not(layer1_outputs(3064)) or (layer1_outputs(1337));
    layer2_outputs(2519) <= (layer1_outputs(2295)) and not (layer1_outputs(4130));
    layer2_outputs(2520) <= not(layer1_outputs(3059));
    layer2_outputs(2521) <= '0';
    layer2_outputs(2522) <= not(layer1_outputs(1370));
    layer2_outputs(2523) <= not((layer1_outputs(2598)) and (layer1_outputs(3507)));
    layer2_outputs(2524) <= not(layer1_outputs(1707));
    layer2_outputs(2525) <= (layer1_outputs(5044)) and not (layer1_outputs(3871));
    layer2_outputs(2526) <= layer1_outputs(4361);
    layer2_outputs(2527) <= not((layer1_outputs(3184)) or (layer1_outputs(657)));
    layer2_outputs(2528) <= layer1_outputs(1593);
    layer2_outputs(2529) <= (layer1_outputs(1640)) and not (layer1_outputs(231));
    layer2_outputs(2530) <= layer1_outputs(999);
    layer2_outputs(2531) <= not((layer1_outputs(4183)) and (layer1_outputs(938)));
    layer2_outputs(2532) <= layer1_outputs(1070);
    layer2_outputs(2533) <= layer1_outputs(1050);
    layer2_outputs(2534) <= not(layer1_outputs(3011)) or (layer1_outputs(5003));
    layer2_outputs(2535) <= not(layer1_outputs(4721));
    layer2_outputs(2536) <= not((layer1_outputs(3796)) or (layer1_outputs(3266)));
    layer2_outputs(2537) <= not((layer1_outputs(4840)) or (layer1_outputs(4841)));
    layer2_outputs(2538) <= not(layer1_outputs(2657)) or (layer1_outputs(1421));
    layer2_outputs(2539) <= not((layer1_outputs(1901)) or (layer1_outputs(4221)));
    layer2_outputs(2540) <= not(layer1_outputs(3715));
    layer2_outputs(2541) <= (layer1_outputs(1460)) and (layer1_outputs(4027));
    layer2_outputs(2542) <= not(layer1_outputs(681));
    layer2_outputs(2543) <= not(layer1_outputs(3376)) or (layer1_outputs(3687));
    layer2_outputs(2544) <= not(layer1_outputs(4013));
    layer2_outputs(2545) <= not((layer1_outputs(5076)) xor (layer1_outputs(5063)));
    layer2_outputs(2546) <= not(layer1_outputs(3992));
    layer2_outputs(2547) <= not(layer1_outputs(4230)) or (layer1_outputs(5054));
    layer2_outputs(2548) <= not(layer1_outputs(674));
    layer2_outputs(2549) <= (layer1_outputs(4937)) and not (layer1_outputs(4278));
    layer2_outputs(2550) <= (layer1_outputs(179)) and not (layer1_outputs(578));
    layer2_outputs(2551) <= (layer1_outputs(3471)) and not (layer1_outputs(1156));
    layer2_outputs(2552) <= layer1_outputs(4728);
    layer2_outputs(2553) <= not(layer1_outputs(3047));
    layer2_outputs(2554) <= layer1_outputs(634);
    layer2_outputs(2555) <= not(layer1_outputs(1664));
    layer2_outputs(2556) <= '0';
    layer2_outputs(2557) <= (layer1_outputs(2303)) and not (layer1_outputs(3326));
    layer2_outputs(2558) <= (layer1_outputs(1080)) or (layer1_outputs(4475));
    layer2_outputs(2559) <= not(layer1_outputs(2385));
    layer2_outputs(2560) <= not(layer1_outputs(1210));
    layer2_outputs(2561) <= not((layer1_outputs(3775)) or (layer1_outputs(675)));
    layer2_outputs(2562) <= not((layer1_outputs(3383)) and (layer1_outputs(96)));
    layer2_outputs(2563) <= layer1_outputs(158);
    layer2_outputs(2564) <= not(layer1_outputs(2623)) or (layer1_outputs(1823));
    layer2_outputs(2565) <= layer1_outputs(5030);
    layer2_outputs(2566) <= (layer1_outputs(2731)) and not (layer1_outputs(1860));
    layer2_outputs(2567) <= not((layer1_outputs(3807)) xor (layer1_outputs(708)));
    layer2_outputs(2568) <= (layer1_outputs(172)) and not (layer1_outputs(807));
    layer2_outputs(2569) <= (layer1_outputs(391)) and not (layer1_outputs(2766));
    layer2_outputs(2570) <= layer1_outputs(4822);
    layer2_outputs(2571) <= (layer1_outputs(632)) xor (layer1_outputs(4330));
    layer2_outputs(2572) <= not(layer1_outputs(776));
    layer2_outputs(2573) <= not((layer1_outputs(458)) xor (layer1_outputs(4402)));
    layer2_outputs(2574) <= not((layer1_outputs(4617)) xor (layer1_outputs(3899)));
    layer2_outputs(2575) <= (layer1_outputs(1368)) and not (layer1_outputs(5047));
    layer2_outputs(2576) <= not(layer1_outputs(2650));
    layer2_outputs(2577) <= not(layer1_outputs(138));
    layer2_outputs(2578) <= (layer1_outputs(774)) and not (layer1_outputs(167));
    layer2_outputs(2579) <= not((layer1_outputs(2468)) or (layer1_outputs(4851)));
    layer2_outputs(2580) <= not(layer1_outputs(1805));
    layer2_outputs(2581) <= (layer1_outputs(4507)) and not (layer1_outputs(4971));
    layer2_outputs(2582) <= (layer1_outputs(806)) and not (layer1_outputs(2640));
    layer2_outputs(2583) <= not(layer1_outputs(1457));
    layer2_outputs(2584) <= not(layer1_outputs(551)) or (layer1_outputs(1519));
    layer2_outputs(2585) <= layer1_outputs(463);
    layer2_outputs(2586) <= (layer1_outputs(3293)) and not (layer1_outputs(640));
    layer2_outputs(2587) <= layer1_outputs(2390);
    layer2_outputs(2588) <= not(layer1_outputs(4627));
    layer2_outputs(2589) <= layer1_outputs(3684);
    layer2_outputs(2590) <= not(layer1_outputs(900));
    layer2_outputs(2591) <= not(layer1_outputs(4182)) or (layer1_outputs(2748));
    layer2_outputs(2592) <= not(layer1_outputs(4006));
    layer2_outputs(2593) <= (layer1_outputs(1972)) and (layer1_outputs(4579));
    layer2_outputs(2594) <= layer1_outputs(1160);
    layer2_outputs(2595) <= layer1_outputs(4838);
    layer2_outputs(2596) <= layer1_outputs(4412);
    layer2_outputs(2597) <= not(layer1_outputs(1799));
    layer2_outputs(2598) <= (layer1_outputs(1891)) or (layer1_outputs(771));
    layer2_outputs(2599) <= not((layer1_outputs(4163)) and (layer1_outputs(3256)));
    layer2_outputs(2600) <= not((layer1_outputs(4910)) or (layer1_outputs(3019)));
    layer2_outputs(2601) <= (layer1_outputs(1701)) or (layer1_outputs(124));
    layer2_outputs(2602) <= not((layer1_outputs(502)) xor (layer1_outputs(4763)));
    layer2_outputs(2603) <= (layer1_outputs(1338)) and (layer1_outputs(2774));
    layer2_outputs(2604) <= (layer1_outputs(814)) and not (layer1_outputs(689));
    layer2_outputs(2605) <= (layer1_outputs(4033)) and not (layer1_outputs(2602));
    layer2_outputs(2606) <= layer1_outputs(2820);
    layer2_outputs(2607) <= layer1_outputs(1471);
    layer2_outputs(2608) <= not(layer1_outputs(2146)) or (layer1_outputs(1844));
    layer2_outputs(2609) <= not((layer1_outputs(3506)) or (layer1_outputs(4590)));
    layer2_outputs(2610) <= not(layer1_outputs(3957));
    layer2_outputs(2611) <= not(layer1_outputs(2818));
    layer2_outputs(2612) <= not((layer1_outputs(751)) and (layer1_outputs(2791)));
    layer2_outputs(2613) <= not((layer1_outputs(182)) xor (layer1_outputs(2594)));
    layer2_outputs(2614) <= layer1_outputs(1395);
    layer2_outputs(2615) <= (layer1_outputs(4452)) and not (layer1_outputs(3340));
    layer2_outputs(2616) <= layer1_outputs(932);
    layer2_outputs(2617) <= not(layer1_outputs(890));
    layer2_outputs(2618) <= (layer1_outputs(2933)) and not (layer1_outputs(2163));
    layer2_outputs(2619) <= layer1_outputs(1797);
    layer2_outputs(2620) <= not((layer1_outputs(2429)) xor (layer1_outputs(5119)));
    layer2_outputs(2621) <= (layer1_outputs(3013)) and not (layer1_outputs(1576));
    layer2_outputs(2622) <= not((layer1_outputs(4098)) and (layer1_outputs(2716)));
    layer2_outputs(2623) <= layer1_outputs(1993);
    layer2_outputs(2624) <= not((layer1_outputs(3808)) xor (layer1_outputs(3722)));
    layer2_outputs(2625) <= not((layer1_outputs(4944)) xor (layer1_outputs(85)));
    layer2_outputs(2626) <= not(layer1_outputs(1183));
    layer2_outputs(2627) <= not(layer1_outputs(1620)) or (layer1_outputs(996));
    layer2_outputs(2628) <= layer1_outputs(3249);
    layer2_outputs(2629) <= not((layer1_outputs(3986)) or (layer1_outputs(2206)));
    layer2_outputs(2630) <= not(layer1_outputs(2453));
    layer2_outputs(2631) <= not(layer1_outputs(4744));
    layer2_outputs(2632) <= layer1_outputs(2762);
    layer2_outputs(2633) <= not(layer1_outputs(5018));
    layer2_outputs(2634) <= not(layer1_outputs(2208));
    layer2_outputs(2635) <= layer1_outputs(2167);
    layer2_outputs(2636) <= layer1_outputs(341);
    layer2_outputs(2637) <= not(layer1_outputs(971));
    layer2_outputs(2638) <= not(layer1_outputs(4249)) or (layer1_outputs(1866));
    layer2_outputs(2639) <= layer1_outputs(4936);
    layer2_outputs(2640) <= layer1_outputs(1430);
    layer2_outputs(2641) <= not(layer1_outputs(4406));
    layer2_outputs(2642) <= (layer1_outputs(953)) and not (layer1_outputs(1151));
    layer2_outputs(2643) <= not((layer1_outputs(4770)) and (layer1_outputs(4783)));
    layer2_outputs(2644) <= (layer1_outputs(2233)) xor (layer1_outputs(1340));
    layer2_outputs(2645) <= layer1_outputs(93);
    layer2_outputs(2646) <= not(layer1_outputs(1711)) or (layer1_outputs(1296));
    layer2_outputs(2647) <= not((layer1_outputs(530)) or (layer1_outputs(181)));
    layer2_outputs(2648) <= layer1_outputs(3636);
    layer2_outputs(2649) <= not(layer1_outputs(1902));
    layer2_outputs(2650) <= not(layer1_outputs(3321));
    layer2_outputs(2651) <= not(layer1_outputs(1052));
    layer2_outputs(2652) <= layer1_outputs(1814);
    layer2_outputs(2653) <= (layer1_outputs(3781)) and not (layer1_outputs(4826));
    layer2_outputs(2654) <= not(layer1_outputs(2690));
    layer2_outputs(2655) <= not((layer1_outputs(688)) or (layer1_outputs(3304)));
    layer2_outputs(2656) <= not(layer1_outputs(1342)) or (layer1_outputs(4705));
    layer2_outputs(2657) <= layer1_outputs(694);
    layer2_outputs(2658) <= '0';
    layer2_outputs(2659) <= layer1_outputs(3325);
    layer2_outputs(2660) <= (layer1_outputs(2735)) xor (layer1_outputs(371));
    layer2_outputs(2661) <= not(layer1_outputs(387)) or (layer1_outputs(3177));
    layer2_outputs(2662) <= (layer1_outputs(608)) and not (layer1_outputs(3742));
    layer2_outputs(2663) <= not(layer1_outputs(66));
    layer2_outputs(2664) <= layer1_outputs(2483);
    layer2_outputs(2665) <= layer1_outputs(4417);
    layer2_outputs(2666) <= layer1_outputs(513);
    layer2_outputs(2667) <= layer1_outputs(3153);
    layer2_outputs(2668) <= layer1_outputs(581);
    layer2_outputs(2669) <= layer1_outputs(705);
    layer2_outputs(2670) <= not(layer1_outputs(357));
    layer2_outputs(2671) <= (layer1_outputs(5052)) and not (layer1_outputs(4068));
    layer2_outputs(2672) <= not(layer1_outputs(2275));
    layer2_outputs(2673) <= not((layer1_outputs(3856)) or (layer1_outputs(2263)));
    layer2_outputs(2674) <= (layer1_outputs(1456)) and not (layer1_outputs(3183));
    layer2_outputs(2675) <= not(layer1_outputs(3782));
    layer2_outputs(2676) <= layer1_outputs(2291);
    layer2_outputs(2677) <= (layer1_outputs(2569)) and not (layer1_outputs(3632));
    layer2_outputs(2678) <= not((layer1_outputs(1037)) and (layer1_outputs(1068)));
    layer2_outputs(2679) <= layer1_outputs(4346);
    layer2_outputs(2680) <= (layer1_outputs(901)) and not (layer1_outputs(4033));
    layer2_outputs(2681) <= not((layer1_outputs(4514)) or (layer1_outputs(893)));
    layer2_outputs(2682) <= not(layer1_outputs(1699));
    layer2_outputs(2683) <= not(layer1_outputs(1485));
    layer2_outputs(2684) <= not((layer1_outputs(1286)) and (layer1_outputs(2520)));
    layer2_outputs(2685) <= layer1_outputs(4089);
    layer2_outputs(2686) <= not(layer1_outputs(4874));
    layer2_outputs(2687) <= layer1_outputs(3678);
    layer2_outputs(2688) <= (layer1_outputs(860)) and not (layer1_outputs(161));
    layer2_outputs(2689) <= not(layer1_outputs(4297));
    layer2_outputs(2690) <= layer1_outputs(2927);
    layer2_outputs(2691) <= (layer1_outputs(3263)) or (layer1_outputs(5073));
    layer2_outputs(2692) <= not(layer1_outputs(908));
    layer2_outputs(2693) <= not(layer1_outputs(2218)) or (layer1_outputs(844));
    layer2_outputs(2694) <= layer1_outputs(4359);
    layer2_outputs(2695) <= layer1_outputs(3298);
    layer2_outputs(2696) <= not(layer1_outputs(4599));
    layer2_outputs(2697) <= (layer1_outputs(4837)) and (layer1_outputs(563));
    layer2_outputs(2698) <= (layer1_outputs(2677)) and (layer1_outputs(2433));
    layer2_outputs(2699) <= not(layer1_outputs(2186));
    layer2_outputs(2700) <= not(layer1_outputs(1671));
    layer2_outputs(2701) <= layer1_outputs(3904);
    layer2_outputs(2702) <= not((layer1_outputs(2172)) and (layer1_outputs(993)));
    layer2_outputs(2703) <= not(layer1_outputs(3207));
    layer2_outputs(2704) <= not(layer1_outputs(4506));
    layer2_outputs(2705) <= (layer1_outputs(4952)) or (layer1_outputs(3976));
    layer2_outputs(2706) <= not(layer1_outputs(5078)) or (layer1_outputs(4331));
    layer2_outputs(2707) <= not((layer1_outputs(2230)) xor (layer1_outputs(2048)));
    layer2_outputs(2708) <= (layer1_outputs(4821)) and not (layer1_outputs(1335));
    layer2_outputs(2709) <= (layer1_outputs(4055)) xor (layer1_outputs(2889));
    layer2_outputs(2710) <= not((layer1_outputs(4874)) xor (layer1_outputs(3771)));
    layer2_outputs(2711) <= (layer1_outputs(3891)) and (layer1_outputs(4559));
    layer2_outputs(2712) <= (layer1_outputs(1019)) and not (layer1_outputs(230));
    layer2_outputs(2713) <= not(layer1_outputs(66));
    layer2_outputs(2714) <= (layer1_outputs(102)) or (layer1_outputs(1741));
    layer2_outputs(2715) <= not((layer1_outputs(3306)) and (layer1_outputs(105)));
    layer2_outputs(2716) <= not(layer1_outputs(4601)) or (layer1_outputs(763));
    layer2_outputs(2717) <= layer1_outputs(292);
    layer2_outputs(2718) <= not(layer1_outputs(2677));
    layer2_outputs(2719) <= layer1_outputs(2684);
    layer2_outputs(2720) <= layer1_outputs(4799);
    layer2_outputs(2721) <= not(layer1_outputs(2259));
    layer2_outputs(2722) <= (layer1_outputs(2638)) xor (layer1_outputs(4968));
    layer2_outputs(2723) <= layer1_outputs(1567);
    layer2_outputs(2724) <= layer1_outputs(4025);
    layer2_outputs(2725) <= not(layer1_outputs(3642)) or (layer1_outputs(2465));
    layer2_outputs(2726) <= not(layer1_outputs(3336)) or (layer1_outputs(851));
    layer2_outputs(2727) <= not((layer1_outputs(2161)) and (layer1_outputs(3498)));
    layer2_outputs(2728) <= (layer1_outputs(2235)) or (layer1_outputs(722));
    layer2_outputs(2729) <= layer1_outputs(4898);
    layer2_outputs(2730) <= layer1_outputs(894);
    layer2_outputs(2731) <= not(layer1_outputs(4219)) or (layer1_outputs(1027));
    layer2_outputs(2732) <= not((layer1_outputs(3378)) or (layer1_outputs(3612)));
    layer2_outputs(2733) <= (layer1_outputs(2196)) and (layer1_outputs(2149));
    layer2_outputs(2734) <= not((layer1_outputs(2732)) and (layer1_outputs(4434)));
    layer2_outputs(2735) <= not(layer1_outputs(1767));
    layer2_outputs(2736) <= layer1_outputs(5113);
    layer2_outputs(2737) <= (layer1_outputs(3239)) and not (layer1_outputs(3194));
    layer2_outputs(2738) <= (layer1_outputs(4300)) and not (layer1_outputs(1546));
    layer2_outputs(2739) <= layer1_outputs(15);
    layer2_outputs(2740) <= layer1_outputs(4273);
    layer2_outputs(2741) <= (layer1_outputs(1830)) and not (layer1_outputs(5093));
    layer2_outputs(2742) <= not((layer1_outputs(4798)) xor (layer1_outputs(2712)));
    layer2_outputs(2743) <= '1';
    layer2_outputs(2744) <= layer1_outputs(4387);
    layer2_outputs(2745) <= not(layer1_outputs(4972));
    layer2_outputs(2746) <= not(layer1_outputs(3238)) or (layer1_outputs(4360));
    layer2_outputs(2747) <= layer1_outputs(933);
    layer2_outputs(2748) <= not(layer1_outputs(3170)) or (layer1_outputs(1105));
    layer2_outputs(2749) <= layer1_outputs(1700);
    layer2_outputs(2750) <= not(layer1_outputs(3056)) or (layer1_outputs(213));
    layer2_outputs(2751) <= layer1_outputs(3012);
    layer2_outputs(2752) <= (layer1_outputs(1126)) and not (layer1_outputs(4771));
    layer2_outputs(2753) <= (layer1_outputs(1283)) xor (layer1_outputs(3195));
    layer2_outputs(2754) <= not(layer1_outputs(4037));
    layer2_outputs(2755) <= not(layer1_outputs(2914));
    layer2_outputs(2756) <= not(layer1_outputs(3732));
    layer2_outputs(2757) <= (layer1_outputs(3189)) xor (layer1_outputs(3212));
    layer2_outputs(2758) <= not(layer1_outputs(3437)) or (layer1_outputs(2588));
    layer2_outputs(2759) <= (layer1_outputs(3653)) and not (layer1_outputs(2564));
    layer2_outputs(2760) <= (layer1_outputs(3605)) and not (layer1_outputs(3756));
    layer2_outputs(2761) <= (layer1_outputs(4998)) and (layer1_outputs(1078));
    layer2_outputs(2762) <= layer1_outputs(2357);
    layer2_outputs(2763) <= layer1_outputs(3267);
    layer2_outputs(2764) <= (layer1_outputs(1813)) and not (layer1_outputs(4980));
    layer2_outputs(2765) <= layer1_outputs(2550);
    layer2_outputs(2766) <= not(layer1_outputs(885));
    layer2_outputs(2767) <= not(layer1_outputs(2391));
    layer2_outputs(2768) <= not(layer1_outputs(318)) or (layer1_outputs(2889));
    layer2_outputs(2769) <= (layer1_outputs(3329)) or (layer1_outputs(644));
    layer2_outputs(2770) <= not(layer1_outputs(62));
    layer2_outputs(2771) <= (layer1_outputs(4597)) and not (layer1_outputs(2718));
    layer2_outputs(2772) <= not(layer1_outputs(3802)) or (layer1_outputs(4857));
    layer2_outputs(2773) <= not(layer1_outputs(3826));
    layer2_outputs(2774) <= not(layer1_outputs(2100));
    layer2_outputs(2775) <= not(layer1_outputs(4931));
    layer2_outputs(2776) <= (layer1_outputs(2041)) and not (layer1_outputs(279));
    layer2_outputs(2777) <= layer1_outputs(2793);
    layer2_outputs(2778) <= layer1_outputs(3707);
    layer2_outputs(2779) <= not(layer1_outputs(1495));
    layer2_outputs(2780) <= not(layer1_outputs(3752));
    layer2_outputs(2781) <= (layer1_outputs(3226)) or (layer1_outputs(297));
    layer2_outputs(2782) <= layer1_outputs(2545);
    layer2_outputs(2783) <= not((layer1_outputs(1329)) and (layer1_outputs(3966)));
    layer2_outputs(2784) <= not(layer1_outputs(4440));
    layer2_outputs(2785) <= layer1_outputs(4208);
    layer2_outputs(2786) <= not((layer1_outputs(1152)) or (layer1_outputs(4494)));
    layer2_outputs(2787) <= not(layer1_outputs(5063));
    layer2_outputs(2788) <= not((layer1_outputs(4844)) or (layer1_outputs(500)));
    layer2_outputs(2789) <= (layer1_outputs(4829)) and not (layer1_outputs(258));
    layer2_outputs(2790) <= layer1_outputs(570);
    layer2_outputs(2791) <= (layer1_outputs(2011)) or (layer1_outputs(4876));
    layer2_outputs(2792) <= layer1_outputs(2389);
    layer2_outputs(2793) <= not(layer1_outputs(3421)) or (layer1_outputs(3432));
    layer2_outputs(2794) <= not(layer1_outputs(3507)) or (layer1_outputs(981));
    layer2_outputs(2795) <= (layer1_outputs(1744)) xor (layer1_outputs(222));
    layer2_outputs(2796) <= not((layer1_outputs(820)) or (layer1_outputs(2541)));
    layer2_outputs(2797) <= layer1_outputs(3695);
    layer2_outputs(2798) <= not(layer1_outputs(2825)) or (layer1_outputs(145));
    layer2_outputs(2799) <= not((layer1_outputs(4180)) xor (layer1_outputs(4451)));
    layer2_outputs(2800) <= '1';
    layer2_outputs(2801) <= not(layer1_outputs(2799));
    layer2_outputs(2802) <= layer1_outputs(3791);
    layer2_outputs(2803) <= not((layer1_outputs(940)) and (layer1_outputs(2493)));
    layer2_outputs(2804) <= not(layer1_outputs(722));
    layer2_outputs(2805) <= not(layer1_outputs(1650)) or (layer1_outputs(2826));
    layer2_outputs(2806) <= not(layer1_outputs(3740));
    layer2_outputs(2807) <= not(layer1_outputs(4345));
    layer2_outputs(2808) <= not(layer1_outputs(403));
    layer2_outputs(2809) <= not(layer1_outputs(593));
    layer2_outputs(2810) <= not(layer1_outputs(4850));
    layer2_outputs(2811) <= (layer1_outputs(898)) xor (layer1_outputs(1960));
    layer2_outputs(2812) <= not(layer1_outputs(2985));
    layer2_outputs(2813) <= not(layer1_outputs(4704));
    layer2_outputs(2814) <= not((layer1_outputs(5049)) or (layer1_outputs(2722)));
    layer2_outputs(2815) <= not(layer1_outputs(4571));
    layer2_outputs(2816) <= not(layer1_outputs(1327));
    layer2_outputs(2817) <= layer1_outputs(3399);
    layer2_outputs(2818) <= not(layer1_outputs(3413));
    layer2_outputs(2819) <= layer1_outputs(5109);
    layer2_outputs(2820) <= not(layer1_outputs(4501));
    layer2_outputs(2821) <= not((layer1_outputs(1064)) and (layer1_outputs(1948)));
    layer2_outputs(2822) <= not((layer1_outputs(2088)) and (layer1_outputs(2104)));
    layer2_outputs(2823) <= (layer1_outputs(750)) and not (layer1_outputs(1079));
    layer2_outputs(2824) <= '1';
    layer2_outputs(2825) <= not(layer1_outputs(988));
    layer2_outputs(2826) <= not(layer1_outputs(3469));
    layer2_outputs(2827) <= not((layer1_outputs(1727)) xor (layer1_outputs(1266)));
    layer2_outputs(2828) <= (layer1_outputs(1216)) and (layer1_outputs(579));
    layer2_outputs(2829) <= layer1_outputs(4992);
    layer2_outputs(2830) <= (layer1_outputs(800)) and not (layer1_outputs(195));
    layer2_outputs(2831) <= (layer1_outputs(2982)) and not (layer1_outputs(4528));
    layer2_outputs(2832) <= layer1_outputs(201);
    layer2_outputs(2833) <= not((layer1_outputs(2732)) or (layer1_outputs(4795)));
    layer2_outputs(2834) <= not(layer1_outputs(4739));
    layer2_outputs(2835) <= not(layer1_outputs(91)) or (layer1_outputs(4505));
    layer2_outputs(2836) <= not(layer1_outputs(992));
    layer2_outputs(2837) <= layer1_outputs(2057);
    layer2_outputs(2838) <= (layer1_outputs(3639)) and not (layer1_outputs(3233));
    layer2_outputs(2839) <= not((layer1_outputs(3531)) and (layer1_outputs(2472)));
    layer2_outputs(2840) <= (layer1_outputs(4303)) and not (layer1_outputs(4370));
    layer2_outputs(2841) <= not((layer1_outputs(2344)) or (layer1_outputs(3703)));
    layer2_outputs(2842) <= not(layer1_outputs(3924));
    layer2_outputs(2843) <= layer1_outputs(3009);
    layer2_outputs(2844) <= not((layer1_outputs(4516)) or (layer1_outputs(3873)));
    layer2_outputs(2845) <= not((layer1_outputs(3043)) xor (layer1_outputs(3006)));
    layer2_outputs(2846) <= not(layer1_outputs(2056));
    layer2_outputs(2847) <= (layer1_outputs(3086)) and not (layer1_outputs(3166));
    layer2_outputs(2848) <= layer1_outputs(4361);
    layer2_outputs(2849) <= not(layer1_outputs(1977));
    layer2_outputs(2850) <= not(layer1_outputs(4713)) or (layer1_outputs(197));
    layer2_outputs(2851) <= layer1_outputs(593);
    layer2_outputs(2852) <= (layer1_outputs(2456)) and not (layer1_outputs(1));
    layer2_outputs(2853) <= (layer1_outputs(4334)) and not (layer1_outputs(588));
    layer2_outputs(2854) <= (layer1_outputs(1577)) and (layer1_outputs(2942));
    layer2_outputs(2855) <= (layer1_outputs(1372)) and not (layer1_outputs(1850));
    layer2_outputs(2856) <= (layer1_outputs(2449)) xor (layer1_outputs(386));
    layer2_outputs(2857) <= layer1_outputs(886);
    layer2_outputs(2858) <= not(layer1_outputs(3316));
    layer2_outputs(2859) <= (layer1_outputs(2733)) and not (layer1_outputs(3252));
    layer2_outputs(2860) <= layer1_outputs(3813);
    layer2_outputs(2861) <= not((layer1_outputs(4431)) or (layer1_outputs(324)));
    layer2_outputs(2862) <= not((layer1_outputs(3708)) or (layer1_outputs(3248)));
    layer2_outputs(2863) <= not(layer1_outputs(3974));
    layer2_outputs(2864) <= (layer1_outputs(4305)) and (layer1_outputs(2947));
    layer2_outputs(2865) <= layer1_outputs(3500);
    layer2_outputs(2866) <= layer1_outputs(3751);
    layer2_outputs(2867) <= layer1_outputs(4049);
    layer2_outputs(2868) <= not((layer1_outputs(2454)) xor (layer1_outputs(3798)));
    layer2_outputs(2869) <= (layer1_outputs(4312)) or (layer1_outputs(3416));
    layer2_outputs(2870) <= layer1_outputs(2859);
    layer2_outputs(2871) <= layer1_outputs(1045);
    layer2_outputs(2872) <= layer1_outputs(2198);
    layer2_outputs(2873) <= not(layer1_outputs(1943)) or (layer1_outputs(5));
    layer2_outputs(2874) <= not((layer1_outputs(1573)) and (layer1_outputs(2526)));
    layer2_outputs(2875) <= (layer1_outputs(3599)) and (layer1_outputs(2581));
    layer2_outputs(2876) <= (layer1_outputs(4541)) and not (layer1_outputs(1833));
    layer2_outputs(2877) <= '1';
    layer2_outputs(2878) <= layer1_outputs(2805);
    layer2_outputs(2879) <= layer1_outputs(4464);
    layer2_outputs(2880) <= layer1_outputs(2707);
    layer2_outputs(2881) <= layer1_outputs(4533);
    layer2_outputs(2882) <= not(layer1_outputs(2351));
    layer2_outputs(2883) <= not((layer1_outputs(4757)) xor (layer1_outputs(3629)));
    layer2_outputs(2884) <= not(layer1_outputs(3003)) or (layer1_outputs(1092));
    layer2_outputs(2885) <= (layer1_outputs(3814)) and not (layer1_outputs(2897));
    layer2_outputs(2886) <= (layer1_outputs(1332)) xor (layer1_outputs(1172));
    layer2_outputs(2887) <= layer1_outputs(1095);
    layer2_outputs(2888) <= (layer1_outputs(3319)) and (layer1_outputs(2610));
    layer2_outputs(2889) <= (layer1_outputs(5066)) and not (layer1_outputs(3280));
    layer2_outputs(2890) <= (layer1_outputs(3324)) or (layer1_outputs(3645));
    layer2_outputs(2891) <= not((layer1_outputs(1003)) or (layer1_outputs(228)));
    layer2_outputs(2892) <= (layer1_outputs(1982)) and not (layer1_outputs(3675));
    layer2_outputs(2893) <= layer1_outputs(4043);
    layer2_outputs(2894) <= (layer1_outputs(2542)) and not (layer1_outputs(3652));
    layer2_outputs(2895) <= layer1_outputs(3499);
    layer2_outputs(2896) <= layer1_outputs(4417);
    layer2_outputs(2897) <= (layer1_outputs(3775)) and not (layer1_outputs(2524));
    layer2_outputs(2898) <= layer1_outputs(2370);
    layer2_outputs(2899) <= not((layer1_outputs(2117)) and (layer1_outputs(1039)));
    layer2_outputs(2900) <= not(layer1_outputs(5118));
    layer2_outputs(2901) <= not(layer1_outputs(243)) or (layer1_outputs(1379));
    layer2_outputs(2902) <= layer1_outputs(3373);
    layer2_outputs(2903) <= not(layer1_outputs(1190)) or (layer1_outputs(4455));
    layer2_outputs(2904) <= layer1_outputs(4109);
    layer2_outputs(2905) <= (layer1_outputs(4483)) and (layer1_outputs(2058));
    layer2_outputs(2906) <= layer1_outputs(2540);
    layer2_outputs(2907) <= (layer1_outputs(2904)) and not (layer1_outputs(3609));
    layer2_outputs(2908) <= (layer1_outputs(4879)) and not (layer1_outputs(4865));
    layer2_outputs(2909) <= layer1_outputs(2961);
    layer2_outputs(2910) <= layer1_outputs(4091);
    layer2_outputs(2911) <= not((layer1_outputs(2047)) or (layer1_outputs(34)));
    layer2_outputs(2912) <= not(layer1_outputs(4762));
    layer2_outputs(2913) <= not(layer1_outputs(216));
    layer2_outputs(2914) <= not(layer1_outputs(1701));
    layer2_outputs(2915) <= layer1_outputs(1715);
    layer2_outputs(2916) <= not(layer1_outputs(4986));
    layer2_outputs(2917) <= layer1_outputs(4050);
    layer2_outputs(2918) <= (layer1_outputs(3914)) or (layer1_outputs(3686));
    layer2_outputs(2919) <= not(layer1_outputs(4515));
    layer2_outputs(2920) <= (layer1_outputs(409)) or (layer1_outputs(2349));
    layer2_outputs(2921) <= layer1_outputs(3339);
    layer2_outputs(2922) <= not(layer1_outputs(754)) or (layer1_outputs(1478));
    layer2_outputs(2923) <= (layer1_outputs(1302)) and (layer1_outputs(1197));
    layer2_outputs(2924) <= not((layer1_outputs(3353)) or (layer1_outputs(1341)));
    layer2_outputs(2925) <= not(layer1_outputs(1517));
    layer2_outputs(2926) <= (layer1_outputs(347)) xor (layer1_outputs(2692));
    layer2_outputs(2927) <= not(layer1_outputs(3984)) or (layer1_outputs(516));
    layer2_outputs(2928) <= layer1_outputs(1369);
    layer2_outputs(2929) <= not(layer1_outputs(2343));
    layer2_outputs(2930) <= (layer1_outputs(4606)) xor (layer1_outputs(2595));
    layer2_outputs(2931) <= not((layer1_outputs(1746)) or (layer1_outputs(499)));
    layer2_outputs(2932) <= layer1_outputs(3561);
    layer2_outputs(2933) <= layer1_outputs(955);
    layer2_outputs(2934) <= (layer1_outputs(669)) xor (layer1_outputs(2093));
    layer2_outputs(2935) <= (layer1_outputs(999)) and not (layer1_outputs(1405));
    layer2_outputs(2936) <= (layer1_outputs(210)) or (layer1_outputs(4019));
    layer2_outputs(2937) <= '1';
    layer2_outputs(2938) <= not(layer1_outputs(2272));
    layer2_outputs(2939) <= not(layer1_outputs(1048)) or (layer1_outputs(4207));
    layer2_outputs(2940) <= not((layer1_outputs(240)) or (layer1_outputs(4642)));
    layer2_outputs(2941) <= (layer1_outputs(3374)) and not (layer1_outputs(2708));
    layer2_outputs(2942) <= layer1_outputs(2472);
    layer2_outputs(2943) <= not(layer1_outputs(2166));
    layer2_outputs(2944) <= layer1_outputs(2744);
    layer2_outputs(2945) <= layer1_outputs(1801);
    layer2_outputs(2946) <= not((layer1_outputs(1199)) xor (layer1_outputs(1952)));
    layer2_outputs(2947) <= '0';
    layer2_outputs(2948) <= not((layer1_outputs(2886)) xor (layer1_outputs(1735)));
    layer2_outputs(2949) <= (layer1_outputs(1000)) and (layer1_outputs(2809));
    layer2_outputs(2950) <= (layer1_outputs(345)) or (layer1_outputs(3980));
    layer2_outputs(2951) <= (layer1_outputs(3965)) or (layer1_outputs(3941));
    layer2_outputs(2952) <= not(layer1_outputs(4724));
    layer2_outputs(2953) <= not(layer1_outputs(2964));
    layer2_outputs(2954) <= layer1_outputs(3188);
    layer2_outputs(2955) <= not(layer1_outputs(3819));
    layer2_outputs(2956) <= (layer1_outputs(733)) xor (layer1_outputs(3502));
    layer2_outputs(2957) <= not(layer1_outputs(327));
    layer2_outputs(2958) <= not(layer1_outputs(103));
    layer2_outputs(2959) <= not(layer1_outputs(2477));
    layer2_outputs(2960) <= not(layer1_outputs(3114));
    layer2_outputs(2961) <= (layer1_outputs(3583)) and not (layer1_outputs(2141));
    layer2_outputs(2962) <= not(layer1_outputs(162));
    layer2_outputs(2963) <= (layer1_outputs(3152)) and (layer1_outputs(2332));
    layer2_outputs(2964) <= (layer1_outputs(4394)) or (layer1_outputs(4895));
    layer2_outputs(2965) <= not((layer1_outputs(835)) and (layer1_outputs(747)));
    layer2_outputs(2966) <= (layer1_outputs(4247)) and (layer1_outputs(306));
    layer2_outputs(2967) <= (layer1_outputs(4952)) and not (layer1_outputs(2314));
    layer2_outputs(2968) <= not(layer1_outputs(975)) or (layer1_outputs(518));
    layer2_outputs(2969) <= not((layer1_outputs(3627)) xor (layer1_outputs(2950)));
    layer2_outputs(2970) <= not(layer1_outputs(1571));
    layer2_outputs(2971) <= layer1_outputs(4211);
    layer2_outputs(2972) <= not(layer1_outputs(1886));
    layer2_outputs(2973) <= not(layer1_outputs(4161));
    layer2_outputs(2974) <= not(layer1_outputs(674));
    layer2_outputs(2975) <= not(layer1_outputs(3138)) or (layer1_outputs(1944));
    layer2_outputs(2976) <= (layer1_outputs(636)) and not (layer1_outputs(3878));
    layer2_outputs(2977) <= not(layer1_outputs(302));
    layer2_outputs(2978) <= (layer1_outputs(264)) and (layer1_outputs(3754));
    layer2_outputs(2979) <= layer1_outputs(3545);
    layer2_outputs(2980) <= not(layer1_outputs(3363));
    layer2_outputs(2981) <= not(layer1_outputs(2589));
    layer2_outputs(2982) <= not(layer1_outputs(3874));
    layer2_outputs(2983) <= not(layer1_outputs(2137));
    layer2_outputs(2984) <= (layer1_outputs(4971)) or (layer1_outputs(175));
    layer2_outputs(2985) <= layer1_outputs(1740);
    layer2_outputs(2986) <= layer1_outputs(4285);
    layer2_outputs(2987) <= not((layer1_outputs(4726)) or (layer1_outputs(3687)));
    layer2_outputs(2988) <= not(layer1_outputs(4189));
    layer2_outputs(2989) <= (layer1_outputs(802)) and not (layer1_outputs(850));
    layer2_outputs(2990) <= layer1_outputs(4545);
    layer2_outputs(2991) <= (layer1_outputs(1042)) and not (layer1_outputs(3461));
    layer2_outputs(2992) <= not(layer1_outputs(434)) or (layer1_outputs(1759));
    layer2_outputs(2993) <= (layer1_outputs(4706)) and not (layer1_outputs(148));
    layer2_outputs(2994) <= (layer1_outputs(624)) and not (layer1_outputs(81));
    layer2_outputs(2995) <= (layer1_outputs(2264)) and not (layer1_outputs(3985));
    layer2_outputs(2996) <= not(layer1_outputs(962));
    layer2_outputs(2997) <= layer1_outputs(207);
    layer2_outputs(2998) <= not(layer1_outputs(3557));
    layer2_outputs(2999) <= not(layer1_outputs(2852)) or (layer1_outputs(5040));
    layer2_outputs(3000) <= not(layer1_outputs(607));
    layer2_outputs(3001) <= not(layer1_outputs(2626));
    layer2_outputs(3002) <= not(layer1_outputs(2452)) or (layer1_outputs(921));
    layer2_outputs(3003) <= not(layer1_outputs(4995));
    layer2_outputs(3004) <= not(layer1_outputs(2816));
    layer2_outputs(3005) <= not((layer1_outputs(998)) or (layer1_outputs(3395)));
    layer2_outputs(3006) <= not((layer1_outputs(4774)) xor (layer1_outputs(456)));
    layer2_outputs(3007) <= not(layer1_outputs(1335));
    layer2_outputs(3008) <= layer1_outputs(183);
    layer2_outputs(3009) <= not(layer1_outputs(2154));
    layer2_outputs(3010) <= not(layer1_outputs(3022));
    layer2_outputs(3011) <= layer1_outputs(1390);
    layer2_outputs(3012) <= layer1_outputs(2242);
    layer2_outputs(3013) <= not((layer1_outputs(4457)) and (layer1_outputs(756)));
    layer2_outputs(3014) <= not((layer1_outputs(3458)) or (layer1_outputs(2600)));
    layer2_outputs(3015) <= layer1_outputs(1488);
    layer2_outputs(3016) <= layer1_outputs(3938);
    layer2_outputs(3017) <= (layer1_outputs(3926)) or (layer1_outputs(928));
    layer2_outputs(3018) <= layer1_outputs(4059);
    layer2_outputs(3019) <= not(layer1_outputs(3478));
    layer2_outputs(3020) <= (layer1_outputs(1762)) and not (layer1_outputs(3224));
    layer2_outputs(3021) <= (layer1_outputs(1280)) xor (layer1_outputs(2723));
    layer2_outputs(3022) <= not(layer1_outputs(1182)) or (layer1_outputs(4588));
    layer2_outputs(3023) <= (layer1_outputs(4667)) xor (layer1_outputs(2515));
    layer2_outputs(3024) <= not(layer1_outputs(1388)) or (layer1_outputs(2278));
    layer2_outputs(3025) <= (layer1_outputs(4820)) and not (layer1_outputs(4959));
    layer2_outputs(3026) <= (layer1_outputs(2231)) or (layer1_outputs(2144));
    layer2_outputs(3027) <= (layer1_outputs(1170)) and not (layer1_outputs(302));
    layer2_outputs(3028) <= not((layer1_outputs(4863)) and (layer1_outputs(723)));
    layer2_outputs(3029) <= not(layer1_outputs(927));
    layer2_outputs(3030) <= not(layer1_outputs(4587));
    layer2_outputs(3031) <= '1';
    layer2_outputs(3032) <= (layer1_outputs(1964)) or (layer1_outputs(276));
    layer2_outputs(3033) <= '0';
    layer2_outputs(3034) <= not(layer1_outputs(3862));
    layer2_outputs(3035) <= (layer1_outputs(4202)) and not (layer1_outputs(633));
    layer2_outputs(3036) <= (layer1_outputs(1047)) xor (layer1_outputs(1924));
    layer2_outputs(3037) <= (layer1_outputs(3566)) and not (layer1_outputs(2835));
    layer2_outputs(3038) <= layer1_outputs(1236);
    layer2_outputs(3039) <= not(layer1_outputs(3442));
    layer2_outputs(3040) <= not(layer1_outputs(2534)) or (layer1_outputs(3962));
    layer2_outputs(3041) <= not((layer1_outputs(4415)) xor (layer1_outputs(3630)));
    layer2_outputs(3042) <= layer1_outputs(3572);
    layer2_outputs(3043) <= not(layer1_outputs(487));
    layer2_outputs(3044) <= not(layer1_outputs(2387));
    layer2_outputs(3045) <= (layer1_outputs(1040)) and not (layer1_outputs(2523));
    layer2_outputs(3046) <= layer1_outputs(4331);
    layer2_outputs(3047) <= not(layer1_outputs(1641));
    layer2_outputs(3048) <= not(layer1_outputs(4703));
    layer2_outputs(3049) <= not(layer1_outputs(4830));
    layer2_outputs(3050) <= (layer1_outputs(1590)) and not (layer1_outputs(1365));
    layer2_outputs(3051) <= (layer1_outputs(252)) and (layer1_outputs(190));
    layer2_outputs(3052) <= '1';
    layer2_outputs(3053) <= layer1_outputs(567);
    layer2_outputs(3054) <= layer1_outputs(1677);
    layer2_outputs(3055) <= layer1_outputs(1322);
    layer2_outputs(3056) <= not((layer1_outputs(423)) xor (layer1_outputs(627)));
    layer2_outputs(3057) <= not(layer1_outputs(4371)) or (layer1_outputs(1929));
    layer2_outputs(3058) <= not(layer1_outputs(1623));
    layer2_outputs(3059) <= (layer1_outputs(828)) and not (layer1_outputs(587));
    layer2_outputs(3060) <= (layer1_outputs(3550)) and not (layer1_outputs(2994));
    layer2_outputs(3061) <= (layer1_outputs(4697)) and not (layer1_outputs(995));
    layer2_outputs(3062) <= not((layer1_outputs(379)) and (layer1_outputs(1671)));
    layer2_outputs(3063) <= not(layer1_outputs(1510)) or (layer1_outputs(2633));
    layer2_outputs(3064) <= (layer1_outputs(4041)) and not (layer1_outputs(471));
    layer2_outputs(3065) <= layer1_outputs(3880);
    layer2_outputs(3066) <= (layer1_outputs(2807)) and (layer1_outputs(4776));
    layer2_outputs(3067) <= layer1_outputs(1760);
    layer2_outputs(3068) <= (layer1_outputs(1175)) and not (layer1_outputs(651));
    layer2_outputs(3069) <= (layer1_outputs(3735)) and not (layer1_outputs(4957));
    layer2_outputs(3070) <= (layer1_outputs(872)) and not (layer1_outputs(229));
    layer2_outputs(3071) <= not(layer1_outputs(3767)) or (layer1_outputs(2067));
    layer2_outputs(3072) <= not(layer1_outputs(2786));
    layer2_outputs(3073) <= layer1_outputs(3074);
    layer2_outputs(3074) <= not((layer1_outputs(2692)) xor (layer1_outputs(526)));
    layer2_outputs(3075) <= not(layer1_outputs(1531)) or (layer1_outputs(2887));
    layer2_outputs(3076) <= (layer1_outputs(2953)) xor (layer1_outputs(1320));
    layer2_outputs(3077) <= (layer1_outputs(2967)) and not (layer1_outputs(4993));
    layer2_outputs(3078) <= (layer1_outputs(2500)) and not (layer1_outputs(973));
    layer2_outputs(3079) <= not(layer1_outputs(126)) or (layer1_outputs(4721));
    layer2_outputs(3080) <= not(layer1_outputs(2277));
    layer2_outputs(3081) <= not(layer1_outputs(3002));
    layer2_outputs(3082) <= not(layer1_outputs(2737));
    layer2_outputs(3083) <= layer1_outputs(5090);
    layer2_outputs(3084) <= not(layer1_outputs(4717));
    layer2_outputs(3085) <= not(layer1_outputs(3786)) or (layer1_outputs(2786));
    layer2_outputs(3086) <= not(layer1_outputs(2393));
    layer2_outputs(3087) <= not(layer1_outputs(414));
    layer2_outputs(3088) <= not(layer1_outputs(623));
    layer2_outputs(3089) <= not(layer1_outputs(2105));
    layer2_outputs(3090) <= not(layer1_outputs(3783));
    layer2_outputs(3091) <= (layer1_outputs(2663)) and not (layer1_outputs(360));
    layer2_outputs(3092) <= not((layer1_outputs(2580)) xor (layer1_outputs(137)));
    layer2_outputs(3093) <= not((layer1_outputs(1805)) or (layer1_outputs(3895)));
    layer2_outputs(3094) <= (layer1_outputs(2375)) and not (layer1_outputs(4104));
    layer2_outputs(3095) <= not((layer1_outputs(4835)) and (layer1_outputs(2579)));
    layer2_outputs(3096) <= (layer1_outputs(1344)) and not (layer1_outputs(2232));
    layer2_outputs(3097) <= not(layer1_outputs(926));
    layer2_outputs(3098) <= layer1_outputs(2333);
    layer2_outputs(3099) <= not((layer1_outputs(724)) xor (layer1_outputs(3157)));
    layer2_outputs(3100) <= not(layer1_outputs(2965)) or (layer1_outputs(740));
    layer2_outputs(3101) <= not(layer1_outputs(2648));
    layer2_outputs(3102) <= not((layer1_outputs(1722)) and (layer1_outputs(5015)));
    layer2_outputs(3103) <= not(layer1_outputs(245)) or (layer1_outputs(2582));
    layer2_outputs(3104) <= not(layer1_outputs(2345));
    layer2_outputs(3105) <= layer1_outputs(4297);
    layer2_outputs(3106) <= (layer1_outputs(4800)) and not (layer1_outputs(1680));
    layer2_outputs(3107) <= not(layer1_outputs(4244));
    layer2_outputs(3108) <= layer1_outputs(1789);
    layer2_outputs(3109) <= layer1_outputs(983);
    layer2_outputs(3110) <= (layer1_outputs(3594)) or (layer1_outputs(1491));
    layer2_outputs(3111) <= (layer1_outputs(2915)) xor (layer1_outputs(1685));
    layer2_outputs(3112) <= not((layer1_outputs(4964)) or (layer1_outputs(72)));
    layer2_outputs(3113) <= not(layer1_outputs(3551)) or (layer1_outputs(2038));
    layer2_outputs(3114) <= not((layer1_outputs(4855)) and (layer1_outputs(4262)));
    layer2_outputs(3115) <= not(layer1_outputs(4488));
    layer2_outputs(3116) <= not((layer1_outputs(4622)) and (layer1_outputs(3361)));
    layer2_outputs(3117) <= not(layer1_outputs(2928)) or (layer1_outputs(2683));
    layer2_outputs(3118) <= not(layer1_outputs(834));
    layer2_outputs(3119) <= not(layer1_outputs(318)) or (layer1_outputs(2674));
    layer2_outputs(3120) <= (layer1_outputs(3098)) or (layer1_outputs(2305));
    layer2_outputs(3121) <= not(layer1_outputs(1083)) or (layer1_outputs(3185));
    layer2_outputs(3122) <= not(layer1_outputs(1502));
    layer2_outputs(3123) <= layer1_outputs(2968);
    layer2_outputs(3124) <= not(layer1_outputs(3020));
    layer2_outputs(3125) <= not(layer1_outputs(268));
    layer2_outputs(3126) <= not((layer1_outputs(3236)) and (layer1_outputs(87)));
    layer2_outputs(3127) <= layer1_outputs(4856);
    layer2_outputs(3128) <= layer1_outputs(5069);
    layer2_outputs(3129) <= not((layer1_outputs(3289)) or (layer1_outputs(1903)));
    layer2_outputs(3130) <= not(layer1_outputs(200));
    layer2_outputs(3131) <= not(layer1_outputs(4141));
    layer2_outputs(3132) <= not(layer1_outputs(3304)) or (layer1_outputs(169));
    layer2_outputs(3133) <= not(layer1_outputs(4156));
    layer2_outputs(3134) <= not(layer1_outputs(4826)) or (layer1_outputs(3066));
    layer2_outputs(3135) <= not(layer1_outputs(3418));
    layer2_outputs(3136) <= not(layer1_outputs(1512));
    layer2_outputs(3137) <= not(layer1_outputs(283));
    layer2_outputs(3138) <= (layer1_outputs(3728)) xor (layer1_outputs(1144));
    layer2_outputs(3139) <= not(layer1_outputs(3121));
    layer2_outputs(3140) <= not((layer1_outputs(721)) and (layer1_outputs(1525)));
    layer2_outputs(3141) <= (layer1_outputs(630)) and not (layer1_outputs(4998));
    layer2_outputs(3142) <= (layer1_outputs(4815)) and not (layer1_outputs(2098));
    layer2_outputs(3143) <= not(layer1_outputs(3951));
    layer2_outputs(3144) <= not((layer1_outputs(3584)) and (layer1_outputs(4032)));
    layer2_outputs(3145) <= not((layer1_outputs(4119)) and (layer1_outputs(3943)));
    layer2_outputs(3146) <= layer1_outputs(5058);
    layer2_outputs(3147) <= not(layer1_outputs(1132)) or (layer1_outputs(2254));
    layer2_outputs(3148) <= not((layer1_outputs(55)) xor (layer1_outputs(4443)));
    layer2_outputs(3149) <= (layer1_outputs(3526)) and (layer1_outputs(4111));
    layer2_outputs(3150) <= not((layer1_outputs(906)) and (layer1_outputs(4718)));
    layer2_outputs(3151) <= (layer1_outputs(2631)) and not (layer1_outputs(737));
    layer2_outputs(3152) <= layer1_outputs(2174);
    layer2_outputs(3153) <= (layer1_outputs(3092)) or (layer1_outputs(3092));
    layer2_outputs(3154) <= not(layer1_outputs(3285)) or (layer1_outputs(1684));
    layer2_outputs(3155) <= not(layer1_outputs(210)) or (layer1_outputs(3931));
    layer2_outputs(3156) <= (layer1_outputs(2342)) and (layer1_outputs(4245));
    layer2_outputs(3157) <= not(layer1_outputs(3369));
    layer2_outputs(3158) <= not(layer1_outputs(1748));
    layer2_outputs(3159) <= not(layer1_outputs(3370));
    layer2_outputs(3160) <= not((layer1_outputs(1597)) xor (layer1_outputs(462)));
    layer2_outputs(3161) <= not(layer1_outputs(543));
    layer2_outputs(3162) <= (layer1_outputs(4151)) and not (layer1_outputs(2420));
    layer2_outputs(3163) <= not(layer1_outputs(247)) or (layer1_outputs(2545));
    layer2_outputs(3164) <= layer1_outputs(215);
    layer2_outputs(3165) <= (layer1_outputs(431)) or (layer1_outputs(363));
    layer2_outputs(3166) <= not((layer1_outputs(346)) or (layer1_outputs(2250)));
    layer2_outputs(3167) <= not(layer1_outputs(10)) or (layer1_outputs(266));
    layer2_outputs(3168) <= not(layer1_outputs(1479));
    layer2_outputs(3169) <= (layer1_outputs(4336)) and not (layer1_outputs(4448));
    layer2_outputs(3170) <= (layer1_outputs(4182)) and (layer1_outputs(1225));
    layer2_outputs(3171) <= not(layer1_outputs(3582));
    layer2_outputs(3172) <= not((layer1_outputs(568)) or (layer1_outputs(3158)));
    layer2_outputs(3173) <= layer1_outputs(1840);
    layer2_outputs(3174) <= not(layer1_outputs(212));
    layer2_outputs(3175) <= not(layer1_outputs(3911));
    layer2_outputs(3176) <= (layer1_outputs(2769)) and (layer1_outputs(1676));
    layer2_outputs(3177) <= not(layer1_outputs(4643));
    layer2_outputs(3178) <= '1';
    layer2_outputs(3179) <= not(layer1_outputs(4957));
    layer2_outputs(3180) <= (layer1_outputs(2358)) and (layer1_outputs(98));
    layer2_outputs(3181) <= not((layer1_outputs(1296)) or (layer1_outputs(1482)));
    layer2_outputs(3182) <= (layer1_outputs(4372)) and (layer1_outputs(4135));
    layer2_outputs(3183) <= layer1_outputs(3117);
    layer2_outputs(3184) <= layer1_outputs(1875);
    layer2_outputs(3185) <= layer1_outputs(4118);
    layer2_outputs(3186) <= not((layer1_outputs(1469)) xor (layer1_outputs(2361)));
    layer2_outputs(3187) <= not(layer1_outputs(2460)) or (layer1_outputs(1775));
    layer2_outputs(3188) <= (layer1_outputs(4540)) or (layer1_outputs(3557));
    layer2_outputs(3189) <= (layer1_outputs(1842)) or (layer1_outputs(3422));
    layer2_outputs(3190) <= (layer1_outputs(1426)) or (layer1_outputs(1194));
    layer2_outputs(3191) <= not((layer1_outputs(4391)) and (layer1_outputs(140)));
    layer2_outputs(3192) <= not(layer1_outputs(2872));
    layer2_outputs(3193) <= layer1_outputs(4662);
    layer2_outputs(3194) <= not(layer1_outputs(270));
    layer2_outputs(3195) <= not(layer1_outputs(3950)) or (layer1_outputs(2559));
    layer2_outputs(3196) <= not(layer1_outputs(3905)) or (layer1_outputs(1927));
    layer2_outputs(3197) <= layer1_outputs(1713);
    layer2_outputs(3198) <= not(layer1_outputs(4272)) or (layer1_outputs(4496));
    layer2_outputs(3199) <= layer1_outputs(1242);
    layer2_outputs(3200) <= layer1_outputs(2430);
    layer2_outputs(3201) <= not(layer1_outputs(2142));
    layer2_outputs(3202) <= layer1_outputs(3408);
    layer2_outputs(3203) <= not((layer1_outputs(3691)) xor (layer1_outputs(642)));
    layer2_outputs(3204) <= (layer1_outputs(2310)) xor (layer1_outputs(2364));
    layer2_outputs(3205) <= not(layer1_outputs(5107));
    layer2_outputs(3206) <= layer1_outputs(1497);
    layer2_outputs(3207) <= layer1_outputs(4938);
    layer2_outputs(3208) <= layer1_outputs(4681);
    layer2_outputs(3209) <= '0';
    layer2_outputs(3210) <= layer1_outputs(4243);
    layer2_outputs(3211) <= (layer1_outputs(1174)) and (layer1_outputs(3518));
    layer2_outputs(3212) <= layer1_outputs(1659);
    layer2_outputs(3213) <= (layer1_outputs(4208)) and not (layer1_outputs(3187));
    layer2_outputs(3214) <= layer1_outputs(1420);
    layer2_outputs(3215) <= layer1_outputs(1227);
    layer2_outputs(3216) <= not((layer1_outputs(4776)) and (layer1_outputs(2377)));
    layer2_outputs(3217) <= (layer1_outputs(422)) xor (layer1_outputs(3083));
    layer2_outputs(3218) <= (layer1_outputs(4211)) and not (layer1_outputs(2503));
    layer2_outputs(3219) <= not(layer1_outputs(1582)) or (layer1_outputs(2070));
    layer2_outputs(3220) <= (layer1_outputs(4641)) and not (layer1_outputs(1858));
    layer2_outputs(3221) <= layer1_outputs(556);
    layer2_outputs(3222) <= not((layer1_outputs(3481)) or (layer1_outputs(3048)));
    layer2_outputs(3223) <= layer1_outputs(2385);
    layer2_outputs(3224) <= not(layer1_outputs(3269)) or (layer1_outputs(4277));
    layer2_outputs(3225) <= (layer1_outputs(3414)) xor (layer1_outputs(4740));
    layer2_outputs(3226) <= layer1_outputs(2043);
    layer2_outputs(3227) <= '1';
    layer2_outputs(3228) <= not(layer1_outputs(4355)) or (layer1_outputs(222));
    layer2_outputs(3229) <= (layer1_outputs(1938)) and not (layer1_outputs(3760));
    layer2_outputs(3230) <= not(layer1_outputs(2033));
    layer2_outputs(3231) <= not(layer1_outputs(5012));
    layer2_outputs(3232) <= not(layer1_outputs(474));
    layer2_outputs(3233) <= (layer1_outputs(1458)) or (layer1_outputs(1378));
    layer2_outputs(3234) <= not(layer1_outputs(256));
    layer2_outputs(3235) <= (layer1_outputs(100)) and not (layer1_outputs(2548));
    layer2_outputs(3236) <= not(layer1_outputs(682));
    layer2_outputs(3237) <= (layer1_outputs(2607)) and not (layer1_outputs(956));
    layer2_outputs(3238) <= not(layer1_outputs(2812));
    layer2_outputs(3239) <= layer1_outputs(4640);
    layer2_outputs(3240) <= (layer1_outputs(3049)) and (layer1_outputs(379));
    layer2_outputs(3241) <= not(layer1_outputs(1728));
    layer2_outputs(3242) <= not((layer1_outputs(4000)) and (layer1_outputs(3235)));
    layer2_outputs(3243) <= not(layer1_outputs(4654));
    layer2_outputs(3244) <= not(layer1_outputs(1285));
    layer2_outputs(3245) <= (layer1_outputs(1521)) or (layer1_outputs(2191));
    layer2_outputs(3246) <= not(layer1_outputs(2269)) or (layer1_outputs(1009));
    layer2_outputs(3247) <= not(layer1_outputs(1864));
    layer2_outputs(3248) <= not(layer1_outputs(2134)) or (layer1_outputs(4038));
    layer2_outputs(3249) <= not(layer1_outputs(2102));
    layer2_outputs(3250) <= not(layer1_outputs(2136));
    layer2_outputs(3251) <= '1';
    layer2_outputs(3252) <= layer1_outputs(332);
    layer2_outputs(3253) <= layer1_outputs(4134);
    layer2_outputs(3254) <= not(layer1_outputs(4518));
    layer2_outputs(3255) <= not(layer1_outputs(1771));
    layer2_outputs(3256) <= (layer1_outputs(903)) and (layer1_outputs(1624));
    layer2_outputs(3257) <= layer1_outputs(1206);
    layer2_outputs(3258) <= layer1_outputs(4142);
    layer2_outputs(3259) <= not(layer1_outputs(129)) or (layer1_outputs(2684));
    layer2_outputs(3260) <= layer1_outputs(2273);
    layer2_outputs(3261) <= not((layer1_outputs(865)) and (layer1_outputs(4522)));
    layer2_outputs(3262) <= (layer1_outputs(1442)) and (layer1_outputs(2698));
    layer2_outputs(3263) <= not(layer1_outputs(2005));
    layer2_outputs(3264) <= not(layer1_outputs(1527)) or (layer1_outputs(3914));
    layer2_outputs(3265) <= not(layer1_outputs(4080));
    layer2_outputs(3266) <= layer1_outputs(472);
    layer2_outputs(3267) <= layer1_outputs(1507);
    layer2_outputs(3268) <= not(layer1_outputs(4472)) or (layer1_outputs(5020));
    layer2_outputs(3269) <= layer1_outputs(4225);
    layer2_outputs(3270) <= layer1_outputs(3854);
    layer2_outputs(3271) <= (layer1_outputs(4387)) and not (layer1_outputs(4738));
    layer2_outputs(3272) <= (layer1_outputs(3349)) and not (layer1_outputs(1779));
    layer2_outputs(3273) <= not(layer1_outputs(1143));
    layer2_outputs(3274) <= layer1_outputs(765);
    layer2_outputs(3275) <= not(layer1_outputs(1578)) or (layer1_outputs(1275));
    layer2_outputs(3276) <= (layer1_outputs(3082)) or (layer1_outputs(1771));
    layer2_outputs(3277) <= layer1_outputs(1334);
    layer2_outputs(3278) <= layer1_outputs(1836);
    layer2_outputs(3279) <= (layer1_outputs(2212)) or (layer1_outputs(1171));
    layer2_outputs(3280) <= layer1_outputs(704);
    layer2_outputs(3281) <= layer1_outputs(4575);
    layer2_outputs(3282) <= (layer1_outputs(1786)) and (layer1_outputs(2874));
    layer2_outputs(3283) <= not(layer1_outputs(4310));
    layer2_outputs(3284) <= (layer1_outputs(3385)) and (layer1_outputs(1290));
    layer2_outputs(3285) <= not(layer1_outputs(2353));
    layer2_outputs(3286) <= layer1_outputs(5114);
    layer2_outputs(3287) <= not(layer1_outputs(3609));
    layer2_outputs(3288) <= not(layer1_outputs(969)) or (layer1_outputs(853));
    layer2_outputs(3289) <= not(layer1_outputs(2415));
    layer2_outputs(3290) <= not((layer1_outputs(3886)) xor (layer1_outputs(4611)));
    layer2_outputs(3291) <= layer1_outputs(4889);
    layer2_outputs(3292) <= not(layer1_outputs(2250));
    layer2_outputs(3293) <= (layer1_outputs(389)) and not (layer1_outputs(5043));
    layer2_outputs(3294) <= (layer1_outputs(1486)) and (layer1_outputs(1453));
    layer2_outputs(3295) <= not(layer1_outputs(2355));
    layer2_outputs(3296) <= (layer1_outputs(1761)) and (layer1_outputs(1923));
    layer2_outputs(3297) <= not((layer1_outputs(4070)) and (layer1_outputs(3318)));
    layer2_outputs(3298) <= not(layer1_outputs(2097));
    layer2_outputs(3299) <= layer1_outputs(4085);
    layer2_outputs(3300) <= not(layer1_outputs(2977));
    layer2_outputs(3301) <= not((layer1_outputs(3928)) or (layer1_outputs(3327)));
    layer2_outputs(3302) <= layer1_outputs(703);
    layer2_outputs(3303) <= not(layer1_outputs(3590)) or (layer1_outputs(4451));
    layer2_outputs(3304) <= not(layer1_outputs(4744));
    layer2_outputs(3305) <= not(layer1_outputs(4712));
    layer2_outputs(3306) <= layer1_outputs(2780);
    layer2_outputs(3307) <= not(layer1_outputs(2551)) or (layer1_outputs(205));
    layer2_outputs(3308) <= not(layer1_outputs(340));
    layer2_outputs(3309) <= (layer1_outputs(2997)) and not (layer1_outputs(4931));
    layer2_outputs(3310) <= not(layer1_outputs(2710)) or (layer1_outputs(4581));
    layer2_outputs(3311) <= not(layer1_outputs(1268));
    layer2_outputs(3312) <= not(layer1_outputs(1044));
    layer2_outputs(3313) <= (layer1_outputs(3703)) or (layer1_outputs(343));
    layer2_outputs(3314) <= not(layer1_outputs(1709));
    layer2_outputs(3315) <= not(layer1_outputs(1351));
    layer2_outputs(3316) <= (layer1_outputs(3124)) and (layer1_outputs(2811));
    layer2_outputs(3317) <= (layer1_outputs(3176)) and (layer1_outputs(289));
    layer2_outputs(3318) <= not(layer1_outputs(4963));
    layer2_outputs(3319) <= (layer1_outputs(1910)) and not (layer1_outputs(1112));
    layer2_outputs(3320) <= layer1_outputs(399);
    layer2_outputs(3321) <= layer1_outputs(156);
    layer2_outputs(3322) <= not(layer1_outputs(2767)) or (layer1_outputs(1452));
    layer2_outputs(3323) <= not((layer1_outputs(4701)) or (layer1_outputs(4268)));
    layer2_outputs(3324) <= layer1_outputs(3572);
    layer2_outputs(3325) <= layer1_outputs(3408);
    layer2_outputs(3326) <= (layer1_outputs(2153)) and not (layer1_outputs(2178));
    layer2_outputs(3327) <= layer1_outputs(2713);
    layer2_outputs(3328) <= not(layer1_outputs(3089)) or (layer1_outputs(4233));
    layer2_outputs(3329) <= not((layer1_outputs(4709)) and (layer1_outputs(549)));
    layer2_outputs(3330) <= not((layer1_outputs(997)) or (layer1_outputs(345)));
    layer2_outputs(3331) <= (layer1_outputs(4607)) and (layer1_outputs(4613));
    layer2_outputs(3332) <= (layer1_outputs(4441)) and not (layer1_outputs(869));
    layer2_outputs(3333) <= (layer1_outputs(4682)) and not (layer1_outputs(1087));
    layer2_outputs(3334) <= not(layer1_outputs(2209));
    layer2_outputs(3335) <= not(layer1_outputs(394)) or (layer1_outputs(3065));
    layer2_outputs(3336) <= layer1_outputs(2376);
    layer2_outputs(3337) <= not((layer1_outputs(2116)) or (layer1_outputs(376)));
    layer2_outputs(3338) <= not(layer1_outputs(753));
    layer2_outputs(3339) <= layer1_outputs(494);
    layer2_outputs(3340) <= layer1_outputs(4352);
    layer2_outputs(3341) <= not(layer1_outputs(3741)) or (layer1_outputs(338));
    layer2_outputs(3342) <= (layer1_outputs(1762)) or (layer1_outputs(899));
    layer2_outputs(3343) <= not(layer1_outputs(4423)) or (layer1_outputs(555));
    layer2_outputs(3344) <= not(layer1_outputs(1654));
    layer2_outputs(3345) <= layer1_outputs(4782);
    layer2_outputs(3346) <= (layer1_outputs(1483)) and (layer1_outputs(1377));
    layer2_outputs(3347) <= not((layer1_outputs(3193)) or (layer1_outputs(4916)));
    layer2_outputs(3348) <= layer1_outputs(3492);
    layer2_outputs(3349) <= layer1_outputs(3555);
    layer2_outputs(3350) <= not(layer1_outputs(1504)) or (layer1_outputs(811));
    layer2_outputs(3351) <= not((layer1_outputs(530)) and (layer1_outputs(2054)));
    layer2_outputs(3352) <= not(layer1_outputs(2446));
    layer2_outputs(3353) <= not(layer1_outputs(2741));
    layer2_outputs(3354) <= (layer1_outputs(1436)) and not (layer1_outputs(3627));
    layer2_outputs(3355) <= not(layer1_outputs(711));
    layer2_outputs(3356) <= not(layer1_outputs(817));
    layer2_outputs(3357) <= not((layer1_outputs(152)) and (layer1_outputs(3973)));
    layer2_outputs(3358) <= not((layer1_outputs(3661)) or (layer1_outputs(4992)));
    layer2_outputs(3359) <= (layer1_outputs(1820)) and (layer1_outputs(2530));
    layer2_outputs(3360) <= layer1_outputs(4311);
    layer2_outputs(3361) <= not(layer1_outputs(2029));
    layer2_outputs(3362) <= (layer1_outputs(79)) and not (layer1_outputs(708));
    layer2_outputs(3363) <= not((layer1_outputs(1066)) xor (layer1_outputs(198)));
    layer2_outputs(3364) <= layer1_outputs(4712);
    layer2_outputs(3365) <= '1';
    layer2_outputs(3366) <= layer1_outputs(791);
    layer2_outputs(3367) <= (layer1_outputs(1909)) and not (layer1_outputs(2074));
    layer2_outputs(3368) <= layer1_outputs(390);
    layer2_outputs(3369) <= not(layer1_outputs(910));
    layer2_outputs(3370) <= not((layer1_outputs(786)) or (layer1_outputs(1155)));
    layer2_outputs(3371) <= (layer1_outputs(3638)) and (layer1_outputs(4906));
    layer2_outputs(3372) <= not(layer1_outputs(2012));
    layer2_outputs(3373) <= not(layer1_outputs(2644));
    layer2_outputs(3374) <= layer1_outputs(2538);
    layer2_outputs(3375) <= not(layer1_outputs(4536));
    layer2_outputs(3376) <= not(layer1_outputs(4226)) or (layer1_outputs(2909));
    layer2_outputs(3377) <= not(layer1_outputs(4909));
    layer2_outputs(3378) <= not(layer1_outputs(878));
    layer2_outputs(3379) <= not(layer1_outputs(73));
    layer2_outputs(3380) <= layer1_outputs(5053);
    layer2_outputs(3381) <= not((layer1_outputs(2673)) or (layer1_outputs(615)));
    layer2_outputs(3382) <= not((layer1_outputs(239)) xor (layer1_outputs(2455)));
    layer2_outputs(3383) <= '1';
    layer2_outputs(3384) <= not(layer1_outputs(1014)) or (layer1_outputs(2797));
    layer2_outputs(3385) <= not((layer1_outputs(1714)) or (layer1_outputs(1097)));
    layer2_outputs(3386) <= not((layer1_outputs(3928)) or (layer1_outputs(3730)));
    layer2_outputs(3387) <= (layer1_outputs(1558)) xor (layer1_outputs(498));
    layer2_outputs(3388) <= not((layer1_outputs(1759)) or (layer1_outputs(4644)));
    layer2_outputs(3389) <= not(layer1_outputs(3411));
    layer2_outputs(3390) <= not(layer1_outputs(1417));
    layer2_outputs(3391) <= not((layer1_outputs(1317)) xor (layer1_outputs(2612)));
    layer2_outputs(3392) <= (layer1_outputs(3313)) or (layer1_outputs(1359));
    layer2_outputs(3393) <= not(layer1_outputs(777));
    layer2_outputs(3394) <= (layer1_outputs(270)) or (layer1_outputs(2050));
    layer2_outputs(3395) <= layer1_outputs(1695);
    layer2_outputs(3396) <= not(layer1_outputs(1522));
    layer2_outputs(3397) <= not(layer1_outputs(2214)) or (layer1_outputs(4231));
    layer2_outputs(3398) <= not(layer1_outputs(2985));
    layer2_outputs(3399) <= not(layer1_outputs(353));
    layer2_outputs(3400) <= layer1_outputs(4342);
    layer2_outputs(3401) <= (layer1_outputs(4261)) and (layer1_outputs(1470));
    layer2_outputs(3402) <= '0';
    layer2_outputs(3403) <= not(layer1_outputs(3514)) or (layer1_outputs(2538));
    layer2_outputs(3404) <= not(layer1_outputs(3684));
    layer2_outputs(3405) <= not((layer1_outputs(952)) or (layer1_outputs(321)));
    layer2_outputs(3406) <= (layer1_outputs(3600)) xor (layer1_outputs(4425));
    layer2_outputs(3407) <= not((layer1_outputs(2239)) xor (layer1_outputs(3465)));
    layer2_outputs(3408) <= (layer1_outputs(3072)) and (layer1_outputs(4598));
    layer2_outputs(3409) <= not((layer1_outputs(3821)) and (layer1_outputs(3280)));
    layer2_outputs(3410) <= not(layer1_outputs(1731));
    layer2_outputs(3411) <= (layer1_outputs(128)) and not (layer1_outputs(620));
    layer2_outputs(3412) <= not(layer1_outputs(3541));
    layer2_outputs(3413) <= (layer1_outputs(2267)) and not (layer1_outputs(2642));
    layer2_outputs(3414) <= not(layer1_outputs(3028));
    layer2_outputs(3415) <= not(layer1_outputs(1630));
    layer2_outputs(3416) <= not(layer1_outputs(4468)) or (layer1_outputs(2166));
    layer2_outputs(3417) <= layer1_outputs(2404);
    layer2_outputs(3418) <= layer1_outputs(5082);
    layer2_outputs(3419) <= not(layer1_outputs(4795)) or (layer1_outputs(882));
    layer2_outputs(3420) <= layer1_outputs(1788);
    layer2_outputs(3421) <= (layer1_outputs(3124)) xor (layer1_outputs(4716));
    layer2_outputs(3422) <= not(layer1_outputs(3501));
    layer2_outputs(3423) <= layer1_outputs(2191);
    layer2_outputs(3424) <= layer1_outputs(617);
    layer2_outputs(3425) <= (layer1_outputs(4075)) or (layer1_outputs(4105));
    layer2_outputs(3426) <= layer1_outputs(4761);
    layer2_outputs(3427) <= not(layer1_outputs(2875));
    layer2_outputs(3428) <= layer1_outputs(2986);
    layer2_outputs(3429) <= not(layer1_outputs(4154)) or (layer1_outputs(1303));
    layer2_outputs(3430) <= not(layer1_outputs(2667)) or (layer1_outputs(1600));
    layer2_outputs(3431) <= not(layer1_outputs(4708));
    layer2_outputs(3432) <= not(layer1_outputs(2397));
    layer2_outputs(3433) <= not(layer1_outputs(3654)) or (layer1_outputs(52));
    layer2_outputs(3434) <= not((layer1_outputs(2746)) or (layer1_outputs(4353)));
    layer2_outputs(3435) <= layer1_outputs(4969);
    layer2_outputs(3436) <= (layer1_outputs(2475)) and not (layer1_outputs(1740));
    layer2_outputs(3437) <= not((layer1_outputs(2743)) and (layer1_outputs(911)));
    layer2_outputs(3438) <= layer1_outputs(3146);
    layer2_outputs(3439) <= (layer1_outputs(424)) xor (layer1_outputs(1548));
    layer2_outputs(3440) <= not(layer1_outputs(2322));
    layer2_outputs(3441) <= not(layer1_outputs(4482));
    layer2_outputs(3442) <= not(layer1_outputs(1703)) or (layer1_outputs(3892));
    layer2_outputs(3443) <= layer1_outputs(457);
    layer2_outputs(3444) <= not((layer1_outputs(4198)) and (layer1_outputs(2796)));
    layer2_outputs(3445) <= not(layer1_outputs(738)) or (layer1_outputs(909));
    layer2_outputs(3446) <= not(layer1_outputs(4702));
    layer2_outputs(3447) <= not(layer1_outputs(1796));
    layer2_outputs(3448) <= (layer1_outputs(4653)) and (layer1_outputs(4509));
    layer2_outputs(3449) <= not(layer1_outputs(4040));
    layer2_outputs(3450) <= not(layer1_outputs(3205));
    layer2_outputs(3451) <= (layer1_outputs(2073)) and (layer1_outputs(2552));
    layer2_outputs(3452) <= layer1_outputs(4718);
    layer2_outputs(3453) <= not(layer1_outputs(1876));
    layer2_outputs(3454) <= not((layer1_outputs(1847)) xor (layer1_outputs(1747)));
    layer2_outputs(3455) <= (layer1_outputs(3134)) and not (layer1_outputs(3589));
    layer2_outputs(3456) <= not(layer1_outputs(3848));
    layer2_outputs(3457) <= not(layer1_outputs(35));
    layer2_outputs(3458) <= not(layer1_outputs(398));
    layer2_outputs(3459) <= not((layer1_outputs(1781)) and (layer1_outputs(1810)));
    layer2_outputs(3460) <= layer1_outputs(227);
    layer2_outputs(3461) <= not(layer1_outputs(4290));
    layer2_outputs(3462) <= layer1_outputs(503);
    layer2_outputs(3463) <= not(layer1_outputs(2925));
    layer2_outputs(3464) <= not(layer1_outputs(1441)) or (layer1_outputs(883));
    layer2_outputs(3465) <= not((layer1_outputs(558)) and (layer1_outputs(3768)));
    layer2_outputs(3466) <= layer1_outputs(348);
    layer2_outputs(3467) <= not(layer1_outputs(2853));
    layer2_outputs(3468) <= not(layer1_outputs(243));
    layer2_outputs(3469) <= not(layer1_outputs(4584));
    layer2_outputs(3470) <= layer1_outputs(3342);
    layer2_outputs(3471) <= not((layer1_outputs(3522)) xor (layer1_outputs(854)));
    layer2_outputs(3472) <= (layer1_outputs(515)) xor (layer1_outputs(5065));
    layer2_outputs(3473) <= (layer1_outputs(2770)) and not (layer1_outputs(2717));
    layer2_outputs(3474) <= not(layer1_outputs(4285));
    layer2_outputs(3475) <= not(layer1_outputs(2937)) or (layer1_outputs(2282));
    layer2_outputs(3476) <= (layer1_outputs(917)) and (layer1_outputs(4899));
    layer2_outputs(3477) <= not(layer1_outputs(3221));
    layer2_outputs(3478) <= layer1_outputs(4583);
    layer2_outputs(3479) <= (layer1_outputs(325)) and not (layer1_outputs(983));
    layer2_outputs(3480) <= (layer1_outputs(5101)) xor (layer1_outputs(3449));
    layer2_outputs(3481) <= layer1_outputs(2454);
    layer2_outputs(3482) <= layer1_outputs(2154);
    layer2_outputs(3483) <= (layer1_outputs(387)) or (layer1_outputs(4447));
    layer2_outputs(3484) <= layer1_outputs(5088);
    layer2_outputs(3485) <= (layer1_outputs(541)) xor (layer1_outputs(1022));
    layer2_outputs(3486) <= (layer1_outputs(2808)) and (layer1_outputs(4774));
    layer2_outputs(3487) <= '1';
    layer2_outputs(3488) <= (layer1_outputs(1458)) and not (layer1_outputs(615));
    layer2_outputs(3489) <= not(layer1_outputs(4731));
    layer2_outputs(3490) <= layer1_outputs(3893);
    layer2_outputs(3491) <= layer1_outputs(4318);
    layer2_outputs(3492) <= not((layer1_outputs(3242)) and (layer1_outputs(4306)));
    layer2_outputs(3493) <= not(layer1_outputs(3690));
    layer2_outputs(3494) <= (layer1_outputs(851)) and (layer1_outputs(734));
    layer2_outputs(3495) <= not(layer1_outputs(51));
    layer2_outputs(3496) <= (layer1_outputs(250)) or (layer1_outputs(2083));
    layer2_outputs(3497) <= layer1_outputs(277);
    layer2_outputs(3498) <= not(layer1_outputs(4562));
    layer2_outputs(3499) <= not((layer1_outputs(1271)) and (layer1_outputs(362)));
    layer2_outputs(3500) <= not(layer1_outputs(3508)) or (layer1_outputs(1077));
    layer2_outputs(3501) <= layer1_outputs(1541);
    layer2_outputs(3502) <= (layer1_outputs(2517)) or (layer1_outputs(4235));
    layer2_outputs(3503) <= layer1_outputs(4238);
    layer2_outputs(3504) <= not((layer1_outputs(2858)) or (layer1_outputs(2165)));
    layer2_outputs(3505) <= (layer1_outputs(4319)) and (layer1_outputs(402));
    layer2_outputs(3506) <= not(layer1_outputs(2857));
    layer2_outputs(3507) <= not(layer1_outputs(737));
    layer2_outputs(3508) <= not(layer1_outputs(450));
    layer2_outputs(3509) <= not(layer1_outputs(3328));
    layer2_outputs(3510) <= not(layer1_outputs(2386)) or (layer1_outputs(1204));
    layer2_outputs(3511) <= (layer1_outputs(3335)) or (layer1_outputs(4008));
    layer2_outputs(3512) <= not((layer1_outputs(4389)) xor (layer1_outputs(2408)));
    layer2_outputs(3513) <= not(layer1_outputs(1955));
    layer2_outputs(3514) <= not(layer1_outputs(2049)) or (layer1_outputs(3907));
    layer2_outputs(3515) <= (layer1_outputs(5053)) and not (layer1_outputs(184));
    layer2_outputs(3516) <= (layer1_outputs(3250)) and (layer1_outputs(1015));
    layer2_outputs(3517) <= (layer1_outputs(1490)) and not (layer1_outputs(1123));
    layer2_outputs(3518) <= not(layer1_outputs(677)) or (layer1_outputs(3049));
    layer2_outputs(3519) <= not(layer1_outputs(787));
    layer2_outputs(3520) <= layer1_outputs(1248);
    layer2_outputs(3521) <= (layer1_outputs(3168)) xor (layer1_outputs(1936));
    layer2_outputs(3522) <= not(layer1_outputs(4270));
    layer2_outputs(3523) <= (layer1_outputs(459)) xor (layer1_outputs(111));
    layer2_outputs(3524) <= not(layer1_outputs(1393));
    layer2_outputs(3525) <= not(layer1_outputs(57));
    layer2_outputs(3526) <= (layer1_outputs(1987)) or (layer1_outputs(2069));
    layer2_outputs(3527) <= not(layer1_outputs(3722)) or (layer1_outputs(4560));
    layer2_outputs(3528) <= not(layer1_outputs(4951)) or (layer1_outputs(712));
    layer2_outputs(3529) <= not(layer1_outputs(2270));
    layer2_outputs(3530) <= '1';
    layer2_outputs(3531) <= not((layer1_outputs(2617)) xor (layer1_outputs(1161)));
    layer2_outputs(3532) <= not(layer1_outputs(3992));
    layer2_outputs(3533) <= not(layer1_outputs(954));
    layer2_outputs(3534) <= not(layer1_outputs(4937)) or (layer1_outputs(1811));
    layer2_outputs(3535) <= not((layer1_outputs(1730)) xor (layer1_outputs(3094)));
    layer2_outputs(3536) <= layer1_outputs(3101);
    layer2_outputs(3537) <= not(layer1_outputs(3819));
    layer2_outputs(3538) <= (layer1_outputs(3355)) and not (layer1_outputs(1234));
    layer2_outputs(3539) <= not(layer1_outputs(690));
    layer2_outputs(3540) <= layer1_outputs(475);
    layer2_outputs(3541) <= layer1_outputs(2372);
    layer2_outputs(3542) <= not(layer1_outputs(1105));
    layer2_outputs(3543) <= not(layer1_outputs(1794));
    layer2_outputs(3544) <= (layer1_outputs(3061)) and (layer1_outputs(2255));
    layer2_outputs(3545) <= not(layer1_outputs(3404));
    layer2_outputs(3546) <= not((layer1_outputs(1280)) and (layer1_outputs(5086)));
    layer2_outputs(3547) <= not(layer1_outputs(3626));
    layer2_outputs(3548) <= (layer1_outputs(1266)) xor (layer1_outputs(3490));
    layer2_outputs(3549) <= (layer1_outputs(1089)) or (layer1_outputs(3598));
    layer2_outputs(3550) <= layer1_outputs(3300);
    layer2_outputs(3551) <= not((layer1_outputs(881)) or (layer1_outputs(2357)));
    layer2_outputs(3552) <= not(layer1_outputs(1752)) or (layer1_outputs(509));
    layer2_outputs(3553) <= layer1_outputs(1290);
    layer2_outputs(3554) <= layer1_outputs(118);
    layer2_outputs(3555) <= (layer1_outputs(1261)) and not (layer1_outputs(4816));
    layer2_outputs(3556) <= (layer1_outputs(1167)) or (layer1_outputs(4878));
    layer2_outputs(3557) <= (layer1_outputs(2450)) xor (layer1_outputs(88));
    layer2_outputs(3558) <= not(layer1_outputs(2145));
    layer2_outputs(3559) <= not((layer1_outputs(822)) and (layer1_outputs(585)));
    layer2_outputs(3560) <= layer1_outputs(4403);
    layer2_outputs(3561) <= layer1_outputs(1522);
    layer2_outputs(3562) <= (layer1_outputs(3344)) or (layer1_outputs(1010));
    layer2_outputs(3563) <= layer1_outputs(3477);
    layer2_outputs(3564) <= (layer1_outputs(2563)) and (layer1_outputs(4275));
    layer2_outputs(3565) <= layer1_outputs(1179);
    layer2_outputs(3566) <= not((layer1_outputs(4188)) and (layer1_outputs(212)));
    layer2_outputs(3567) <= not(layer1_outputs(4682));
    layer2_outputs(3568) <= not(layer1_outputs(2606));
    layer2_outputs(3569) <= not(layer1_outputs(2031));
    layer2_outputs(3570) <= layer1_outputs(4407);
    layer2_outputs(3571) <= not(layer1_outputs(1088));
    layer2_outputs(3572) <= (layer1_outputs(4573)) and not (layer1_outputs(789));
    layer2_outputs(3573) <= layer1_outputs(4461);
    layer2_outputs(3574) <= not(layer1_outputs(4604)) or (layer1_outputs(4640));
    layer2_outputs(3575) <= (layer1_outputs(1103)) and not (layer1_outputs(4462));
    layer2_outputs(3576) <= not((layer1_outputs(1322)) and (layer1_outputs(1440)));
    layer2_outputs(3577) <= (layer1_outputs(4075)) or (layer1_outputs(784));
    layer2_outputs(3578) <= (layer1_outputs(4548)) and (layer1_outputs(1635));
    layer2_outputs(3579) <= layer1_outputs(3208);
    layer2_outputs(3580) <= (layer1_outputs(741)) and not (layer1_outputs(5034));
    layer2_outputs(3581) <= '1';
    layer2_outputs(3582) <= (layer1_outputs(1871)) or (layer1_outputs(1563));
    layer2_outputs(3583) <= not(layer1_outputs(4096));
    layer2_outputs(3584) <= not(layer1_outputs(3118)) or (layer1_outputs(3317));
    layer2_outputs(3585) <= not((layer1_outputs(590)) or (layer1_outputs(1708)));
    layer2_outputs(3586) <= not(layer1_outputs(5061)) or (layer1_outputs(336));
    layer2_outputs(3587) <= (layer1_outputs(439)) and not (layer1_outputs(1566));
    layer2_outputs(3588) <= not(layer1_outputs(2048));
    layer2_outputs(3589) <= (layer1_outputs(15)) or (layer1_outputs(354));
    layer2_outputs(3590) <= not(layer1_outputs(4946));
    layer2_outputs(3591) <= (layer1_outputs(4175)) or (layer1_outputs(2563));
    layer2_outputs(3592) <= not(layer1_outputs(3568));
    layer2_outputs(3593) <= not(layer1_outputs(383)) or (layer1_outputs(280));
    layer2_outputs(3594) <= not((layer1_outputs(4986)) or (layer1_outputs(206)));
    layer2_outputs(3595) <= (layer1_outputs(914)) or (layer1_outputs(1043));
    layer2_outputs(3596) <= not(layer1_outputs(3025));
    layer2_outputs(3597) <= not(layer1_outputs(2764));
    layer2_outputs(3598) <= not(layer1_outputs(863));
    layer2_outputs(3599) <= layer1_outputs(702);
    layer2_outputs(3600) <= not((layer1_outputs(4054)) or (layer1_outputs(4093)));
    layer2_outputs(3601) <= not((layer1_outputs(2607)) and (layer1_outputs(3857)));
    layer2_outputs(3602) <= not((layer1_outputs(822)) and (layer1_outputs(4883)));
    layer2_outputs(3603) <= not(layer1_outputs(888));
    layer2_outputs(3604) <= '0';
    layer2_outputs(3605) <= '0';
    layer2_outputs(3606) <= '0';
    layer2_outputs(3607) <= not(layer1_outputs(4225)) or (layer1_outputs(369));
    layer2_outputs(3608) <= (layer1_outputs(4772)) xor (layer1_outputs(4351));
    layer2_outputs(3609) <= (layer1_outputs(5039)) and not (layer1_outputs(1618));
    layer2_outputs(3610) <= (layer1_outputs(4386)) or (layer1_outputs(2130));
    layer2_outputs(3611) <= (layer1_outputs(1711)) and not (layer1_outputs(3437));
    layer2_outputs(3612) <= not((layer1_outputs(3039)) xor (layer1_outputs(799)));
    layer2_outputs(3613) <= '1';
    layer2_outputs(3614) <= layer1_outputs(3672);
    layer2_outputs(3615) <= layer1_outputs(4175);
    layer2_outputs(3616) <= not((layer1_outputs(4259)) or (layer1_outputs(3440)));
    layer2_outputs(3617) <= not(layer1_outputs(1926));
    layer2_outputs(3618) <= not(layer1_outputs(1655));
    layer2_outputs(3619) <= not(layer1_outputs(1225)) or (layer1_outputs(3915));
    layer2_outputs(3620) <= not((layer1_outputs(1544)) xor (layer1_outputs(4137)));
    layer2_outputs(3621) <= (layer1_outputs(590)) or (layer1_outputs(510));
    layer2_outputs(3622) <= layer1_outputs(1314);
    layer2_outputs(3623) <= (layer1_outputs(2558)) and not (layer1_outputs(284));
    layer2_outputs(3624) <= not((layer1_outputs(4548)) or (layer1_outputs(3543)));
    layer2_outputs(3625) <= layer1_outputs(3269);
    layer2_outputs(3626) <= (layer1_outputs(3798)) and not (layer1_outputs(3376));
    layer2_outputs(3627) <= layer1_outputs(276);
    layer2_outputs(3628) <= (layer1_outputs(3516)) and not (layer1_outputs(1694));
    layer2_outputs(3629) <= (layer1_outputs(3357)) and not (layer1_outputs(553));
    layer2_outputs(3630) <= not(layer1_outputs(447));
    layer2_outputs(3631) <= not(layer1_outputs(3590));
    layer2_outputs(3632) <= (layer1_outputs(1292)) or (layer1_outputs(467));
    layer2_outputs(3633) <= layer1_outputs(3031);
    layer2_outputs(3634) <= not(layer1_outputs(3152));
    layer2_outputs(3635) <= layer1_outputs(3088);
    layer2_outputs(3636) <= layer1_outputs(926);
    layer2_outputs(3637) <= (layer1_outputs(3030)) and not (layer1_outputs(3824));
    layer2_outputs(3638) <= not(layer1_outputs(286));
    layer2_outputs(3639) <= layer1_outputs(3150);
    layer2_outputs(3640) <= (layer1_outputs(1457)) and not (layer1_outputs(3698));
    layer2_outputs(3641) <= not((layer1_outputs(3394)) or (layer1_outputs(3285)));
    layer2_outputs(3642) <= not(layer1_outputs(974)) or (layer1_outputs(1533));
    layer2_outputs(3643) <= not(layer1_outputs(524));
    layer2_outputs(3644) <= not(layer1_outputs(4280));
    layer2_outputs(3645) <= layer1_outputs(2658);
    layer2_outputs(3646) <= layer1_outputs(2519);
    layer2_outputs(3647) <= not(layer1_outputs(366));
    layer2_outputs(3648) <= not(layer1_outputs(204));
    layer2_outputs(3649) <= (layer1_outputs(2880)) or (layer1_outputs(328));
    layer2_outputs(3650) <= not(layer1_outputs(1295));
    layer2_outputs(3651) <= not(layer1_outputs(1743));
    layer2_outputs(3652) <= not(layer1_outputs(1059));
    layer2_outputs(3653) <= not(layer1_outputs(1305));
    layer2_outputs(3654) <= '1';
    layer2_outputs(3655) <= layer1_outputs(3970);
    layer2_outputs(3656) <= not((layer1_outputs(2542)) and (layer1_outputs(406)));
    layer2_outputs(3657) <= not(layer1_outputs(1424));
    layer2_outputs(3658) <= '1';
    layer2_outputs(3659) <= not((layer1_outputs(3333)) and (layer1_outputs(1972)));
    layer2_outputs(3660) <= layer1_outputs(391);
    layer2_outputs(3661) <= (layer1_outputs(4051)) and not (layer1_outputs(630));
    layer2_outputs(3662) <= not(layer1_outputs(2073));
    layer2_outputs(3663) <= not((layer1_outputs(893)) and (layer1_outputs(3127)));
    layer2_outputs(3664) <= layer1_outputs(3409);
    layer2_outputs(3665) <= not(layer1_outputs(3863));
    layer2_outputs(3666) <= (layer1_outputs(4600)) and not (layer1_outputs(2495));
    layer2_outputs(3667) <= not((layer1_outputs(782)) or (layer1_outputs(4859)));
    layer2_outputs(3668) <= not(layer1_outputs(168));
    layer2_outputs(3669) <= not(layer1_outputs(2514));
    layer2_outputs(3670) <= not((layer1_outputs(3643)) xor (layer1_outputs(818)));
    layer2_outputs(3671) <= (layer1_outputs(3389)) and not (layer1_outputs(4070));
    layer2_outputs(3672) <= layer1_outputs(660);
    layer2_outputs(3673) <= (layer1_outputs(2661)) and not (layer1_outputs(4707));
    layer2_outputs(3674) <= (layer1_outputs(4960)) xor (layer1_outputs(209));
    layer2_outputs(3675) <= layer1_outputs(3740);
    layer2_outputs(3676) <= not(layer1_outputs(2805));
    layer2_outputs(3677) <= not((layer1_outputs(3876)) and (layer1_outputs(3890)));
    layer2_outputs(3678) <= (layer1_outputs(118)) or (layer1_outputs(2991));
    layer2_outputs(3679) <= not(layer1_outputs(1882));
    layer2_outputs(3680) <= layer1_outputs(4181);
    layer2_outputs(3681) <= not(layer1_outputs(4279));
    layer2_outputs(3682) <= not(layer1_outputs(858));
    layer2_outputs(3683) <= not((layer1_outputs(2100)) or (layer1_outputs(4433)));
    layer2_outputs(3684) <= (layer1_outputs(4485)) and (layer1_outputs(4106));
    layer2_outputs(3685) <= layer1_outputs(1055);
    layer2_outputs(3686) <= layer1_outputs(2431);
    layer2_outputs(3687) <= (layer1_outputs(3621)) or (layer1_outputs(1602));
    layer2_outputs(3688) <= (layer1_outputs(3922)) or (layer1_outputs(560));
    layer2_outputs(3689) <= (layer1_outputs(1957)) and (layer1_outputs(2863));
    layer2_outputs(3690) <= not(layer1_outputs(1455));
    layer2_outputs(3691) <= layer1_outputs(2970);
    layer2_outputs(3692) <= not((layer1_outputs(2574)) and (layer1_outputs(2260)));
    layer2_outputs(3693) <= (layer1_outputs(1461)) xor (layer1_outputs(3840));
    layer2_outputs(3694) <= (layer1_outputs(121)) or (layer1_outputs(1724));
    layer2_outputs(3695) <= layer1_outputs(2908);
    layer2_outputs(3696) <= layer1_outputs(2648);
    layer2_outputs(3697) <= not(layer1_outputs(428));
    layer2_outputs(3698) <= not(layer1_outputs(2244)) or (layer1_outputs(2470));
    layer2_outputs(3699) <= not(layer1_outputs(1394));
    layer2_outputs(3700) <= layer1_outputs(3358);
    layer2_outputs(3701) <= layer1_outputs(435);
    layer2_outputs(3702) <= '1';
    layer2_outputs(3703) <= not(layer1_outputs(2678));
    layer2_outputs(3704) <= not(layer1_outputs(2283));
    layer2_outputs(3705) <= not(layer1_outputs(3994)) or (layer1_outputs(2253));
    layer2_outputs(3706) <= not(layer1_outputs(2616));
    layer2_outputs(3707) <= not(layer1_outputs(682));
    layer2_outputs(3708) <= layer1_outputs(1215);
    layer2_outputs(3709) <= not(layer1_outputs(5097));
    layer2_outputs(3710) <= not(layer1_outputs(2618));
    layer2_outputs(3711) <= not(layer1_outputs(5091)) or (layer1_outputs(2469));
    layer2_outputs(3712) <= layer1_outputs(2425);
    layer2_outputs(3713) <= layer1_outputs(5109);
    layer2_outputs(3714) <= not(layer1_outputs(4980));
    layer2_outputs(3715) <= '0';
    layer2_outputs(3716) <= layer1_outputs(2724);
    layer2_outputs(3717) <= not(layer1_outputs(862));
    layer2_outputs(3718) <= not(layer1_outputs(3340)) or (layer1_outputs(1947));
    layer2_outputs(3719) <= not(layer1_outputs(2940));
    layer2_outputs(3720) <= not(layer1_outputs(4089));
    layer2_outputs(3721) <= (layer1_outputs(4367)) and (layer1_outputs(3623));
    layer2_outputs(3722) <= not(layer1_outputs(1846));
    layer2_outputs(3723) <= not(layer1_outputs(2161));
    layer2_outputs(3724) <= (layer1_outputs(2057)) xor (layer1_outputs(3016));
    layer2_outputs(3725) <= not((layer1_outputs(2742)) and (layer1_outputs(2589)));
    layer2_outputs(3726) <= not(layer1_outputs(2885));
    layer2_outputs(3727) <= layer1_outputs(3379);
    layer2_outputs(3728) <= (layer1_outputs(1284)) and (layer1_outputs(1851));
    layer2_outputs(3729) <= not(layer1_outputs(434)) or (layer1_outputs(4480));
    layer2_outputs(3730) <= (layer1_outputs(2885)) xor (layer1_outputs(3278));
    layer2_outputs(3731) <= not((layer1_outputs(4683)) xor (layer1_outputs(735)));
    layer2_outputs(3732) <= layer1_outputs(1649);
    layer2_outputs(3733) <= not(layer1_outputs(3957));
    layer2_outputs(3734) <= (layer1_outputs(2149)) and not (layer1_outputs(494));
    layer2_outputs(3735) <= (layer1_outputs(2754)) and not (layer1_outputs(235));
    layer2_outputs(3736) <= (layer1_outputs(4039)) and (layer1_outputs(4533));
    layer2_outputs(3737) <= layer1_outputs(1217);
    layer2_outputs(3738) <= layer1_outputs(3038);
    layer2_outputs(3739) <= (layer1_outputs(1819)) and (layer1_outputs(1616));
    layer2_outputs(3740) <= not(layer1_outputs(1135));
    layer2_outputs(3741) <= not(layer1_outputs(3434));
    layer2_outputs(3742) <= not(layer1_outputs(4087));
    layer2_outputs(3743) <= layer1_outputs(4347);
    layer2_outputs(3744) <= not(layer1_outputs(4426));
    layer2_outputs(3745) <= layer1_outputs(3511);
    layer2_outputs(3746) <= (layer1_outputs(1895)) and not (layer1_outputs(2535));
    layer2_outputs(3747) <= (layer1_outputs(3916)) and (layer1_outputs(268));
    layer2_outputs(3748) <= (layer1_outputs(512)) and (layer1_outputs(3217));
    layer2_outputs(3749) <= (layer1_outputs(4390)) or (layer1_outputs(1435));
    layer2_outputs(3750) <= layer1_outputs(2005);
    layer2_outputs(3751) <= layer1_outputs(4450);
    layer2_outputs(3752) <= layer1_outputs(2911);
    layer2_outputs(3753) <= '0';
    layer2_outputs(3754) <= (layer1_outputs(4756)) xor (layer1_outputs(4570));
    layer2_outputs(3755) <= not(layer1_outputs(888));
    layer2_outputs(3756) <= (layer1_outputs(3599)) or (layer1_outputs(4930));
    layer2_outputs(3757) <= (layer1_outputs(2911)) and not (layer1_outputs(2634));
    layer2_outputs(3758) <= not((layer1_outputs(31)) or (layer1_outputs(4093)));
    layer2_outputs(3759) <= not(layer1_outputs(3644));
    layer2_outputs(3760) <= (layer1_outputs(4456)) and not (layer1_outputs(798));
    layer2_outputs(3761) <= layer1_outputs(1248);
    layer2_outputs(3762) <= not(layer1_outputs(4812));
    layer2_outputs(3763) <= (layer1_outputs(3787)) xor (layer1_outputs(1364));
    layer2_outputs(3764) <= not(layer1_outputs(213));
    layer2_outputs(3765) <= not((layer1_outputs(2745)) or (layer1_outputs(4809)));
    layer2_outputs(3766) <= not(layer1_outputs(1072)) or (layer1_outputs(431));
    layer2_outputs(3767) <= layer1_outputs(4845);
    layer2_outputs(3768) <= not((layer1_outputs(4928)) xor (layer1_outputs(1025)));
    layer2_outputs(3769) <= not(layer1_outputs(3327));
    layer2_outputs(3770) <= (layer1_outputs(3664)) and (layer1_outputs(720));
    layer2_outputs(3771) <= layer1_outputs(1160);
    layer2_outputs(3772) <= not(layer1_outputs(375));
    layer2_outputs(3773) <= layer1_outputs(2660);
    layer2_outputs(3774) <= not((layer1_outputs(1588)) and (layer1_outputs(2248)));
    layer2_outputs(3775) <= layer1_outputs(2032);
    layer2_outputs(3776) <= not(layer1_outputs(739));
    layer2_outputs(3777) <= (layer1_outputs(1767)) and not (layer1_outputs(1526));
    layer2_outputs(3778) <= not((layer1_outputs(3175)) and (layer1_outputs(2366)));
    layer2_outputs(3779) <= layer1_outputs(3944);
    layer2_outputs(3780) <= not(layer1_outputs(2929)) or (layer1_outputs(4766));
    layer2_outputs(3781) <= not(layer1_outputs(5050));
    layer2_outputs(3782) <= not(layer1_outputs(3923));
    layer2_outputs(3783) <= layer1_outputs(3816);
    layer2_outputs(3784) <= layer1_outputs(3516);
    layer2_outputs(3785) <= (layer1_outputs(4722)) or (layer1_outputs(2014));
    layer2_outputs(3786) <= layer1_outputs(658);
    layer2_outputs(3787) <= not(layer1_outputs(2207));
    layer2_outputs(3788) <= '0';
    layer2_outputs(3789) <= not(layer1_outputs(1774));
    layer2_outputs(3790) <= (layer1_outputs(1975)) or (layer1_outputs(2119));
    layer2_outputs(3791) <= layer1_outputs(3784);
    layer2_outputs(3792) <= not(layer1_outputs(3560));
    layer2_outputs(3793) <= (layer1_outputs(1221)) or (layer1_outputs(4916));
    layer2_outputs(3794) <= not(layer1_outputs(4667));
    layer2_outputs(3795) <= layer1_outputs(1175);
    layer2_outputs(3796) <= (layer1_outputs(1139)) and (layer1_outputs(3955));
    layer2_outputs(3797) <= not((layer1_outputs(2703)) and (layer1_outputs(4543)));
    layer2_outputs(3798) <= (layer1_outputs(2974)) or (layer1_outputs(2480));
    layer2_outputs(3799) <= layer1_outputs(333);
    layer2_outputs(3800) <= not((layer1_outputs(2415)) and (layer1_outputs(2252)));
    layer2_outputs(3801) <= not(layer1_outputs(4320));
    layer2_outputs(3802) <= not(layer1_outputs(4877));
    layer2_outputs(3803) <= layer1_outputs(2850);
    layer2_outputs(3804) <= not(layer1_outputs(1176));
    layer2_outputs(3805) <= (layer1_outputs(3459)) xor (layer1_outputs(2939));
    layer2_outputs(3806) <= not(layer1_outputs(1121));
    layer2_outputs(3807) <= not(layer1_outputs(910)) or (layer1_outputs(4187));
    layer2_outputs(3808) <= not(layer1_outputs(1150)) or (layer1_outputs(3443));
    layer2_outputs(3809) <= not((layer1_outputs(1204)) and (layer1_outputs(53)));
    layer2_outputs(3810) <= '1';
    layer2_outputs(3811) <= not(layer1_outputs(558));
    layer2_outputs(3812) <= (layer1_outputs(2476)) and (layer1_outputs(3439));
    layer2_outputs(3813) <= (layer1_outputs(312)) or (layer1_outputs(1136));
    layer2_outputs(3814) <= not(layer1_outputs(5040)) or (layer1_outputs(3691));
    layer2_outputs(3815) <= layer1_outputs(4913);
    layer2_outputs(3816) <= not(layer1_outputs(2749));
    layer2_outputs(3817) <= (layer1_outputs(3638)) xor (layer1_outputs(2750));
    layer2_outputs(3818) <= (layer1_outputs(1400)) and (layer1_outputs(4808));
    layer2_outputs(3819) <= (layer1_outputs(2883)) or (layer1_outputs(1133));
    layer2_outputs(3820) <= not(layer1_outputs(3523));
    layer2_outputs(3821) <= '1';
    layer2_outputs(3822) <= '1';
    layer2_outputs(3823) <= layer1_outputs(2582);
    layer2_outputs(3824) <= not(layer1_outputs(3396));
    layer2_outputs(3825) <= not(layer1_outputs(1953)) or (layer1_outputs(2844));
    layer2_outputs(3826) <= layer1_outputs(3658);
    layer2_outputs(3827) <= not(layer1_outputs(4646)) or (layer1_outputs(4078));
    layer2_outputs(3828) <= (layer1_outputs(843)) and (layer1_outputs(149));
    layer2_outputs(3829) <= '0';
    layer2_outputs(3830) <= not(layer1_outputs(2315));
    layer2_outputs(3831) <= not(layer1_outputs(717)) or (layer1_outputs(3483));
    layer2_outputs(3832) <= layer1_outputs(3776);
    layer2_outputs(3833) <= not(layer1_outputs(426));
    layer2_outputs(3834) <= layer1_outputs(1904);
    layer2_outputs(3835) <= layer1_outputs(330);
    layer2_outputs(3836) <= not(layer1_outputs(2226));
    layer2_outputs(3837) <= layer1_outputs(381);
    layer2_outputs(3838) <= layer1_outputs(2559);
    layer2_outputs(3839) <= layer1_outputs(1029);
    layer2_outputs(3840) <= not(layer1_outputs(3394));
    layer2_outputs(3841) <= not(layer1_outputs(919));
    layer2_outputs(3842) <= not((layer1_outputs(5108)) or (layer1_outputs(249)));
    layer2_outputs(3843) <= layer1_outputs(4519);
    layer2_outputs(3844) <= (layer1_outputs(295)) and (layer1_outputs(2627));
    layer2_outputs(3845) <= not(layer1_outputs(1688)) or (layer1_outputs(892));
    layer2_outputs(3846) <= not((layer1_outputs(2260)) or (layer1_outputs(1916)));
    layer2_outputs(3847) <= not(layer1_outputs(3621));
    layer2_outputs(3848) <= (layer1_outputs(372)) and not (layer1_outputs(612));
    layer2_outputs(3849) <= not(layer1_outputs(4349)) or (layer1_outputs(4586));
    layer2_outputs(3850) <= '0';
    layer2_outputs(3851) <= not(layer1_outputs(1223));
    layer2_outputs(3852) <= layer1_outputs(897);
    layer2_outputs(3853) <= not(layer1_outputs(4309));
    layer2_outputs(3854) <= not((layer1_outputs(4922)) and (layer1_outputs(5099)));
    layer2_outputs(3855) <= (layer1_outputs(1118)) xor (layer1_outputs(1727));
    layer2_outputs(3856) <= layer1_outputs(2785);
    layer2_outputs(3857) <= (layer1_outputs(4507)) xor (layer1_outputs(1908));
    layer2_outputs(3858) <= (layer1_outputs(3683)) and not (layer1_outputs(3128));
    layer2_outputs(3859) <= not(layer1_outputs(1254));
    layer2_outputs(3860) <= not(layer1_outputs(4258));
    layer2_outputs(3861) <= layer1_outputs(3877);
    layer2_outputs(3862) <= layer1_outputs(1907);
    layer2_outputs(3863) <= (layer1_outputs(3932)) xor (layer1_outputs(3906));
    layer2_outputs(3864) <= not(layer1_outputs(1468));
    layer2_outputs(3865) <= not(layer1_outputs(3171));
    layer2_outputs(3866) <= not(layer1_outputs(3113)) or (layer1_outputs(86));
    layer2_outputs(3867) <= (layer1_outputs(3810)) and not (layer1_outputs(4487));
    layer2_outputs(3868) <= layer1_outputs(4580);
    layer2_outputs(3869) <= not(layer1_outputs(3659));
    layer2_outputs(3870) <= not((layer1_outputs(3855)) and (layer1_outputs(2182)));
    layer2_outputs(3871) <= layer1_outputs(3218);
    layer2_outputs(3872) <= not(layer1_outputs(3738));
    layer2_outputs(3873) <= layer1_outputs(1276);
    layer2_outputs(3874) <= layer1_outputs(3875);
    layer2_outputs(3875) <= layer1_outputs(1289);
    layer2_outputs(3876) <= not(layer1_outputs(1538));
    layer2_outputs(3877) <= not(layer1_outputs(460));
    layer2_outputs(3878) <= not((layer1_outputs(3952)) xor (layer1_outputs(3624)));
    layer2_outputs(3879) <= not(layer1_outputs(2992));
    layer2_outputs(3880) <= not((layer1_outputs(1998)) or (layer1_outputs(1249)));
    layer2_outputs(3881) <= not(layer1_outputs(1361));
    layer2_outputs(3882) <= layer1_outputs(2862);
    layer2_outputs(3883) <= not(layer1_outputs(625));
    layer2_outputs(3884) <= not(layer1_outputs(1107));
    layer2_outputs(3885) <= (layer1_outputs(3887)) or (layer1_outputs(238));
    layer2_outputs(3886) <= (layer1_outputs(1568)) and (layer1_outputs(3420));
    layer2_outputs(3887) <= not(layer1_outputs(672));
    layer2_outputs(3888) <= not(layer1_outputs(4130)) or (layer1_outputs(984));
    layer2_outputs(3889) <= not((layer1_outputs(553)) and (layer1_outputs(779)));
    layer2_outputs(3890) <= not(layer1_outputs(330));
    layer2_outputs(3891) <= not(layer1_outputs(4914));
    layer2_outputs(3892) <= layer1_outputs(1845);
    layer2_outputs(3893) <= not(layer1_outputs(616));
    layer2_outputs(3894) <= not(layer1_outputs(2671));
    layer2_outputs(3895) <= not(layer1_outputs(1137));
    layer2_outputs(3896) <= layer1_outputs(3353);
    layer2_outputs(3897) <= not((layer1_outputs(611)) xor (layer1_outputs(3973)));
    layer2_outputs(3898) <= not((layer1_outputs(4339)) and (layer1_outputs(2770)));
    layer2_outputs(3899) <= not(layer1_outputs(193));
    layer2_outputs(3900) <= layer1_outputs(5047);
    layer2_outputs(3901) <= layer1_outputs(2004);
    layer2_outputs(3902) <= not((layer1_outputs(162)) xor (layer1_outputs(1646)));
    layer2_outputs(3903) <= not((layer1_outputs(3126)) or (layer1_outputs(731)));
    layer2_outputs(3904) <= (layer1_outputs(2848)) and not (layer1_outputs(3504));
    layer2_outputs(3905) <= not((layer1_outputs(2906)) and (layer1_outputs(3926)));
    layer2_outputs(3906) <= not(layer1_outputs(473));
    layer2_outputs(3907) <= layer1_outputs(3244);
    layer2_outputs(3908) <= not(layer1_outputs(1632));
    layer2_outputs(3909) <= (layer1_outputs(1114)) and not (layer1_outputs(3692));
    layer2_outputs(3910) <= not(layer1_outputs(1487)) or (layer1_outputs(4764));
    layer2_outputs(3911) <= layer1_outputs(1262);
    layer2_outputs(3912) <= not((layer1_outputs(341)) or (layer1_outputs(114)));
    layer2_outputs(3913) <= not(layer1_outputs(2765));
    layer2_outputs(3914) <= (layer1_outputs(1242)) xor (layer1_outputs(3903));
    layer2_outputs(3915) <= not((layer1_outputs(4864)) or (layer1_outputs(2614)));
    layer2_outputs(3916) <= (layer1_outputs(71)) and (layer1_outputs(2113));
    layer2_outputs(3917) <= not(layer1_outputs(967));
    layer2_outputs(3918) <= layer1_outputs(4484);
    layer2_outputs(3919) <= not(layer1_outputs(4221));
    layer2_outputs(3920) <= '1';
    layer2_outputs(3921) <= not((layer1_outputs(4616)) xor (layer1_outputs(4423)));
    layer2_outputs(3922) <= layer1_outputs(1720);
    layer2_outputs(3923) <= layer1_outputs(1062);
    layer2_outputs(3924) <= not(layer1_outputs(3630)) or (layer1_outputs(3840));
    layer2_outputs(3925) <= layer1_outputs(3864);
    layer2_outputs(3926) <= (layer1_outputs(2524)) xor (layer1_outputs(807));
    layer2_outputs(3927) <= layer1_outputs(1274);
    layer2_outputs(3928) <= layer1_outputs(4036);
    layer2_outputs(3929) <= not(layer1_outputs(3956)) or (layer1_outputs(4190));
    layer2_outputs(3930) <= not(layer1_outputs(1364));
    layer2_outputs(3931) <= layer1_outputs(3518);
    layer2_outputs(3932) <= not(layer1_outputs(4503));
    layer2_outputs(3933) <= not(layer1_outputs(2041));
    layer2_outputs(3934) <= layer1_outputs(4929);
    layer2_outputs(3935) <= layer1_outputs(4811);
    layer2_outputs(3936) <= (layer1_outputs(315)) or (layer1_outputs(1669));
    layer2_outputs(3937) <= (layer1_outputs(4979)) and not (layer1_outputs(3723));
    layer2_outputs(3938) <= (layer1_outputs(2455)) and not (layer1_outputs(781));
    layer2_outputs(3939) <= not(layer1_outputs(4305));
    layer2_outputs(3940) <= not(layer1_outputs(1098));
    layer2_outputs(3941) <= layer1_outputs(3828);
    layer2_outputs(3942) <= not(layer1_outputs(1622));
    layer2_outputs(3943) <= not(layer1_outputs(4729));
    layer2_outputs(3944) <= (layer1_outputs(2011)) or (layer1_outputs(396));
    layer2_outputs(3945) <= (layer1_outputs(3231)) and not (layer1_outputs(4932));
    layer2_outputs(3946) <= not((layer1_outputs(1595)) or (layer1_outputs(3888)));
    layer2_outputs(3947) <= not(layer1_outputs(5051));
    layer2_outputs(3948) <= not(layer1_outputs(4234));
    layer2_outputs(3949) <= layer1_outputs(1307);
    layer2_outputs(3950) <= not((layer1_outputs(788)) or (layer1_outputs(2993)));
    layer2_outputs(3951) <= not(layer1_outputs(679)) or (layer1_outputs(1841));
    layer2_outputs(3952) <= not(layer1_outputs(2995));
    layer2_outputs(3953) <= (layer1_outputs(2409)) or (layer1_outputs(1387));
    layer2_outputs(3954) <= (layer1_outputs(4125)) xor (layer1_outputs(4393));
    layer2_outputs(3955) <= layer1_outputs(490);
    layer2_outputs(3956) <= layer1_outputs(2907);
    layer2_outputs(3957) <= (layer1_outputs(1969)) and not (layer1_outputs(1584));
    layer2_outputs(3958) <= (layer1_outputs(3116)) and not (layer1_outputs(916));
    layer2_outputs(3959) <= not(layer1_outputs(1591));
    layer2_outputs(3960) <= (layer1_outputs(2129)) and not (layer1_outputs(2778));
    layer2_outputs(3961) <= not(layer1_outputs(1793));
    layer2_outputs(3962) <= not(layer1_outputs(804));
    layer2_outputs(3963) <= not(layer1_outputs(2373));
    layer2_outputs(3964) <= layer1_outputs(3352);
    layer2_outputs(3965) <= (layer1_outputs(1287)) and not (layer1_outputs(605));
    layer2_outputs(3966) <= not((layer1_outputs(4329)) and (layer1_outputs(2494)));
    layer2_outputs(3967) <= '0';
    layer2_outputs(3968) <= not((layer1_outputs(4077)) xor (layer1_outputs(3823)));
    layer2_outputs(3969) <= not(layer1_outputs(4834));
    layer2_outputs(3970) <= not(layer1_outputs(3181)) or (layer1_outputs(3699));
    layer2_outputs(3971) <= layer1_outputs(4112);
    layer2_outputs(3972) <= not(layer1_outputs(261));
    layer2_outputs(3973) <= (layer1_outputs(1330)) and (layer1_outputs(4371));
    layer2_outputs(3974) <= not(layer1_outputs(1789));
    layer2_outputs(3975) <= layer1_outputs(9);
    layer2_outputs(3976) <= (layer1_outputs(1825)) or (layer1_outputs(5023));
    layer2_outputs(3977) <= not((layer1_outputs(1353)) and (layer1_outputs(2558)));
    layer2_outputs(3978) <= layer1_outputs(1342);
    layer2_outputs(3979) <= not((layer1_outputs(1506)) and (layer1_outputs(2550)));
    layer2_outputs(3980) <= layer1_outputs(4268);
    layer2_outputs(3981) <= not(layer1_outputs(2003));
    layer2_outputs(3982) <= not(layer1_outputs(556)) or (layer1_outputs(2173));
    layer2_outputs(3983) <= layer1_outputs(7);
    layer2_outputs(3984) <= not(layer1_outputs(1317));
    layer2_outputs(3985) <= layer1_outputs(604);
    layer2_outputs(3986) <= not(layer1_outputs(943)) or (layer1_outputs(4558));
    layer2_outputs(3987) <= not(layer1_outputs(4308));
    layer2_outputs(3988) <= not(layer1_outputs(2873));
    layer2_outputs(3989) <= layer1_outputs(2686);
    layer2_outputs(3990) <= layer1_outputs(4831);
    layer2_outputs(3991) <= layer1_outputs(1553);
    layer2_outputs(3992) <= not(layer1_outputs(326)) or (layer1_outputs(1339));
    layer2_outputs(3993) <= (layer1_outputs(3472)) and not (layer1_outputs(3999));
    layer2_outputs(3994) <= not(layer1_outputs(3035));
    layer2_outputs(3995) <= layer1_outputs(3167);
    layer2_outputs(3996) <= not(layer1_outputs(3755));
    layer2_outputs(3997) <= (layer1_outputs(1404)) xor (layer1_outputs(2497));
    layer2_outputs(3998) <= layer1_outputs(1270);
    layer2_outputs(3999) <= not(layer1_outputs(2068));
    layer2_outputs(4000) <= layer1_outputs(4428);
    layer2_outputs(4001) <= not(layer1_outputs(1950)) or (layer1_outputs(5077));
    layer2_outputs(4002) <= not(layer1_outputs(4274)) or (layer1_outputs(3151));
    layer2_outputs(4003) <= not(layer1_outputs(4378)) or (layer1_outputs(94));
    layer2_outputs(4004) <= layer1_outputs(4502);
    layer2_outputs(4005) <= (layer1_outputs(2876)) and (layer1_outputs(4380));
    layer2_outputs(4006) <= not(layer1_outputs(104));
    layer2_outputs(4007) <= layer1_outputs(4425);
    layer2_outputs(4008) <= not(layer1_outputs(1010));
    layer2_outputs(4009) <= layer1_outputs(1102);
    layer2_outputs(4010) <= layer1_outputs(4967);
    layer2_outputs(4011) <= (layer1_outputs(3484)) and (layer1_outputs(3764));
    layer2_outputs(4012) <= layer1_outputs(1825);
    layer2_outputs(4013) <= not(layer1_outputs(1131));
    layer2_outputs(4014) <= not((layer1_outputs(4953)) or (layer1_outputs(3170)));
    layer2_outputs(4015) <= layer1_outputs(1039);
    layer2_outputs(4016) <= not(layer1_outputs(3234)) or (layer1_outputs(691));
    layer2_outputs(4017) <= (layer1_outputs(2502)) and not (layer1_outputs(3867));
    layer2_outputs(4018) <= layer1_outputs(2520);
    layer2_outputs(4019) <= not((layer1_outputs(2652)) and (layer1_outputs(2413)));
    layer2_outputs(4020) <= layer1_outputs(1653);
    layer2_outputs(4021) <= (layer1_outputs(196)) xor (layer1_outputs(4691));
    layer2_outputs(4022) <= not(layer1_outputs(4593));
    layer2_outputs(4023) <= not((layer1_outputs(2671)) and (layer1_outputs(233)));
    layer2_outputs(4024) <= '0';
    layer2_outputs(4025) <= not((layer1_outputs(375)) or (layer1_outputs(3115)));
    layer2_outputs(4026) <= not(layer1_outputs(4775)) or (layer1_outputs(2556));
    layer2_outputs(4027) <= not((layer1_outputs(2490)) and (layer1_outputs(1476)));
    layer2_outputs(4028) <= not(layer1_outputs(2020));
    layer2_outputs(4029) <= not((layer1_outputs(4337)) xor (layer1_outputs(4200)));
    layer2_outputs(4030) <= (layer1_outputs(3110)) and not (layer1_outputs(3442));
    layer2_outputs(4031) <= layer1_outputs(517);
    layer2_outputs(4032) <= not(layer1_outputs(4280)) or (layer1_outputs(2009));
    layer2_outputs(4033) <= not((layer1_outputs(1256)) and (layer1_outputs(4940)));
    layer2_outputs(4034) <= (layer1_outputs(4252)) xor (layer1_outputs(1096));
    layer2_outputs(4035) <= not(layer1_outputs(3305));
    layer2_outputs(4036) <= (layer1_outputs(4374)) and not (layer1_outputs(43));
    layer2_outputs(4037) <= not(layer1_outputs(1258)) or (layer1_outputs(2965));
    layer2_outputs(4038) <= not(layer1_outputs(1769));
    layer2_outputs(4039) <= not(layer1_outputs(4571));
    layer2_outputs(4040) <= layer1_outputs(1377);
    layer2_outputs(4041) <= not(layer1_outputs(2236));
    layer2_outputs(4042) <= layer1_outputs(792);
    layer2_outputs(4043) <= not(layer1_outputs(4194));
    layer2_outputs(4044) <= (layer1_outputs(4445)) and not (layer1_outputs(4232));
    layer2_outputs(4045) <= (layer1_outputs(1893)) and not (layer1_outputs(4898));
    layer2_outputs(4046) <= not((layer1_outputs(4747)) or (layer1_outputs(4018)));
    layer2_outputs(4047) <= not(layer1_outputs(150));
    layer2_outputs(4048) <= not(layer1_outputs(3));
    layer2_outputs(4049) <= not(layer1_outputs(3287)) or (layer1_outputs(2197));
    layer2_outputs(4050) <= not(layer1_outputs(449));
    layer2_outputs(4051) <= (layer1_outputs(1608)) or (layer1_outputs(3206));
    layer2_outputs(4052) <= not(layer1_outputs(3111));
    layer2_outputs(4053) <= not(layer1_outputs(3365)) or (layer1_outputs(4861));
    layer2_outputs(4054) <= not(layer1_outputs(3136));
    layer2_outputs(4055) <= not((layer1_outputs(1367)) xor (layer1_outputs(3211)));
    layer2_outputs(4056) <= (layer1_outputs(4003)) and (layer1_outputs(3864));
    layer2_outputs(4057) <= (layer1_outputs(1547)) and not (layer1_outputs(3172));
    layer2_outputs(4058) <= layer1_outputs(1386);
    layer2_outputs(4059) <= not(layer1_outputs(3682));
    layer2_outputs(4060) <= '0';
    layer2_outputs(4061) <= (layer1_outputs(1863)) or (layer1_outputs(2845));
    layer2_outputs(4062) <= layer1_outputs(122);
    layer2_outputs(4063) <= not(layer1_outputs(4804));
    layer2_outputs(4064) <= not((layer1_outputs(1670)) and (layer1_outputs(1156)));
    layer2_outputs(4065) <= not(layer1_outputs(2661));
    layer2_outputs(4066) <= not(layer1_outputs(1011));
    layer2_outputs(4067) <= not(layer1_outputs(4022)) or (layer1_outputs(1189));
    layer2_outputs(4068) <= layer1_outputs(1850);
    layer2_outputs(4069) <= (layer1_outputs(3758)) or (layer1_outputs(4385));
    layer2_outputs(4070) <= not(layer1_outputs(96));
    layer2_outputs(4071) <= not(layer1_outputs(2082)) or (layer1_outputs(4702));
    layer2_outputs(4072) <= (layer1_outputs(1907)) or (layer1_outputs(5062));
    layer2_outputs(4073) <= (layer1_outputs(4234)) and not (layer1_outputs(3721));
    layer2_outputs(4074) <= (layer1_outputs(4484)) and (layer1_outputs(444));
    layer2_outputs(4075) <= not((layer1_outputs(25)) or (layer1_outputs(2508)));
    layer2_outputs(4076) <= layer1_outputs(319);
    layer2_outputs(4077) <= layer1_outputs(2789);
    layer2_outputs(4078) <= (layer1_outputs(4053)) and (layer1_outputs(3855));
    layer2_outputs(4079) <= not(layer1_outputs(3270));
    layer2_outputs(4080) <= layer1_outputs(1841);
    layer2_outputs(4081) <= not((layer1_outputs(36)) xor (layer1_outputs(2773)));
    layer2_outputs(4082) <= not((layer1_outputs(4286)) or (layer1_outputs(4845)));
    layer2_outputs(4083) <= not((layer1_outputs(2089)) and (layer1_outputs(4837)));
    layer2_outputs(4084) <= not(layer1_outputs(2649));
    layer2_outputs(4085) <= (layer1_outputs(1541)) or (layer1_outputs(2446));
    layer2_outputs(4086) <= (layer1_outputs(1733)) or (layer1_outputs(1050));
    layer2_outputs(4087) <= not(layer1_outputs(2467));
    layer2_outputs(4088) <= not((layer1_outputs(296)) and (layer1_outputs(1660)));
    layer2_outputs(4089) <= (layer1_outputs(1826)) and not (layer1_outputs(4415));
    layer2_outputs(4090) <= layer1_outputs(3024);
    layer2_outputs(4091) <= not(layer1_outputs(4072));
    layer2_outputs(4092) <= layer1_outputs(2821);
    layer2_outputs(4093) <= not(layer1_outputs(1583)) or (layer1_outputs(1877));
    layer2_outputs(4094) <= not(layer1_outputs(4184));
    layer2_outputs(4095) <= (layer1_outputs(59)) or (layer1_outputs(1237));
    layer2_outputs(4096) <= (layer1_outputs(788)) xor (layer1_outputs(2094));
    layer2_outputs(4097) <= not(layer1_outputs(41));
    layer2_outputs(4098) <= (layer1_outputs(3446)) and not (layer1_outputs(609));
    layer2_outputs(4099) <= layer1_outputs(968);
    layer2_outputs(4100) <= layer1_outputs(1241);
    layer2_outputs(4101) <= not(layer1_outputs(127)) or (layer1_outputs(3581));
    layer2_outputs(4102) <= not(layer1_outputs(2897)) or (layer1_outputs(4377));
    layer2_outputs(4103) <= not(layer1_outputs(2851)) or (layer1_outputs(3306));
    layer2_outputs(4104) <= not(layer1_outputs(854));
    layer2_outputs(4105) <= layer1_outputs(1932);
    layer2_outputs(4106) <= layer1_outputs(2867);
    layer2_outputs(4107) <= layer1_outputs(1534);
    layer2_outputs(4108) <= layer1_outputs(1086);
    layer2_outputs(4109) <= layer1_outputs(4969);
    layer2_outputs(4110) <= not((layer1_outputs(1491)) or (layer1_outputs(4869)));
    layer2_outputs(4111) <= not((layer1_outputs(3946)) and (layer1_outputs(859)));
    layer2_outputs(4112) <= not(layer1_outputs(821)) or (layer1_outputs(1424));
    layer2_outputs(4113) <= not((layer1_outputs(2758)) and (layer1_outputs(2021)));
    layer2_outputs(4114) <= layer1_outputs(2036);
    layer2_outputs(4115) <= not(layer1_outputs(2103));
    layer2_outputs(4116) <= layer1_outputs(1075);
    layer2_outputs(4117) <= not(layer1_outputs(3046)) or (layer1_outputs(3080));
    layer2_outputs(4118) <= (layer1_outputs(3263)) and not (layer1_outputs(3844));
    layer2_outputs(4119) <= layer1_outputs(4801);
    layer2_outputs(4120) <= not(layer1_outputs(2870));
    layer2_outputs(4121) <= (layer1_outputs(993)) and (layer1_outputs(1933));
    layer2_outputs(4122) <= layer1_outputs(4355);
    layer2_outputs(4123) <= not(layer1_outputs(461));
    layer2_outputs(4124) <= not(layer1_outputs(4081));
    layer2_outputs(4125) <= (layer1_outputs(1128)) and not (layer1_outputs(601));
    layer2_outputs(4126) <= not(layer1_outputs(1679)) or (layer1_outputs(2262));
    layer2_outputs(4127) <= '0';
    layer2_outputs(4128) <= '0';
    layer2_outputs(4129) <= not((layer1_outputs(3286)) and (layer1_outputs(216)));
    layer2_outputs(4130) <= not(layer1_outputs(2842));
    layer2_outputs(4131) <= (layer1_outputs(3299)) and (layer1_outputs(1557));
    layer2_outputs(4132) <= (layer1_outputs(2695)) or (layer1_outputs(348));
    layer2_outputs(4133) <= not(layer1_outputs(920));
    layer2_outputs(4134) <= not(layer1_outputs(4785)) or (layer1_outputs(1167));
    layer2_outputs(4135) <= not(layer1_outputs(4655));
    layer2_outputs(4136) <= not(layer1_outputs(126));
    layer2_outputs(4137) <= (layer1_outputs(1108)) or (layer1_outputs(183));
    layer2_outputs(4138) <= layer1_outputs(1999);
    layer2_outputs(4139) <= layer1_outputs(3168);
    layer2_outputs(4140) <= (layer1_outputs(700)) xor (layer1_outputs(1207));
    layer2_outputs(4141) <= not(layer1_outputs(2598));
    layer2_outputs(4142) <= layer1_outputs(742);
    layer2_outputs(4143) <= (layer1_outputs(4588)) and not (layer1_outputs(3222));
    layer2_outputs(4144) <= (layer1_outputs(2828)) and not (layer1_outputs(920));
    layer2_outputs(4145) <= not(layer1_outputs(244)) or (layer1_outputs(4491));
    layer2_outputs(4146) <= (layer1_outputs(1970)) or (layer1_outputs(3709));
    layer2_outputs(4147) <= layer1_outputs(1472);
    layer2_outputs(4148) <= not(layer1_outputs(1946));
    layer2_outputs(4149) <= not(layer1_outputs(4014));
    layer2_outputs(4150) <= (layer1_outputs(1093)) or (layer1_outputs(626));
    layer2_outputs(4151) <= not(layer1_outputs(472));
    layer2_outputs(4152) <= not(layer1_outputs(1053));
    layer2_outputs(4153) <= layer1_outputs(2776);
    layer2_outputs(4154) <= (layer1_outputs(2084)) and not (layer1_outputs(637));
    layer2_outputs(4155) <= not(layer1_outputs(2176));
    layer2_outputs(4156) <= not((layer1_outputs(4836)) or (layer1_outputs(1440)));
    layer2_outputs(4157) <= not(layer1_outputs(1325)) or (layer1_outputs(344));
    layer2_outputs(4158) <= (layer1_outputs(673)) and not (layer1_outputs(5110));
    layer2_outputs(4159) <= not(layer1_outputs(2521));
    layer2_outputs(4160) <= layer1_outputs(4162);
    layer2_outputs(4161) <= not(layer1_outputs(4421)) or (layer1_outputs(1246));
    layer2_outputs(4162) <= not(layer1_outputs(1477)) or (layer1_outputs(4584));
    layer2_outputs(4163) <= (layer1_outputs(522)) and (layer1_outputs(2604));
    layer2_outputs(4164) <= layer1_outputs(2601);
    layer2_outputs(4165) <= not((layer1_outputs(3147)) or (layer1_outputs(1891)));
    layer2_outputs(4166) <= layer1_outputs(3910);
    layer2_outputs(4167) <= not(layer1_outputs(2903));
    layer2_outputs(4168) <= '0';
    layer2_outputs(4169) <= layer1_outputs(3766);
    layer2_outputs(4170) <= not(layer1_outputs(3448));
    layer2_outputs(4171) <= not(layer1_outputs(464));
    layer2_outputs(4172) <= not((layer1_outputs(2512)) or (layer1_outputs(121)));
    layer2_outputs(4173) <= not(layer1_outputs(841));
    layer2_outputs(4174) <= not(layer1_outputs(1775));
    layer2_outputs(4175) <= not(layer1_outputs(725)) or (layer1_outputs(2711));
    layer2_outputs(4176) <= layer1_outputs(527);
    layer2_outputs(4177) <= not(layer1_outputs(947));
    layer2_outputs(4178) <= not(layer1_outputs(4778)) or (layer1_outputs(2510));
    layer2_outputs(4179) <= (layer1_outputs(4453)) xor (layer1_outputs(397));
    layer2_outputs(4180) <= (layer1_outputs(801)) or (layer1_outputs(3159));
    layer2_outputs(4181) <= not((layer1_outputs(1627)) and (layer1_outputs(2376)));
    layer2_outputs(4182) <= not((layer1_outputs(4482)) xor (layer1_outputs(833)));
    layer2_outputs(4183) <= not(layer1_outputs(1707));
    layer2_outputs(4184) <= (layer1_outputs(1617)) and not (layer1_outputs(144));
    layer2_outputs(4185) <= layer1_outputs(2467);
    layer2_outputs(4186) <= layer1_outputs(550);
    layer2_outputs(4187) <= '1';
    layer2_outputs(4188) <= layer1_outputs(2277);
    layer2_outputs(4189) <= layer1_outputs(479);
    layer2_outputs(4190) <= layer1_outputs(2854);
    layer2_outputs(4191) <= (layer1_outputs(193)) and not (layer1_outputs(4674));
    layer2_outputs(4192) <= not(layer1_outputs(288));
    layer2_outputs(4193) <= layer1_outputs(3385);
    layer2_outputs(4194) <= layer1_outputs(3793);
    layer2_outputs(4195) <= layer1_outputs(1619);
    layer2_outputs(4196) <= not(layer1_outputs(1764));
    layer2_outputs(4197) <= (layer1_outputs(1269)) or (layer1_outputs(3238));
    layer2_outputs(4198) <= not(layer1_outputs(1949));
    layer2_outputs(4199) <= (layer1_outputs(987)) and not (layer1_outputs(1246));
    layer2_outputs(4200) <= (layer1_outputs(2111)) and not (layer1_outputs(4526));
    layer2_outputs(4201) <= (layer1_outputs(2505)) or (layer1_outputs(5062));
    layer2_outputs(4202) <= (layer1_outputs(1461)) and not (layer1_outputs(1679));
    layer2_outputs(4203) <= not(layer1_outputs(3196));
    layer2_outputs(4204) <= layer1_outputs(2796);
    layer2_outputs(4205) <= layer1_outputs(4987);
    layer2_outputs(4206) <= (layer1_outputs(1433)) and not (layer1_outputs(1674));
    layer2_outputs(4207) <= layer1_outputs(3450);
    layer2_outputs(4208) <= not((layer1_outputs(5103)) xor (layer1_outputs(1770)));
    layer2_outputs(4209) <= not(layer1_outputs(232));
    layer2_outputs(4210) <= layer1_outputs(1116);
    layer2_outputs(4211) <= layer1_outputs(5093);
    layer2_outputs(4212) <= not((layer1_outputs(869)) and (layer1_outputs(1403)));
    layer2_outputs(4213) <= (layer1_outputs(1226)) and not (layer1_outputs(3227));
    layer2_outputs(4214) <= (layer1_outputs(618)) and not (layer1_outputs(2139));
    layer2_outputs(4215) <= layer1_outputs(2219);
    layer2_outputs(4216) <= not(layer1_outputs(480));
    layer2_outputs(4217) <= not(layer1_outputs(3941));
    layer2_outputs(4218) <= layer1_outputs(3650);
    layer2_outputs(4219) <= not((layer1_outputs(484)) or (layer1_outputs(3832)));
    layer2_outputs(4220) <= not(layer1_outputs(1888));
    layer2_outputs(4221) <= layer1_outputs(1921);
    layer2_outputs(4222) <= not(layer1_outputs(1308));
    layer2_outputs(4223) <= layer1_outputs(3281);
    layer2_outputs(4224) <= not(layer1_outputs(1220));
    layer2_outputs(4225) <= not(layer1_outputs(2181));
    layer2_outputs(4226) <= (layer1_outputs(3234)) and (layer1_outputs(2841));
    layer2_outputs(4227) <= layer1_outputs(4138);
    layer2_outputs(4228) <= layer1_outputs(4953);
    layer2_outputs(4229) <= not(layer1_outputs(3720));
    layer2_outputs(4230) <= layer1_outputs(3308);
    layer2_outputs(4231) <= layer1_outputs(1943);
    layer2_outputs(4232) <= layer1_outputs(1006);
    layer2_outputs(4233) <= (layer1_outputs(1940)) and not (layer1_outputs(4958));
    layer2_outputs(4234) <= '1';
    layer2_outputs(4235) <= (layer1_outputs(4330)) and (layer1_outputs(683));
    layer2_outputs(4236) <= not(layer1_outputs(4901));
    layer2_outputs(4237) <= not(layer1_outputs(4271)) or (layer1_outputs(290));
    layer2_outputs(4238) <= '0';
    layer2_outputs(4239) <= (layer1_outputs(4250)) or (layer1_outputs(5027));
    layer2_outputs(4240) <= not(layer1_outputs(4696)) or (layer1_outputs(3784));
    layer2_outputs(4241) <= (layer1_outputs(4508)) and (layer1_outputs(1400));
    layer2_outputs(4242) <= not(layer1_outputs(1544));
    layer2_outputs(4243) <= layer1_outputs(2026);
    layer2_outputs(4244) <= layer1_outputs(2272);
    layer2_outputs(4245) <= (layer1_outputs(1511)) xor (layer1_outputs(4687));
    layer2_outputs(4246) <= not((layer1_outputs(1802)) xor (layer1_outputs(3318)));
    layer2_outputs(4247) <= (layer1_outputs(1783)) and not (layer1_outputs(745));
    layer2_outputs(4248) <= not(layer1_outputs(3503));
    layer2_outputs(4249) <= not((layer1_outputs(1524)) and (layer1_outputs(2635)));
    layer2_outputs(4250) <= not(layer1_outputs(1988));
    layer2_outputs(4251) <= not(layer1_outputs(3227)) or (layer1_outputs(2587));
    layer2_outputs(4252) <= layer1_outputs(1559);
    layer2_outputs(4253) <= not(layer1_outputs(3096));
    layer2_outputs(4254) <= layer1_outputs(4817);
    layer2_outputs(4255) <= layer1_outputs(1253);
    layer2_outputs(4256) <= (layer1_outputs(4363)) xor (layer1_outputs(2934));
    layer2_outputs(4257) <= layer1_outputs(2616);
    layer2_outputs(4258) <= not(layer1_outputs(2654));
    layer2_outputs(4259) <= not(layer1_outputs(3456));
    layer2_outputs(4260) <= not(layer1_outputs(2466)) or (layer1_outputs(5021));
    layer2_outputs(4261) <= layer1_outputs(3478);
    layer2_outputs(4262) <= (layer1_outputs(3071)) and not (layer1_outputs(3381));
    layer2_outputs(4263) <= not(layer1_outputs(28));
    layer2_outputs(4264) <= not(layer1_outputs(724));
    layer2_outputs(4265) <= not(layer1_outputs(154));
    layer2_outputs(4266) <= (layer1_outputs(871)) and not (layer1_outputs(4763));
    layer2_outputs(4267) <= not(layer1_outputs(982)) or (layer1_outputs(1562));
    layer2_outputs(4268) <= layer1_outputs(2536);
    layer2_outputs(4269) <= (layer1_outputs(3403)) and not (layer1_outputs(2453));
    layer2_outputs(4270) <= '0';
    layer2_outputs(4271) <= not(layer1_outputs(2931)) or (layer1_outputs(4449));
    layer2_outputs(4272) <= (layer1_outputs(5024)) and (layer1_outputs(3940));
    layer2_outputs(4273) <= (layer1_outputs(1297)) or (layer1_outputs(1966));
    layer2_outputs(4274) <= not(layer1_outputs(1363));
    layer2_outputs(4275) <= layer1_outputs(3191);
    layer2_outputs(4276) <= not(layer1_outputs(1438));
    layer2_outputs(4277) <= layer1_outputs(4839);
    layer2_outputs(4278) <= not(layer1_outputs(4204));
    layer2_outputs(4279) <= (layer1_outputs(4858)) and not (layer1_outputs(259));
    layer2_outputs(4280) <= layer1_outputs(1806);
    layer2_outputs(4281) <= not(layer1_outputs(3078)) or (layer1_outputs(3921));
    layer2_outputs(4282) <= not(layer1_outputs(3375));
    layer2_outputs(4283) <= not((layer1_outputs(2700)) xor (layer1_outputs(1071)));
    layer2_outputs(4284) <= not(layer1_outputs(1980));
    layer2_outputs(4285) <= (layer1_outputs(1614)) xor (layer1_outputs(3967));
    layer2_outputs(4286) <= layer1_outputs(464);
    layer2_outputs(4287) <= layer1_outputs(899);
    layer2_outputs(4288) <= not(layer1_outputs(2038));
    layer2_outputs(4289) <= layer1_outputs(1325);
    layer2_outputs(4290) <= '1';
    layer2_outputs(4291) <= (layer1_outputs(2619)) or (layer1_outputs(3078));
    layer2_outputs(4292) <= not((layer1_outputs(3445)) and (layer1_outputs(2193)));
    layer2_outputs(4293) <= layer1_outputs(3198);
    layer2_outputs(4294) <= (layer1_outputs(3835)) or (layer1_outputs(4344));
    layer2_outputs(4295) <= not((layer1_outputs(749)) and (layer1_outputs(2623)));
    layer2_outputs(4296) <= not((layer1_outputs(2076)) and (layer1_outputs(532)));
    layer2_outputs(4297) <= (layer1_outputs(3397)) xor (layer1_outputs(5034));
    layer2_outputs(4298) <= (layer1_outputs(1538)) xor (layer1_outputs(1111));
    layer2_outputs(4299) <= not((layer1_outputs(1673)) and (layer1_outputs(254)));
    layer2_outputs(4300) <= (layer1_outputs(3192)) and (layer1_outputs(274));
    layer2_outputs(4301) <= not(layer1_outputs(3094));
    layer2_outputs(4302) <= layer1_outputs(3743);
    layer2_outputs(4303) <= not((layer1_outputs(1038)) and (layer1_outputs(3483)));
    layer2_outputs(4304) <= (layer1_outputs(3148)) xor (layer1_outputs(3213));
    layer2_outputs(4305) <= not((layer1_outputs(2593)) and (layer1_outputs(3698)));
    layer2_outputs(4306) <= not(layer1_outputs(5048)) or (layer1_outputs(436));
    layer2_outputs(4307) <= not(layer1_outputs(4021)) or (layer1_outputs(4201));
    layer2_outputs(4308) <= '0';
    layer2_outputs(4309) <= not(layer1_outputs(535));
    layer2_outputs(4310) <= not(layer1_outputs(1606));
    layer2_outputs(4311) <= not((layer1_outputs(552)) xor (layer1_outputs(3842)));
    layer2_outputs(4312) <= layer1_outputs(1545);
    layer2_outputs(4313) <= layer1_outputs(2656);
    layer2_outputs(4314) <= (layer1_outputs(169)) and not (layer1_outputs(760));
    layer2_outputs(4315) <= layer1_outputs(635);
    layer2_outputs(4316) <= layer1_outputs(170);
    layer2_outputs(4317) <= (layer1_outputs(4750)) xor (layer1_outputs(3392));
    layer2_outputs(4318) <= not(layer1_outputs(3802));
    layer2_outputs(4319) <= layer1_outputs(3257);
    layer2_outputs(4320) <= layer1_outputs(5083);
    layer2_outputs(4321) <= (layer1_outputs(4040)) and not (layer1_outputs(1381));
    layer2_outputs(4322) <= (layer1_outputs(2177)) and not (layer1_outputs(1489));
    layer2_outputs(4323) <= (layer1_outputs(3071)) or (layer1_outputs(2398));
    layer2_outputs(4324) <= layer1_outputs(2778);
    layer2_outputs(4325) <= not(layer1_outputs(4493));
    layer2_outputs(4326) <= not(layer1_outputs(11));
    layer2_outputs(4327) <= not(layer1_outputs(4000));
    layer2_outputs(4328) <= layer1_outputs(4688);
    layer2_outputs(4329) <= (layer1_outputs(1436)) and not (layer1_outputs(3975));
    layer2_outputs(4330) <= not(layer1_outputs(2827));
    layer2_outputs(4331) <= not(layer1_outputs(3642)) or (layer1_outputs(3993));
    layer2_outputs(4332) <= layer1_outputs(2921);
    layer2_outputs(4333) <= not(layer1_outputs(2026));
    layer2_outputs(4334) <= layer1_outputs(1607);
    layer2_outputs(4335) <= not(layer1_outputs(4560));
    layer2_outputs(4336) <= (layer1_outputs(1777)) and (layer1_outputs(3861));
    layer2_outputs(4337) <= not(layer1_outputs(2335));
    layer2_outputs(4338) <= layer1_outputs(4770);
    layer2_outputs(4339) <= not(layer1_outputs(405));
    layer2_outputs(4340) <= not(layer1_outputs(383)) or (layer1_outputs(2797));
    layer2_outputs(4341) <= (layer1_outputs(407)) and not (layer1_outputs(4469));
    layer2_outputs(4342) <= layer1_outputs(4370);
    layer2_outputs(4343) <= (layer1_outputs(743)) and not (layer1_outputs(386));
    layer2_outputs(4344) <= not(layer1_outputs(3797)) or (layer1_outputs(1125));
    layer2_outputs(4345) <= not((layer1_outputs(1887)) or (layer1_outputs(1600)));
    layer2_outputs(4346) <= not(layer1_outputs(2603));
    layer2_outputs(4347) <= (layer1_outputs(4517)) and not (layer1_outputs(3054));
    layer2_outputs(4348) <= (layer1_outputs(552)) and not (layer1_outputs(232));
    layer2_outputs(4349) <= (layer1_outputs(4903)) or (layer1_outputs(1360));
    layer2_outputs(4350) <= (layer1_outputs(974)) and not (layer1_outputs(4893));
    layer2_outputs(4351) <= not(layer1_outputs(2955));
    layer2_outputs(4352) <= not(layer1_outputs(2091)) or (layer1_outputs(744));
    layer2_outputs(4353) <= (layer1_outputs(4541)) and (layer1_outputs(4785));
    layer2_outputs(4354) <= not(layer1_outputs(165));
    layer2_outputs(4355) <= layer1_outputs(416);
    layer2_outputs(4356) <= (layer1_outputs(1033)) or (layer1_outputs(367));
    layer2_outputs(4357) <= layer1_outputs(4473);
    layer2_outputs(4358) <= not(layer1_outputs(4858)) or (layer1_outputs(196));
    layer2_outputs(4359) <= not(layer1_outputs(1976));
    layer2_outputs(4360) <= not(layer1_outputs(3201)) or (layer1_outputs(2013));
    layer2_outputs(4361) <= (layer1_outputs(4259)) and (layer1_outputs(5115));
    layer2_outputs(4362) <= not(layer1_outputs(3083));
    layer2_outputs(4363) <= not(layer1_outputs(1525));
    layer2_outputs(4364) <= layer1_outputs(4526);
    layer2_outputs(4365) <= not(layer1_outputs(1));
    layer2_outputs(4366) <= not(layer1_outputs(717));
    layer2_outputs(4367) <= layer1_outputs(4050);
    layer2_outputs(4368) <= '1';
    layer2_outputs(4369) <= layer1_outputs(4542);
    layer2_outputs(4370) <= not((layer1_outputs(1807)) or (layer1_outputs(4073)));
    layer2_outputs(4371) <= not((layer1_outputs(32)) and (layer1_outputs(965)));
    layer2_outputs(4372) <= layer1_outputs(1595);
    layer2_outputs(4373) <= layer1_outputs(3109);
    layer2_outputs(4374) <= layer1_outputs(2203);
    layer2_outputs(4375) <= (layer1_outputs(2544)) and (layer1_outputs(4680));
    layer2_outputs(4376) <= not(layer1_outputs(1316));
    layer2_outputs(4377) <= layer1_outputs(4164);
    layer2_outputs(4378) <= not(layer1_outputs(1587)) or (layer1_outputs(4689));
    layer2_outputs(4379) <= layer1_outputs(3165);
    layer2_outputs(4380) <= not(layer1_outputs(581)) or (layer1_outputs(4849));
    layer2_outputs(4381) <= layer1_outputs(2066);
    layer2_outputs(4382) <= not(layer1_outputs(3700));
    layer2_outputs(4383) <= not(layer1_outputs(34)) or (layer1_outputs(4001));
    layer2_outputs(4384) <= (layer1_outputs(2094)) xor (layer1_outputs(3763));
    layer2_outputs(4385) <= (layer1_outputs(3849)) xor (layer1_outputs(1682));
    layer2_outputs(4386) <= (layer1_outputs(4076)) or (layer1_outputs(1051));
    layer2_outputs(4387) <= (layer1_outputs(1661)) and (layer1_outputs(372));
    layer2_outputs(4388) <= '0';
    layer2_outputs(4389) <= not(layer1_outputs(4046));
    layer2_outputs(4390) <= layer1_outputs(2794);
    layer2_outputs(4391) <= not(layer1_outputs(976)) or (layer1_outputs(588));
    layer2_outputs(4392) <= not(layer1_outputs(2006));
    layer2_outputs(4393) <= (layer1_outputs(2405)) and not (layer1_outputs(292));
    layer2_outputs(4394) <= not((layer1_outputs(1159)) xor (layer1_outputs(1120)));
    layer2_outputs(4395) <= (layer1_outputs(3800)) and (layer1_outputs(2823));
    layer2_outputs(4396) <= (layer1_outputs(1983)) or (layer1_outputs(17));
    layer2_outputs(4397) <= (layer1_outputs(2236)) and (layer1_outputs(4240));
    layer2_outputs(4398) <= not((layer1_outputs(1308)) or (layer1_outputs(1030)));
    layer2_outputs(4399) <= (layer1_outputs(1331)) and (layer1_outputs(4974));
    layer2_outputs(4400) <= layer1_outputs(0);
    layer2_outputs(4401) <= layer1_outputs(4253);
    layer2_outputs(4402) <= layer1_outputs(554);
    layer2_outputs(4403) <= not((layer1_outputs(1912)) and (layer1_outputs(1141)));
    layer2_outputs(4404) <= not(layer1_outputs(4072));
    layer2_outputs(4405) <= layer1_outputs(1514);
    layer2_outputs(4406) <= (layer1_outputs(1168)) and (layer1_outputs(1467));
    layer2_outputs(4407) <= layer1_outputs(3865);
    layer2_outputs(4408) <= not((layer1_outputs(181)) and (layer1_outputs(2780)));
    layer2_outputs(4409) <= (layer1_outputs(1742)) and (layer1_outputs(3293));
    layer2_outputs(4410) <= not(layer1_outputs(2507));
    layer2_outputs(4411) <= layer1_outputs(2403);
    layer2_outputs(4412) <= not((layer1_outputs(2585)) and (layer1_outputs(5011)));
    layer2_outputs(4413) <= not(layer1_outputs(1519));
    layer2_outputs(4414) <= not(layer1_outputs(1659));
    layer2_outputs(4415) <= layer1_outputs(4853);
    layer2_outputs(4416) <= layer1_outputs(4178);
    layer2_outputs(4417) <= not(layer1_outputs(978));
    layer2_outputs(4418) <= not((layer1_outputs(1247)) or (layer1_outputs(709)));
    layer2_outputs(4419) <= not(layer1_outputs(2302));
    layer2_outputs(4420) <= not((layer1_outputs(844)) and (layer1_outputs(4699)));
    layer2_outputs(4421) <= not((layer1_outputs(3051)) and (layer1_outputs(1902)));
    layer2_outputs(4422) <= layer1_outputs(1725);
    layer2_outputs(4423) <= (layer1_outputs(1489)) and not (layer1_outputs(358));
    layer2_outputs(4424) <= not(layer1_outputs(1675));
    layer2_outputs(4425) <= not(layer1_outputs(905));
    layer2_outputs(4426) <= (layer1_outputs(3050)) or (layer1_outputs(3491));
    layer2_outputs(4427) <= not((layer1_outputs(39)) and (layer1_outputs(4663)));
    layer2_outputs(4428) <= not(layer1_outputs(884));
    layer2_outputs(4429) <= not(layer1_outputs(3748));
    layer2_outputs(4430) <= not((layer1_outputs(52)) and (layer1_outputs(3905)));
    layer2_outputs(4431) <= not((layer1_outputs(3834)) or (layer1_outputs(3702)));
    layer2_outputs(4432) <= (layer1_outputs(499)) and (layer1_outputs(3451));
    layer2_outputs(4433) <= layer1_outputs(2584);
    layer2_outputs(4434) <= layer1_outputs(2813);
    layer2_outputs(4435) <= not(layer1_outputs(2367));
    layer2_outputs(4436) <= not(layer1_outputs(3413));
    layer2_outputs(4437) <= '0';
    layer2_outputs(4438) <= not(layer1_outputs(4741)) or (layer1_outputs(3575));
    layer2_outputs(4439) <= not(layer1_outputs(37));
    layer2_outputs(4440) <= (layer1_outputs(4996)) and not (layer1_outputs(48));
    layer2_outputs(4441) <= (layer1_outputs(4394)) and not (layer1_outputs(2640));
    layer2_outputs(4442) <= not(layer1_outputs(3309)) or (layer1_outputs(1127));
    layer2_outputs(4443) <= not(layer1_outputs(2022)) or (layer1_outputs(3438));
    layer2_outputs(4444) <= not((layer1_outputs(2817)) and (layer1_outputs(1221)));
    layer2_outputs(4445) <= not(layer1_outputs(600));
    layer2_outputs(4446) <= not((layer1_outputs(3912)) xor (layer1_outputs(4217)));
    layer2_outputs(4447) <= not(layer1_outputs(1653));
    layer2_outputs(4448) <= '1';
    layer2_outputs(4449) <= (layer1_outputs(1004)) and (layer1_outputs(1095));
    layer2_outputs(4450) <= not(layer1_outputs(4317));
    layer2_outputs(4451) <= layer1_outputs(2025);
    layer2_outputs(4452) <= layer1_outputs(3644);
    layer2_outputs(4453) <= layer1_outputs(44);
    layer2_outputs(4454) <= layer1_outputs(3329);
    layer2_outputs(4455) <= '1';
    layer2_outputs(4456) <= not(layer1_outputs(2739));
    layer2_outputs(4457) <= not(layer1_outputs(2888));
    layer2_outputs(4458) <= (layer1_outputs(3539)) and not (layer1_outputs(4647));
    layer2_outputs(4459) <= not((layer1_outputs(1867)) or (layer1_outputs(4345)));
    layer2_outputs(4460) <= (layer1_outputs(1462)) and not (layer1_outputs(665));
    layer2_outputs(4461) <= (layer1_outputs(2167)) and (layer1_outputs(3922));
    layer2_outputs(4462) <= not((layer1_outputs(2585)) or (layer1_outputs(3452)));
    layer2_outputs(4463) <= not((layer1_outputs(1437)) or (layer1_outputs(2777)));
    layer2_outputs(4464) <= layer1_outputs(835);
    layer2_outputs(4465) <= not(layer1_outputs(4658));
    layer2_outputs(4466) <= layer1_outputs(4401);
    layer2_outputs(4467) <= (layer1_outputs(4589)) or (layer1_outputs(3140));
    layer2_outputs(4468) <= not(layer1_outputs(4010)) or (layer1_outputs(136));
    layer2_outputs(4469) <= not(layer1_outputs(3319));
    layer2_outputs(4470) <= not(layer1_outputs(498)) or (layer1_outputs(2560));
    layer2_outputs(4471) <= (layer1_outputs(939)) xor (layer1_outputs(4884));
    layer2_outputs(4472) <= layer1_outputs(3279);
    layer2_outputs(4473) <= not((layer1_outputs(4694)) and (layer1_outputs(2233)));
    layer2_outputs(4474) <= layer1_outputs(4714);
    layer2_outputs(4475) <= layer1_outputs(272);
    layer2_outputs(4476) <= not(layer1_outputs(1905)) or (layer1_outputs(1718));
    layer2_outputs(4477) <= not(layer1_outputs(4223));
    layer2_outputs(4478) <= not(layer1_outputs(224));
    layer2_outputs(4479) <= not((layer1_outputs(2893)) or (layer1_outputs(2650)));
    layer2_outputs(4480) <= '0';
    layer2_outputs(4481) <= not(layer1_outputs(448));
    layer2_outputs(4482) <= not(layer1_outputs(3975)) or (layer1_outputs(1008));
    layer2_outputs(4483) <= (layer1_outputs(3898)) or (layer1_outputs(1999));
    layer2_outputs(4484) <= (layer1_outputs(4535)) xor (layer1_outputs(2615));
    layer2_outputs(4485) <= layer1_outputs(5029);
    layer2_outputs(4486) <= layer1_outputs(393);
    layer2_outputs(4487) <= not(layer1_outputs(4229));
    layer2_outputs(4488) <= layer1_outputs(3149);
    layer2_outputs(4489) <= '0';
    layer2_outputs(4490) <= '1';
    layer2_outputs(4491) <= layer1_outputs(3247);
    layer2_outputs(4492) <= layer1_outputs(3426);
    layer2_outputs(4493) <= not(layer1_outputs(4620));
    layer2_outputs(4494) <= not(layer1_outputs(970)) or (layer1_outputs(424));
    layer2_outputs(4495) <= not(layer1_outputs(3130)) or (layer1_outputs(2107));
    layer2_outputs(4496) <= layer1_outputs(1673);
    layer2_outputs(4497) <= layer1_outputs(1196);
    layer2_outputs(4498) <= not(layer1_outputs(1475));
    layer2_outputs(4499) <= (layer1_outputs(2668)) and not (layer1_outputs(3995));
    layer2_outputs(4500) <= layer1_outputs(3155);
    layer2_outputs(4501) <= not(layer1_outputs(2869)) or (layer1_outputs(4242));
    layer2_outputs(4502) <= not(layer1_outputs(4269));
    layer2_outputs(4503) <= (layer1_outputs(643)) or (layer1_outputs(224));
    layer2_outputs(4504) <= not(layer1_outputs(4843));
    layer2_outputs(4505) <= not((layer1_outputs(4071)) or (layer1_outputs(1598)));
    layer2_outputs(4506) <= layer1_outputs(632);
    layer2_outputs(4507) <= not(layer1_outputs(3933));
    layer2_outputs(4508) <= (layer1_outputs(1861)) or (layer1_outputs(594));
    layer2_outputs(4509) <= layer1_outputs(2291);
    layer2_outputs(4510) <= (layer1_outputs(1373)) and not (layer1_outputs(1498));
    layer2_outputs(4511) <= (layer1_outputs(3870)) or (layer1_outputs(3291));
    layer2_outputs(4512) <= (layer1_outputs(8)) and (layer1_outputs(3508));
    layer2_outputs(4513) <= (layer1_outputs(4888)) and not (layer1_outputs(4340));
    layer2_outputs(4514) <= (layer1_outputs(757)) and not (layer1_outputs(2503));
    layer2_outputs(4515) <= layer1_outputs(2529);
    layer2_outputs(4516) <= layer1_outputs(4460);
    layer2_outputs(4517) <= not(layer1_outputs(4711));
    layer2_outputs(4518) <= not((layer1_outputs(1581)) or (layer1_outputs(577)));
    layer2_outputs(4519) <= not(layer1_outputs(5038));
    layer2_outputs(4520) <= not(layer1_outputs(2362));
    layer2_outputs(4521) <= (layer1_outputs(2394)) and not (layer1_outputs(275));
    layer2_outputs(4522) <= (layer1_outputs(1592)) and not (layer1_outputs(3002));
    layer2_outputs(4523) <= not(layer1_outputs(3441));
    layer2_outputs(4524) <= not(layer1_outputs(2938));
    layer2_outputs(4525) <= (layer1_outputs(2682)) and (layer1_outputs(2838));
    layer2_outputs(4526) <= (layer1_outputs(919)) and not (layer1_outputs(1945));
    layer2_outputs(4527) <= not((layer1_outputs(465)) or (layer1_outputs(2471)));
    layer2_outputs(4528) <= (layer1_outputs(1751)) or (layer1_outputs(4891));
    layer2_outputs(4529) <= not(layer1_outputs(1580));
    layer2_outputs(4530) <= not((layer1_outputs(4649)) and (layer1_outputs(4601)));
    layer2_outputs(4531) <= layer1_outputs(4664);
    layer2_outputs(4532) <= layer1_outputs(3770);
    layer2_outputs(4533) <= not(layer1_outputs(4789));
    layer2_outputs(4534) <= '1';
    layer2_outputs(4535) <= (layer1_outputs(2922)) and (layer1_outputs(3311));
    layer2_outputs(4536) <= layer1_outputs(1628);
    layer2_outputs(4537) <= (layer1_outputs(359)) and not (layer1_outputs(2400));
    layer2_outputs(4538) <= (layer1_outputs(3789)) and not (layer1_outputs(78));
    layer2_outputs(4539) <= not(layer1_outputs(1410));
    layer2_outputs(4540) <= not(layer1_outputs(4220));
    layer2_outputs(4541) <= (layer1_outputs(246)) or (layer1_outputs(819));
    layer2_outputs(4542) <= not((layer1_outputs(5083)) xor (layer1_outputs(3711)));
    layer2_outputs(4543) <= not(layer1_outputs(3307));
    layer2_outputs(4544) <= not((layer1_outputs(373)) and (layer1_outputs(845)));
    layer2_outputs(4545) <= not((layer1_outputs(2611)) and (layer1_outputs(3013)));
    layer2_outputs(4546) <= '1';
    layer2_outputs(4547) <= not((layer1_outputs(548)) xor (layer1_outputs(2294)));
    layer2_outputs(4548) <= (layer1_outputs(4083)) and not (layer1_outputs(3076));
    layer2_outputs(4549) <= layer1_outputs(3024);
    layer2_outputs(4550) <= not(layer1_outputs(3135));
    layer2_outputs(4551) <= not(layer1_outputs(2756)) or (layer1_outputs(157));
    layer2_outputs(4552) <= layer1_outputs(1667);
    layer2_outputs(4553) <= not(layer1_outputs(715)) or (layer1_outputs(2613));
    layer2_outputs(4554) <= layer1_outputs(1849);
    layer2_outputs(4555) <= (layer1_outputs(2108)) and not (layer1_outputs(922));
    layer2_outputs(4556) <= layer1_outputs(5097);
    layer2_outputs(4557) <= not(layer1_outputs(3920));
    layer2_outputs(4558) <= layer1_outputs(857);
    layer2_outputs(4559) <= (layer1_outputs(2181)) and not (layer1_outputs(4382));
    layer2_outputs(4560) <= not(layer1_outputs(1706));
    layer2_outputs(4561) <= layer1_outputs(1629);
    layer2_outputs(4562) <= (layer1_outputs(4444)) or (layer1_outputs(203));
    layer2_outputs(4563) <= (layer1_outputs(3060)) and (layer1_outputs(5084));
    layer2_outputs(4564) <= not(layer1_outputs(2645));
    layer2_outputs(4565) <= not(layer1_outputs(3537));
    layer2_outputs(4566) <= (layer1_outputs(3894)) xor (layer1_outputs(4981));
    layer2_outputs(4567) <= layer1_outputs(2706);
    layer2_outputs(4568) <= layer1_outputs(176);
    layer2_outputs(4569) <= not((layer1_outputs(1816)) or (layer1_outputs(848)));
    layer2_outputs(4570) <= not(layer1_outputs(4446));
    layer2_outputs(4571) <= (layer1_outputs(2002)) and not (layer1_outputs(4732));
    layer2_outputs(4572) <= layer1_outputs(704);
    layer2_outputs(4573) <= (layer1_outputs(5071)) or (layer1_outputs(4933));
    layer2_outputs(4574) <= layer1_outputs(2459);
    layer2_outputs(4575) <= layer1_outputs(3303);
    layer2_outputs(4576) <= not((layer1_outputs(4781)) and (layer1_outputs(2942)));
    layer2_outputs(4577) <= not(layer1_outputs(2685));
    layer2_outputs(4578) <= layer1_outputs(3488);
    layer2_outputs(4579) <= not((layer1_outputs(374)) and (layer1_outputs(1726)));
    layer2_outputs(4580) <= layer1_outputs(4408);
    layer2_outputs(4581) <= (layer1_outputs(2410)) and (layer1_outputs(1327));
    layer2_outputs(4582) <= layer1_outputs(4186);
    layer2_outputs(4583) <= '0';
    layer2_outputs(4584) <= not(layer1_outputs(934));
    layer2_outputs(4585) <= not(layer1_outputs(3824));
    layer2_outputs(4586) <= not((layer1_outputs(3188)) and (layer1_outputs(258)));
    layer2_outputs(4587) <= (layer1_outputs(2565)) and (layer1_outputs(535));
    layer2_outputs(4588) <= (layer1_outputs(648)) and not (layer1_outputs(4592));
    layer2_outputs(4589) <= not(layer1_outputs(2739));
    layer2_outputs(4590) <= not((layer1_outputs(4097)) or (layer1_outputs(101)));
    layer2_outputs(4591) <= '1';
    layer2_outputs(4592) <= (layer1_outputs(2176)) and not (layer1_outputs(3278));
    layer2_outputs(4593) <= layer1_outputs(4111);
    layer2_outputs(4594) <= (layer1_outputs(1853)) or (layer1_outputs(3746));
    layer2_outputs(4595) <= not(layer1_outputs(3173));
    layer2_outputs(4596) <= not(layer1_outputs(1352));
    layer2_outputs(4597) <= not(layer1_outputs(3332));
    layer2_outputs(4598) <= layer1_outputs(5114);
    layer2_outputs(4599) <= layer1_outputs(4203);
    layer2_outputs(4600) <= (layer1_outputs(1928)) or (layer1_outputs(4580));
    layer2_outputs(4601) <= (layer1_outputs(3882)) xor (layer1_outputs(3677));
    layer2_outputs(4602) <= not(layer1_outputs(214));
    layer2_outputs(4603) <= not(layer1_outputs(4975));
    layer2_outputs(4604) <= not(layer1_outputs(1433));
    layer2_outputs(4605) <= (layer1_outputs(559)) and (layer1_outputs(3718));
    layer2_outputs(4606) <= layer1_outputs(4680);
    layer2_outputs(4607) <= not(layer1_outputs(4020));
    layer2_outputs(4608) <= layer1_outputs(320);
    layer2_outputs(4609) <= (layer1_outputs(1959)) or (layer1_outputs(3424));
    layer2_outputs(4610) <= not((layer1_outputs(4736)) xor (layer1_outputs(1200)));
    layer2_outputs(4611) <= (layer1_outputs(4201)) or (layer1_outputs(849));
    layer2_outputs(4612) <= not(layer1_outputs(2783));
    layer2_outputs(4613) <= layer1_outputs(1480);
    layer2_outputs(4614) <= not(layer1_outputs(3021));
    layer2_outputs(4615) <= not(layer1_outputs(4327));
    layer2_outputs(4616) <= not(layer1_outputs(1251));
    layer2_outputs(4617) <= not((layer1_outputs(4263)) and (layer1_outputs(564)));
    layer2_outputs(4618) <= (layer1_outputs(298)) and (layer1_outputs(4678));
    layer2_outputs(4619) <= (layer1_outputs(2348)) and not (layer1_outputs(1745));
    layer2_outputs(4620) <= (layer1_outputs(2744)) and (layer1_outputs(5013));
    layer2_outputs(4621) <= (layer1_outputs(2662)) and not (layer1_outputs(2373));
    layer2_outputs(4622) <= not(layer1_outputs(3607));
    layer2_outputs(4623) <= not(layer1_outputs(4779));
    layer2_outputs(4624) <= not(layer1_outputs(2086)) or (layer1_outputs(905));
    layer2_outputs(4625) <= (layer1_outputs(4440)) or (layer1_outputs(5087));
    layer2_outputs(4626) <= (layer1_outputs(3610)) xor (layer1_outputs(449));
    layer2_outputs(4627) <= not((layer1_outputs(1118)) and (layer1_outputs(489)));
    layer2_outputs(4628) <= (layer1_outputs(5096)) and not (layer1_outputs(4187));
    layer2_outputs(4629) <= not(layer1_outputs(4176));
    layer2_outputs(4630) <= layer1_outputs(65);
    layer2_outputs(4631) <= not((layer1_outputs(2104)) and (layer1_outputs(1636)));
    layer2_outputs(4632) <= not(layer1_outputs(4218));
    layer2_outputs(4633) <= not((layer1_outputs(4797)) or (layer1_outputs(4860)));
    layer2_outputs(4634) <= (layer1_outputs(977)) or (layer1_outputs(2905));
    layer2_outputs(4635) <= layer1_outputs(4202);
    layer2_outputs(4636) <= not((layer1_outputs(470)) and (layer1_outputs(189)));
    layer2_outputs(4637) <= layer1_outputs(1618);
    layer2_outputs(4638) <= not(layer1_outputs(5006));
    layer2_outputs(4639) <= (layer1_outputs(1056)) or (layer1_outputs(3811));
    layer2_outputs(4640) <= not(layer1_outputs(4518));
    layer2_outputs(4641) <= not((layer1_outputs(1860)) or (layer1_outputs(3707)));
    layer2_outputs(4642) <= not(layer1_outputs(49));
    layer2_outputs(4643) <= layer1_outputs(47);
    layer2_outputs(4644) <= '0';
    layer2_outputs(4645) <= (layer1_outputs(4666)) and not (layer1_outputs(4167));
    layer2_outputs(4646) <= layer1_outputs(365);
    layer2_outputs(4647) <= layer1_outputs(3753);
    layer2_outputs(4648) <= not(layer1_outputs(2317));
    layer2_outputs(4649) <= not(layer1_outputs(4222)) or (layer1_outputs(1723));
    layer2_outputs(4650) <= layer1_outputs(4508);
    layer2_outputs(4651) <= layer1_outputs(3597);
    layer2_outputs(4652) <= (layer1_outputs(2435)) xor (layer1_outputs(3582));
    layer2_outputs(4653) <= (layer1_outputs(2380)) and not (layer1_outputs(944));
    layer2_outputs(4654) <= not(layer1_outputs(1201)) or (layer1_outputs(4042));
    layer2_outputs(4655) <= not(layer1_outputs(5015));
    layer2_outputs(4656) <= not(layer1_outputs(4195)) or (layer1_outputs(2141));
    layer2_outputs(4657) <= layer1_outputs(3618);
    layer2_outputs(4658) <= not(layer1_outputs(3029));
    layer2_outputs(4659) <= not(layer1_outputs(735));
    layer2_outputs(4660) <= layer1_outputs(3229);
    layer2_outputs(4661) <= not(layer1_outputs(267)) or (layer1_outputs(226));
    layer2_outputs(4662) <= layer1_outputs(602);
    layer2_outputs(4663) <= layer1_outputs(1765);
    layer2_outputs(4664) <= layer1_outputs(2395);
    layer2_outputs(4665) <= layer1_outputs(4045);
    layer2_outputs(4666) <= not((layer1_outputs(3073)) or (layer1_outputs(810)));
    layer2_outputs(4667) <= not((layer1_outputs(2080)) and (layer1_outputs(766)));
    layer2_outputs(4668) <= (layer1_outputs(3586)) and not (layer1_outputs(2087));
    layer2_outputs(4669) <= layer1_outputs(3616);
    layer2_outputs(4670) <= not(layer1_outputs(310));
    layer2_outputs(4671) <= not((layer1_outputs(443)) and (layer1_outputs(4140)));
    layer2_outputs(4672) <= layer1_outputs(1465);
    layer2_outputs(4673) <= (layer1_outputs(2865)) xor (layer1_outputs(4561));
    layer2_outputs(4674) <= layer1_outputs(4870);
    layer2_outputs(4675) <= layer1_outputs(1697);
    layer2_outputs(4676) <= not(layer1_outputs(2327)) or (layer1_outputs(861));
    layer2_outputs(4677) <= not(layer1_outputs(2402));
    layer2_outputs(4678) <= not((layer1_outputs(4818)) or (layer1_outputs(1074)));
    layer2_outputs(4679) <= not(layer1_outputs(3303));
    layer2_outputs(4680) <= layer1_outputs(3592);
    layer2_outputs(4681) <= layer1_outputs(3511);
    layer2_outputs(4682) <= (layer1_outputs(1883)) and not (layer1_outputs(4216));
    layer2_outputs(4683) <= not((layer1_outputs(1138)) or (layer1_outputs(331)));
    layer2_outputs(4684) <= (layer1_outputs(71)) or (layer1_outputs(4880));
    layer2_outputs(4685) <= layer1_outputs(1985);
    layer2_outputs(4686) <= not(layer1_outputs(2668)) or (layer1_outputs(501));
    layer2_outputs(4687) <= (layer1_outputs(1721)) or (layer1_outputs(536));
    layer2_outputs(4688) <= layer1_outputs(1791);
    layer2_outputs(4689) <= not((layer1_outputs(4364)) xor (layer1_outputs(4798)));
    layer2_outputs(4690) <= (layer1_outputs(2159)) and not (layer1_outputs(1572));
    layer2_outputs(4691) <= not(layer1_outputs(4772));
    layer2_outputs(4692) <= layer1_outputs(3267);
    layer2_outputs(4693) <= layer1_outputs(160);
    layer2_outputs(4694) <= (layer1_outputs(4761)) xor (layer1_outputs(1890));
    layer2_outputs(4695) <= (layer1_outputs(1177)) and not (layer1_outputs(957));
    layer2_outputs(4696) <= (layer1_outputs(958)) and (layer1_outputs(3070));
    layer2_outputs(4697) <= not(layer1_outputs(2156));
    layer2_outputs(4698) <= (layer1_outputs(4730)) and not (layer1_outputs(752));
    layer2_outputs(4699) <= layer1_outputs(1142);
    layer2_outputs(4700) <= (layer1_outputs(3743)) xor (layer1_outputs(2093));
    layer2_outputs(4701) <= not((layer1_outputs(1527)) and (layer1_outputs(2567)));
    layer2_outputs(4702) <= not(layer1_outputs(3277));
    layer2_outputs(4703) <= not(layer1_outputs(1376));
    layer2_outputs(4704) <= not(layer1_outputs(359));
    layer2_outputs(4705) <= layer1_outputs(3982);
    layer2_outputs(4706) <= layer1_outputs(166);
    layer2_outputs(4707) <= not((layer1_outputs(1359)) or (layer1_outputs(192)));
    layer2_outputs(4708) <= layer1_outputs(4001);
    layer2_outputs(4709) <= (layer1_outputs(481)) or (layer1_outputs(3391));
    layer2_outputs(4710) <= not(layer1_outputs(1281)) or (layer1_outputs(4148));
    layer2_outputs(4711) <= not(layer1_outputs(3135));
    layer2_outputs(4712) <= not(layer1_outputs(1336)) or (layer1_outputs(3123));
    layer2_outputs(4713) <= (layer1_outputs(4656)) and not (layer1_outputs(2551));
    layer2_outputs(4714) <= '1';
    layer2_outputs(4715) <= (layer1_outputs(467)) and not (layer1_outputs(672));
    layer2_outputs(4716) <= (layer1_outputs(2399)) and not (layer1_outputs(1962));
    layer2_outputs(4717) <= layer1_outputs(4701);
    layer2_outputs(4718) <= not(layer1_outputs(16)) or (layer1_outputs(5099));
    layer2_outputs(4719) <= (layer1_outputs(2099)) and not (layer1_outputs(2918));
    layer2_outputs(4720) <= layer1_outputs(3244);
    layer2_outputs(4721) <= (layer1_outputs(3257)) and not (layer1_outputs(247));
    layer2_outputs(4722) <= (layer1_outputs(707)) and not (layer1_outputs(1512));
    layer2_outputs(4723) <= not(layer1_outputs(2820));
    layer2_outputs(4724) <= not(layer1_outputs(3045)) or (layer1_outputs(3726));
    layer2_outputs(4725) <= (layer1_outputs(1826)) and not (layer1_outputs(4811));
    layer2_outputs(4726) <= not(layer1_outputs(3977));
    layer2_outputs(4727) <= (layer1_outputs(3998)) and not (layer1_outputs(2292));
    layer2_outputs(4728) <= not(layer1_outputs(1277)) or (layer1_outputs(2720));
    layer2_outputs(4729) <= not(layer1_outputs(4438)) or (layer1_outputs(2039));
    layer2_outputs(4730) <= not(layer1_outputs(525));
    layer2_outputs(4731) <= not(layer1_outputs(369)) or (layer1_outputs(1251));
    layer2_outputs(4732) <= not((layer1_outputs(3584)) xor (layer1_outputs(907)));
    layer2_outputs(4733) <= not(layer1_outputs(1471));
    layer2_outputs(4734) <= layer1_outputs(3291);
    layer2_outputs(4735) <= not(layer1_outputs(2226)) or (layer1_outputs(3945));
    layer2_outputs(4736) <= not(layer1_outputs(2037)) or (layer1_outputs(2789));
    layer2_outputs(4737) <= (layer1_outputs(1613)) xor (layer1_outputs(3881));
    layer2_outputs(4738) <= layer1_outputs(2101);
    layer2_outputs(4739) <= layer1_outputs(2383);
    layer2_outputs(4740) <= not(layer1_outputs(2813));
    layer2_outputs(4741) <= (layer1_outputs(4479)) and not (layer1_outputs(490));
    layer2_outputs(4742) <= (layer1_outputs(4965)) or (layer1_outputs(3717));
    layer2_outputs(4743) <= not(layer1_outputs(4463));
    layer2_outputs(4744) <= '1';
    layer2_outputs(4745) <= not(layer1_outputs(3822));
    layer2_outputs(4746) <= (layer1_outputs(4348)) and not (layer1_outputs(437));
    layer2_outputs(4747) <= layer1_outputs(1796);
    layer2_outputs(4748) <= layer1_outputs(912);
    layer2_outputs(4749) <= (layer1_outputs(1459)) or (layer1_outputs(191));
    layer2_outputs(4750) <= layer1_outputs(2211);
    layer2_outputs(4751) <= layer1_outputs(4200);
    layer2_outputs(4752) <= not((layer1_outputs(873)) and (layer1_outputs(4637)));
    layer2_outputs(4753) <= not((layer1_outputs(1913)) and (layer1_outputs(2727)));
    layer2_outputs(4754) <= (layer1_outputs(4881)) and not (layer1_outputs(583));
    layer2_outputs(4755) <= not(layer1_outputs(2213));
    layer2_outputs(4756) <= not((layer1_outputs(2762)) and (layer1_outputs(4314)));
    layer2_outputs(4757) <= (layer1_outputs(1369)) xor (layer1_outputs(4589));
    layer2_outputs(4758) <= (layer1_outputs(2757)) and not (layer1_outputs(3364));
    layer2_outputs(4759) <= (layer1_outputs(3643)) and not (layer1_outputs(2288));
    layer2_outputs(4760) <= (layer1_outputs(2275)) xor (layer1_outputs(2247));
    layer2_outputs(4761) <= not(layer1_outputs(1817));
    layer2_outputs(4762) <= layer1_outputs(2807);
    layer2_outputs(4763) <= layer1_outputs(4461);
    layer2_outputs(4764) <= not((layer1_outputs(771)) xor (layer1_outputs(4135)));
    layer2_outputs(4765) <= (layer1_outputs(4129)) or (layer1_outputs(2879));
    layer2_outputs(4766) <= layer1_outputs(421);
    layer2_outputs(4767) <= layer1_outputs(3937);
    layer2_outputs(4768) <= not(layer1_outputs(1399));
    layer2_outputs(4769) <= layer1_outputs(3144);
    layer2_outputs(4770) <= (layer1_outputs(3764)) xor (layer1_outputs(3121));
    layer2_outputs(4771) <= layer1_outputs(3313);
    layer2_outputs(4772) <= (layer1_outputs(4121)) or (layer1_outputs(4612));
    layer2_outputs(4773) <= not(layer1_outputs(1205));
    layer2_outputs(4774) <= not((layer1_outputs(3422)) xor (layer1_outputs(655)));
    layer2_outputs(4775) <= not((layer1_outputs(1261)) or (layer1_outputs(4511)));
    layer2_outputs(4776) <= (layer1_outputs(3991)) and (layer1_outputs(1154));
    layer2_outputs(4777) <= layer1_outputs(1162);
    layer2_outputs(4778) <= layer1_outputs(2706);
    layer2_outputs(4779) <= not(layer1_outputs(1158));
    layer2_outputs(4780) <= not(layer1_outputs(2984)) or (layer1_outputs(4397));
    layer2_outputs(4781) <= (layer1_outputs(401)) and (layer1_outputs(4758));
    layer2_outputs(4782) <= not(layer1_outputs(4945));
    layer2_outputs(4783) <= '1';
    layer2_outputs(4784) <= layer1_outputs(376);
    layer2_outputs(4785) <= (layer1_outputs(2323)) and (layer1_outputs(2678));
    layer2_outputs(4786) <= not(layer1_outputs(4470)) or (layer1_outputs(4030));
    layer2_outputs(4787) <= (layer1_outputs(3120)) and not (layer1_outputs(2629));
    layer2_outputs(4788) <= not(layer1_outputs(3504)) or (layer1_outputs(1615));
    layer2_outputs(4789) <= not(layer1_outputs(2223)) or (layer1_outputs(4406));
    layer2_outputs(4790) <= (layer1_outputs(477)) and not (layer1_outputs(2952));
    layer2_outputs(4791) <= not((layer1_outputs(1108)) and (layer1_outputs(3589)));
    layer2_outputs(4792) <= layer1_outputs(637);
    layer2_outputs(4793) <= not((layer1_outputs(4563)) or (layer1_outputs(4489)));
    layer2_outputs(4794) <= layer1_outputs(3868);
    layer2_outputs(4795) <= layer1_outputs(803);
    layer2_outputs(4796) <= (layer1_outputs(240)) xor (layer1_outputs(3519));
    layer2_outputs(4797) <= (layer1_outputs(3111)) or (layer1_outputs(551));
    layer2_outputs(4798) <= not(layer1_outputs(1732)) or (layer1_outputs(3275));
    layer2_outputs(4799) <= not(layer1_outputs(4492));
    layer2_outputs(4800) <= not(layer1_outputs(5002));
    layer2_outputs(4801) <= (layer1_outputs(393)) or (layer1_outputs(1310));
    layer2_outputs(4802) <= layer1_outputs(743);
    layer2_outputs(4803) <= '1';
    layer2_outputs(4804) <= (layer1_outputs(3044)) and (layer1_outputs(2205));
    layer2_outputs(4805) <= (layer1_outputs(3418)) and (layer1_outputs(3548));
    layer2_outputs(4806) <= layer1_outputs(4822);
    layer2_outputs(4807) <= (layer1_outputs(3361)) xor (layer1_outputs(2015));
    layer2_outputs(4808) <= layer1_outputs(5051);
    layer2_outputs(4809) <= (layer1_outputs(3509)) and (layer1_outputs(1592));
    layer2_outputs(4810) <= (layer1_outputs(1181)) and not (layer1_outputs(4547));
    layer2_outputs(4811) <= not(layer1_outputs(3825));
    layer2_outputs(4812) <= not((layer1_outputs(3473)) xor (layer1_outputs(2620)));
    layer2_outputs(4813) <= (layer1_outputs(3597)) xor (layer1_outputs(1367));
    layer2_outputs(4814) <= not(layer1_outputs(5019));
    layer2_outputs(4815) <= not(layer1_outputs(2628));
    layer2_outputs(4816) <= not(layer1_outputs(5102));
    layer2_outputs(4817) <= layer1_outputs(2478);
    layer2_outputs(4818) <= layer1_outputs(1319);
    layer2_outputs(4819) <= not(layer1_outputs(837));
    layer2_outputs(4820) <= layer1_outputs(2961);
    layer2_outputs(4821) <= (layer1_outputs(2307)) xor (layer1_outputs(2474));
    layer2_outputs(4822) <= not(layer1_outputs(2718));
    layer2_outputs(4823) <= not(layer1_outputs(3219)) or (layer1_outputs(816));
    layer2_outputs(4824) <= not(layer1_outputs(3132));
    layer2_outputs(4825) <= '0';
    layer2_outputs(4826) <= '0';
    layer2_outputs(4827) <= layer1_outputs(3610);
    layer2_outputs(4828) <= not(layer1_outputs(2354));
    layer2_outputs(4829) <= not(layer1_outputs(4690)) or (layer1_outputs(2966));
    layer2_outputs(4830) <= not(layer1_outputs(2899)) or (layer1_outputs(4860));
    layer2_outputs(4831) <= layer1_outputs(1449);
    layer2_outputs(4832) <= not((layer1_outputs(4707)) or (layer1_outputs(3009)));
    layer2_outputs(4833) <= not(layer1_outputs(1757)) or (layer1_outputs(331));
    layer2_outputs(4834) <= not(layer1_outputs(1764));
    layer2_outputs(4835) <= '0';
    layer2_outputs(4836) <= not(layer1_outputs(2259)) or (layer1_outputs(3174));
    layer2_outputs(4837) <= (layer1_outputs(2024)) xor (layer1_outputs(4847));
    layer2_outputs(4838) <= layer1_outputs(794);
    layer2_outputs(4839) <= layer1_outputs(2764);
    layer2_outputs(4840) <= layer1_outputs(1333);
    layer2_outputs(4841) <= (layer1_outputs(1532)) and not (layer1_outputs(2892));
    layer2_outputs(4842) <= layer1_outputs(2760);
    layer2_outputs(4843) <= not(layer1_outputs(1905));
    layer2_outputs(4844) <= not(layer1_outputs(4769));
    layer2_outputs(4845) <= not(layer1_outputs(2847));
    layer2_outputs(4846) <= layer1_outputs(2621);
    layer2_outputs(4847) <= layer1_outputs(4198);
    layer2_outputs(4848) <= not(layer1_outputs(728));
    layer2_outputs(4849) <= layer1_outputs(17);
    layer2_outputs(4850) <= (layer1_outputs(2486)) and not (layer1_outputs(157));
    layer2_outputs(4851) <= (layer1_outputs(1847)) and not (layer1_outputs(1040));
    layer2_outputs(4852) <= layer1_outputs(3279);
    layer2_outputs(4853) <= not(layer1_outputs(1856));
    layer2_outputs(4854) <= layer1_outputs(4597);
    layer2_outputs(4855) <= layer1_outputs(4612);
    layer2_outputs(4856) <= not(layer1_outputs(1152));
    layer2_outputs(4857) <= not(layer1_outputs(1633));
    layer2_outputs(4858) <= layer1_outputs(4333);
    layer2_outputs(4859) <= not(layer1_outputs(3872)) or (layer1_outputs(1264));
    layer2_outputs(4860) <= layer1_outputs(4214);
    layer2_outputs(4861) <= not(layer1_outputs(1717));
    layer2_outputs(4862) <= not(layer1_outputs(809)) or (layer1_outputs(4537));
    layer2_outputs(4863) <= layer1_outputs(982);
    layer2_outputs(4864) <= not(layer1_outputs(2356));
    layer2_outputs(4865) <= not((layer1_outputs(3852)) xor (layer1_outputs(1511)));
    layer2_outputs(4866) <= (layer1_outputs(2544)) or (layer1_outputs(4949));
    layer2_outputs(4867) <= not((layer1_outputs(4185)) or (layer1_outputs(4521)));
    layer2_outputs(4868) <= (layer1_outputs(4740)) and (layer1_outputs(4888));
    layer2_outputs(4869) <= layer1_outputs(1757);
    layer2_outputs(4870) <= layer1_outputs(272);
    layer2_outputs(4871) <= not(layer1_outputs(1870));
    layer2_outputs(4872) <= not(layer1_outputs(3990)) or (layer1_outputs(3052));
    layer2_outputs(4873) <= layer1_outputs(4103);
    layer2_outputs(4874) <= layer1_outputs(4007);
    layer2_outputs(4875) <= layer1_outputs(3520);
    layer2_outputs(4876) <= not(layer1_outputs(317));
    layer2_outputs(4877) <= not(layer1_outputs(2869));
    layer2_outputs(4878) <= (layer1_outputs(2469)) and not (layer1_outputs(4794));
    layer2_outputs(4879) <= (layer1_outputs(2687)) and not (layer1_outputs(1081));
    layer2_outputs(4880) <= not(layer1_outputs(3718));
    layer2_outputs(4881) <= not((layer1_outputs(3446)) and (layer1_outputs(3611)));
    layer2_outputs(4882) <= (layer1_outputs(4260)) and not (layer1_outputs(4024));
    layer2_outputs(4883) <= not((layer1_outputs(1615)) or (layer1_outputs(1056)));
    layer2_outputs(4884) <= not(layer1_outputs(2484));
    layer2_outputs(4885) <= not(layer1_outputs(4132)) or (layer1_outputs(4460));
    layer2_outputs(4886) <= not(layer1_outputs(5007)) or (layer1_outputs(876));
    layer2_outputs(4887) <= not(layer1_outputs(2125));
    layer2_outputs(4888) <= layer1_outputs(3499);
    layer2_outputs(4889) <= (layer1_outputs(217)) and not (layer1_outputs(2407));
    layer2_outputs(4890) <= not((layer1_outputs(3031)) and (layer1_outputs(2923)));
    layer2_outputs(4891) <= not(layer1_outputs(4041));
    layer2_outputs(4892) <= not(layer1_outputs(3023)) or (layer1_outputs(5020));
    layer2_outputs(4893) <= not(layer1_outputs(1297));
    layer2_outputs(4894) <= layer1_outputs(2345);
    layer2_outputs(4895) <= not(layer1_outputs(234));
    layer2_outputs(4896) <= layer1_outputs(42);
    layer2_outputs(4897) <= not(layer1_outputs(2728)) or (layer1_outputs(1041));
    layer2_outputs(4898) <= (layer1_outputs(5105)) xor (layer1_outputs(562));
    layer2_outputs(4899) <= '1';
    layer2_outputs(4900) <= not((layer1_outputs(2622)) xor (layer1_outputs(136)));
    layer2_outputs(4901) <= not((layer1_outputs(4611)) and (layer1_outputs(1001)));
    layer2_outputs(4902) <= (layer1_outputs(569)) and (layer1_outputs(2018));
    layer2_outputs(4903) <= not(layer1_outputs(2416)) or (layer1_outputs(575));
    layer2_outputs(4904) <= (layer1_outputs(480)) and not (layer1_outputs(5091));
    layer2_outputs(4905) <= (layer1_outputs(2261)) and not (layer1_outputs(4685));
    layer2_outputs(4906) <= not(layer1_outputs(2185)) or (layer1_outputs(112));
    layer2_outputs(4907) <= layer1_outputs(2027);
    layer2_outputs(4908) <= not((layer1_outputs(461)) and (layer1_outputs(1316)));
    layer2_outputs(4909) <= not(layer1_outputs(408));
    layer2_outputs(4910) <= (layer1_outputs(3749)) and not (layer1_outputs(1768));
    layer2_outputs(4911) <= not(layer1_outputs(4166));
    layer2_outputs(4912) <= not(layer1_outputs(4493));
    layer2_outputs(4913) <= layer1_outputs(4900);
    layer2_outputs(4914) <= not((layer1_outputs(2120)) and (layer1_outputs(3262)));
    layer2_outputs(4915) <= not((layer1_outputs(4349)) and (layer1_outputs(734)));
    layer2_outputs(4916) <= layer1_outputs(4120);
    layer2_outputs(4917) <= not(layer1_outputs(1564));
    layer2_outputs(4918) <= (layer1_outputs(357)) and (layer1_outputs(3640));
    layer2_outputs(4919) <= not(layer1_outputs(2405));
    layer2_outputs(4920) <= not(layer1_outputs(4278));
    layer2_outputs(4921) <= not(layer1_outputs(2313));
    layer2_outputs(4922) <= not(layer1_outputs(3289)) or (layer1_outputs(2050));
    layer2_outputs(4923) <= not((layer1_outputs(2504)) and (layer1_outputs(4100)));
    layer2_outputs(4924) <= layer1_outputs(4501);
    layer2_outputs(4925) <= not((layer1_outputs(3836)) xor (layer1_outputs(3381)));
    layer2_outputs(4926) <= layer1_outputs(1668);
    layer2_outputs(4927) <= not(layer1_outputs(3338));
    layer2_outputs(4928) <= not(layer1_outputs(1174));
    layer2_outputs(4929) <= not((layer1_outputs(4236)) xor (layer1_outputs(963)));
    layer2_outputs(4930) <= (layer1_outputs(1734)) and not (layer1_outputs(4868));
    layer2_outputs(4931) <= layer1_outputs(4399);
    layer2_outputs(4932) <= layer1_outputs(5001);
    layer2_outputs(4933) <= not(layer1_outputs(2245));
    layer2_outputs(4934) <= not(layer1_outputs(1086));
    layer2_outputs(4935) <= (layer1_outputs(3064)) and not (layer1_outputs(1375));
    layer2_outputs(4936) <= (layer1_outputs(933)) and (layer1_outputs(1227));
    layer2_outputs(4937) <= not(layer1_outputs(4648));
    layer2_outputs(4938) <= layer1_outputs(4209);
    layer2_outputs(4939) <= not(layer1_outputs(334)) or (layer1_outputs(1918));
    layer2_outputs(4940) <= layer1_outputs(496);
    layer2_outputs(4941) <= not((layer1_outputs(4941)) and (layer1_outputs(4303)));
    layer2_outputs(4942) <= not(layer1_outputs(5094));
    layer2_outputs(4943) <= layer1_outputs(1620);
    layer2_outputs(4944) <= not(layer1_outputs(2610)) or (layer1_outputs(3209));
    layer2_outputs(4945) <= not(layer1_outputs(1586));
    layer2_outputs(4946) <= (layer1_outputs(3570)) or (layer1_outputs(1744));
    layer2_outputs(4947) <= (layer1_outputs(4633)) and not (layer1_outputs(2329));
    layer2_outputs(4948) <= layer1_outputs(1495);
    layer2_outputs(4949) <= layer1_outputs(1117);
    layer2_outputs(4950) <= not((layer1_outputs(1084)) xor (layer1_outputs(2244)));
    layer2_outputs(4951) <= (layer1_outputs(381)) and not (layer1_outputs(519));
    layer2_outputs(4952) <= layer1_outputs(2243);
    layer2_outputs(4953) <= not(layer1_outputs(205));
    layer2_outputs(4954) <= (layer1_outputs(4537)) and (layer1_outputs(3401));
    layer2_outputs(4955) <= layer1_outputs(2061);
    layer2_outputs(4956) <= not(layer1_outputs(3742)) or (layer1_outputs(772));
    layer2_outputs(4957) <= not(layer1_outputs(904));
    layer2_outputs(4958) <= not(layer1_outputs(2564));
    layer2_outputs(4959) <= not(layer1_outputs(3043)) or (layer1_outputs(3240));
    layer2_outputs(4960) <= not(layer1_outputs(2369)) or (layer1_outputs(133));
    layer2_outputs(4961) <= not((layer1_outputs(4802)) and (layer1_outputs(5055)));
    layer2_outputs(4962) <= (layer1_outputs(4088)) or (layer1_outputs(1694));
    layer2_outputs(4963) <= (layer1_outputs(23)) and not (layer1_outputs(2448));
    layer2_outputs(4964) <= layer1_outputs(343);
    layer2_outputs(4965) <= (layer1_outputs(400)) or (layer1_outputs(3416));
    layer2_outputs(4966) <= not(layer1_outputs(2359));
    layer2_outputs(4967) <= (layer1_outputs(959)) and not (layer1_outputs(4114));
    layer2_outputs(4968) <= layer1_outputs(2274);
    layer2_outputs(4969) <= (layer1_outputs(286)) and not (layer1_outputs(2081));
    layer2_outputs(4970) <= not((layer1_outputs(2572)) and (layer1_outputs(1715)));
    layer2_outputs(4971) <= not(layer1_outputs(2133));
    layer2_outputs(4972) <= layer1_outputs(4261);
    layer2_outputs(4973) <= layer1_outputs(3038);
    layer2_outputs(4974) <= not(layer1_outputs(644));
    layer2_outputs(4975) <= (layer1_outputs(1710)) and (layer1_outputs(4169));
    layer2_outputs(4976) <= not((layer1_outputs(4544)) or (layer1_outputs(3780)));
    layer2_outputs(4977) <= layer1_outputs(2440);
    layer2_outputs(4978) <= '1';
    layer2_outputs(4979) <= not(layer1_outputs(1192));
    layer2_outputs(4980) <= not((layer1_outputs(3808)) and (layer1_outputs(1398)));
    layer2_outputs(4981) <= not(layer1_outputs(2830)) or (layer1_outputs(3817));
    layer2_outputs(4982) <= not((layer1_outputs(1416)) or (layer1_outputs(2120)));
    layer2_outputs(4983) <= not(layer1_outputs(4498));
    layer2_outputs(4984) <= (layer1_outputs(3586)) and not (layer1_outputs(2450));
    layer2_outputs(4985) <= not((layer1_outputs(2124)) and (layer1_outputs(4764)));
    layer2_outputs(4986) <= not(layer1_outputs(1609));
    layer2_outputs(4987) <= not(layer1_outputs(1988));
    layer2_outputs(4988) <= (layer1_outputs(3843)) and not (layer1_outputs(901));
    layer2_outputs(4989) <= layer1_outputs(131);
    layer2_outputs(4990) <= (layer1_outputs(1621)) or (layer1_outputs(3772));
    layer2_outputs(4991) <= layer1_outputs(4256);
    layer2_outputs(4992) <= (layer1_outputs(3258)) and (layer1_outputs(1948));
    layer2_outputs(4993) <= not(layer1_outputs(3311));
    layer2_outputs(4994) <= not(layer1_outputs(2667));
    layer2_outputs(4995) <= layer1_outputs(3246);
    layer2_outputs(4996) <= '1';
    layer2_outputs(4997) <= not(layer1_outputs(281));
    layer2_outputs(4998) <= not(layer1_outputs(4753));
    layer2_outputs(4999) <= not(layer1_outputs(4351));
    layer2_outputs(5000) <= (layer1_outputs(4057)) and not (layer1_outputs(892));
    layer2_outputs(5001) <= not(layer1_outputs(4108));
    layer2_outputs(5002) <= (layer1_outputs(342)) and not (layer1_outputs(3297));
    layer2_outputs(5003) <= not(layer1_outputs(4133));
    layer2_outputs(5004) <= layer1_outputs(934);
    layer2_outputs(5005) <= (layer1_outputs(1651)) and (layer1_outputs(4452));
    layer2_outputs(5006) <= not(layer1_outputs(1404));
    layer2_outputs(5007) <= not(layer1_outputs(296));
    layer2_outputs(5008) <= not(layer1_outputs(4357));
    layer2_outputs(5009) <= not(layer1_outputs(689));
    layer2_outputs(5010) <= (layer1_outputs(2935)) xor (layer1_outputs(1617));
    layer2_outputs(5011) <= not(layer1_outputs(1046)) or (layer1_outputs(4012));
    layer2_outputs(5012) <= (layer1_outputs(2676)) or (layer1_outputs(25));
    layer2_outputs(5013) <= not((layer1_outputs(3606)) and (layer1_outputs(3934)));
    layer2_outputs(5014) <= not(layer1_outputs(2966));
    layer2_outputs(5015) <= '1';
    layer2_outputs(5016) <= layer1_outputs(561);
    layer2_outputs(5017) <= not(layer1_outputs(3169)) or (layer1_outputs(943));
    layer2_outputs(5018) <= (layer1_outputs(915)) and not (layer1_outputs(4193));
    layer2_outputs(5019) <= not(layer1_outputs(3618)) or (layer1_outputs(85));
    layer2_outputs(5020) <= not(layer1_outputs(842)) or (layer1_outputs(3175));
    layer2_outputs(5021) <= layer1_outputs(2715);
    layer2_outputs(5022) <= layer1_outputs(3601);
    layer2_outputs(5023) <= layer1_outputs(4557);
    layer2_outputs(5024) <= not(layer1_outputs(3677));
    layer2_outputs(5025) <= not((layer1_outputs(3869)) or (layer1_outputs(3463)));
    layer2_outputs(5026) <= layer1_outputs(1996);
    layer2_outputs(5027) <= (layer1_outputs(1363)) or (layer1_outputs(3412));
    layer2_outputs(5028) <= (layer1_outputs(4777)) or (layer1_outputs(604));
    layer2_outputs(5029) <= (layer1_outputs(4825)) and not (layer1_outputs(1073));
    layer2_outputs(5030) <= (layer1_outputs(1140)) or (layer1_outputs(2688));
    layer2_outputs(5031) <= not(layer1_outputs(860)) or (layer1_outputs(4017));
    layer2_outputs(5032) <= not((layer1_outputs(3915)) or (layer1_outputs(2703)));
    layer2_outputs(5033) <= (layer1_outputs(1178)) and (layer1_outputs(932));
    layer2_outputs(5034) <= not(layer1_outputs(3788));
    layer2_outputs(5035) <= (layer1_outputs(940)) and (layer1_outputs(3659));
    layer2_outputs(5036) <= layer1_outputs(3195);
    layer2_outputs(5037) <= (layer1_outputs(852)) xor (layer1_outputs(1878));
    layer2_outputs(5038) <= not(layer1_outputs(2040)) or (layer1_outputs(2325));
    layer2_outputs(5039) <= layer1_outputs(2884);
    layer2_outputs(5040) <= layer1_outputs(4743);
    layer2_outputs(5041) <= (layer1_outputs(598)) and (layer1_outputs(913));
    layer2_outputs(5042) <= not(layer1_outputs(442)) or (layer1_outputs(2792));
    layer2_outputs(5043) <= layer1_outputs(4754);
    layer2_outputs(5044) <= (layer1_outputs(505)) xor (layer1_outputs(1478));
    layer2_outputs(5045) <= not(layer1_outputs(1500));
    layer2_outputs(5046) <= '0';
    layer2_outputs(5047) <= layer1_outputs(3594);
    layer2_outputs(5048) <= not(layer1_outputs(4458));
    layer2_outputs(5049) <= not((layer1_outputs(436)) xor (layer1_outputs(3512)));
    layer2_outputs(5050) <= layer1_outputs(1173);
    layer2_outputs(5051) <= not(layer1_outputs(1900));
    layer2_outputs(5052) <= layer1_outputs(199);
    layer2_outputs(5053) <= not(layer1_outputs(3322));
    layer2_outputs(5054) <= layer1_outputs(1654);
    layer2_outputs(5055) <= not(layer1_outputs(840)) or (layer1_outputs(3021));
    layer2_outputs(5056) <= not(layer1_outputs(3270)) or (layer1_outputs(561));
    layer2_outputs(5057) <= (layer1_outputs(3676)) and not (layer1_outputs(793));
    layer2_outputs(5058) <= not((layer1_outputs(1220)) or (layer1_outputs(4538)));
    layer2_outputs(5059) <= layer1_outputs(1876);
    layer2_outputs(5060) <= layer1_outputs(2341);
    layer2_outputs(5061) <= (layer1_outputs(2933)) and not (layer1_outputs(4129));
    layer2_outputs(5062) <= '1';
    layer2_outputs(5063) <= not(layer1_outputs(1554));
    layer2_outputs(5064) <= not(layer1_outputs(3720));
    layer2_outputs(5065) <= layer1_outputs(309);
    layer2_outputs(5066) <= not((layer1_outputs(4002)) and (layer1_outputs(4194)));
    layer2_outputs(5067) <= layer1_outputs(825);
    layer2_outputs(5068) <= (layer1_outputs(1655)) xor (layer1_outputs(4411));
    layer2_outputs(5069) <= (layer1_outputs(2855)) or (layer1_outputs(3667));
    layer2_outputs(5070) <= layer1_outputs(1063);
    layer2_outputs(5071) <= (layer1_outputs(3419)) and not (layer1_outputs(2875));
    layer2_outputs(5072) <= not((layer1_outputs(53)) or (layer1_outputs(463)));
    layer2_outputs(5073) <= (layer1_outputs(866)) and not (layer1_outputs(3919));
    layer2_outputs(5074) <= (layer1_outputs(1983)) and (layer1_outputs(2361));
    layer2_outputs(5075) <= (layer1_outputs(248)) and not (layer1_outputs(4823));
    layer2_outputs(5076) <= (layer1_outputs(4471)) and not (layer1_outputs(285));
    layer2_outputs(5077) <= layer1_outputs(2458);
    layer2_outputs(5078) <= (layer1_outputs(1231)) or (layer1_outputs(4500));
    layer2_outputs(5079) <= not(layer1_outputs(3149));
    layer2_outputs(5080) <= not(layer1_outputs(2952));
    layer2_outputs(5081) <= not(layer1_outputs(540));
    layer2_outputs(5082) <= layer1_outputs(2491);
    layer2_outputs(5083) <= (layer1_outputs(3773)) and not (layer1_outputs(2363));
    layer2_outputs(5084) <= not(layer1_outputs(2222));
    layer2_outputs(5085) <= not(layer1_outputs(3069));
    layer2_outputs(5086) <= (layer1_outputs(964)) and not (layer1_outputs(1920));
    layer2_outputs(5087) <= layer1_outputs(3849);
    layer2_outputs(5088) <= layer1_outputs(2526);
    layer2_outputs(5089) <= layer1_outputs(2511);
    layer2_outputs(5090) <= not(layer1_outputs(4101));
    layer2_outputs(5091) <= (layer1_outputs(1464)) and (layer1_outputs(451));
    layer2_outputs(5092) <= (layer1_outputs(3147)) or (layer1_outputs(3971));
    layer2_outputs(5093) <= not(layer1_outputs(2079)) or (layer1_outputs(596));
    layer2_outputs(5094) <= not((layer1_outputs(956)) or (layer1_outputs(5087)));
    layer2_outputs(5095) <= (layer1_outputs(4793)) and not (layer1_outputs(3503));
    layer2_outputs(5096) <= not(layer1_outputs(838));
    layer2_outputs(5097) <= not(layer1_outputs(2782)) or (layer1_outputs(1398));
    layer2_outputs(5098) <= layer1_outputs(897);
    layer2_outputs(5099) <= layer1_outputs(175);
    layer2_outputs(5100) <= layer1_outputs(2427);
    layer2_outputs(5101) <= not(layer1_outputs(1945)) or (layer1_outputs(4299));
    layer2_outputs(5102) <= layer1_outputs(2600);
    layer2_outputs(5103) <= not(layer1_outputs(3312));
    layer2_outputs(5104) <= not(layer1_outputs(2268));
    layer2_outputs(5105) <= (layer1_outputs(1949)) or (layer1_outputs(3585));
    layer2_outputs(5106) <= not((layer1_outputs(3133)) or (layer1_outputs(4977)));
    layer2_outputs(5107) <= not((layer1_outputs(1198)) or (layer1_outputs(2781)));
    layer2_outputs(5108) <= not(layer1_outputs(3214));
    layer2_outputs(5109) <= '0';
    layer2_outputs(5110) <= not((layer1_outputs(4864)) or (layer1_outputs(4291)));
    layer2_outputs(5111) <= (layer1_outputs(3563)) and not (layer1_outputs(4843));
    layer2_outputs(5112) <= (layer1_outputs(2170)) and not (layer1_outputs(1323));
    layer2_outputs(5113) <= layer1_outputs(857);
    layer2_outputs(5114) <= (layer1_outputs(3186)) or (layer1_outputs(4354));
    layer2_outputs(5115) <= layer1_outputs(2576);
    layer2_outputs(5116) <= (layer1_outputs(2701)) or (layer1_outputs(4427));
    layer2_outputs(5117) <= '1';
    layer2_outputs(5118) <= (layer1_outputs(4636)) or (layer1_outputs(656));
    layer2_outputs(5119) <= not(layer1_outputs(3614));
    outputs(0) <= layer2_outputs(3578);
    outputs(1) <= (layer2_outputs(3377)) and (layer2_outputs(4976));
    outputs(2) <= not(layer2_outputs(4593));
    outputs(3) <= layer2_outputs(538);
    outputs(4) <= layer2_outputs(1322);
    outputs(5) <= not((layer2_outputs(938)) or (layer2_outputs(968)));
    outputs(6) <= (layer2_outputs(983)) and not (layer2_outputs(917));
    outputs(7) <= not(layer2_outputs(2769));
    outputs(8) <= layer2_outputs(2396);
    outputs(9) <= (layer2_outputs(753)) and (layer2_outputs(3508));
    outputs(10) <= not(layer2_outputs(4663));
    outputs(11) <= layer2_outputs(3506);
    outputs(12) <= not(layer2_outputs(642));
    outputs(13) <= not(layer2_outputs(3692));
    outputs(14) <= (layer2_outputs(256)) and (layer2_outputs(1658));
    outputs(15) <= (layer2_outputs(1000)) xor (layer2_outputs(3276));
    outputs(16) <= layer2_outputs(4475);
    outputs(17) <= (layer2_outputs(3154)) xor (layer2_outputs(2968));
    outputs(18) <= not(layer2_outputs(4474));
    outputs(19) <= not(layer2_outputs(3299));
    outputs(20) <= (layer2_outputs(685)) and not (layer2_outputs(4943));
    outputs(21) <= not(layer2_outputs(4909));
    outputs(22) <= not(layer2_outputs(4487));
    outputs(23) <= not(layer2_outputs(2517));
    outputs(24) <= not(layer2_outputs(2033));
    outputs(25) <= layer2_outputs(4325);
    outputs(26) <= layer2_outputs(3664);
    outputs(27) <= layer2_outputs(2761);
    outputs(28) <= not(layer2_outputs(1223));
    outputs(29) <= layer2_outputs(1699);
    outputs(30) <= layer2_outputs(1656);
    outputs(31) <= layer2_outputs(1356);
    outputs(32) <= not(layer2_outputs(1897));
    outputs(33) <= (layer2_outputs(1588)) and not (layer2_outputs(2547));
    outputs(34) <= not(layer2_outputs(3807));
    outputs(35) <= not((layer2_outputs(1594)) xor (layer2_outputs(4869)));
    outputs(36) <= layer2_outputs(677);
    outputs(37) <= layer2_outputs(413);
    outputs(38) <= layer2_outputs(4842);
    outputs(39) <= (layer2_outputs(926)) xor (layer2_outputs(3570));
    outputs(40) <= not(layer2_outputs(2895));
    outputs(41) <= not((layer2_outputs(1702)) or (layer2_outputs(694)));
    outputs(42) <= (layer2_outputs(865)) and (layer2_outputs(4742));
    outputs(43) <= layer2_outputs(445);
    outputs(44) <= (layer2_outputs(3308)) and not (layer2_outputs(3887));
    outputs(45) <= not(layer2_outputs(4549)) or (layer2_outputs(4029));
    outputs(46) <= layer2_outputs(3696);
    outputs(47) <= layer2_outputs(4283);
    outputs(48) <= (layer2_outputs(2251)) and not (layer2_outputs(3414));
    outputs(49) <= layer2_outputs(965);
    outputs(50) <= not((layer2_outputs(4814)) and (layer2_outputs(3986)));
    outputs(51) <= (layer2_outputs(412)) and (layer2_outputs(1911));
    outputs(52) <= layer2_outputs(1697);
    outputs(53) <= (layer2_outputs(1084)) and (layer2_outputs(2767));
    outputs(54) <= (layer2_outputs(1029)) and not (layer2_outputs(528));
    outputs(55) <= not(layer2_outputs(3963));
    outputs(56) <= layer2_outputs(4405);
    outputs(57) <= not(layer2_outputs(1794));
    outputs(58) <= layer2_outputs(4582);
    outputs(59) <= (layer2_outputs(2231)) and (layer2_outputs(2839));
    outputs(60) <= layer2_outputs(4482);
    outputs(61) <= layer2_outputs(1630);
    outputs(62) <= layer2_outputs(3059);
    outputs(63) <= layer2_outputs(3349);
    outputs(64) <= not((layer2_outputs(4902)) xor (layer2_outputs(1015)));
    outputs(65) <= (layer2_outputs(2269)) and not (layer2_outputs(390));
    outputs(66) <= not(layer2_outputs(559));
    outputs(67) <= not(layer2_outputs(285));
    outputs(68) <= not(layer2_outputs(626));
    outputs(69) <= not((layer2_outputs(1080)) and (layer2_outputs(4150)));
    outputs(70) <= not(layer2_outputs(931));
    outputs(71) <= (layer2_outputs(4508)) and (layer2_outputs(2806));
    outputs(72) <= layer2_outputs(4842);
    outputs(73) <= not(layer2_outputs(2126));
    outputs(74) <= not(layer2_outputs(3572));
    outputs(75) <= not(layer2_outputs(2545));
    outputs(76) <= layer2_outputs(257);
    outputs(77) <= layer2_outputs(1138);
    outputs(78) <= (layer2_outputs(1680)) and (layer2_outputs(4783));
    outputs(79) <= layer2_outputs(797);
    outputs(80) <= layer2_outputs(2109);
    outputs(81) <= layer2_outputs(4240);
    outputs(82) <= not(layer2_outputs(3131));
    outputs(83) <= not((layer2_outputs(3055)) and (layer2_outputs(4280)));
    outputs(84) <= not(layer2_outputs(2121));
    outputs(85) <= layer2_outputs(2986);
    outputs(86) <= not(layer2_outputs(231));
    outputs(87) <= not(layer2_outputs(4911)) or (layer2_outputs(4338));
    outputs(88) <= not(layer2_outputs(441));
    outputs(89) <= not(layer2_outputs(3404)) or (layer2_outputs(1106));
    outputs(90) <= layer2_outputs(3039);
    outputs(91) <= layer2_outputs(350);
    outputs(92) <= layer2_outputs(363);
    outputs(93) <= not((layer2_outputs(4016)) and (layer2_outputs(1874)));
    outputs(94) <= layer2_outputs(510);
    outputs(95) <= not(layer2_outputs(1617));
    outputs(96) <= layer2_outputs(1433);
    outputs(97) <= not(layer2_outputs(4812));
    outputs(98) <= not(layer2_outputs(1706));
    outputs(99) <= not(layer2_outputs(1249));
    outputs(100) <= layer2_outputs(969);
    outputs(101) <= (layer2_outputs(2255)) and (layer2_outputs(371));
    outputs(102) <= not(layer2_outputs(1133));
    outputs(103) <= layer2_outputs(2972);
    outputs(104) <= layer2_outputs(4013);
    outputs(105) <= layer2_outputs(4256);
    outputs(106) <= (layer2_outputs(541)) and not (layer2_outputs(3962));
    outputs(107) <= (layer2_outputs(3064)) or (layer2_outputs(2581));
    outputs(108) <= layer2_outputs(4976);
    outputs(109) <= (layer2_outputs(1178)) and not (layer2_outputs(64));
    outputs(110) <= not(layer2_outputs(661));
    outputs(111) <= not(layer2_outputs(1309));
    outputs(112) <= not(layer2_outputs(3321));
    outputs(113) <= not((layer2_outputs(2233)) xor (layer2_outputs(431)));
    outputs(114) <= layer2_outputs(2788);
    outputs(115) <= (layer2_outputs(4272)) and not (layer2_outputs(4498));
    outputs(116) <= not(layer2_outputs(5119));
    outputs(117) <= not(layer2_outputs(2702)) or (layer2_outputs(2065));
    outputs(118) <= layer2_outputs(4787);
    outputs(119) <= layer2_outputs(4030);
    outputs(120) <= layer2_outputs(2890);
    outputs(121) <= not(layer2_outputs(2979)) or (layer2_outputs(3836));
    outputs(122) <= not(layer2_outputs(2075));
    outputs(123) <= not(layer2_outputs(3072));
    outputs(124) <= (layer2_outputs(1107)) xor (layer2_outputs(3357));
    outputs(125) <= layer2_outputs(221);
    outputs(126) <= (layer2_outputs(505)) or (layer2_outputs(4305));
    outputs(127) <= not(layer2_outputs(3527));
    outputs(128) <= not(layer2_outputs(791));
    outputs(129) <= not(layer2_outputs(2769));
    outputs(130) <= layer2_outputs(4193);
    outputs(131) <= not(layer2_outputs(4821)) or (layer2_outputs(4952));
    outputs(132) <= not((layer2_outputs(923)) or (layer2_outputs(1443)));
    outputs(133) <= not(layer2_outputs(775));
    outputs(134) <= not(layer2_outputs(2910));
    outputs(135) <= (layer2_outputs(2733)) xor (layer2_outputs(1190));
    outputs(136) <= not(layer2_outputs(3028));
    outputs(137) <= not(layer2_outputs(1728));
    outputs(138) <= (layer2_outputs(305)) or (layer2_outputs(11));
    outputs(139) <= layer2_outputs(4866);
    outputs(140) <= not(layer2_outputs(532));
    outputs(141) <= not((layer2_outputs(945)) or (layer2_outputs(1816)));
    outputs(142) <= not((layer2_outputs(2939)) and (layer2_outputs(1487)));
    outputs(143) <= layer2_outputs(117);
    outputs(144) <= not(layer2_outputs(2422));
    outputs(145) <= not((layer2_outputs(478)) or (layer2_outputs(2450)));
    outputs(146) <= not(layer2_outputs(5013)) or (layer2_outputs(4746));
    outputs(147) <= layer2_outputs(145);
    outputs(148) <= not(layer2_outputs(1452));
    outputs(149) <= not(layer2_outputs(3245));
    outputs(150) <= not(layer2_outputs(2497));
    outputs(151) <= not(layer2_outputs(4802));
    outputs(152) <= layer2_outputs(1473);
    outputs(153) <= layer2_outputs(133);
    outputs(154) <= layer2_outputs(2553);
    outputs(155) <= (layer2_outputs(4149)) and not (layer2_outputs(3858));
    outputs(156) <= not(layer2_outputs(4027));
    outputs(157) <= not(layer2_outputs(1994));
    outputs(158) <= not(layer2_outputs(4982));
    outputs(159) <= not(layer2_outputs(4888));
    outputs(160) <= not(layer2_outputs(3183));
    outputs(161) <= not(layer2_outputs(4421));
    outputs(162) <= not(layer2_outputs(4712));
    outputs(163) <= not(layer2_outputs(2284));
    outputs(164) <= layer2_outputs(3968);
    outputs(165) <= not(layer2_outputs(3007));
    outputs(166) <= not(layer2_outputs(1046));
    outputs(167) <= not(layer2_outputs(3093)) or (layer2_outputs(4038));
    outputs(168) <= not(layer2_outputs(434));
    outputs(169) <= not(layer2_outputs(1437));
    outputs(170) <= layer2_outputs(1363);
    outputs(171) <= not((layer2_outputs(3354)) or (layer2_outputs(4209)));
    outputs(172) <= (layer2_outputs(1472)) and not (layer2_outputs(355));
    outputs(173) <= not(layer2_outputs(5060));
    outputs(174) <= layer2_outputs(3242);
    outputs(175) <= not(layer2_outputs(3784));
    outputs(176) <= (layer2_outputs(4211)) and not (layer2_outputs(2665));
    outputs(177) <= layer2_outputs(3417);
    outputs(178) <= (layer2_outputs(93)) and (layer2_outputs(4263));
    outputs(179) <= not((layer2_outputs(2870)) or (layer2_outputs(2996)));
    outputs(180) <= not((layer2_outputs(1641)) xor (layer2_outputs(2032)));
    outputs(181) <= layer2_outputs(3849);
    outputs(182) <= (layer2_outputs(1475)) xor (layer2_outputs(32));
    outputs(183) <= (layer2_outputs(379)) and not (layer2_outputs(3996));
    outputs(184) <= not((layer2_outputs(2962)) xor (layer2_outputs(4983)));
    outputs(185) <= not(layer2_outputs(846));
    outputs(186) <= not((layer2_outputs(1422)) xor (layer2_outputs(238)));
    outputs(187) <= layer2_outputs(1759);
    outputs(188) <= not(layer2_outputs(884));
    outputs(189) <= not((layer2_outputs(4088)) xor (layer2_outputs(3744)));
    outputs(190) <= layer2_outputs(658);
    outputs(191) <= not(layer2_outputs(3983));
    outputs(192) <= layer2_outputs(2502);
    outputs(193) <= not(layer2_outputs(3364));
    outputs(194) <= layer2_outputs(5075);
    outputs(195) <= not(layer2_outputs(1554));
    outputs(196) <= not((layer2_outputs(1485)) or (layer2_outputs(4365)));
    outputs(197) <= layer2_outputs(116);
    outputs(198) <= layer2_outputs(2091);
    outputs(199) <= layer2_outputs(4239);
    outputs(200) <= (layer2_outputs(4923)) and not (layer2_outputs(3668));
    outputs(201) <= not(layer2_outputs(4950));
    outputs(202) <= layer2_outputs(2042);
    outputs(203) <= (layer2_outputs(958)) and not (layer2_outputs(4075));
    outputs(204) <= layer2_outputs(895);
    outputs(205) <= layer2_outputs(4750);
    outputs(206) <= layer2_outputs(4859);
    outputs(207) <= (layer2_outputs(3403)) xor (layer2_outputs(3660));
    outputs(208) <= not(layer2_outputs(2052));
    outputs(209) <= not((layer2_outputs(4456)) and (layer2_outputs(3062)));
    outputs(210) <= layer2_outputs(3794);
    outputs(211) <= not(layer2_outputs(3935));
    outputs(212) <= layer2_outputs(191);
    outputs(213) <= not(layer2_outputs(3026)) or (layer2_outputs(4121));
    outputs(214) <= layer2_outputs(3398);
    outputs(215) <= not(layer2_outputs(4739));
    outputs(216) <= not((layer2_outputs(4989)) and (layer2_outputs(425)));
    outputs(217) <= not(layer2_outputs(4105));
    outputs(218) <= not(layer2_outputs(1544));
    outputs(219) <= not(layer2_outputs(4829));
    outputs(220) <= layer2_outputs(2901);
    outputs(221) <= layer2_outputs(2248);
    outputs(222) <= not(layer2_outputs(2118));
    outputs(223) <= layer2_outputs(1377);
    outputs(224) <= not(layer2_outputs(866));
    outputs(225) <= not(layer2_outputs(2100));
    outputs(226) <= layer2_outputs(4628);
    outputs(227) <= not((layer2_outputs(3206)) xor (layer2_outputs(1305)));
    outputs(228) <= layer2_outputs(4535);
    outputs(229) <= layer2_outputs(3461);
    outputs(230) <= not(layer2_outputs(3243));
    outputs(231) <= layer2_outputs(490);
    outputs(232) <= not(layer2_outputs(4949));
    outputs(233) <= layer2_outputs(2578);
    outputs(234) <= not(layer2_outputs(3212)) or (layer2_outputs(2718));
    outputs(235) <= not(layer2_outputs(3799)) or (layer2_outputs(4795));
    outputs(236) <= not(layer2_outputs(651));
    outputs(237) <= layer2_outputs(3099);
    outputs(238) <= (layer2_outputs(4886)) and not (layer2_outputs(137));
    outputs(239) <= not((layer2_outputs(1932)) xor (layer2_outputs(4825)));
    outputs(240) <= not(layer2_outputs(2996));
    outputs(241) <= not(layer2_outputs(4484));
    outputs(242) <= not(layer2_outputs(1461)) or (layer2_outputs(1117));
    outputs(243) <= (layer2_outputs(3508)) and not (layer2_outputs(4049));
    outputs(244) <= not(layer2_outputs(2628));
    outputs(245) <= layer2_outputs(3166);
    outputs(246) <= layer2_outputs(3420);
    outputs(247) <= (layer2_outputs(4284)) or (layer2_outputs(1017));
    outputs(248) <= layer2_outputs(1623);
    outputs(249) <= layer2_outputs(2098);
    outputs(250) <= not(layer2_outputs(2316));
    outputs(251) <= not((layer2_outputs(1706)) or (layer2_outputs(2182)));
    outputs(252) <= not(layer2_outputs(3057));
    outputs(253) <= layer2_outputs(4086);
    outputs(254) <= layer2_outputs(4535);
    outputs(255) <= not(layer2_outputs(3809));
    outputs(256) <= (layer2_outputs(5004)) and (layer2_outputs(2148));
    outputs(257) <= layer2_outputs(1881);
    outputs(258) <= not(layer2_outputs(3617)) or (layer2_outputs(1587));
    outputs(259) <= not(layer2_outputs(3725));
    outputs(260) <= (layer2_outputs(1773)) and not (layer2_outputs(454));
    outputs(261) <= not((layer2_outputs(3983)) or (layer2_outputs(3782)));
    outputs(262) <= not(layer2_outputs(3896));
    outputs(263) <= layer2_outputs(4885);
    outputs(264) <= not(layer2_outputs(694));
    outputs(265) <= (layer2_outputs(2304)) xor (layer2_outputs(1210));
    outputs(266) <= not(layer2_outputs(2703));
    outputs(267) <= layer2_outputs(2034);
    outputs(268) <= layer2_outputs(699);
    outputs(269) <= (layer2_outputs(4658)) or (layer2_outputs(937));
    outputs(270) <= layer2_outputs(1810);
    outputs(271) <= not(layer2_outputs(3042)) or (layer2_outputs(2362));
    outputs(272) <= layer2_outputs(574);
    outputs(273) <= layer2_outputs(542);
    outputs(274) <= (layer2_outputs(1615)) or (layer2_outputs(4884));
    outputs(275) <= not(layer2_outputs(2708));
    outputs(276) <= not(layer2_outputs(4602));
    outputs(277) <= layer2_outputs(1199);
    outputs(278) <= not((layer2_outputs(1908)) and (layer2_outputs(3405)));
    outputs(279) <= layer2_outputs(599);
    outputs(280) <= layer2_outputs(3785);
    outputs(281) <= layer2_outputs(2566);
    outputs(282) <= layer2_outputs(103);
    outputs(283) <= not(layer2_outputs(2908));
    outputs(284) <= layer2_outputs(4755);
    outputs(285) <= layer2_outputs(2468);
    outputs(286) <= not(layer2_outputs(719));
    outputs(287) <= (layer2_outputs(271)) and not (layer2_outputs(3750));
    outputs(288) <= (layer2_outputs(4673)) and not (layer2_outputs(4664));
    outputs(289) <= not(layer2_outputs(2825));
    outputs(290) <= not(layer2_outputs(3063));
    outputs(291) <= not((layer2_outputs(414)) and (layer2_outputs(851)));
    outputs(292) <= not(layer2_outputs(3304));
    outputs(293) <= not((layer2_outputs(3585)) xor (layer2_outputs(1427)));
    outputs(294) <= layer2_outputs(3985);
    outputs(295) <= (layer2_outputs(3800)) and (layer2_outputs(1221));
    outputs(296) <= not((layer2_outputs(4421)) or (layer2_outputs(4261)));
    outputs(297) <= (layer2_outputs(4899)) and not (layer2_outputs(2779));
    outputs(298) <= layer2_outputs(4000);
    outputs(299) <= layer2_outputs(3490);
    outputs(300) <= layer2_outputs(3452);
    outputs(301) <= not(layer2_outputs(4998)) or (layer2_outputs(4545));
    outputs(302) <= not(layer2_outputs(1741));
    outputs(303) <= layer2_outputs(1424);
    outputs(304) <= not(layer2_outputs(349)) or (layer2_outputs(2006));
    outputs(305) <= layer2_outputs(4222);
    outputs(306) <= (layer2_outputs(3273)) or (layer2_outputs(1153));
    outputs(307) <= not(layer2_outputs(3731));
    outputs(308) <= not((layer2_outputs(3297)) and (layer2_outputs(4251)));
    outputs(309) <= not((layer2_outputs(3924)) xor (layer2_outputs(501)));
    outputs(310) <= not((layer2_outputs(1230)) xor (layer2_outputs(1072)));
    outputs(311) <= layer2_outputs(4808);
    outputs(312) <= (layer2_outputs(3083)) and not (layer2_outputs(2683));
    outputs(313) <= not(layer2_outputs(512));
    outputs(314) <= not((layer2_outputs(3869)) or (layer2_outputs(892)));
    outputs(315) <= not((layer2_outputs(3432)) xor (layer2_outputs(391)));
    outputs(316) <= layer2_outputs(2220);
    outputs(317) <= not(layer2_outputs(1969));
    outputs(318) <= not(layer2_outputs(2431));
    outputs(319) <= (layer2_outputs(4948)) and not (layer2_outputs(1057));
    outputs(320) <= not(layer2_outputs(1457));
    outputs(321) <= (layer2_outputs(1495)) xor (layer2_outputs(1220));
    outputs(322) <= not(layer2_outputs(4592));
    outputs(323) <= (layer2_outputs(2920)) and not (layer2_outputs(4072));
    outputs(324) <= not(layer2_outputs(4401));
    outputs(325) <= not(layer2_outputs(2379));
    outputs(326) <= layer2_outputs(1355);
    outputs(327) <= not((layer2_outputs(2169)) or (layer2_outputs(400)));
    outputs(328) <= layer2_outputs(1700);
    outputs(329) <= (layer2_outputs(465)) xor (layer2_outputs(2445));
    outputs(330) <= (layer2_outputs(4282)) and not (layer2_outputs(2778));
    outputs(331) <= not(layer2_outputs(803));
    outputs(332) <= not((layer2_outputs(4386)) xor (layer2_outputs(3960)));
    outputs(333) <= layer2_outputs(1927);
    outputs(334) <= not(layer2_outputs(2357));
    outputs(335) <= not(layer2_outputs(1108));
    outputs(336) <= not(layer2_outputs(4587));
    outputs(337) <= not(layer2_outputs(1873));
    outputs(338) <= not(layer2_outputs(452));
    outputs(339) <= not(layer2_outputs(4957));
    outputs(340) <= not(layer2_outputs(2150));
    outputs(341) <= layer2_outputs(4221);
    outputs(342) <= not(layer2_outputs(244));
    outputs(343) <= (layer2_outputs(1626)) and not (layer2_outputs(4933));
    outputs(344) <= not(layer2_outputs(3136));
    outputs(345) <= not(layer2_outputs(2471));
    outputs(346) <= (layer2_outputs(1746)) xor (layer2_outputs(2016));
    outputs(347) <= not((layer2_outputs(4635)) or (layer2_outputs(1205)));
    outputs(348) <= (layer2_outputs(3648)) and not (layer2_outputs(1339));
    outputs(349) <= not(layer2_outputs(4965));
    outputs(350) <= (layer2_outputs(364)) xor (layer2_outputs(2579));
    outputs(351) <= layer2_outputs(3039);
    outputs(352) <= not(layer2_outputs(3132));
    outputs(353) <= not(layer2_outputs(4663));
    outputs(354) <= not((layer2_outputs(4736)) xor (layer2_outputs(2345)));
    outputs(355) <= (layer2_outputs(3646)) and not (layer2_outputs(4154));
    outputs(356) <= (layer2_outputs(1479)) and not (layer2_outputs(3935));
    outputs(357) <= layer2_outputs(748);
    outputs(358) <= layer2_outputs(3795);
    outputs(359) <= layer2_outputs(3953);
    outputs(360) <= layer2_outputs(3467);
    outputs(361) <= layer2_outputs(2551);
    outputs(362) <= not(layer2_outputs(1115));
    outputs(363) <= not(layer2_outputs(3659)) or (layer2_outputs(3034));
    outputs(364) <= not(layer2_outputs(4090));
    outputs(365) <= (layer2_outputs(3260)) and (layer2_outputs(847));
    outputs(366) <= layer2_outputs(3463);
    outputs(367) <= layer2_outputs(1881);
    outputs(368) <= not(layer2_outputs(671));
    outputs(369) <= (layer2_outputs(5079)) and not (layer2_outputs(4231));
    outputs(370) <= not(layer2_outputs(543));
    outputs(371) <= layer2_outputs(970);
    outputs(372) <= not(layer2_outputs(1613));
    outputs(373) <= layer2_outputs(3348);
    outputs(374) <= not(layer2_outputs(2486));
    outputs(375) <= layer2_outputs(3945);
    outputs(376) <= not(layer2_outputs(2159));
    outputs(377) <= not((layer2_outputs(783)) or (layer2_outputs(2911)));
    outputs(378) <= (layer2_outputs(3196)) xor (layer2_outputs(1670));
    outputs(379) <= layer2_outputs(2386);
    outputs(380) <= not(layer2_outputs(1514));
    outputs(381) <= layer2_outputs(19);
    outputs(382) <= layer2_outputs(944);
    outputs(383) <= layer2_outputs(4725);
    outputs(384) <= layer2_outputs(839);
    outputs(385) <= not(layer2_outputs(3189));
    outputs(386) <= layer2_outputs(1882);
    outputs(387) <= (layer2_outputs(1055)) and (layer2_outputs(57));
    outputs(388) <= not(layer2_outputs(1660));
    outputs(389) <= not((layer2_outputs(1733)) or (layer2_outputs(1504)));
    outputs(390) <= layer2_outputs(4822);
    outputs(391) <= layer2_outputs(1500);
    outputs(392) <= layer2_outputs(191);
    outputs(393) <= not(layer2_outputs(1379));
    outputs(394) <= not(layer2_outputs(635));
    outputs(395) <= not(layer2_outputs(1769));
    outputs(396) <= layer2_outputs(2385);
    outputs(397) <= (layer2_outputs(1549)) and not (layer2_outputs(4623));
    outputs(398) <= not(layer2_outputs(4102)) or (layer2_outputs(3140));
    outputs(399) <= not(layer2_outputs(2279));
    outputs(400) <= not(layer2_outputs(5119));
    outputs(401) <= (layer2_outputs(2222)) and not (layer2_outputs(3401));
    outputs(402) <= not(layer2_outputs(4249));
    outputs(403) <= not((layer2_outputs(4861)) and (layer2_outputs(2648)));
    outputs(404) <= layer2_outputs(777);
    outputs(405) <= layer2_outputs(39);
    outputs(406) <= layer2_outputs(4232);
    outputs(407) <= not(layer2_outputs(2170));
    outputs(408) <= not(layer2_outputs(199));
    outputs(409) <= (layer2_outputs(4028)) and not (layer2_outputs(4935));
    outputs(410) <= layer2_outputs(249);
    outputs(411) <= not(layer2_outputs(4053));
    outputs(412) <= not(layer2_outputs(975));
    outputs(413) <= layer2_outputs(2529);
    outputs(414) <= not(layer2_outputs(3675));
    outputs(415) <= not((layer2_outputs(2942)) and (layer2_outputs(2167)));
    outputs(416) <= not(layer2_outputs(1051)) or (layer2_outputs(527));
    outputs(417) <= layer2_outputs(2887);
    outputs(418) <= not(layer2_outputs(2366));
    outputs(419) <= not((layer2_outputs(3824)) xor (layer2_outputs(4709)));
    outputs(420) <= layer2_outputs(828);
    outputs(421) <= not(layer2_outputs(4595));
    outputs(422) <= not((layer2_outputs(2742)) and (layer2_outputs(2640)));
    outputs(423) <= not(layer2_outputs(2784));
    outputs(424) <= not(layer2_outputs(5077));
    outputs(425) <= (layer2_outputs(2540)) and not (layer2_outputs(3788));
    outputs(426) <= layer2_outputs(472);
    outputs(427) <= not((layer2_outputs(4782)) or (layer2_outputs(4258)));
    outputs(428) <= layer2_outputs(2565);
    outputs(429) <= not(layer2_outputs(4940));
    outputs(430) <= not(layer2_outputs(104));
    outputs(431) <= layer2_outputs(293);
    outputs(432) <= layer2_outputs(2985);
    outputs(433) <= not(layer2_outputs(2092));
    outputs(434) <= not(layer2_outputs(882));
    outputs(435) <= layer2_outputs(1011);
    outputs(436) <= layer2_outputs(4705);
    outputs(437) <= layer2_outputs(1625);
    outputs(438) <= (layer2_outputs(4458)) and not (layer2_outputs(3091));
    outputs(439) <= not(layer2_outputs(4225));
    outputs(440) <= not((layer2_outputs(2149)) xor (layer2_outputs(1038)));
    outputs(441) <= not(layer2_outputs(2224));
    outputs(442) <= not(layer2_outputs(4328));
    outputs(443) <= layer2_outputs(4966);
    outputs(444) <= layer2_outputs(857);
    outputs(445) <= (layer2_outputs(3293)) and not (layer2_outputs(3413));
    outputs(446) <= layer2_outputs(1836);
    outputs(447) <= not(layer2_outputs(606));
    outputs(448) <= (layer2_outputs(2269)) xor (layer2_outputs(2789));
    outputs(449) <= not((layer2_outputs(3171)) or (layer2_outputs(2400)));
    outputs(450) <= (layer2_outputs(638)) and not (layer2_outputs(3330));
    outputs(451) <= layer2_outputs(3137);
    outputs(452) <= (layer2_outputs(4847)) xor (layer2_outputs(5029));
    outputs(453) <= not((layer2_outputs(3362)) or (layer2_outputs(1547)));
    outputs(454) <= layer2_outputs(1575);
    outputs(455) <= (layer2_outputs(2393)) and not (layer2_outputs(3788));
    outputs(456) <= not((layer2_outputs(967)) xor (layer2_outputs(166)));
    outputs(457) <= (layer2_outputs(4137)) xor (layer2_outputs(268));
    outputs(458) <= layer2_outputs(3568);
    outputs(459) <= layer2_outputs(3210);
    outputs(460) <= not(layer2_outputs(4498));
    outputs(461) <= not(layer2_outputs(2616));
    outputs(462) <= (layer2_outputs(4619)) xor (layer2_outputs(3580));
    outputs(463) <= not(layer2_outputs(2365));
    outputs(464) <= layer2_outputs(4228);
    outputs(465) <= not(layer2_outputs(1411));
    outputs(466) <= not(layer2_outputs(1393));
    outputs(467) <= layer2_outputs(4449);
    outputs(468) <= layer2_outputs(933);
    outputs(469) <= layer2_outputs(4947);
    outputs(470) <= not(layer2_outputs(3932));
    outputs(471) <= (layer2_outputs(206)) xor (layer2_outputs(4199));
    outputs(472) <= (layer2_outputs(3494)) and (layer2_outputs(2098));
    outputs(473) <= layer2_outputs(840);
    outputs(474) <= layer2_outputs(3065);
    outputs(475) <= not((layer2_outputs(2146)) or (layer2_outputs(3655)));
    outputs(476) <= not(layer2_outputs(1578));
    outputs(477) <= (layer2_outputs(2505)) and (layer2_outputs(3648));
    outputs(478) <= layer2_outputs(427);
    outputs(479) <= layer2_outputs(1473);
    outputs(480) <= not(layer2_outputs(3500));
    outputs(481) <= (layer2_outputs(3961)) and not (layer2_outputs(3554));
    outputs(482) <= layer2_outputs(1773);
    outputs(483) <= (layer2_outputs(4612)) and not (layer2_outputs(5058));
    outputs(484) <= layer2_outputs(1127);
    outputs(485) <= not(layer2_outputs(2453)) or (layer2_outputs(2332));
    outputs(486) <= (layer2_outputs(524)) and not (layer2_outputs(2432));
    outputs(487) <= not(layer2_outputs(3150));
    outputs(488) <= (layer2_outputs(2790)) and not (layer2_outputs(4229));
    outputs(489) <= layer2_outputs(1017);
    outputs(490) <= layer2_outputs(433);
    outputs(491) <= not(layer2_outputs(1618));
    outputs(492) <= not((layer2_outputs(2101)) xor (layer2_outputs(4647)));
    outputs(493) <= (layer2_outputs(2165)) and not (layer2_outputs(182));
    outputs(494) <= not((layer2_outputs(3007)) and (layer2_outputs(2660)));
    outputs(495) <= layer2_outputs(443);
    outputs(496) <= not(layer2_outputs(999));
    outputs(497) <= layer2_outputs(2899);
    outputs(498) <= not(layer2_outputs(4788));
    outputs(499) <= (layer2_outputs(3573)) and (layer2_outputs(3199));
    outputs(500) <= layer2_outputs(211);
    outputs(501) <= layer2_outputs(3852);
    outputs(502) <= not(layer2_outputs(1545));
    outputs(503) <= not(layer2_outputs(1663));
    outputs(504) <= not(layer2_outputs(771));
    outputs(505) <= not(layer2_outputs(2004));
    outputs(506) <= not((layer2_outputs(4220)) or (layer2_outputs(2216)));
    outputs(507) <= not(layer2_outputs(3811));
    outputs(508) <= layer2_outputs(514);
    outputs(509) <= not((layer2_outputs(955)) xor (layer2_outputs(3851)));
    outputs(510) <= '1';
    outputs(511) <= not(layer2_outputs(2819));
    outputs(512) <= not(layer2_outputs(4881));
    outputs(513) <= layer2_outputs(2649);
    outputs(514) <= not((layer2_outputs(2796)) xor (layer2_outputs(699)));
    outputs(515) <= layer2_outputs(4776);
    outputs(516) <= not(layer2_outputs(2473));
    outputs(517) <= (layer2_outputs(2592)) and (layer2_outputs(488));
    outputs(518) <= layer2_outputs(2316);
    outputs(519) <= layer2_outputs(1025);
    outputs(520) <= (layer2_outputs(3306)) and (layer2_outputs(767));
    outputs(521) <= (layer2_outputs(1391)) and (layer2_outputs(686));
    outputs(522) <= layer2_outputs(3237);
    outputs(523) <= (layer2_outputs(1906)) or (layer2_outputs(3911));
    outputs(524) <= not(layer2_outputs(1023));
    outputs(525) <= not(layer2_outputs(616));
    outputs(526) <= not((layer2_outputs(2171)) or (layer2_outputs(832)));
    outputs(527) <= (layer2_outputs(608)) and not (layer2_outputs(2374));
    outputs(528) <= (layer2_outputs(3062)) xor (layer2_outputs(4058));
    outputs(529) <= '0';
    outputs(530) <= (layer2_outputs(724)) and not (layer2_outputs(1410));
    outputs(531) <= (layer2_outputs(2071)) and not (layer2_outputs(1202));
    outputs(532) <= layer2_outputs(471);
    outputs(533) <= (layer2_outputs(1744)) and not (layer2_outputs(925));
    outputs(534) <= not(layer2_outputs(2375));
    outputs(535) <= not(layer2_outputs(162));
    outputs(536) <= (layer2_outputs(21)) and (layer2_outputs(1242));
    outputs(537) <= (layer2_outputs(4311)) and not (layer2_outputs(4632));
    outputs(538) <= layer2_outputs(3948);
    outputs(539) <= not(layer2_outputs(875));
    outputs(540) <= not((layer2_outputs(4551)) or (layer2_outputs(272)));
    outputs(541) <= layer2_outputs(3466);
    outputs(542) <= not(layer2_outputs(2501));
    outputs(543) <= layer2_outputs(4879);
    outputs(544) <= (layer2_outputs(741)) or (layer2_outputs(4538));
    outputs(545) <= not(layer2_outputs(4780));
    outputs(546) <= (layer2_outputs(4727)) and (layer2_outputs(2614));
    outputs(547) <= layer2_outputs(4816);
    outputs(548) <= (layer2_outputs(4218)) and (layer2_outputs(972));
    outputs(549) <= not(layer2_outputs(2438)) or (layer2_outputs(3904));
    outputs(550) <= (layer2_outputs(1001)) and not (layer2_outputs(660));
    outputs(551) <= layer2_outputs(4717);
    outputs(552) <= layer2_outputs(452);
    outputs(553) <= not(layer2_outputs(4457));
    outputs(554) <= not((layer2_outputs(3840)) or (layer2_outputs(1088)));
    outputs(555) <= (layer2_outputs(4022)) and (layer2_outputs(4420));
    outputs(556) <= layer2_outputs(217);
    outputs(557) <= layer2_outputs(3436);
    outputs(558) <= (layer2_outputs(4112)) and (layer2_outputs(4790));
    outputs(559) <= not((layer2_outputs(1035)) or (layer2_outputs(157)));
    outputs(560) <= not(layer2_outputs(969));
    outputs(561) <= not(layer2_outputs(4001));
    outputs(562) <= layer2_outputs(4647);
    outputs(563) <= not(layer2_outputs(2127));
    outputs(564) <= not((layer2_outputs(2585)) xor (layer2_outputs(2198)));
    outputs(565) <= not(layer2_outputs(4322));
    outputs(566) <= (layer2_outputs(388)) and (layer2_outputs(1616));
    outputs(567) <= (layer2_outputs(5007)) and (layer2_outputs(900));
    outputs(568) <= (layer2_outputs(3378)) and not (layer2_outputs(723));
    outputs(569) <= (layer2_outputs(3351)) and (layer2_outputs(1442));
    outputs(570) <= (layer2_outputs(2259)) and (layer2_outputs(3891));
    outputs(571) <= not(layer2_outputs(36));
    outputs(572) <= layer2_outputs(3035);
    outputs(573) <= not((layer2_outputs(1281)) xor (layer2_outputs(3361)));
    outputs(574) <= not(layer2_outputs(4901));
    outputs(575) <= (layer2_outputs(4008)) and not (layer2_outputs(4476));
    outputs(576) <= layer2_outputs(2207);
    outputs(577) <= not((layer2_outputs(4089)) or (layer2_outputs(1713)));
    outputs(578) <= layer2_outputs(413);
    outputs(579) <= (layer2_outputs(2757)) and not (layer2_outputs(654));
    outputs(580) <= layer2_outputs(2208);
    outputs(581) <= (layer2_outputs(5105)) and not (layer2_outputs(4916));
    outputs(582) <= (layer2_outputs(1198)) and (layer2_outputs(3654));
    outputs(583) <= not(layer2_outputs(4296));
    outputs(584) <= not((layer2_outputs(989)) xor (layer2_outputs(5006)));
    outputs(585) <= not(layer2_outputs(2951));
    outputs(586) <= layer2_outputs(3093);
    outputs(587) <= not((layer2_outputs(4649)) or (layer2_outputs(1265)));
    outputs(588) <= layer2_outputs(4261);
    outputs(589) <= not(layer2_outputs(4371));
    outputs(590) <= not(layer2_outputs(4516));
    outputs(591) <= not((layer2_outputs(4373)) or (layer2_outputs(2129)));
    outputs(592) <= (layer2_outputs(3646)) and (layer2_outputs(4110));
    outputs(593) <= layer2_outputs(4424);
    outputs(594) <= layer2_outputs(4366);
    outputs(595) <= (layer2_outputs(265)) and not (layer2_outputs(1123));
    outputs(596) <= (layer2_outputs(5078)) and not (layer2_outputs(1170));
    outputs(597) <= (layer2_outputs(3912)) and not (layer2_outputs(1225));
    outputs(598) <= (layer2_outputs(4908)) and not (layer2_outputs(664));
    outputs(599) <= not((layer2_outputs(4143)) or (layer2_outputs(3872)));
    outputs(600) <= not((layer2_outputs(2198)) or (layer2_outputs(735)));
    outputs(601) <= not((layer2_outputs(4391)) xor (layer2_outputs(4487)));
    outputs(602) <= (layer2_outputs(2351)) and not (layer2_outputs(624));
    outputs(603) <= not(layer2_outputs(1200));
    outputs(604) <= (layer2_outputs(1506)) and (layer2_outputs(4078));
    outputs(605) <= (layer2_outputs(841)) and not (layer2_outputs(340));
    outputs(606) <= (layer2_outputs(2116)) and not (layer2_outputs(5071));
    outputs(607) <= not((layer2_outputs(3799)) or (layer2_outputs(4135)));
    outputs(608) <= (layer2_outputs(2817)) and not (layer2_outputs(4467));
    outputs(609) <= not(layer2_outputs(4854));
    outputs(610) <= (layer2_outputs(1981)) and (layer2_outputs(999));
    outputs(611) <= not(layer2_outputs(3529));
    outputs(612) <= not((layer2_outputs(1877)) or (layer2_outputs(2361)));
    outputs(613) <= not((layer2_outputs(3878)) or (layer2_outputs(2875)));
    outputs(614) <= (layer2_outputs(3892)) and (layer2_outputs(3136));
    outputs(615) <= not(layer2_outputs(1195));
    outputs(616) <= not((layer2_outputs(2606)) xor (layer2_outputs(4011)));
    outputs(617) <= layer2_outputs(209);
    outputs(618) <= (layer2_outputs(4061)) and (layer2_outputs(4992));
    outputs(619) <= (layer2_outputs(3692)) and not (layer2_outputs(3434));
    outputs(620) <= layer2_outputs(4775);
    outputs(621) <= (layer2_outputs(2173)) and (layer2_outputs(2590));
    outputs(622) <= (layer2_outputs(1527)) and not (layer2_outputs(2906));
    outputs(623) <= not(layer2_outputs(4916));
    outputs(624) <= not(layer2_outputs(4858));
    outputs(625) <= not(layer2_outputs(4793));
    outputs(626) <= not((layer2_outputs(1194)) or (layer2_outputs(3780)));
    outputs(627) <= not(layer2_outputs(1082));
    outputs(628) <= (layer2_outputs(623)) and (layer2_outputs(2997));
    outputs(629) <= not(layer2_outputs(364));
    outputs(630) <= not((layer2_outputs(5016)) or (layer2_outputs(4068)));
    outputs(631) <= not(layer2_outputs(1962));
    outputs(632) <= layer2_outputs(4838);
    outputs(633) <= layer2_outputs(3319);
    outputs(634) <= (layer2_outputs(702)) and not (layer2_outputs(2808));
    outputs(635) <= (layer2_outputs(328)) and not (layer2_outputs(495));
    outputs(636) <= (layer2_outputs(2119)) and not (layer2_outputs(14));
    outputs(637) <= (layer2_outputs(2582)) and (layer2_outputs(4395));
    outputs(638) <= (layer2_outputs(2241)) and not (layer2_outputs(928));
    outputs(639) <= (layer2_outputs(2891)) and not (layer2_outputs(2227));
    outputs(640) <= (layer2_outputs(2482)) and not (layer2_outputs(4450));
    outputs(641) <= not(layer2_outputs(4529));
    outputs(642) <= not(layer2_outputs(3977));
    outputs(643) <= (layer2_outputs(2125)) and (layer2_outputs(1943));
    outputs(644) <= (layer2_outputs(1987)) and (layer2_outputs(4295));
    outputs(645) <= layer2_outputs(947);
    outputs(646) <= (layer2_outputs(1833)) and (layer2_outputs(2491));
    outputs(647) <= (layer2_outputs(4766)) and not (layer2_outputs(4398));
    outputs(648) <= (layer2_outputs(2130)) and not (layer2_outputs(4586));
    outputs(649) <= (layer2_outputs(672)) and not (layer2_outputs(1385));
    outputs(650) <= (layer2_outputs(3672)) and not (layer2_outputs(5080));
    outputs(651) <= (layer2_outputs(4223)) and not (layer2_outputs(97));
    outputs(652) <= not(layer2_outputs(2916));
    outputs(653) <= (layer2_outputs(1767)) and not (layer2_outputs(4891));
    outputs(654) <= (layer2_outputs(4689)) xor (layer2_outputs(2271));
    outputs(655) <= (layer2_outputs(4386)) and not (layer2_outputs(2733));
    outputs(656) <= not(layer2_outputs(4103));
    outputs(657) <= (layer2_outputs(607)) and not (layer2_outputs(1344));
    outputs(658) <= (layer2_outputs(1550)) and not (layer2_outputs(4667));
    outputs(659) <= (layer2_outputs(2741)) and not (layer2_outputs(2879));
    outputs(660) <= not((layer2_outputs(1395)) or (layer2_outputs(3543)));
    outputs(661) <= (layer2_outputs(3574)) and (layer2_outputs(4832));
    outputs(662) <= not(layer2_outputs(1312));
    outputs(663) <= not((layer2_outputs(833)) xor (layer2_outputs(1242)));
    outputs(664) <= (layer2_outputs(2456)) and not (layer2_outputs(127));
    outputs(665) <= not(layer2_outputs(1703));
    outputs(666) <= not((layer2_outputs(3272)) or (layer2_outputs(2843)));
    outputs(667) <= (layer2_outputs(2543)) and (layer2_outputs(390));
    outputs(668) <= (layer2_outputs(818)) and not (layer2_outputs(3808));
    outputs(669) <= (layer2_outputs(4)) and not (layer2_outputs(3019));
    outputs(670) <= not(layer2_outputs(3966));
    outputs(671) <= (layer2_outputs(3236)) and (layer2_outputs(4666));
    outputs(672) <= layer2_outputs(2149);
    outputs(673) <= layer2_outputs(3880);
    outputs(674) <= (layer2_outputs(3320)) and (layer2_outputs(3512));
    outputs(675) <= layer2_outputs(4484);
    outputs(676) <= not((layer2_outputs(4542)) or (layer2_outputs(495)));
    outputs(677) <= layer2_outputs(4070);
    outputs(678) <= (layer2_outputs(869)) and not (layer2_outputs(3088));
    outputs(679) <= layer2_outputs(4686);
    outputs(680) <= (layer2_outputs(79)) xor (layer2_outputs(4762));
    outputs(681) <= (layer2_outputs(4820)) and not (layer2_outputs(4227));
    outputs(682) <= (layer2_outputs(3516)) and not (layer2_outputs(733));
    outputs(683) <= (layer2_outputs(1309)) and not (layer2_outputs(1267));
    outputs(684) <= layer2_outputs(2794);
    outputs(685) <= layer2_outputs(2378);
    outputs(686) <= not(layer2_outputs(3916));
    outputs(687) <= not(layer2_outputs(1089));
    outputs(688) <= layer2_outputs(4390);
    outputs(689) <= not((layer2_outputs(1219)) or (layer2_outputs(2205)));
    outputs(690) <= (layer2_outputs(1528)) xor (layer2_outputs(1972));
    outputs(691) <= (layer2_outputs(3758)) and (layer2_outputs(3801));
    outputs(692) <= layer2_outputs(518);
    outputs(693) <= not(layer2_outputs(1579));
    outputs(694) <= (layer2_outputs(218)) xor (layer2_outputs(278));
    outputs(695) <= not((layer2_outputs(4814)) xor (layer2_outputs(3561)));
    outputs(696) <= not((layer2_outputs(4685)) xor (layer2_outputs(1879)));
    outputs(697) <= not((layer2_outputs(236)) or (layer2_outputs(4012)));
    outputs(698) <= layer2_outputs(25);
    outputs(699) <= (layer2_outputs(720)) xor (layer2_outputs(3988));
    outputs(700) <= (layer2_outputs(763)) and not (layer2_outputs(423));
    outputs(701) <= (layer2_outputs(3318)) and not (layer2_outputs(2750));
    outputs(702) <= layer2_outputs(3277);
    outputs(703) <= not((layer2_outputs(103)) or (layer2_outputs(4372)));
    outputs(704) <= layer2_outputs(3502);
    outputs(705) <= layer2_outputs(4144);
    outputs(706) <= not(layer2_outputs(22));
    outputs(707) <= not(layer2_outputs(2288));
    outputs(708) <= (layer2_outputs(2035)) and not (layer2_outputs(50));
    outputs(709) <= (layer2_outputs(3748)) and (layer2_outputs(2007));
    outputs(710) <= (layer2_outputs(2561)) and not (layer2_outputs(4939));
    outputs(711) <= not(layer2_outputs(4831));
    outputs(712) <= not(layer2_outputs(4648));
    outputs(713) <= layer2_outputs(2993);
    outputs(714) <= layer2_outputs(4431);
    outputs(715) <= (layer2_outputs(2487)) and (layer2_outputs(1169));
    outputs(716) <= not((layer2_outputs(1)) or (layer2_outputs(4026)));
    outputs(717) <= (layer2_outputs(1593)) and not (layer2_outputs(508));
    outputs(718) <= layer2_outputs(462);
    outputs(719) <= layer2_outputs(4017);
    outputs(720) <= (layer2_outputs(47)) and not (layer2_outputs(1596));
    outputs(721) <= not(layer2_outputs(5089));
    outputs(722) <= not(layer2_outputs(15));
    outputs(723) <= not((layer2_outputs(3885)) or (layer2_outputs(1716)));
    outputs(724) <= (layer2_outputs(289)) and (layer2_outputs(519));
    outputs(725) <= (layer2_outputs(2791)) and (layer2_outputs(3649));
    outputs(726) <= not(layer2_outputs(3884));
    outputs(727) <= (layer2_outputs(2660)) and (layer2_outputs(1486));
    outputs(728) <= (layer2_outputs(3326)) xor (layer2_outputs(3682));
    outputs(729) <= not(layer2_outputs(481));
    outputs(730) <= (layer2_outputs(49)) and not (layer2_outputs(50));
    outputs(731) <= (layer2_outputs(3055)) and not (layer2_outputs(3374));
    outputs(732) <= not(layer2_outputs(2848)) or (layer2_outputs(5095));
    outputs(733) <= (layer2_outputs(2075)) and not (layer2_outputs(2227));
    outputs(734) <= (layer2_outputs(2264)) and (layer2_outputs(4121));
    outputs(735) <= (layer2_outputs(114)) and (layer2_outputs(3830));
    outputs(736) <= (layer2_outputs(1768)) xor (layer2_outputs(3035));
    outputs(737) <= not(layer2_outputs(2873));
    outputs(738) <= (layer2_outputs(1545)) xor (layer2_outputs(2140));
    outputs(739) <= not((layer2_outputs(4368)) and (layer2_outputs(961)));
    outputs(740) <= not(layer2_outputs(1468));
    outputs(741) <= (layer2_outputs(2360)) and not (layer2_outputs(2345));
    outputs(742) <= (layer2_outputs(2595)) and not (layer2_outputs(2002));
    outputs(743) <= (layer2_outputs(4992)) and not (layer2_outputs(233));
    outputs(744) <= layer2_outputs(1378);
    outputs(745) <= not(layer2_outputs(1386));
    outputs(746) <= (layer2_outputs(2768)) and not (layer2_outputs(5086));
    outputs(747) <= layer2_outputs(666);
    outputs(748) <= layer2_outputs(518);
    outputs(749) <= not(layer2_outputs(4953));
    outputs(750) <= not((layer2_outputs(4656)) or (layer2_outputs(3595)));
    outputs(751) <= not(layer2_outputs(730));
    outputs(752) <= not(layer2_outputs(2190));
    outputs(753) <= not(layer2_outputs(3023));
    outputs(754) <= not(layer2_outputs(1915));
    outputs(755) <= (layer2_outputs(2086)) and (layer2_outputs(5064));
    outputs(756) <= not(layer2_outputs(3219));
    outputs(757) <= not(layer2_outputs(489));
    outputs(758) <= not(layer2_outputs(1467));
    outputs(759) <= (layer2_outputs(2324)) and not (layer2_outputs(5086));
    outputs(760) <= layer2_outputs(4241);
    outputs(761) <= layer2_outputs(820);
    outputs(762) <= not((layer2_outputs(1905)) or (layer2_outputs(3133)));
    outputs(763) <= (layer2_outputs(2781)) xor (layer2_outputs(86));
    outputs(764) <= not(layer2_outputs(2236));
    outputs(765) <= (layer2_outputs(5011)) and (layer2_outputs(1250));
    outputs(766) <= not(layer2_outputs(2436));
    outputs(767) <= (layer2_outputs(2925)) and (layer2_outputs(5088));
    outputs(768) <= (layer2_outputs(736)) xor (layer2_outputs(3564));
    outputs(769) <= not((layer2_outputs(684)) or (layer2_outputs(1739)));
    outputs(770) <= not((layer2_outputs(3447)) or (layer2_outputs(2565)));
    outputs(771) <= not((layer2_outputs(2010)) or (layer2_outputs(1035)));
    outputs(772) <= not(layer2_outputs(250));
    outputs(773) <= layer2_outputs(2940);
    outputs(774) <= (layer2_outputs(1317)) and (layer2_outputs(1340));
    outputs(775) <= layer2_outputs(2339);
    outputs(776) <= (layer2_outputs(3026)) xor (layer2_outputs(2911));
    outputs(777) <= not((layer2_outputs(4863)) or (layer2_outputs(1475)));
    outputs(778) <= (layer2_outputs(2185)) and not (layer2_outputs(4928));
    outputs(779) <= not((layer2_outputs(2906)) or (layer2_outputs(1417)));
    outputs(780) <= (layer2_outputs(2134)) and (layer2_outputs(2758));
    outputs(781) <= layer2_outputs(3875);
    outputs(782) <= layer2_outputs(2191);
    outputs(783) <= (layer2_outputs(2929)) and (layer2_outputs(1478));
    outputs(784) <= (layer2_outputs(3559)) and (layer2_outputs(628));
    outputs(785) <= layer2_outputs(3937);
    outputs(786) <= (layer2_outputs(2747)) and not (layer2_outputs(2459));
    outputs(787) <= (layer2_outputs(3175)) and not (layer2_outputs(1362));
    outputs(788) <= not((layer2_outputs(5033)) or (layer2_outputs(1858)));
    outputs(789) <= not((layer2_outputs(2435)) or (layer2_outputs(2546)));
    outputs(790) <= (layer2_outputs(3138)) and (layer2_outputs(4514));
    outputs(791) <= not((layer2_outputs(1939)) or (layer2_outputs(334)));
    outputs(792) <= layer2_outputs(4158);
    outputs(793) <= not(layer2_outputs(1720)) or (layer2_outputs(990));
    outputs(794) <= (layer2_outputs(3321)) and not (layer2_outputs(619));
    outputs(795) <= not((layer2_outputs(2342)) or (layer2_outputs(1488)));
    outputs(796) <= (layer2_outputs(4313)) and (layer2_outputs(672));
    outputs(797) <= (layer2_outputs(859)) xor (layer2_outputs(842));
    outputs(798) <= not(layer2_outputs(2480));
    outputs(799) <= (layer2_outputs(1324)) and (layer2_outputs(4770));
    outputs(800) <= not(layer2_outputs(1308));
    outputs(801) <= not(layer2_outputs(1811));
    outputs(802) <= (layer2_outputs(613)) and not (layer2_outputs(1122));
    outputs(803) <= (layer2_outputs(3965)) and (layer2_outputs(2991));
    outputs(804) <= not(layer2_outputs(4378));
    outputs(805) <= (layer2_outputs(2266)) and (layer2_outputs(2404));
    outputs(806) <= not(layer2_outputs(2448));
    outputs(807) <= '0';
    outputs(808) <= layer2_outputs(160);
    outputs(809) <= layer2_outputs(4882);
    outputs(810) <= layer2_outputs(3742);
    outputs(811) <= (layer2_outputs(1926)) and (layer2_outputs(425));
    outputs(812) <= (layer2_outputs(614)) and not (layer2_outputs(457));
    outputs(813) <= not(layer2_outputs(5113));
    outputs(814) <= (layer2_outputs(1360)) and not (layer2_outputs(82));
    outputs(815) <= not((layer2_outputs(3106)) xor (layer2_outputs(1873)));
    outputs(816) <= (layer2_outputs(964)) and not (layer2_outputs(589));
    outputs(817) <= layer2_outputs(3066);
    outputs(818) <= not((layer2_outputs(156)) or (layer2_outputs(3100)));
    outputs(819) <= layer2_outputs(5075);
    outputs(820) <= (layer2_outputs(3161)) and (layer2_outputs(353));
    outputs(821) <= not((layer2_outputs(3166)) xor (layer2_outputs(3876)));
    outputs(822) <= layer2_outputs(1691);
    outputs(823) <= (layer2_outputs(3513)) and not (layer2_outputs(473));
    outputs(824) <= (layer2_outputs(3584)) and not (layer2_outputs(1447));
    outputs(825) <= not((layer2_outputs(4146)) or (layer2_outputs(1383)));
    outputs(826) <= (layer2_outputs(2854)) xor (layer2_outputs(1796));
    outputs(827) <= not(layer2_outputs(3428));
    outputs(828) <= (layer2_outputs(240)) and (layer2_outputs(3697));
    outputs(829) <= not(layer2_outputs(3198));
    outputs(830) <= (layer2_outputs(1021)) and not (layer2_outputs(3793));
    outputs(831) <= layer2_outputs(2008);
    outputs(832) <= (layer2_outputs(1683)) and not (layer2_outputs(1351));
    outputs(833) <= (layer2_outputs(4118)) and not (layer2_outputs(1273));
    outputs(834) <= (layer2_outputs(3664)) and (layer2_outputs(3235));
    outputs(835) <= (layer2_outputs(1141)) and not (layer2_outputs(4646));
    outputs(836) <= (layer2_outputs(3814)) and not (layer2_outputs(333));
    outputs(837) <= (layer2_outputs(2681)) and not (layer2_outputs(3426));
    outputs(838) <= (layer2_outputs(305)) and not (layer2_outputs(3527));
    outputs(839) <= (layer2_outputs(2352)) and not (layer2_outputs(716));
    outputs(840) <= (layer2_outputs(1636)) and not (layer2_outputs(1907));
    outputs(841) <= layer2_outputs(183);
    outputs(842) <= not(layer2_outputs(1050));
    outputs(843) <= not(layer2_outputs(2160));
    outputs(844) <= not(layer2_outputs(460));
    outputs(845) <= (layer2_outputs(2796)) and not (layer2_outputs(1465));
    outputs(846) <= (layer2_outputs(2178)) and not (layer2_outputs(427));
    outputs(847) <= (layer2_outputs(2779)) and (layer2_outputs(3607));
    outputs(848) <= layer2_outputs(509);
    outputs(849) <= not((layer2_outputs(4801)) or (layer2_outputs(1591)));
    outputs(850) <= not(layer2_outputs(2355));
    outputs(851) <= layer2_outputs(4664);
    outputs(852) <= not(layer2_outputs(3987));
    outputs(853) <= (layer2_outputs(3344)) and not (layer2_outputs(2372));
    outputs(854) <= layer2_outputs(1420);
    outputs(855) <= not((layer2_outputs(277)) or (layer2_outputs(128)));
    outputs(856) <= not(layer2_outputs(3500));
    outputs(857) <= (layer2_outputs(3722)) and not (layer2_outputs(1293));
    outputs(858) <= (layer2_outputs(1373)) and not (layer2_outputs(65));
    outputs(859) <= layer2_outputs(4020);
    outputs(860) <= layer2_outputs(3501);
    outputs(861) <= (layer2_outputs(6)) and (layer2_outputs(263));
    outputs(862) <= not(layer2_outputs(4501));
    outputs(863) <= (layer2_outputs(3848)) and not (layer2_outputs(2693));
    outputs(864) <= not((layer2_outputs(1519)) or (layer2_outputs(2950)));
    outputs(865) <= (layer2_outputs(3874)) and not (layer2_outputs(2210));
    outputs(866) <= not(layer2_outputs(2972));
    outputs(867) <= not((layer2_outputs(4655)) or (layer2_outputs(3092)));
    outputs(868) <= not(layer2_outputs(4263));
    outputs(869) <= not(layer2_outputs(3632));
    outputs(870) <= not((layer2_outputs(3144)) or (layer2_outputs(3899)));
    outputs(871) <= not(layer2_outputs(3110));
    outputs(872) <= not(layer2_outputs(2274));
    outputs(873) <= not(layer2_outputs(556));
    outputs(874) <= (layer2_outputs(883)) and not (layer2_outputs(2836));
    outputs(875) <= layer2_outputs(3415);
    outputs(876) <= (layer2_outputs(4927)) and not (layer2_outputs(2380));
    outputs(877) <= not(layer2_outputs(333));
    outputs(878) <= not((layer2_outputs(2505)) xor (layer2_outputs(4163)));
    outputs(879) <= not(layer2_outputs(1344));
    outputs(880) <= layer2_outputs(4406);
    outputs(881) <= layer2_outputs(3662);
    outputs(882) <= layer2_outputs(3893);
    outputs(883) <= (layer2_outputs(1087)) and not (layer2_outputs(113));
    outputs(884) <= not(layer2_outputs(3651));
    outputs(885) <= not(layer2_outputs(2644));
    outputs(886) <= layer2_outputs(4767);
    outputs(887) <= layer2_outputs(3423);
    outputs(888) <= layer2_outputs(4967);
    outputs(889) <= not(layer2_outputs(1564));
    outputs(890) <= not(layer2_outputs(1966));
    outputs(891) <= layer2_outputs(4597);
    outputs(892) <= (layer2_outputs(4234)) and (layer2_outputs(1076));
    outputs(893) <= not(layer2_outputs(2964)) or (layer2_outputs(2136));
    outputs(894) <= not(layer2_outputs(982));
    outputs(895) <= (layer2_outputs(3829)) xor (layer2_outputs(622));
    outputs(896) <= not(layer2_outputs(3103));
    outputs(897) <= not(layer2_outputs(2657));
    outputs(898) <= layer2_outputs(172);
    outputs(899) <= not(layer2_outputs(3475));
    outputs(900) <= (layer2_outputs(3005)) and (layer2_outputs(1548));
    outputs(901) <= (layer2_outputs(1131)) and not (layer2_outputs(723));
    outputs(902) <= (layer2_outputs(494)) or (layer2_outputs(4375));
    outputs(903) <= (layer2_outputs(1968)) or (layer2_outputs(134));
    outputs(904) <= not(layer2_outputs(1785));
    outputs(905) <= not(layer2_outputs(1397));
    outputs(906) <= not(layer2_outputs(4577));
    outputs(907) <= (layer2_outputs(4455)) and not (layer2_outputs(4752));
    outputs(908) <= not(layer2_outputs(2956));
    outputs(909) <= (layer2_outputs(3609)) xor (layer2_outputs(1870));
    outputs(910) <= not((layer2_outputs(4862)) or (layer2_outputs(3191)));
    outputs(911) <= not((layer2_outputs(3264)) or (layer2_outputs(2965)));
    outputs(912) <= not(layer2_outputs(2230));
    outputs(913) <= layer2_outputs(3436);
    outputs(914) <= not(layer2_outputs(2673));
    outputs(915) <= not(layer2_outputs(4859));
    outputs(916) <= layer2_outputs(1738);
    outputs(917) <= (layer2_outputs(4243)) and (layer2_outputs(2834));
    outputs(918) <= not(layer2_outputs(1336));
    outputs(919) <= not(layer2_outputs(3457));
    outputs(920) <= layer2_outputs(4191);
    outputs(921) <= layer2_outputs(1586);
    outputs(922) <= layer2_outputs(3252);
    outputs(923) <= not(layer2_outputs(2626));
    outputs(924) <= (layer2_outputs(4336)) and not (layer2_outputs(84));
    outputs(925) <= (layer2_outputs(4316)) and not (layer2_outputs(2314));
    outputs(926) <= layer2_outputs(2275);
    outputs(927) <= not((layer2_outputs(560)) or (layer2_outputs(3256)));
    outputs(928) <= not(layer2_outputs(2236));
    outputs(929) <= layer2_outputs(2987);
    outputs(930) <= (layer2_outputs(3048)) and not (layer2_outputs(4903));
    outputs(931) <= (layer2_outputs(1478)) and not (layer2_outputs(3870));
    outputs(932) <= (layer2_outputs(1870)) xor (layer2_outputs(4359));
    outputs(933) <= not(layer2_outputs(4763));
    outputs(934) <= not(layer2_outputs(2212));
    outputs(935) <= not((layer2_outputs(4146)) or (layer2_outputs(4126)));
    outputs(936) <= layer2_outputs(3689);
    outputs(937) <= (layer2_outputs(843)) and (layer2_outputs(737));
    outputs(938) <= not(layer2_outputs(2632));
    outputs(939) <= (layer2_outputs(3944)) and not (layer2_outputs(4557));
    outputs(940) <= not(layer2_outputs(3190));
    outputs(941) <= not((layer2_outputs(3623)) xor (layer2_outputs(4959)));
    outputs(942) <= not(layer2_outputs(2421));
    outputs(943) <= not(layer2_outputs(484));
    outputs(944) <= (layer2_outputs(4388)) or (layer2_outputs(3295));
    outputs(945) <= (layer2_outputs(3742)) and (layer2_outputs(515));
    outputs(946) <= (layer2_outputs(960)) and not (layer2_outputs(2607));
    outputs(947) <= (layer2_outputs(2162)) and not (layer2_outputs(2633));
    outputs(948) <= not((layer2_outputs(2212)) or (layer2_outputs(560)));
    outputs(949) <= not(layer2_outputs(1180));
    outputs(950) <= (layer2_outputs(1470)) and not (layer2_outputs(4034));
    outputs(951) <= layer2_outputs(3699);
    outputs(952) <= layer2_outputs(5095);
    outputs(953) <= not(layer2_outputs(1771));
    outputs(954) <= layer2_outputs(3802);
    outputs(955) <= layer2_outputs(1381);
    outputs(956) <= layer2_outputs(3564);
    outputs(957) <= not(layer2_outputs(1842));
    outputs(958) <= not(layer2_outputs(2858));
    outputs(959) <= layer2_outputs(2629);
    outputs(960) <= layer2_outputs(916);
    outputs(961) <= not((layer2_outputs(4945)) or (layer2_outputs(2788)));
    outputs(962) <= not((layer2_outputs(1299)) or (layer2_outputs(755)));
    outputs(963) <= not((layer2_outputs(2094)) and (layer2_outputs(5019)));
    outputs(964) <= layer2_outputs(3280);
    outputs(965) <= not(layer2_outputs(2890));
    outputs(966) <= not(layer2_outputs(3392));
    outputs(967) <= (layer2_outputs(819)) xor (layer2_outputs(549));
    outputs(968) <= layer2_outputs(3142);
    outputs(969) <= not(layer2_outputs(5056));
    outputs(970) <= (layer2_outputs(2823)) and (layer2_outputs(2605));
    outputs(971) <= not((layer2_outputs(1428)) xor (layer2_outputs(1435)));
    outputs(972) <= (layer2_outputs(2400)) and (layer2_outputs(4495));
    outputs(973) <= not((layer2_outputs(4044)) or (layer2_outputs(1113)));
    outputs(974) <= not(layer2_outputs(2538));
    outputs(975) <= not(layer2_outputs(487));
    outputs(976) <= not((layer2_outputs(2831)) xor (layer2_outputs(3176)));
    outputs(977) <= layer2_outputs(4344);
    outputs(978) <= layer2_outputs(4738);
    outputs(979) <= not(layer2_outputs(5101));
    outputs(980) <= not(layer2_outputs(1736));
    outputs(981) <= (layer2_outputs(3319)) and not (layer2_outputs(4555));
    outputs(982) <= layer2_outputs(3665);
    outputs(983) <= not(layer2_outputs(1429));
    outputs(984) <= not((layer2_outputs(2535)) xor (layer2_outputs(468)));
    outputs(985) <= layer2_outputs(2519);
    outputs(986) <= layer2_outputs(2341);
    outputs(987) <= layer2_outputs(2816);
    outputs(988) <= not((layer2_outputs(3793)) or (layer2_outputs(3531)));
    outputs(989) <= layer2_outputs(2153);
    outputs(990) <= (layer2_outputs(3143)) or (layer2_outputs(4393));
    outputs(991) <= not(layer2_outputs(987));
    outputs(992) <= (layer2_outputs(4604)) and (layer2_outputs(2162));
    outputs(993) <= layer2_outputs(520);
    outputs(994) <= layer2_outputs(3181);
    outputs(995) <= not(layer2_outputs(4201));
    outputs(996) <= not((layer2_outputs(4656)) or (layer2_outputs(1832)));
    outputs(997) <= not((layer2_outputs(836)) xor (layer2_outputs(156)));
    outputs(998) <= (layer2_outputs(2940)) and not (layer2_outputs(2081));
    outputs(999) <= not(layer2_outputs(1463)) or (layer2_outputs(4314));
    outputs(1000) <= not(layer2_outputs(1713));
    outputs(1001) <= (layer2_outputs(210)) and (layer2_outputs(702));
    outputs(1002) <= not((layer2_outputs(3100)) or (layer2_outputs(760)));
    outputs(1003) <= (layer2_outputs(3237)) and not (layer2_outputs(4060));
    outputs(1004) <= (layer2_outputs(3615)) or (layer2_outputs(2732));
    outputs(1005) <= layer2_outputs(491);
    outputs(1006) <= (layer2_outputs(2674)) and not (layer2_outputs(3269));
    outputs(1007) <= not(layer2_outputs(1688));
    outputs(1008) <= not(layer2_outputs(410));
    outputs(1009) <= (layer2_outputs(1325)) and (layer2_outputs(1284));
    outputs(1010) <= layer2_outputs(2025);
    outputs(1011) <= (layer2_outputs(4827)) and not (layer2_outputs(41));
    outputs(1012) <= (layer2_outputs(3422)) and not (layer2_outputs(4174));
    outputs(1013) <= (layer2_outputs(2437)) and not (layer2_outputs(254));
    outputs(1014) <= (layer2_outputs(3758)) and (layer2_outputs(1571));
    outputs(1015) <= layer2_outputs(2337);
    outputs(1016) <= not(layer2_outputs(2903));
    outputs(1017) <= layer2_outputs(1659);
    outputs(1018) <= layer2_outputs(4440);
    outputs(1019) <= not((layer2_outputs(599)) xor (layer2_outputs(1676)));
    outputs(1020) <= (layer2_outputs(1435)) and (layer2_outputs(4124));
    outputs(1021) <= layer2_outputs(2381);
    outputs(1022) <= (layer2_outputs(2389)) and (layer2_outputs(4909));
    outputs(1023) <= layer2_outputs(4880);
    outputs(1024) <= not((layer2_outputs(4035)) and (layer2_outputs(3474)));
    outputs(1025) <= layer2_outputs(591);
    outputs(1026) <= (layer2_outputs(2770)) and not (layer2_outputs(3504));
    outputs(1027) <= (layer2_outputs(3861)) and not (layer2_outputs(4226));
    outputs(1028) <= not(layer2_outputs(1177));
    outputs(1029) <= not((layer2_outputs(438)) xor (layer2_outputs(4849)));
    outputs(1030) <= not(layer2_outputs(2004));
    outputs(1031) <= layer2_outputs(4765);
    outputs(1032) <= not(layer2_outputs(3222));
    outputs(1033) <= layer2_outputs(4056);
    outputs(1034) <= not(layer2_outputs(1786));
    outputs(1035) <= layer2_outputs(1744);
    outputs(1036) <= not((layer2_outputs(3153)) and (layer2_outputs(3779)));
    outputs(1037) <= layer2_outputs(1420);
    outputs(1038) <= layer2_outputs(1265);
    outputs(1039) <= not(layer2_outputs(1576));
    outputs(1040) <= not(layer2_outputs(4392));
    outputs(1041) <= not(layer2_outputs(738));
    outputs(1042) <= not(layer2_outputs(1027));
    outputs(1043) <= not(layer2_outputs(412));
    outputs(1044) <= layer2_outputs(2328);
    outputs(1045) <= not(layer2_outputs(3092));
    outputs(1046) <= not(layer2_outputs(976));
    outputs(1047) <= not(layer2_outputs(3060)) or (layer2_outputs(2018));
    outputs(1048) <= not((layer2_outputs(1541)) xor (layer2_outputs(4168)));
    outputs(1049) <= (layer2_outputs(350)) and not (layer2_outputs(1822));
    outputs(1050) <= not(layer2_outputs(3687)) or (layer2_outputs(4556));
    outputs(1051) <= layer2_outputs(3625);
    outputs(1052) <= layer2_outputs(1020);
    outputs(1053) <= layer2_outputs(1946);
    outputs(1054) <= not((layer2_outputs(246)) xor (layer2_outputs(4065)));
    outputs(1055) <= layer2_outputs(4289);
    outputs(1056) <= (layer2_outputs(2464)) and (layer2_outputs(159));
    outputs(1057) <= not(layer2_outputs(2699));
    outputs(1058) <= not(layer2_outputs(372));
    outputs(1059) <= layer2_outputs(2710);
    outputs(1060) <= not((layer2_outputs(1052)) xor (layer2_outputs(2891)));
    outputs(1061) <= not(layer2_outputs(1814));
    outputs(1062) <= layer2_outputs(4374);
    outputs(1063) <= not(layer2_outputs(3427));
    outputs(1064) <= layer2_outputs(4874);
    outputs(1065) <= layer2_outputs(867);
    outputs(1066) <= not((layer2_outputs(2423)) xor (layer2_outputs(2145)));
    outputs(1067) <= layer2_outputs(3050);
    outputs(1068) <= not(layer2_outputs(1594)) or (layer2_outputs(3477));
    outputs(1069) <= not(layer2_outputs(3489)) or (layer2_outputs(3359));
    outputs(1070) <= not(layer2_outputs(4135));
    outputs(1071) <= layer2_outputs(119);
    outputs(1072) <= layer2_outputs(622);
    outputs(1073) <= layer2_outputs(842);
    outputs(1074) <= not(layer2_outputs(4820));
    outputs(1075) <= layer2_outputs(3534);
    outputs(1076) <= layer2_outputs(2806);
    outputs(1077) <= (layer2_outputs(2462)) and (layer2_outputs(0));
    outputs(1078) <= (layer2_outputs(3496)) and not (layer2_outputs(3887));
    outputs(1079) <= not(layer2_outputs(3201));
    outputs(1080) <= layer2_outputs(3230);
    outputs(1081) <= not(layer2_outputs(3803));
    outputs(1082) <= not(layer2_outputs(4575));
    outputs(1083) <= not(layer2_outputs(1786));
    outputs(1084) <= (layer2_outputs(943)) and not (layer2_outputs(4063));
    outputs(1085) <= not(layer2_outputs(2248));
    outputs(1086) <= (layer2_outputs(3726)) and not (layer2_outputs(1068));
    outputs(1087) <= layer2_outputs(2971);
    outputs(1088) <= layer2_outputs(4009);
    outputs(1089) <= layer2_outputs(40);
    outputs(1090) <= layer2_outputs(3806);
    outputs(1091) <= layer2_outputs(547);
    outputs(1092) <= layer2_outputs(769);
    outputs(1093) <= not((layer2_outputs(4943)) xor (layer2_outputs(2814)));
    outputs(1094) <= not(layer2_outputs(4094));
    outputs(1095) <= not((layer2_outputs(3307)) xor (layer2_outputs(1655)));
    outputs(1096) <= not(layer2_outputs(1167));
    outputs(1097) <= not(layer2_outputs(612));
    outputs(1098) <= layer2_outputs(3022);
    outputs(1099) <= layer2_outputs(2284);
    outputs(1100) <= layer2_outputs(4378);
    outputs(1101) <= (layer2_outputs(4152)) and not (layer2_outputs(1272));
    outputs(1102) <= layer2_outputs(3809);
    outputs(1103) <= not(layer2_outputs(1012));
    outputs(1104) <= (layer2_outputs(1520)) xor (layer2_outputs(4092));
    outputs(1105) <= not(layer2_outputs(1362)) or (layer2_outputs(706));
    outputs(1106) <= layer2_outputs(1116);
    outputs(1107) <= not(layer2_outputs(5035));
    outputs(1108) <= not(layer2_outputs(1177)) or (layer2_outputs(2647));
    outputs(1109) <= layer2_outputs(1516);
    outputs(1110) <= not(layer2_outputs(2614));
    outputs(1111) <= (layer2_outputs(4713)) or (layer2_outputs(3651));
    outputs(1112) <= layer2_outputs(4760);
    outputs(1113) <= not(layer2_outputs(1761));
    outputs(1114) <= layer2_outputs(1145);
    outputs(1115) <= (layer2_outputs(1577)) and (layer2_outputs(344));
    outputs(1116) <= (layer2_outputs(1991)) xor (layer2_outputs(384));
    outputs(1117) <= (layer2_outputs(4237)) and not (layer2_outputs(3428));
    outputs(1118) <= not(layer2_outputs(2231));
    outputs(1119) <= layer2_outputs(1189);
    outputs(1120) <= layer2_outputs(2291);
    outputs(1121) <= (layer2_outputs(2452)) or (layer2_outputs(3540));
    outputs(1122) <= not((layer2_outputs(131)) xor (layer2_outputs(1253)));
    outputs(1123) <= layer2_outputs(3425);
    outputs(1124) <= layer2_outputs(463);
    outputs(1125) <= layer2_outputs(1780);
    outputs(1126) <= not((layer2_outputs(3098)) and (layer2_outputs(1165)));
    outputs(1127) <= layer2_outputs(3653);
    outputs(1128) <= layer2_outputs(1402);
    outputs(1129) <= not((layer2_outputs(1649)) or (layer2_outputs(2136)));
    outputs(1130) <= layer2_outputs(2910);
    outputs(1131) <= layer2_outputs(3649);
    outputs(1132) <= not(layer2_outputs(2564));
    outputs(1133) <= not(layer2_outputs(4620));
    outputs(1134) <= (layer2_outputs(1661)) and not (layer2_outputs(796));
    outputs(1135) <= layer2_outputs(4485);
    outputs(1136) <= not(layer2_outputs(3326));
    outputs(1137) <= layer2_outputs(1532);
    outputs(1138) <= layer2_outputs(4592);
    outputs(1139) <= not((layer2_outputs(2123)) xor (layer2_outputs(2726)));
    outputs(1140) <= (layer2_outputs(2145)) xor (layer2_outputs(1672));
    outputs(1141) <= layer2_outputs(4506);
    outputs(1142) <= not(layer2_outputs(3271));
    outputs(1143) <= layer2_outputs(4441);
    outputs(1144) <= not(layer2_outputs(2441));
    outputs(1145) <= not((layer2_outputs(2393)) xor (layer2_outputs(4553)));
    outputs(1146) <= (layer2_outputs(4361)) xor (layer2_outputs(2956));
    outputs(1147) <= layer2_outputs(4276);
    outputs(1148) <= layer2_outputs(2760);
    outputs(1149) <= layer2_outputs(5036);
    outputs(1150) <= layer2_outputs(3381);
    outputs(1151) <= not(layer2_outputs(1636));
    outputs(1152) <= not(layer2_outputs(1569));
    outputs(1153) <= layer2_outputs(3542);
    outputs(1154) <= not(layer2_outputs(4667));
    outputs(1155) <= layer2_outputs(4760);
    outputs(1156) <= (layer2_outputs(522)) xor (layer2_outputs(3141));
    outputs(1157) <= not(layer2_outputs(588));
    outputs(1158) <= layer2_outputs(1457);
    outputs(1159) <= layer2_outputs(1754);
    outputs(1160) <= layer2_outputs(2675);
    outputs(1161) <= not(layer2_outputs(4442));
    outputs(1162) <= layer2_outputs(1154);
    outputs(1163) <= not(layer2_outputs(567)) or (layer2_outputs(2188));
    outputs(1164) <= not((layer2_outputs(2607)) xor (layer2_outputs(1850)));
    outputs(1165) <= not(layer2_outputs(4674));
    outputs(1166) <= not(layer2_outputs(3834));
    outputs(1167) <= not(layer2_outputs(3430));
    outputs(1168) <= not(layer2_outputs(251)) or (layer2_outputs(572));
    outputs(1169) <= not(layer2_outputs(614));
    outputs(1170) <= not((layer2_outputs(744)) and (layer2_outputs(843)));
    outputs(1171) <= layer2_outputs(4202);
    outputs(1172) <= not(layer2_outputs(3333));
    outputs(1173) <= not(layer2_outputs(111));
    outputs(1174) <= layer2_outputs(3264);
    outputs(1175) <= not(layer2_outputs(4856));
    outputs(1176) <= layer2_outputs(1341);
    outputs(1177) <= not(layer2_outputs(4563));
    outputs(1178) <= not((layer2_outputs(169)) xor (layer2_outputs(3537)));
    outputs(1179) <= not((layer2_outputs(4903)) xor (layer2_outputs(2114)));
    outputs(1180) <= (layer2_outputs(170)) and (layer2_outputs(119));
    outputs(1181) <= layer2_outputs(2292);
    outputs(1182) <= (layer2_outputs(2876)) and (layer2_outputs(285));
    outputs(1183) <= not((layer2_outputs(5076)) or (layer2_outputs(4870)));
    outputs(1184) <= layer2_outputs(2474);
    outputs(1185) <= layer2_outputs(4603);
    outputs(1186) <= not(layer2_outputs(2029));
    outputs(1187) <= layer2_outputs(5030);
    outputs(1188) <= layer2_outputs(3089);
    outputs(1189) <= layer2_outputs(1980);
    outputs(1190) <= not(layer2_outputs(3024));
    outputs(1191) <= not((layer2_outputs(1281)) or (layer2_outputs(3129)));
    outputs(1192) <= not(layer2_outputs(744));
    outputs(1193) <= (layer2_outputs(1720)) and (layer2_outputs(1168));
    outputs(1194) <= not(layer2_outputs(2696)) or (layer2_outputs(3225));
    outputs(1195) <= layer2_outputs(4590);
    outputs(1196) <= not(layer2_outputs(4117)) or (layer2_outputs(3536));
    outputs(1197) <= not(layer2_outputs(4481));
    outputs(1198) <= layer2_outputs(1417);
    outputs(1199) <= layer2_outputs(1895);
    outputs(1200) <= layer2_outputs(3634);
    outputs(1201) <= (layer2_outputs(1434)) xor (layer2_outputs(3713));
    outputs(1202) <= not(layer2_outputs(4290)) or (layer2_outputs(90));
    outputs(1203) <= (layer2_outputs(4258)) or (layer2_outputs(2006));
    outputs(1204) <= layer2_outputs(3438);
    outputs(1205) <= not(layer2_outputs(3011)) or (layer2_outputs(1322));
    outputs(1206) <= layer2_outputs(343);
    outputs(1207) <= not(layer2_outputs(4296));
    outputs(1208) <= not(layer2_outputs(910)) or (layer2_outputs(1682));
    outputs(1209) <= layer2_outputs(1098);
    outputs(1210) <= not((layer2_outputs(1608)) xor (layer2_outputs(3943)));
    outputs(1211) <= layer2_outputs(1001);
    outputs(1212) <= layer2_outputs(3188);
    outputs(1213) <= layer2_outputs(4905);
    outputs(1214) <= not(layer2_outputs(1994));
    outputs(1215) <= not((layer2_outputs(558)) or (layer2_outputs(2197)));
    outputs(1216) <= layer2_outputs(1148);
    outputs(1217) <= layer2_outputs(1936);
    outputs(1218) <= not(layer2_outputs(939));
    outputs(1219) <= not((layer2_outputs(1181)) and (layer2_outputs(3709)));
    outputs(1220) <= not((layer2_outputs(3485)) xor (layer2_outputs(4304)));
    outputs(1221) <= not((layer2_outputs(1089)) or (layer2_outputs(3736)));
    outputs(1222) <= (layer2_outputs(2898)) and not (layer2_outputs(3640));
    outputs(1223) <= not(layer2_outputs(3820));
    outputs(1224) <= not(layer2_outputs(4411));
    outputs(1225) <= not(layer2_outputs(442));
    outputs(1226) <= layer2_outputs(2002);
    outputs(1227) <= not(layer2_outputs(4070));
    outputs(1228) <= (layer2_outputs(499)) xor (layer2_outputs(2070));
    outputs(1229) <= layer2_outputs(4105);
    outputs(1230) <= not(layer2_outputs(3601));
    outputs(1231) <= not(layer2_outputs(2619)) or (layer2_outputs(881));
    outputs(1232) <= (layer2_outputs(988)) xor (layer2_outputs(629));
    outputs(1233) <= layer2_outputs(4408);
    outputs(1234) <= layer2_outputs(3919);
    outputs(1235) <= layer2_outputs(1848);
    outputs(1236) <= not(layer2_outputs(2301));
    outputs(1237) <= not((layer2_outputs(2674)) xor (layer2_outputs(455)));
    outputs(1238) <= layer2_outputs(725);
    outputs(1239) <= layer2_outputs(618);
    outputs(1240) <= not(layer2_outputs(2944));
    outputs(1241) <= (layer2_outputs(3513)) and not (layer2_outputs(4309));
    outputs(1242) <= not(layer2_outputs(2463));
    outputs(1243) <= not(layer2_outputs(5032));
    outputs(1244) <= layer2_outputs(1461);
    outputs(1245) <= not(layer2_outputs(2055));
    outputs(1246) <= not(layer2_outputs(1776));
    outputs(1247) <= layer2_outputs(5037);
    outputs(1248) <= not(layer2_outputs(4494));
    outputs(1249) <= not(layer2_outputs(2544));
    outputs(1250) <= not(layer2_outputs(143));
    outputs(1251) <= not((layer2_outputs(4491)) or (layer2_outputs(2356)));
    outputs(1252) <= layer2_outputs(2395);
    outputs(1253) <= layer2_outputs(2817);
    outputs(1254) <= not(layer2_outputs(314));
    outputs(1255) <= (layer2_outputs(1522)) xor (layer2_outputs(196));
    outputs(1256) <= layer2_outputs(2211);
    outputs(1257) <= not((layer2_outputs(53)) xor (layer2_outputs(3178)));
    outputs(1258) <= layer2_outputs(4360);
    outputs(1259) <= layer2_outputs(1007);
    outputs(1260) <= layer2_outputs(362);
    outputs(1261) <= layer2_outputs(521);
    outputs(1262) <= (layer2_outputs(513)) and not (layer2_outputs(4302));
    outputs(1263) <= not(layer2_outputs(3957));
    outputs(1264) <= (layer2_outputs(4098)) and (layer2_outputs(1108));
    outputs(1265) <= layer2_outputs(4100);
    outputs(1266) <= layer2_outputs(4964);
    outputs(1267) <= not(layer2_outputs(3353));
    outputs(1268) <= layer2_outputs(3519);
    outputs(1269) <= not(layer2_outputs(3015));
    outputs(1270) <= not((layer2_outputs(4591)) and (layer2_outputs(1208)));
    outputs(1271) <= not(layer2_outputs(2745));
    outputs(1272) <= not(layer2_outputs(3070));
    outputs(1273) <= (layer2_outputs(3263)) and (layer2_outputs(2243));
    outputs(1274) <= not(layer2_outputs(2021)) or (layer2_outputs(3332));
    outputs(1275) <= (layer2_outputs(3539)) xor (layer2_outputs(949));
    outputs(1276) <= (layer2_outputs(1213)) and not (layer2_outputs(1528));
    outputs(1277) <= not((layer2_outputs(3435)) xor (layer2_outputs(577)));
    outputs(1278) <= not(layer2_outputs(3278));
    outputs(1279) <= not(layer2_outputs(29));
    outputs(1280) <= not(layer2_outputs(733));
    outputs(1281) <= not((layer2_outputs(1694)) or (layer2_outputs(3323)));
    outputs(1282) <= not(layer2_outputs(4558)) or (layer2_outputs(1846));
    outputs(1283) <= layer2_outputs(1551);
    outputs(1284) <= (layer2_outputs(259)) and not (layer2_outputs(4197));
    outputs(1285) <= layer2_outputs(1214);
    outputs(1286) <= layer2_outputs(4003);
    outputs(1287) <= not(layer2_outputs(1564));
    outputs(1288) <= layer2_outputs(4253);
    outputs(1289) <= layer2_outputs(2451);
    outputs(1290) <= not((layer2_outputs(3767)) or (layer2_outputs(757)));
    outputs(1291) <= not((layer2_outputs(2174)) xor (layer2_outputs(929)));
    outputs(1292) <= not((layer2_outputs(1006)) or (layer2_outputs(2500)));
    outputs(1293) <= layer2_outputs(1816);
    outputs(1294) <= layer2_outputs(1524);
    outputs(1295) <= not(layer2_outputs(2228));
    outputs(1296) <= (layer2_outputs(4600)) xor (layer2_outputs(1010));
    outputs(1297) <= layer2_outputs(1331);
    outputs(1298) <= (layer2_outputs(328)) and not (layer2_outputs(4413));
    outputs(1299) <= layer2_outputs(2452);
    outputs(1300) <= not(layer2_outputs(4166));
    outputs(1301) <= (layer2_outputs(1353)) or (layer2_outputs(3492));
    outputs(1302) <= not(layer2_outputs(3430));
    outputs(1303) <= layer2_outputs(3358);
    outputs(1304) <= (layer2_outputs(653)) and (layer2_outputs(743));
    outputs(1305) <= (layer2_outputs(1766)) xor (layer2_outputs(2418));
    outputs(1306) <= layer2_outputs(213);
    outputs(1307) <= (layer2_outputs(336)) and not (layer2_outputs(813));
    outputs(1308) <= layer2_outputs(3003);
    outputs(1309) <= layer2_outputs(1848);
    outputs(1310) <= layer2_outputs(4082);
    outputs(1311) <= layer2_outputs(1893);
    outputs(1312) <= not(layer2_outputs(3892));
    outputs(1313) <= not(layer2_outputs(2429));
    outputs(1314) <= layer2_outputs(4265);
    outputs(1315) <= layer2_outputs(4625);
    outputs(1316) <= not(layer2_outputs(1006));
    outputs(1317) <= layer2_outputs(5002);
    outputs(1318) <= (layer2_outputs(4152)) and not (layer2_outputs(656));
    outputs(1319) <= not(layer2_outputs(1369));
    outputs(1320) <= not(layer2_outputs(4866));
    outputs(1321) <= not(layer2_outputs(387));
    outputs(1322) <= not(layer2_outputs(2871));
    outputs(1323) <= layer2_outputs(3655);
    outputs(1324) <= layer2_outputs(4749);
    outputs(1325) <= layer2_outputs(2513);
    outputs(1326) <= layer2_outputs(1827);
    outputs(1327) <= not(layer2_outputs(3613)) or (layer2_outputs(520));
    outputs(1328) <= (layer2_outputs(4253)) and not (layer2_outputs(2225));
    outputs(1329) <= not(layer2_outputs(4684)) or (layer2_outputs(1904));
    outputs(1330) <= layer2_outputs(525);
    outputs(1331) <= layer2_outputs(2314);
    outputs(1332) <= not(layer2_outputs(2865));
    outputs(1333) <= not(layer2_outputs(2572));
    outputs(1334) <= layer2_outputs(774);
    outputs(1335) <= not(layer2_outputs(1252));
    outputs(1336) <= not(layer2_outputs(2577));
    outputs(1337) <= layer2_outputs(4069);
    outputs(1338) <= (layer2_outputs(2492)) or (layer2_outputs(303));
    outputs(1339) <= (layer2_outputs(4060)) or (layer2_outputs(493));
    outputs(1340) <= not((layer2_outputs(4452)) xor (layer2_outputs(2436)));
    outputs(1341) <= not((layer2_outputs(332)) xor (layer2_outputs(2303)));
    outputs(1342) <= not((layer2_outputs(2530)) xor (layer2_outputs(4375)));
    outputs(1343) <= not(layer2_outputs(4591)) or (layer2_outputs(2579));
    outputs(1344) <= layer2_outputs(3281);
    outputs(1345) <= (layer2_outputs(3388)) xor (layer2_outputs(216));
    outputs(1346) <= not((layer2_outputs(402)) xor (layer2_outputs(4295)));
    outputs(1347) <= layer2_outputs(86);
    outputs(1348) <= layer2_outputs(1861);
    outputs(1349) <= not((layer2_outputs(2527)) and (layer2_outputs(1207)));
    outputs(1350) <= not(layer2_outputs(4972));
    outputs(1351) <= not(layer2_outputs(1542));
    outputs(1352) <= not(layer2_outputs(2685)) or (layer2_outputs(1094));
    outputs(1353) <= layer2_outputs(4346);
    outputs(1354) <= not(layer2_outputs(2142)) or (layer2_outputs(2862));
    outputs(1355) <= not(layer2_outputs(280));
    outputs(1356) <= not(layer2_outputs(1540));
    outputs(1357) <= not(layer2_outputs(942));
    outputs(1358) <= not((layer2_outputs(5074)) or (layer2_outputs(1191)));
    outputs(1359) <= not(layer2_outputs(273));
    outputs(1360) <= not(layer2_outputs(3340));
    outputs(1361) <= not(layer2_outputs(2354));
    outputs(1362) <= not(layer2_outputs(1523));
    outputs(1363) <= not(layer2_outputs(4547)) or (layer2_outputs(1103));
    outputs(1364) <= not(layer2_outputs(831)) or (layer2_outputs(1504));
    outputs(1365) <= not(layer2_outputs(1432));
    outputs(1366) <= layer2_outputs(1114);
    outputs(1367) <= (layer2_outputs(3090)) and not (layer2_outputs(4188));
    outputs(1368) <= layer2_outputs(4936);
    outputs(1369) <= layer2_outputs(1682);
    outputs(1370) <= not((layer2_outputs(766)) or (layer2_outputs(1328)));
    outputs(1371) <= layer2_outputs(3204);
    outputs(1372) <= layer2_outputs(1020);
    outputs(1373) <= layer2_outputs(2117);
    outputs(1374) <= not(layer2_outputs(1617));
    outputs(1375) <= not(layer2_outputs(4299));
    outputs(1376) <= not(layer2_outputs(4638));
    outputs(1377) <= (layer2_outputs(3714)) xor (layer2_outputs(4125));
    outputs(1378) <= not((layer2_outputs(121)) xor (layer2_outputs(3402)));
    outputs(1379) <= not(layer2_outputs(4293));
    outputs(1380) <= not(layer2_outputs(2536));
    outputs(1381) <= layer2_outputs(4254);
    outputs(1382) <= layer2_outputs(4500);
    outputs(1383) <= layer2_outputs(1557);
    outputs(1384) <= not(layer2_outputs(1675));
    outputs(1385) <= (layer2_outputs(4740)) or (layer2_outputs(3091));
    outputs(1386) <= not((layer2_outputs(1622)) and (layer2_outputs(4475)));
    outputs(1387) <= layer2_outputs(161);
    outputs(1388) <= (layer2_outputs(4409)) xor (layer2_outputs(1159));
    outputs(1389) <= layer2_outputs(3915);
    outputs(1390) <= layer2_outputs(1494);
    outputs(1391) <= not(layer2_outputs(2245));
    outputs(1392) <= not(layer2_outputs(2544));
    outputs(1393) <= not(layer2_outputs(2591)) or (layer2_outputs(4504));
    outputs(1394) <= not(layer2_outputs(4990)) or (layer2_outputs(4381));
    outputs(1395) <= not(layer2_outputs(1633));
    outputs(1396) <= (layer2_outputs(3258)) and (layer2_outputs(3396));
    outputs(1397) <= layer2_outputs(4931);
    outputs(1398) <= layer2_outputs(3999);
    outputs(1399) <= not((layer2_outputs(4837)) xor (layer2_outputs(4260)));
    outputs(1400) <= layer2_outputs(1818);
    outputs(1401) <= not(layer2_outputs(4438));
    outputs(1402) <= layer2_outputs(1367);
    outputs(1403) <= (layer2_outputs(636)) xor (layer2_outputs(166));
    outputs(1404) <= (layer2_outputs(4789)) xor (layer2_outputs(886));
    outputs(1405) <= layer2_outputs(2571);
    outputs(1406) <= not(layer2_outputs(1521));
    outputs(1407) <= not((layer2_outputs(2528)) xor (layer2_outputs(893)));
    outputs(1408) <= not(layer2_outputs(3103));
    outputs(1409) <= not(layer2_outputs(1009));
    outputs(1410) <= not(layer2_outputs(894));
    outputs(1411) <= not(layer2_outputs(2087));
    outputs(1412) <= layer2_outputs(2168);
    outputs(1413) <= layer2_outputs(4526);
    outputs(1414) <= layer2_outputs(63);
    outputs(1415) <= not(layer2_outputs(1948));
    outputs(1416) <= not(layer2_outputs(1287)) or (layer2_outputs(3720));
    outputs(1417) <= not(layer2_outputs(1027));
    outputs(1418) <= not(layer2_outputs(3906));
    outputs(1419) <= not(layer2_outputs(4394));
    outputs(1420) <= (layer2_outputs(3048)) xor (layer2_outputs(3643));
    outputs(1421) <= layer2_outputs(3399);
    outputs(1422) <= not(layer2_outputs(1470));
    outputs(1423) <= not(layer2_outputs(4674));
    outputs(1424) <= layer2_outputs(891);
    outputs(1425) <= layer2_outputs(601);
    outputs(1426) <= not(layer2_outputs(4120));
    outputs(1427) <= (layer2_outputs(3140)) and not (layer2_outputs(5099));
    outputs(1428) <= (layer2_outputs(799)) xor (layer2_outputs(546));
    outputs(1429) <= not((layer2_outputs(1484)) xor (layer2_outputs(4156)));
    outputs(1430) <= layer2_outputs(4594);
    outputs(1431) <= (layer2_outputs(459)) and not (layer2_outputs(2172));
    outputs(1432) <= not(layer2_outputs(2049));
    outputs(1433) <= layer2_outputs(959);
    outputs(1434) <= not((layer2_outputs(2482)) and (layer2_outputs(192)));
    outputs(1435) <= (layer2_outputs(354)) xor (layer2_outputs(4519));
    outputs(1436) <= not((layer2_outputs(2840)) or (layer2_outputs(3600)));
    outputs(1437) <= layer2_outputs(3412);
    outputs(1438) <= layer2_outputs(1358);
    outputs(1439) <= (layer2_outputs(2960)) and (layer2_outputs(1635));
    outputs(1440) <= layer2_outputs(3444);
    outputs(1441) <= layer2_outputs(4649);
    outputs(1442) <= layer2_outputs(2897);
    outputs(1443) <= not(layer2_outputs(3657));
    outputs(1444) <= layer2_outputs(3230);
    outputs(1445) <= layer2_outputs(3936);
    outputs(1446) <= layer2_outputs(502);
    outputs(1447) <= not((layer2_outputs(1160)) or (layer2_outputs(4984)));
    outputs(1448) <= not(layer2_outputs(5038));
    outputs(1449) <= (layer2_outputs(3719)) xor (layer2_outputs(2009));
    outputs(1450) <= not(layer2_outputs(2913));
    outputs(1451) <= not(layer2_outputs(3015));
    outputs(1452) <= not((layer2_outputs(93)) and (layer2_outputs(1899)));
    outputs(1453) <= not(layer2_outputs(4305));
    outputs(1454) <= layer2_outputs(1003);
    outputs(1455) <= layer2_outputs(951);
    outputs(1456) <= layer2_outputs(2239);
    outputs(1457) <= not(layer2_outputs(2718));
    outputs(1458) <= not(layer2_outputs(927));
    outputs(1459) <= not((layer2_outputs(3773)) xor (layer2_outputs(4412)));
    outputs(1460) <= layer2_outputs(4173);
    outputs(1461) <= (layer2_outputs(204)) or (layer2_outputs(822));
    outputs(1462) <= not(layer2_outputs(4751));
    outputs(1463) <= not(layer2_outputs(4259));
    outputs(1464) <= not(layer2_outputs(2137));
    outputs(1465) <= layer2_outputs(4858);
    outputs(1466) <= (layer2_outputs(5064)) xor (layer2_outputs(1919));
    outputs(1467) <= layer2_outputs(2552);
    outputs(1468) <= not(layer2_outputs(492));
    outputs(1469) <= layer2_outputs(2073);
    outputs(1470) <= (layer2_outputs(1787)) and not (layer2_outputs(1012));
    outputs(1471) <= not(layer2_outputs(3897));
    outputs(1472) <= (layer2_outputs(4450)) and (layer2_outputs(1940));
    outputs(1473) <= not(layer2_outputs(3591)) or (layer2_outputs(3786));
    outputs(1474) <= layer2_outputs(4529);
    outputs(1475) <= layer2_outputs(3067);
    outputs(1476) <= not(layer2_outputs(4768));
    outputs(1477) <= (layer2_outputs(1546)) or (layer2_outputs(1793));
    outputs(1478) <= not((layer2_outputs(2390)) xor (layer2_outputs(1048)));
    outputs(1479) <= layer2_outputs(4626);
    outputs(1480) <= not(layer2_outputs(544));
    outputs(1481) <= not(layer2_outputs(879));
    outputs(1482) <= not((layer2_outputs(920)) xor (layer2_outputs(2173)));
    outputs(1483) <= (layer2_outputs(4262)) and (layer2_outputs(810));
    outputs(1484) <= (layer2_outputs(3223)) or (layer2_outputs(2970));
    outputs(1485) <= layer2_outputs(4938);
    outputs(1486) <= not(layer2_outputs(3212));
    outputs(1487) <= not(layer2_outputs(2822));
    outputs(1488) <= not(layer2_outputs(4399));
    outputs(1489) <= not(layer2_outputs(2967));
    outputs(1490) <= layer2_outputs(1916);
    outputs(1491) <= layer2_outputs(2524);
    outputs(1492) <= not(layer2_outputs(3484));
    outputs(1493) <= not(layer2_outputs(1835));
    outputs(1494) <= layer2_outputs(4660);
    outputs(1495) <= not(layer2_outputs(4476));
    outputs(1496) <= not((layer2_outputs(2536)) xor (layer2_outputs(3647)));
    outputs(1497) <= not(layer2_outputs(4438));
    outputs(1498) <= not(layer2_outputs(2915));
    outputs(1499) <= not((layer2_outputs(4293)) and (layer2_outputs(1451)));
    outputs(1500) <= not(layer2_outputs(537));
    outputs(1501) <= layer2_outputs(549);
    outputs(1502) <= not(layer2_outputs(2861));
    outputs(1503) <= not((layer2_outputs(717)) xor (layer2_outputs(557)));
    outputs(1504) <= (layer2_outputs(2841)) or (layer2_outputs(4143));
    outputs(1505) <= not(layer2_outputs(1634));
    outputs(1506) <= (layer2_outputs(320)) and not (layer2_outputs(2598));
    outputs(1507) <= not(layer2_outputs(2893));
    outputs(1508) <= not(layer2_outputs(2195));
    outputs(1509) <= (layer2_outputs(665)) or (layer2_outputs(2639));
    outputs(1510) <= not(layer2_outputs(4025));
    outputs(1511) <= (layer2_outputs(1926)) and not (layer2_outputs(3604));
    outputs(1512) <= not(layer2_outputs(1258));
    outputs(1513) <= not(layer2_outputs(2965));
    outputs(1514) <= not(layer2_outputs(3385));
    outputs(1515) <= not(layer2_outputs(3012));
    outputs(1516) <= layer2_outputs(4680);
    outputs(1517) <= not((layer2_outputs(958)) and (layer2_outputs(1480)));
    outputs(1518) <= not((layer2_outputs(762)) xor (layer2_outputs(300)));
    outputs(1519) <= (layer2_outputs(2608)) and not (layer2_outputs(3674));
    outputs(1520) <= (layer2_outputs(3851)) and (layer2_outputs(1307));
    outputs(1521) <= not(layer2_outputs(265));
    outputs(1522) <= layer2_outputs(1436);
    outputs(1523) <= (layer2_outputs(3115)) and not (layer2_outputs(2922));
    outputs(1524) <= layer2_outputs(2135);
    outputs(1525) <= layer2_outputs(772);
    outputs(1526) <= not(layer2_outputs(287));
    outputs(1527) <= not(layer2_outputs(436));
    outputs(1528) <= not(layer2_outputs(4054));
    outputs(1529) <= (layer2_outputs(1231)) xor (layer2_outputs(3285));
    outputs(1530) <= layer2_outputs(1950);
    outputs(1531) <= not(layer2_outputs(194)) or (layer2_outputs(1202));
    outputs(1532) <= not(layer2_outputs(4563));
    outputs(1533) <= not(layer2_outputs(1126)) or (layer2_outputs(3627));
    outputs(1534) <= not(layer2_outputs(130));
    outputs(1535) <= not(layer2_outputs(3268));
    outputs(1536) <= not(layer2_outputs(2919));
    outputs(1537) <= not((layer2_outputs(4884)) or (layer2_outputs(178)));
    outputs(1538) <= not(layer2_outputs(1028));
    outputs(1539) <= layer2_outputs(3441);
    outputs(1540) <= layer2_outputs(3740);
    outputs(1541) <= layer2_outputs(2203);
    outputs(1542) <= layer2_outputs(477);
    outputs(1543) <= layer2_outputs(3313);
    outputs(1544) <= not(layer2_outputs(1963));
    outputs(1545) <= not(layer2_outputs(1217));
    outputs(1546) <= layer2_outputs(3294);
    outputs(1547) <= layer2_outputs(5073);
    outputs(1548) <= (layer2_outputs(4437)) xor (layer2_outputs(865));
    outputs(1549) <= not(layer2_outputs(4268));
    outputs(1550) <= not((layer2_outputs(675)) xor (layer2_outputs(4712)));
    outputs(1551) <= not(layer2_outputs(4257));
    outputs(1552) <= not(layer2_outputs(3045));
    outputs(1553) <= (layer2_outputs(4360)) and (layer2_outputs(2680));
    outputs(1554) <= not(layer2_outputs(1146));
    outputs(1555) <= layer2_outputs(2140);
    outputs(1556) <= layer2_outputs(3265);
    outputs(1557) <= layer2_outputs(2195);
    outputs(1558) <= not(layer2_outputs(4629));
    outputs(1559) <= layer2_outputs(2318);
    outputs(1560) <= layer2_outputs(1831);
    outputs(1561) <= layer2_outputs(3625);
    outputs(1562) <= layer2_outputs(1285);
    outputs(1563) <= not(layer2_outputs(5077));
    outputs(1564) <= not(layer2_outputs(4104)) or (layer2_outputs(4819));
    outputs(1565) <= (layer2_outputs(3018)) xor (layer2_outputs(4007));
    outputs(1566) <= layer2_outputs(2479);
    outputs(1567) <= layer2_outputs(4165);
    outputs(1568) <= not((layer2_outputs(4773)) or (layer2_outputs(1462)));
    outputs(1569) <= (layer2_outputs(1460)) and not (layer2_outputs(4659));
    outputs(1570) <= (layer2_outputs(627)) and (layer2_outputs(457));
    outputs(1571) <= layer2_outputs(1314);
    outputs(1572) <= (layer2_outputs(2354)) and not (layer2_outputs(1930));
    outputs(1573) <= not(layer2_outputs(4731));
    outputs(1574) <= layer2_outputs(42);
    outputs(1575) <= layer2_outputs(856);
    outputs(1576) <= (layer2_outputs(1842)) and not (layer2_outputs(2708));
    outputs(1577) <= not(layer2_outputs(200));
    outputs(1578) <= not(layer2_outputs(2376));
    outputs(1579) <= not(layer2_outputs(1104));
    outputs(1580) <= (layer2_outputs(2518)) and not (layer2_outputs(4536));
    outputs(1581) <= (layer2_outputs(3002)) and (layer2_outputs(617));
    outputs(1582) <= not(layer2_outputs(4559));
    outputs(1583) <= layer2_outputs(2457);
    outputs(1584) <= (layer2_outputs(4294)) and (layer2_outputs(3972));
    outputs(1585) <= not((layer2_outputs(1291)) or (layer2_outputs(4640)));
    outputs(1586) <= (layer2_outputs(3764)) and not (layer2_outputs(4815));
    outputs(1587) <= layer2_outputs(2618);
    outputs(1588) <= not((layer2_outputs(2847)) xor (layer2_outputs(824)));
    outputs(1589) <= (layer2_outputs(4568)) and not (layer2_outputs(1956));
    outputs(1590) <= not(layer2_outputs(3231));
    outputs(1591) <= layer2_outputs(3439);
    outputs(1592) <= layer2_outputs(4777);
    outputs(1593) <= not(layer2_outputs(3918));
    outputs(1594) <= not((layer2_outputs(4074)) or (layer2_outputs(3218)));
    outputs(1595) <= (layer2_outputs(2062)) and (layer2_outputs(4429));
    outputs(1596) <= layer2_outputs(2747);
    outputs(1597) <= not(layer2_outputs(2576));
    outputs(1598) <= not(layer2_outputs(4809)) or (layer2_outputs(4758));
    outputs(1599) <= not(layer2_outputs(3167));
    outputs(1600) <= not(layer2_outputs(1466)) or (layer2_outputs(4045));
    outputs(1601) <= not(layer2_outputs(3224));
    outputs(1602) <= not((layer2_outputs(2653)) or (layer2_outputs(1559)));
    outputs(1603) <= layer2_outputs(373);
    outputs(1604) <= not(layer2_outputs(35));
    outputs(1605) <= not((layer2_outputs(4918)) xor (layer2_outputs(889)));
    outputs(1606) <= layer2_outputs(1738);
    outputs(1607) <= layer2_outputs(678);
    outputs(1608) <= not(layer2_outputs(3855));
    outputs(1609) <= layer2_outputs(1433);
    outputs(1610) <= not((layer2_outputs(1152)) or (layer2_outputs(3087)));
    outputs(1611) <= (layer2_outputs(2743)) and not (layer2_outputs(1274));
    outputs(1612) <= not((layer2_outputs(1656)) or (layer2_outputs(2237)));
    outputs(1613) <= not((layer2_outputs(4855)) xor (layer2_outputs(4300)));
    outputs(1614) <= layer2_outputs(2116);
    outputs(1615) <= (layer2_outputs(1314)) and not (layer2_outputs(176));
    outputs(1616) <= (layer2_outputs(1807)) and not (layer2_outputs(1548));
    outputs(1617) <= not(layer2_outputs(107));
    outputs(1618) <= not(layer2_outputs(284));
    outputs(1619) <= not(layer2_outputs(5049));
    outputs(1620) <= layer2_outputs(2618);
    outputs(1621) <= layer2_outputs(2872);
    outputs(1622) <= (layer2_outputs(377)) and (layer2_outputs(2744));
    outputs(1623) <= not((layer2_outputs(2560)) or (layer2_outputs(1028)));
    outputs(1624) <= not(layer2_outputs(996));
    outputs(1625) <= layer2_outputs(4963);
    outputs(1626) <= not(layer2_outputs(1726));
    outputs(1627) <= (layer2_outputs(5003)) and not (layer2_outputs(881));
    outputs(1628) <= layer2_outputs(2630);
    outputs(1629) <= not(layer2_outputs(45));
    outputs(1630) <= layer2_outputs(2738);
    outputs(1631) <= (layer2_outputs(854)) and (layer2_outputs(1517));
    outputs(1632) <= not(layer2_outputs(1399));
    outputs(1633) <= layer2_outputs(1803);
    outputs(1634) <= not(layer2_outputs(3030));
    outputs(1635) <= not(layer2_outputs(210));
    outputs(1636) <= layer2_outputs(198);
    outputs(1637) <= (layer2_outputs(4749)) and (layer2_outputs(3822));
    outputs(1638) <= (layer2_outputs(1116)) and not (layer2_outputs(1199));
    outputs(1639) <= layer2_outputs(1690);
    outputs(1640) <= (layer2_outputs(3384)) and not (layer2_outputs(1376));
    outputs(1641) <= (layer2_outputs(3247)) xor (layer2_outputs(2487));
    outputs(1642) <= layer2_outputs(3818);
    outputs(1643) <= layer2_outputs(311);
    outputs(1644) <= not((layer2_outputs(568)) or (layer2_outputs(4694)));
    outputs(1645) <= not(layer2_outputs(800));
    outputs(1646) <= (layer2_outputs(4952)) xor (layer2_outputs(3730));
    outputs(1647) <= not((layer2_outputs(361)) or (layer2_outputs(1710)));
    outputs(1648) <= not(layer2_outputs(2656));
    outputs(1649) <= layer2_outputs(76);
    outputs(1650) <= not((layer2_outputs(3410)) xor (layer2_outputs(4716)));
    outputs(1651) <= not(layer2_outputs(2701));
    outputs(1652) <= (layer2_outputs(4873)) and (layer2_outputs(1065));
    outputs(1653) <= layer2_outputs(2961);
    outputs(1654) <= (layer2_outputs(1498)) and not (layer2_outputs(3691));
    outputs(1655) <= layer2_outputs(2558);
    outputs(1656) <= layer2_outputs(2763);
    outputs(1657) <= not((layer2_outputs(1041)) or (layer2_outputs(480)));
    outputs(1658) <= (layer2_outputs(5080)) and not (layer2_outputs(1968));
    outputs(1659) <= layer2_outputs(4012);
    outputs(1660) <= (layer2_outputs(1895)) and not (layer2_outputs(1732));
    outputs(1661) <= not(layer2_outputs(1541));
    outputs(1662) <= (layer2_outputs(1977)) and (layer2_outputs(1933));
    outputs(1663) <= not((layer2_outputs(1071)) xor (layer2_outputs(2712)));
    outputs(1664) <= layer2_outputs(4801);
    outputs(1665) <= not((layer2_outputs(1440)) xor (layer2_outputs(3064)));
    outputs(1666) <= layer2_outputs(3717);
    outputs(1667) <= not(layer2_outputs(3898));
    outputs(1668) <= layer2_outputs(1681);
    outputs(1669) <= (layer2_outputs(3517)) xor (layer2_outputs(4222));
    outputs(1670) <= layer2_outputs(223);
    outputs(1671) <= not(layer2_outputs(4892));
    outputs(1672) <= not(layer2_outputs(3027));
    outputs(1673) <= (layer2_outputs(1133)) and not (layer2_outputs(250));
    outputs(1674) <= (layer2_outputs(1659)) and not (layer2_outputs(2785));
    outputs(1675) <= (layer2_outputs(1751)) and (layer2_outputs(4587));
    outputs(1676) <= layer2_outputs(4322);
    outputs(1677) <= not((layer2_outputs(2390)) xor (layer2_outputs(2124)));
    outputs(1678) <= not(layer2_outputs(4210));
    outputs(1679) <= (layer2_outputs(4176)) and (layer2_outputs(1212));
    outputs(1680) <= not((layer2_outputs(5051)) or (layer2_outputs(1352)));
    outputs(1681) <= not(layer2_outputs(1249));
    outputs(1682) <= not(layer2_outputs(2575));
    outputs(1683) <= not(layer2_outputs(2924));
    outputs(1684) <= layer2_outputs(3903);
    outputs(1685) <= layer2_outputs(2610);
    outputs(1686) <= not(layer2_outputs(3053));
    outputs(1687) <= not(layer2_outputs(4312));
    outputs(1688) <= layer2_outputs(3735);
    outputs(1689) <= (layer2_outputs(432)) and not (layer2_outputs(4161));
    outputs(1690) <= (layer2_outputs(1951)) and not (layer2_outputs(3600));
    outputs(1691) <= layer2_outputs(3683);
    outputs(1692) <= (layer2_outputs(2667)) and not (layer2_outputs(2209));
    outputs(1693) <= not(layer2_outputs(483));
    outputs(1694) <= layer2_outputs(4641);
    outputs(1695) <= not((layer2_outputs(1784)) xor (layer2_outputs(5087)));
    outputs(1696) <= layer2_outputs(3005);
    outputs(1697) <= not(layer2_outputs(530));
    outputs(1698) <= not(layer2_outputs(1318));
    outputs(1699) <= (layer2_outputs(1327)) or (layer2_outputs(1311));
    outputs(1700) <= layer2_outputs(2776);
    outputs(1701) <= layer2_outputs(2903);
    outputs(1702) <= layer2_outputs(3545);
    outputs(1703) <= not((layer2_outputs(2156)) or (layer2_outputs(2086)));
    outputs(1704) <= (layer2_outputs(4496)) and (layer2_outputs(3014));
    outputs(1705) <= not((layer2_outputs(1213)) xor (layer2_outputs(4915)));
    outputs(1706) <= not(layer2_outputs(355));
    outputs(1707) <= (layer2_outputs(0)) xor (layer2_outputs(2930));
    outputs(1708) <= not((layer2_outputs(2238)) or (layer2_outputs(3481)));
    outputs(1709) <= not((layer2_outputs(4913)) or (layer2_outputs(2112)));
    outputs(1710) <= (layer2_outputs(1231)) and not (layer2_outputs(2394));
    outputs(1711) <= layer2_outputs(2916);
    outputs(1712) <= layer2_outputs(1792);
    outputs(1713) <= (layer2_outputs(3503)) and not (layer2_outputs(3714));
    outputs(1714) <= layer2_outputs(4343);
    outputs(1715) <= layer2_outputs(315);
    outputs(1716) <= not(layer2_outputs(4439));
    outputs(1717) <= not(layer2_outputs(2977));
    outputs(1718) <= (layer2_outputs(1197)) and (layer2_outputs(4733));
    outputs(1719) <= not(layer2_outputs(2243));
    outputs(1720) <= (layer2_outputs(4777)) or (layer2_outputs(2045));
    outputs(1721) <= not(layer2_outputs(2721));
    outputs(1722) <= not((layer2_outputs(2397)) xor (layer2_outputs(2650)));
    outputs(1723) <= not(layer2_outputs(3396));
    outputs(1724) <= not((layer2_outputs(3883)) or (layer2_outputs(2102)));
    outputs(1725) <= not(layer2_outputs(4107));
    outputs(1726) <= layer2_outputs(315);
    outputs(1727) <= (layer2_outputs(4480)) xor (layer2_outputs(1477));
    outputs(1728) <= not(layer2_outputs(4639)) or (layer2_outputs(4080));
    outputs(1729) <= not(layer2_outputs(385)) or (layer2_outputs(4480));
    outputs(1730) <= layer2_outputs(2080);
    outputs(1731) <= not(layer2_outputs(45));
    outputs(1732) <= not(layer2_outputs(695));
    outputs(1733) <= (layer2_outputs(2067)) xor (layer2_outputs(383));
    outputs(1734) <= layer2_outputs(941);
    outputs(1735) <= not(layer2_outputs(2797));
    outputs(1736) <= layer2_outputs(4266);
    outputs(1737) <= not(layer2_outputs(2881));
    outputs(1738) <= not(layer2_outputs(1230)) or (layer2_outputs(654));
    outputs(1739) <= layer2_outputs(2668);
    outputs(1740) <= layer2_outputs(353);
    outputs(1741) <= not(layer2_outputs(773));
    outputs(1742) <= not(layer2_outputs(2466));
    outputs(1743) <= (layer2_outputs(3479)) and not (layer2_outputs(3490));
    outputs(1744) <= layer2_outputs(3755);
    outputs(1745) <= layer2_outputs(745);
    outputs(1746) <= not(layer2_outputs(288));
    outputs(1747) <= not(layer2_outputs(4541));
    outputs(1748) <= (layer2_outputs(4492)) and not (layer2_outputs(2583));
    outputs(1749) <= layer2_outputs(229);
    outputs(1750) <= (layer2_outputs(149)) xor (layer2_outputs(2372));
    outputs(1751) <= layer2_outputs(1955);
    outputs(1752) <= not(layer2_outputs(489));
    outputs(1753) <= (layer2_outputs(5118)) and not (layer2_outputs(3588));
    outputs(1754) <= layer2_outputs(3763);
    outputs(1755) <= layer2_outputs(3542);
    outputs(1756) <= not(layer2_outputs(3030));
    outputs(1757) <= layer2_outputs(4400);
    outputs(1758) <= (layer2_outputs(1690)) and not (layer2_outputs(462));
    outputs(1759) <= not(layer2_outputs(2532));
    outputs(1760) <= layer2_outputs(1171);
    outputs(1761) <= not(layer2_outputs(4639));
    outputs(1762) <= layer2_outputs(371);
    outputs(1763) <= (layer2_outputs(2438)) and (layer2_outputs(1058));
    outputs(1764) <= layer2_outputs(17);
    outputs(1765) <= (layer2_outputs(798)) and not (layer2_outputs(3477));
    outputs(1766) <= not(layer2_outputs(2245));
    outputs(1767) <= layer2_outputs(4367);
    outputs(1768) <= not(layer2_outputs(1132));
    outputs(1769) <= (layer2_outputs(4026)) xor (layer2_outputs(1374));
    outputs(1770) <= not(layer2_outputs(1566));
    outputs(1771) <= not(layer2_outputs(1486));
    outputs(1772) <= not(layer2_outputs(3830));
    outputs(1773) <= layer2_outputs(3783);
    outputs(1774) <= not(layer2_outputs(3110));
    outputs(1775) <= layer2_outputs(4552);
    outputs(1776) <= (layer2_outputs(3406)) and (layer2_outputs(3615));
    outputs(1777) <= not(layer2_outputs(4380));
    outputs(1778) <= not(layer2_outputs(4836)) or (layer2_outputs(5111));
    outputs(1779) <= layer2_outputs(3903);
    outputs(1780) <= (layer2_outputs(552)) and not (layer2_outputs(1458));
    outputs(1781) <= layer2_outputs(2776);
    outputs(1782) <= (layer2_outputs(860)) and not (layer2_outputs(1796));
    outputs(1783) <= not(layer2_outputs(2783));
    outputs(1784) <= layer2_outputs(1570);
    outputs(1785) <= (layer2_outputs(4190)) and not (layer2_outputs(2653));
    outputs(1786) <= layer2_outputs(5052);
    outputs(1787) <= not(layer2_outputs(3463));
    outputs(1788) <= layer2_outputs(2670);
    outputs(1789) <= not(layer2_outputs(4806));
    outputs(1790) <= not((layer2_outputs(57)) or (layer2_outputs(3151)));
    outputs(1791) <= not(layer2_outputs(230)) or (layer2_outputs(877));
    outputs(1792) <= (layer2_outputs(55)) and not (layer2_outputs(645));
    outputs(1793) <= not(layer2_outputs(4928));
    outputs(1794) <= (layer2_outputs(1960)) and not (layer2_outputs(1388));
    outputs(1795) <= not(layer2_outputs(3971)) or (layer2_outputs(70));
    outputs(1796) <= not((layer2_outputs(4588)) or (layer2_outputs(3235)));
    outputs(1797) <= not(layer2_outputs(3660));
    outputs(1798) <= (layer2_outputs(4805)) xor (layer2_outputs(3631));
    outputs(1799) <= not((layer2_outputs(1798)) xor (layer2_outputs(930)));
    outputs(1800) <= layer2_outputs(3372);
    outputs(1801) <= layer2_outputs(2147);
    outputs(1802) <= layer2_outputs(807);
    outputs(1803) <= not(layer2_outputs(1805));
    outputs(1804) <= not(layer2_outputs(2583));
    outputs(1805) <= not(layer2_outputs(4077));
    outputs(1806) <= not(layer2_outputs(1650));
    outputs(1807) <= not((layer2_outputs(347)) xor (layer2_outputs(1033)));
    outputs(1808) <= not(layer2_outputs(1996));
    outputs(1809) <= not(layer2_outputs(4875));
    outputs(1810) <= not((layer2_outputs(3693)) xor (layer2_outputs(3610)));
    outputs(1811) <= layer2_outputs(804);
    outputs(1812) <= layer2_outputs(4298);
    outputs(1813) <= not(layer2_outputs(2920));
    outputs(1814) <= (layer2_outputs(5020)) and not (layer2_outputs(1423));
    outputs(1815) <= not(layer2_outputs(706));
    outputs(1816) <= not(layer2_outputs(4853)) or (layer2_outputs(85));
    outputs(1817) <= layer2_outputs(4824);
    outputs(1818) <= not(layer2_outputs(3996));
    outputs(1819) <= not(layer2_outputs(3922));
    outputs(1820) <= (layer2_outputs(4847)) and not (layer2_outputs(1729));
    outputs(1821) <= not(layer2_outputs(1728));
    outputs(1822) <= not(layer2_outputs(62));
    outputs(1823) <= not((layer2_outputs(3426)) or (layer2_outputs(770)));
    outputs(1824) <= not(layer2_outputs(2175));
    outputs(1825) <= layer2_outputs(1446);
    outputs(1826) <= not(layer2_outputs(4772));
    outputs(1827) <= not((layer2_outputs(790)) or (layer2_outputs(2425)));
    outputs(1828) <= not((layer2_outputs(3086)) xor (layer2_outputs(4887)));
    outputs(1829) <= not((layer2_outputs(66)) and (layer2_outputs(983)));
    outputs(1830) <= not(layer2_outputs(1268));
    outputs(1831) <= (layer2_outputs(1295)) xor (layer2_outputs(4732));
    outputs(1832) <= (layer2_outputs(2989)) and (layer2_outputs(4001));
    outputs(1833) <= layer2_outputs(4819);
    outputs(1834) <= not((layer2_outputs(2683)) and (layer2_outputs(1216)));
    outputs(1835) <= (layer2_outputs(438)) xor (layer2_outputs(1742));
    outputs(1836) <= layer2_outputs(2554);
    outputs(1837) <= layer2_outputs(1405);
    outputs(1838) <= not(layer2_outputs(4679));
    outputs(1839) <= not(layer2_outputs(3652)) or (layer2_outputs(3346));
    outputs(1840) <= (layer2_outputs(2793)) xor (layer2_outputs(2672));
    outputs(1841) <= not(layer2_outputs(708)) or (layer2_outputs(1639));
    outputs(1842) <= (layer2_outputs(725)) and not (layer2_outputs(2555));
    outputs(1843) <= layer2_outputs(1389);
    outputs(1844) <= not(layer2_outputs(3185));
    outputs(1845) <= not(layer2_outputs(4341));
    outputs(1846) <= (layer2_outputs(5040)) and (layer2_outputs(4281));
    outputs(1847) <= not((layer2_outputs(2441)) xor (layer2_outputs(437)));
    outputs(1848) <= not(layer2_outputs(2832));
    outputs(1849) <= not((layer2_outputs(517)) xor (layer2_outputs(651)));
    outputs(1850) <= layer2_outputs(3759);
    outputs(1851) <= not(layer2_outputs(2383));
    outputs(1852) <= (layer2_outputs(1183)) and (layer2_outputs(1901));
    outputs(1853) <= not(layer2_outputs(4164));
    outputs(1854) <= layer2_outputs(4543);
    outputs(1855) <= not((layer2_outputs(2346)) xor (layer2_outputs(237)));
    outputs(1856) <= not(layer2_outputs(426));
    outputs(1857) <= (layer2_outputs(4288)) and (layer2_outputs(925));
    outputs(1858) <= not(layer2_outputs(301));
    outputs(1859) <= layer2_outputs(4366);
    outputs(1860) <= not(layer2_outputs(2689));
    outputs(1861) <= not(layer2_outputs(3010)) or (layer2_outputs(1666));
    outputs(1862) <= layer2_outputs(4766);
    outputs(1863) <= (layer2_outputs(3705)) and (layer2_outputs(4441));
    outputs(1864) <= (layer2_outputs(4443)) and (layer2_outputs(1062));
    outputs(1865) <= not(layer2_outputs(3898));
    outputs(1866) <= (layer2_outputs(4119)) and not (layer2_outputs(1412));
    outputs(1867) <= layer2_outputs(4138);
    outputs(1868) <= layer2_outputs(2680);
    outputs(1869) <= not(layer2_outputs(113));
    outputs(1870) <= layer2_outputs(2011);
    outputs(1871) <= (layer2_outputs(3727)) and (layer2_outputs(1338));
    outputs(1872) <= not(layer2_outputs(4528));
    outputs(1873) <= not(layer2_outputs(2860));
    outputs(1874) <= layer2_outputs(4377);
    outputs(1875) <= (layer2_outputs(2710)) and (layer2_outputs(1700));
    outputs(1876) <= not(layer2_outputs(3497));
    outputs(1877) <= (layer2_outputs(3013)) and (layer2_outputs(2072));
    outputs(1878) <= not(layer2_outputs(1559));
    outputs(1879) <= (layer2_outputs(3886)) xor (layer2_outputs(262));
    outputs(1880) <= (layer2_outputs(3843)) and not (layer2_outputs(3418));
    outputs(1881) <= not(layer2_outputs(646));
    outputs(1882) <= not(layer2_outputs(4417));
    outputs(1883) <= not(layer2_outputs(303));
    outputs(1884) <= (layer2_outputs(3051)) xor (layer2_outputs(4735));
    outputs(1885) <= not(layer2_outputs(4419));
    outputs(1886) <= (layer2_outputs(705)) and not (layer2_outputs(3533));
    outputs(1887) <= not(layer2_outputs(1747));
    outputs(1888) <= not(layer2_outputs(3601));
    outputs(1889) <= (layer2_outputs(2835)) and not (layer2_outputs(2899));
    outputs(1890) <= not(layer2_outputs(4424));
    outputs(1891) <= not((layer2_outputs(3296)) xor (layer2_outputs(1502)));
    outputs(1892) <= layer2_outputs(4570);
    outputs(1893) <= not((layer2_outputs(994)) or (layer2_outputs(1496)));
    outputs(1894) <= not((layer2_outputs(3004)) or (layer2_outputs(2762)));
    outputs(1895) <= layer2_outputs(4584);
    outputs(1896) <= layer2_outputs(2080);
    outputs(1897) <= not((layer2_outputs(4363)) or (layer2_outputs(2792)));
    outputs(1898) <= layer2_outputs(955);
    outputs(1899) <= layer2_outputs(4050);
    outputs(1900) <= not((layer2_outputs(4141)) or (layer2_outputs(1931)));
    outputs(1901) <= (layer2_outputs(5061)) and (layer2_outputs(3976));
    outputs(1902) <= not(layer2_outputs(4547)) or (layer2_outputs(2712));
    outputs(1903) <= not(layer2_outputs(4521));
    outputs(1904) <= (layer2_outputs(3711)) and not (layer2_outputs(2445));
    outputs(1905) <= (layer2_outputs(3779)) and not (layer2_outputs(2321));
    outputs(1906) <= (layer2_outputs(1130)) and (layer2_outputs(609));
    outputs(1907) <= layer2_outputs(4831);
    outputs(1908) <= layer2_outputs(28);
    outputs(1909) <= layer2_outputs(1389);
    outputs(1910) <= not(layer2_outputs(4524));
    outputs(1911) <= not(layer2_outputs(3123));
    outputs(1912) <= not((layer2_outputs(4091)) or (layer2_outputs(396)));
    outputs(1913) <= not(layer2_outputs(2907));
    outputs(1914) <= layer2_outputs(522);
    outputs(1915) <= layer2_outputs(3310);
    outputs(1916) <= not(layer2_outputs(1734));
    outputs(1917) <= layer2_outputs(2737);
    outputs(1918) <= (layer2_outputs(88)) and not (layer2_outputs(4808));
    outputs(1919) <= '0';
    outputs(1920) <= (layer2_outputs(3790)) and not (layer2_outputs(276));
    outputs(1921) <= not(layer2_outputs(2570));
    outputs(1922) <= layer2_outputs(293);
    outputs(1923) <= (layer2_outputs(2882)) and not (layer2_outputs(1441));
    outputs(1924) <= (layer2_outputs(1648)) and (layer2_outputs(3187));
    outputs(1925) <= not(layer2_outputs(1331)) or (layer2_outputs(4804));
    outputs(1926) <= not(layer2_outputs(4772));
    outputs(1927) <= layer2_outputs(496);
    outputs(1928) <= (layer2_outputs(2247)) and not (layer2_outputs(2468));
    outputs(1929) <= not(layer2_outputs(4161));
    outputs(1930) <= not(layer2_outputs(1141));
    outputs(1931) <= layer2_outputs(4306);
    outputs(1932) <= (layer2_outputs(3236)) and not (layer2_outputs(261));
    outputs(1933) <= layer2_outputs(1727);
    outputs(1934) <= layer2_outputs(217);
    outputs(1935) <= not(layer2_outputs(4122)) or (layer2_outputs(2692));
    outputs(1936) <= not(layer2_outputs(1746));
    outputs(1937) <= (layer2_outputs(5027)) and not (layer2_outputs(255));
    outputs(1938) <= layer2_outputs(4723);
    outputs(1939) <= (layer2_outputs(4015)) and not (layer2_outputs(201));
    outputs(1940) <= (layer2_outputs(838)) and (layer2_outputs(3406));
    outputs(1941) <= not((layer2_outputs(2820)) or (layer2_outputs(2054)));
    outputs(1942) <= not(layer2_outputs(1947));
    outputs(1943) <= not(layer2_outputs(1275));
    outputs(1944) <= layer2_outputs(3375);
    outputs(1945) <= layer2_outputs(1953);
    outputs(1946) <= not(layer2_outputs(2456));
    outputs(1947) <= not((layer2_outputs(56)) and (layer2_outputs(2285)));
    outputs(1948) <= not(layer2_outputs(3839));
    outputs(1949) <= not(layer2_outputs(3845));
    outputs(1950) <= not(layer2_outputs(4479));
    outputs(1951) <= not((layer2_outputs(2987)) or (layer2_outputs(32)));
    outputs(1952) <= layer2_outputs(2549);
    outputs(1953) <= not(layer2_outputs(2395));
    outputs(1954) <= not(layer2_outputs(2180));
    outputs(1955) <= (layer2_outputs(3118)) xor (layer2_outputs(2820));
    outputs(1956) <= (layer2_outputs(2189)) and not (layer2_outputs(3743));
    outputs(1957) <= not(layer2_outputs(871));
    outputs(1958) <= layer2_outputs(4870);
    outputs(1959) <= layer2_outputs(2765);
    outputs(1960) <= (layer2_outputs(3238)) and (layer2_outputs(1220));
    outputs(1961) <= not((layer2_outputs(1385)) xor (layer2_outputs(3530)));
    outputs(1962) <= layer2_outputs(3200);
    outputs(1963) <= layer2_outputs(1536);
    outputs(1964) <= not(layer2_outputs(3815));
    outputs(1965) <= not(layer2_outputs(4467));
    outputs(1966) <= (layer2_outputs(1644)) and (layer2_outputs(718));
    outputs(1967) <= layer2_outputs(4022);
    outputs(1968) <= not((layer2_outputs(3000)) and (layer2_outputs(4242)));
    outputs(1969) <= layer2_outputs(4593);
    outputs(1970) <= not((layer2_outputs(3645)) or (layer2_outputs(3546)));
    outputs(1971) <= not(layer2_outputs(2520));
    outputs(1972) <= (layer2_outputs(4306)) and (layer2_outputs(3107));
    outputs(1973) <= not(layer2_outputs(2648));
    outputs(1974) <= (layer2_outputs(3890)) xor (layer2_outputs(1784));
    outputs(1975) <= not(layer2_outputs(1121));
    outputs(1976) <= (layer2_outputs(2517)) and not (layer2_outputs(1350));
    outputs(1977) <= not((layer2_outputs(3863)) and (layer2_outputs(4290)));
    outputs(1978) <= (layer2_outputs(1904)) xor (layer2_outputs(4238));
    outputs(1979) <= layer2_outputs(1431);
    outputs(1980) <= not((layer2_outputs(2281)) or (layer2_outputs(3087)));
    outputs(1981) <= not(layer2_outputs(1620)) or (layer2_outputs(445));
    outputs(1982) <= (layer2_outputs(2533)) and (layer2_outputs(1284));
    outputs(1983) <= layer2_outputs(2408);
    outputs(1984) <= not(layer2_outputs(3739));
    outputs(1985) <= layer2_outputs(3951);
    outputs(1986) <= layer2_outputs(3826);
    outputs(1987) <= (layer2_outputs(2272)) xor (layer2_outputs(3207));
    outputs(1988) <= layer2_outputs(4219);
    outputs(1989) <= layer2_outputs(746);
    outputs(1990) <= not(layer2_outputs(2798));
    outputs(1991) <= not(layer2_outputs(1862));
    outputs(1992) <= layer2_outputs(3997);
    outputs(1993) <= layer2_outputs(2253);
    outputs(1994) <= (layer2_outputs(232)) xor (layer2_outputs(3710));
    outputs(1995) <= layer2_outputs(2133);
    outputs(1996) <= layer2_outputs(533);
    outputs(1997) <= not((layer2_outputs(2281)) or (layer2_outputs(1740)));
    outputs(1998) <= not(layer2_outputs(2858));
    outputs(1999) <= not(layer2_outputs(4564));
    outputs(2000) <= (layer2_outputs(2036)) and (layer2_outputs(4556));
    outputs(2001) <= not((layer2_outputs(4072)) and (layer2_outputs(2300)));
    outputs(2002) <= not(layer2_outputs(3075));
    outputs(2003) <= (layer2_outputs(621)) and not (layer2_outputs(1124));
    outputs(2004) <= layer2_outputs(3936);
    outputs(2005) <= layer2_outputs(430);
    outputs(2006) <= not(layer2_outputs(3024));
    outputs(2007) <= (layer2_outputs(650)) and (layer2_outputs(868));
    outputs(2008) <= not(layer2_outputs(3728));
    outputs(2009) <= not(layer2_outputs(2319));
    outputs(2010) <= layer2_outputs(4818);
    outputs(2011) <= not((layer2_outputs(3695)) or (layer2_outputs(700)));
    outputs(2012) <= (layer2_outputs(3591)) and not (layer2_outputs(213));
    outputs(2013) <= not(layer2_outputs(3038));
    outputs(2014) <= layer2_outputs(1187);
    outputs(2015) <= not(layer2_outputs(3341));
    outputs(2016) <= not((layer2_outputs(4423)) or (layer2_outputs(4739)));
    outputs(2017) <= not(layer2_outputs(3368));
    outputs(2018) <= layer2_outputs(2509);
    outputs(2019) <= layer2_outputs(440);
    outputs(2020) <= (layer2_outputs(4874)) and not (layer2_outputs(1366));
    outputs(2021) <= not(layer2_outputs(2875));
    outputs(2022) <= not((layer2_outputs(1808)) xor (layer2_outputs(3640)));
    outputs(2023) <= not(layer2_outputs(1610));
    outputs(2024) <= (layer2_outputs(4298)) and not (layer2_outputs(1471));
    outputs(2025) <= layer2_outputs(3538);
    outputs(2026) <= not(layer2_outputs(4147));
    outputs(2027) <= not(layer2_outputs(98));
    outputs(2028) <= not(layer2_outputs(1204));
    outputs(2029) <= (layer2_outputs(1421)) and (layer2_outputs(4281));
    outputs(2030) <= (layer2_outputs(1898)) and (layer2_outputs(840));
    outputs(2031) <= not(layer2_outputs(2752));
    outputs(2032) <= not((layer2_outputs(2352)) xor (layer2_outputs(4923)));
    outputs(2033) <= not(layer2_outputs(3834));
    outputs(2034) <= not((layer2_outputs(606)) or (layer2_outputs(1845)));
    outputs(2035) <= (layer2_outputs(324)) and not (layer2_outputs(3841));
    outputs(2036) <= not(layer2_outputs(4116));
    outputs(2037) <= not(layer2_outputs(4180));
    outputs(2038) <= (layer2_outputs(234)) and (layer2_outputs(3762));
    outputs(2039) <= not((layer2_outputs(4550)) or (layer2_outputs(3438)));
    outputs(2040) <= layer2_outputs(2588);
    outputs(2041) <= (layer2_outputs(4609)) and (layer2_outputs(2933));
    outputs(2042) <= layer2_outputs(4526);
    outputs(2043) <= not((layer2_outputs(4731)) and (layer2_outputs(4107)));
    outputs(2044) <= layer2_outputs(1658);
    outputs(2045) <= not(layer2_outputs(501)) or (layer2_outputs(1292));
    outputs(2046) <= (layer2_outputs(380)) and not (layer2_outputs(2924));
    outputs(2047) <= layer2_outputs(2433);
    outputs(2048) <= not(layer2_outputs(3634));
    outputs(2049) <= (layer2_outputs(1886)) or (layer2_outputs(243));
    outputs(2050) <= layer2_outputs(3666);
    outputs(2051) <= not(layer2_outputs(1075));
    outputs(2052) <= (layer2_outputs(2051)) and (layer2_outputs(1849));
    outputs(2053) <= not(layer2_outputs(242));
    outputs(2054) <= layer2_outputs(5069);
    outputs(2055) <= layer2_outputs(2904);
    outputs(2056) <= layer2_outputs(1239);
    outputs(2057) <= not(layer2_outputs(896));
    outputs(2058) <= layer2_outputs(3884);
    outputs(2059) <= layer2_outputs(4595);
    outputs(2060) <= not((layer2_outputs(1621)) xor (layer2_outputs(802)));
    outputs(2061) <= not(layer2_outputs(5063));
    outputs(2062) <= not(layer2_outputs(4560));
    outputs(2063) <= not(layer2_outputs(4678));
    outputs(2064) <= layer2_outputs(443);
    outputs(2065) <= not(layer2_outputs(2625));
    outputs(2066) <= not(layer2_outputs(1159)) or (layer2_outputs(4018));
    outputs(2067) <= (layer2_outputs(124)) and not (layer2_outputs(1228));
    outputs(2068) <= not(layer2_outputs(3583));
    outputs(2069) <= (layer2_outputs(1253)) or (layer2_outputs(1063));
    outputs(2070) <= not(layer2_outputs(2765)) or (layer2_outputs(7));
    outputs(2071) <= layer2_outputs(2205);
    outputs(2072) <= (layer2_outputs(1481)) and (layer2_outputs(5094));
    outputs(2073) <= (layer2_outputs(3421)) and (layer2_outputs(2550));
    outputs(2074) <= not(layer2_outputs(1588));
    outputs(2075) <= not(layer2_outputs(838));
    outputs(2076) <= not((layer2_outputs(3205)) and (layer2_outputs(4444)));
    outputs(2077) <= (layer2_outputs(609)) and (layer2_outputs(4204));
    outputs(2078) <= not(layer2_outputs(2610));
    outputs(2079) <= (layer2_outputs(2331)) and not (layer2_outputs(1686));
    outputs(2080) <= not((layer2_outputs(1014)) xor (layer2_outputs(2331)));
    outputs(2081) <= (layer2_outputs(4821)) and (layer2_outputs(3525));
    outputs(2082) <= not(layer2_outputs(275));
    outputs(2083) <= not((layer2_outputs(168)) xor (layer2_outputs(4569)));
    outputs(2084) <= not(layer2_outputs(4195));
    outputs(2085) <= not((layer2_outputs(1614)) xor (layer2_outputs(3116)));
    outputs(2086) <= not((layer2_outputs(565)) xor (layer2_outputs(5083)));
    outputs(2087) <= (layer2_outputs(179)) or (layer2_outputs(3806));
    outputs(2088) <= not((layer2_outputs(83)) xor (layer2_outputs(2043)));
    outputs(2089) <= not(layer2_outputs(394));
    outputs(2090) <= layer2_outputs(389);
    outputs(2091) <= not((layer2_outputs(3590)) xor (layer2_outputs(1936)));
    outputs(2092) <= not(layer2_outputs(868));
    outputs(2093) <= (layer2_outputs(4113)) and not (layer2_outputs(114));
    outputs(2094) <= layer2_outputs(3916);
    outputs(2095) <= layer2_outputs(4720);
    outputs(2096) <= layer2_outputs(1448);
    outputs(2097) <= layer2_outputs(2077);
    outputs(2098) <= (layer2_outputs(4718)) xor (layer2_outputs(431));
    outputs(2099) <= not(layer2_outputs(2696));
    outputs(2100) <= layer2_outputs(3548);
    outputs(2101) <= not(layer2_outputs(317));
    outputs(2102) <= not(layer2_outputs(3745));
    outputs(2103) <= (layer2_outputs(1)) and (layer2_outputs(3549));
    outputs(2104) <= not((layer2_outputs(2865)) xor (layer2_outputs(2201)));
    outputs(2105) <= layer2_outputs(2881);
    outputs(2106) <= (layer2_outputs(1567)) and (layer2_outputs(1944));
    outputs(2107) <= layer2_outputs(2428);
    outputs(2108) <= not((layer2_outputs(4585)) and (layer2_outputs(1065)));
    outputs(2109) <= not(layer2_outputs(3919));
    outputs(2110) <= layer2_outputs(2896);
    outputs(2111) <= not(layer2_outputs(4912));
    outputs(2112) <= layer2_outputs(3337);
    outputs(2113) <= not(layer2_outputs(611));
    outputs(2114) <= layer2_outputs(5107);
    outputs(2115) <= not(layer2_outputs(1931));
    outputs(2116) <= not(layer2_outputs(4590));
    outputs(2117) <= not(layer2_outputs(4148));
    outputs(2118) <= not((layer2_outputs(4397)) xor (layer2_outputs(1326)));
    outputs(2119) <= (layer2_outputs(3216)) and (layer2_outputs(3277));
    outputs(2120) <= not(layer2_outputs(4532));
    outputs(2121) <= not(layer2_outputs(1294));
    outputs(2122) <= (layer2_outputs(844)) and (layer2_outputs(4488));
    outputs(2123) <= layer2_outputs(2250);
    outputs(2124) <= (layer2_outputs(2272)) and (layer2_outputs(1874));
    outputs(2125) <= not(layer2_outputs(1240));
    outputs(2126) <= not(layer2_outputs(2901)) or (layer2_outputs(4757));
    outputs(2127) <= not(layer2_outputs(1664));
    outputs(2128) <= (layer2_outputs(1520)) xor (layer2_outputs(1553));
    outputs(2129) <= not(layer2_outputs(59));
    outputs(2130) <= (layer2_outputs(482)) xor (layer2_outputs(3347));
    outputs(2131) <= (layer2_outputs(2818)) and not (layer2_outputs(1889));
    outputs(2132) <= not(layer2_outputs(1654));
    outputs(2133) <= (layer2_outputs(1029)) and not (layer2_outputs(3332));
    outputs(2134) <= not((layer2_outputs(4437)) xor (layer2_outputs(3017)));
    outputs(2135) <= not(layer2_outputs(1152));
    outputs(2136) <= (layer2_outputs(2268)) and not (layer2_outputs(2815));
    outputs(2137) <= not(layer2_outputs(2155));
    outputs(2138) <= layer2_outputs(3521);
    outputs(2139) <= not(layer2_outputs(1179));
    outputs(2140) <= not(layer2_outputs(135)) or (layer2_outputs(3102));
    outputs(2141) <= (layer2_outputs(1178)) xor (layer2_outputs(407));
    outputs(2142) <= layer2_outputs(4512);
    outputs(2143) <= layer2_outputs(3221);
    outputs(2144) <= not(layer2_outputs(1084)) or (layer2_outputs(3543));
    outputs(2145) <= not((layer2_outputs(3325)) or (layer2_outputs(3578)));
    outputs(2146) <= layer2_outputs(1379);
    outputs(2147) <= not((layer2_outputs(207)) or (layer2_outputs(5005)));
    outputs(2148) <= layer2_outputs(4524);
    outputs(2149) <= layer2_outputs(586);
    outputs(2150) <= not(layer2_outputs(4665)) or (layer2_outputs(1191));
    outputs(2151) <= (layer2_outputs(4825)) xor (layer2_outputs(3222));
    outputs(2152) <= (layer2_outputs(3287)) and (layer2_outputs(4114));
    outputs(2153) <= layer2_outputs(2263);
    outputs(2154) <= (layer2_outputs(2682)) and (layer2_outputs(4743));
    outputs(2155) <= layer2_outputs(110);
    outputs(2156) <= not(layer2_outputs(572));
    outputs(2157) <= not(layer2_outputs(1778));
    outputs(2158) <= not((layer2_outputs(49)) xor (layer2_outputs(2640)));
    outputs(2159) <= not(layer2_outputs(155));
    outputs(2160) <= not((layer2_outputs(4643)) or (layer2_outputs(2410)));
    outputs(2161) <= layer2_outputs(1771);
    outputs(2162) <= layer2_outputs(1522);
    outputs(2163) <= (layer2_outputs(2828)) and not (layer2_outputs(3301));
    outputs(2164) <= not((layer2_outputs(1503)) or (layer2_outputs(2577)));
    outputs(2165) <= not(layer2_outputs(4945));
    outputs(2166) <= not(layer2_outputs(2902));
    outputs(2167) <= layer2_outputs(2040);
    outputs(2168) <= (layer2_outputs(2999)) and not (layer2_outputs(4968));
    outputs(2169) <= layer2_outputs(104);
    outputs(2170) <= (layer2_outputs(1093)) and (layer2_outputs(4990));
    outputs(2171) <= not((layer2_outputs(1264)) xor (layer2_outputs(1691)));
    outputs(2172) <= not(layer2_outputs(713));
    outputs(2173) <= (layer2_outputs(3888)) and (layer2_outputs(2810));
    outputs(2174) <= not(layer2_outputs(3121));
    outputs(2175) <= not(layer2_outputs(3061));
    outputs(2176) <= not(layer2_outputs(322)) or (layer2_outputs(2642));
    outputs(2177) <= not(layer2_outputs(4069));
    outputs(2178) <= not(layer2_outputs(4334));
    outputs(2179) <= not((layer2_outputs(4519)) and (layer2_outputs(4193)));
    outputs(2180) <= not(layer2_outputs(43));
    outputs(2181) <= layer2_outputs(255);
    outputs(2182) <= (layer2_outputs(4919)) xor (layer2_outputs(1657));
    outputs(2183) <= layer2_outputs(4478);
    outputs(2184) <= layer2_outputs(1039);
    outputs(2185) <= not(layer2_outputs(1665));
    outputs(2186) <= layer2_outputs(1355);
    outputs(2187) <= layer2_outputs(3180);
    outputs(2188) <= layer2_outputs(1057);
    outputs(2189) <= not((layer2_outputs(934)) or (layer2_outputs(106)));
    outputs(2190) <= layer2_outputs(4994);
    outputs(2191) <= (layer2_outputs(4907)) xor (layer2_outputs(1571));
    outputs(2192) <= not(layer2_outputs(222));
    outputs(2193) <= layer2_outputs(3117);
    outputs(2194) <= not(layer2_outputs(68));
    outputs(2195) <= not(layer2_outputs(2443));
    outputs(2196) <= not(layer2_outputs(3529));
    outputs(2197) <= (layer2_outputs(2654)) and not (layer2_outputs(1142));
    outputs(2198) <= layer2_outputs(1286);
    outputs(2199) <= layer2_outputs(1612);
    outputs(2200) <= (layer2_outputs(649)) and not (layer2_outputs(2529));
    outputs(2201) <= layer2_outputs(3250);
    outputs(2202) <= not(layer2_outputs(2827));
    outputs(2203) <= not(layer2_outputs(1511));
    outputs(2204) <= not(layer2_outputs(1359));
    outputs(2205) <= not(layer2_outputs(2011));
    outputs(2206) <= not(layer2_outputs(4960)) or (layer2_outputs(2990));
    outputs(2207) <= not(layer2_outputs(1140));
    outputs(2208) <= not(layer2_outputs(1293));
    outputs(2209) <= layer2_outputs(1709);
    outputs(2210) <= not(layer2_outputs(3202));
    outputs(2211) <= layer2_outputs(4659);
    outputs(2212) <= not(layer2_outputs(2042));
    outputs(2213) <= not(layer2_outputs(5108)) or (layer2_outputs(3478));
    outputs(2214) <= (layer2_outputs(2411)) xor (layer2_outputs(4330));
    outputs(2215) <= not(layer2_outputs(3050));
    outputs(2216) <= not(layer2_outputs(2804));
    outputs(2217) <= (layer2_outputs(4215)) and not (layer2_outputs(1019));
    outputs(2218) <= layer2_outputs(252);
    outputs(2219) <= (layer2_outputs(400)) and not (layer2_outputs(226));
    outputs(2220) <= layer2_outputs(4844);
    outputs(2221) <= not((layer2_outputs(5059)) xor (layer2_outputs(2201)));
    outputs(2222) <= layer2_outputs(2131);
    outputs(2223) <= layer2_outputs(4843);
    outputs(2224) <= not(layer2_outputs(3978));
    outputs(2225) <= not(layer2_outputs(5061)) or (layer2_outputs(2432));
    outputs(2226) <= layer2_outputs(5112);
    outputs(2227) <= (layer2_outputs(3083)) and not (layer2_outputs(4428));
    outputs(2228) <= not(layer2_outputs(2247)) or (layer2_outputs(4279));
    outputs(2229) <= (layer2_outputs(991)) and not (layer2_outputs(2371));
    outputs(2230) <= layer2_outputs(578);
    outputs(2231) <= not((layer2_outputs(4792)) and (layer2_outputs(3288)));
    outputs(2232) <= layer2_outputs(3707);
    outputs(2233) <= not((layer2_outputs(1906)) xor (layer2_outputs(3606)));
    outputs(2234) <= layer2_outputs(985);
    outputs(2235) <= layer2_outputs(3257);
    outputs(2236) <= layer2_outputs(1984);
    outputs(2237) <= layer2_outputs(2350);
    outputs(2238) <= not(layer2_outputs(4352));
    outputs(2239) <= not(layer2_outputs(4004));
    outputs(2240) <= layer2_outputs(4355);
    outputs(2241) <= not(layer2_outputs(207));
    outputs(2242) <= (layer2_outputs(3157)) or (layer2_outputs(778));
    outputs(2243) <= not(layer2_outputs(2277));
    outputs(2244) <= not((layer2_outputs(4011)) xor (layer2_outputs(630)));
    outputs(2245) <= layer2_outputs(4937);
    outputs(2246) <= (layer2_outputs(1266)) and (layer2_outputs(5116));
    outputs(2247) <= layer2_outputs(3421);
    outputs(2248) <= not((layer2_outputs(3316)) xor (layer2_outputs(4042)));
    outputs(2249) <= layer2_outputs(4230);
    outputs(2250) <= not(layer2_outputs(339)) or (layer2_outputs(171));
    outputs(2251) <= not(layer2_outputs(470));
    outputs(2252) <= not(layer2_outputs(4962));
    outputs(2253) <= (layer2_outputs(4457)) and (layer2_outputs(200));
    outputs(2254) <= (layer2_outputs(2547)) and not (layer2_outputs(1106));
    outputs(2255) <= not(layer2_outputs(3877));
    outputs(2256) <= not(layer2_outputs(470));
    outputs(2257) <= layer2_outputs(1346);
    outputs(2258) <= layer2_outputs(4975);
    outputs(2259) <= layer2_outputs(1584);
    outputs(2260) <= not((layer2_outputs(3369)) xor (layer2_outputs(4518)));
    outputs(2261) <= not(layer2_outputs(1503));
    outputs(2262) <= layer2_outputs(3614);
    outputs(2263) <= layer2_outputs(2070);
    outputs(2264) <= (layer2_outputs(3794)) and (layer2_outputs(3567));
    outputs(2265) <= layer2_outputs(5016);
    outputs(2266) <= (layer2_outputs(4655)) xor (layer2_outputs(833));
    outputs(2267) <= not(layer2_outputs(1609));
    outputs(2268) <= not(layer2_outputs(4481));
    outputs(2269) <= not((layer2_outputs(4369)) and (layer2_outputs(5093)));
    outputs(2270) <= not(layer2_outputs(240));
    outputs(2271) <= not(layer2_outputs(575));
    outputs(2272) <= (layer2_outputs(1860)) and (layer2_outputs(3756));
    outputs(2273) <= layer2_outputs(1556);
    outputs(2274) <= layer2_outputs(4122);
    outputs(2275) <= not(layer2_outputs(860));
    outputs(2276) <= not((layer2_outputs(4560)) or (layer2_outputs(926)));
    outputs(2277) <= not(layer2_outputs(1894));
    outputs(2278) <= (layer2_outputs(1399)) and not (layer2_outputs(2668));
    outputs(2279) <= not(layer2_outputs(4846));
    outputs(2280) <= layer2_outputs(2208);
    outputs(2281) <= not((layer2_outputs(27)) and (layer2_outputs(2030)));
    outputs(2282) <= layer2_outputs(749);
    outputs(2283) <= layer2_outputs(1059);
    outputs(2284) <= not(layer2_outputs(4101));
    outputs(2285) <= layer2_outputs(3780);
    outputs(2286) <= layer2_outputs(2621);
    outputs(2287) <= not(layer2_outputs(4132));
    outputs(2288) <= (layer2_outputs(424)) and not (layer2_outputs(834));
    outputs(2289) <= layer2_outputs(3768);
    outputs(2290) <= not((layer2_outputs(3453)) or (layer2_outputs(3314)));
    outputs(2291) <= (layer2_outputs(4922)) xor (layer2_outputs(3562));
    outputs(2292) <= not(layer2_outputs(66));
    outputs(2293) <= not(layer2_outputs(4020));
    outputs(2294) <= (layer2_outputs(964)) and not (layer2_outputs(2387));
    outputs(2295) <= layer2_outputs(4863);
    outputs(2296) <= not(layer2_outputs(2684));
    outputs(2297) <= (layer2_outputs(3681)) xor (layer2_outputs(407));
    outputs(2298) <= layer2_outputs(2378);
    outputs(2299) <= layer2_outputs(2719);
    outputs(2300) <= layer2_outputs(3620);
    outputs(2301) <= layer2_outputs(801);
    outputs(2302) <= not(layer2_outputs(4327));
    outputs(2303) <= not(layer2_outputs(1023));
    outputs(2304) <= not(layer2_outputs(4796));
    outputs(2305) <= (layer2_outputs(1717)) and not (layer2_outputs(4125));
    outputs(2306) <= (layer2_outputs(3577)) xor (layer2_outputs(3586));
    outputs(2307) <= not(layer2_outputs(3485));
    outputs(2308) <= not(layer2_outputs(3619));
    outputs(2309) <= not(layer2_outputs(3229));
    outputs(2310) <= layer2_outputs(2092);
    outputs(2311) <= not(layer2_outputs(4551));
    outputs(2312) <= not(layer2_outputs(2511));
    outputs(2313) <= not(layer2_outputs(2069));
    outputs(2314) <= layer2_outputs(596);
    outputs(2315) <= (layer2_outputs(3314)) xor (layer2_outputs(2908));
    outputs(2316) <= (layer2_outputs(1319)) and not (layer2_outputs(53));
    outputs(2317) <= (layer2_outputs(2973)) or (layer2_outputs(1537));
    outputs(2318) <= layer2_outputs(3750);
    outputs(2319) <= (layer2_outputs(2542)) and (layer2_outputs(1222));
    outputs(2320) <= layer2_outputs(4286);
    outputs(2321) <= not(layer2_outputs(1136));
    outputs(2322) <= not(layer2_outputs(2475));
    outputs(2323) <= layer2_outputs(3506);
    outputs(2324) <= (layer2_outputs(4788)) and not (layer2_outputs(2443));
    outputs(2325) <= layer2_outputs(3098);
    outputs(2326) <= not((layer2_outputs(512)) xor (layer2_outputs(3614)));
    outputs(2327) <= layer2_outputs(4977);
    outputs(2328) <= layer2_outputs(153);
    outputs(2329) <= not(layer2_outputs(5018)) or (layer2_outputs(51));
    outputs(2330) <= not(layer2_outputs(4511));
    outputs(2331) <= not((layer2_outputs(2068)) xor (layer2_outputs(351)));
    outputs(2332) <= not(layer2_outputs(1188));
    outputs(2333) <= layer2_outputs(3993);
    outputs(2334) <= not(layer2_outputs(4727));
    outputs(2335) <= layer2_outputs(1776);
    outputs(2336) <= (layer2_outputs(3658)) and (layer2_outputs(1971));
    outputs(2337) <= (layer2_outputs(568)) and (layer2_outputs(1756));
    outputs(2338) <= not(layer2_outputs(2802));
    outputs(2339) <= not(layer2_outputs(2276));
    outputs(2340) <= not(layer2_outputs(1245)) or (layer2_outputs(1212));
    outputs(2341) <= layer2_outputs(190);
    outputs(2342) <= (layer2_outputs(3678)) and (layer2_outputs(1884));
    outputs(2343) <= layer2_outputs(3474);
    outputs(2344) <= not(layer2_outputs(826));
    outputs(2345) <= (layer2_outputs(3033)) xor (layer2_outputs(3803));
    outputs(2346) <= layer2_outputs(1170);
    outputs(2347) <= not(layer2_outputs(3339)) or (layer2_outputs(1102));
    outputs(2348) <= layer2_outputs(2522);
    outputs(2349) <= layer2_outputs(2687);
    outputs(2350) <= layer2_outputs(2268);
    outputs(2351) <= not(layer2_outputs(1423));
    outputs(2352) <= not(layer2_outputs(4882));
    outputs(2353) <= (layer2_outputs(691)) and not (layer2_outputs(5007));
    outputs(2354) <= (layer2_outputs(4608)) and not (layer2_outputs(5079));
    outputs(2355) <= layer2_outputs(816);
    outputs(2356) <= not(layer2_outputs(793));
    outputs(2357) <= layer2_outputs(1164);
    outputs(2358) <= layer2_outputs(3734);
    outputs(2359) <= (layer2_outputs(4244)) and (layer2_outputs(3741));
    outputs(2360) <= (layer2_outputs(189)) and (layer2_outputs(2060));
    outputs(2361) <= (layer2_outputs(4955)) and not (layer2_outputs(2276));
    outputs(2362) <= not((layer2_outputs(2590)) xor (layer2_outputs(1166)));
    outputs(2363) <= (layer2_outputs(1708)) xor (layer2_outputs(3227));
    outputs(2364) <= layer2_outputs(2559);
    outputs(2365) <= (layer2_outputs(2923)) xor (layer2_outputs(570));
    outputs(2366) <= not(layer2_outputs(1280));
    outputs(2367) <= layer2_outputs(708);
    outputs(2368) <= (layer2_outputs(757)) and not (layer2_outputs(608));
    outputs(2369) <= not(layer2_outputs(28));
    outputs(2370) <= not(layer2_outputs(4410));
    outputs(2371) <= not((layer2_outputs(1256)) and (layer2_outputs(2270)));
    outputs(2372) <= not((layer2_outputs(4531)) xor (layer2_outputs(2929)));
    outputs(2373) <= not(layer2_outputs(2057));
    outputs(2374) <= not(layer2_outputs(331));
    outputs(2375) <= layer2_outputs(2573);
    outputs(2376) <= not(layer2_outputs(2516));
    outputs(2377) <= layer2_outputs(3837);
    outputs(2378) <= layer2_outputs(1527);
    outputs(2379) <= layer2_outputs(1497);
    outputs(2380) <= not(layer2_outputs(4282));
    outputs(2381) <= not(layer2_outputs(4813));
    outputs(2382) <= not(layer2_outputs(1354));
    outputs(2383) <= layer2_outputs(1610);
    outputs(2384) <= layer2_outputs(3959);
    outputs(2385) <= not((layer2_outputs(326)) or (layer2_outputs(1555)));
    outputs(2386) <= (layer2_outputs(551)) xor (layer2_outputs(678));
    outputs(2387) <= layer2_outputs(2267);
    outputs(2388) <= not((layer2_outputs(3153)) xor (layer2_outputs(129)));
    outputs(2389) <= layer2_outputs(3492);
    outputs(2390) <= (layer2_outputs(2046)) xor (layer2_outputs(4187));
    outputs(2391) <= not(layer2_outputs(3532));
    outputs(2392) <= layer2_outputs(3169);
    outputs(2393) <= not(layer2_outputs(684));
    outputs(2394) <= not(layer2_outputs(1524));
    outputs(2395) <= not((layer2_outputs(4160)) xor (layer2_outputs(1086)));
    outputs(2396) <= not(layer2_outputs(1494));
    outputs(2397) <= layer2_outputs(418);
    outputs(2398) <= not(layer2_outputs(4123));
    outputs(2399) <= not(layer2_outputs(713));
    outputs(2400) <= not((layer2_outputs(1416)) or (layer2_outputs(4335)));
    outputs(2401) <= (layer2_outputs(2258)) xor (layer2_outputs(876));
    outputs(2402) <= not(layer2_outputs(4725));
    outputs(2403) <= layer2_outputs(3942);
    outputs(2404) <= layer2_outputs(2022);
    outputs(2405) <= layer2_outputs(5089);
    outputs(2406) <= (layer2_outputs(3342)) xor (layer2_outputs(4251));
    outputs(2407) <= (layer2_outputs(1989)) and not (layer2_outputs(2470));
    outputs(2408) <= layer2_outputs(596);
    outputs(2409) <= (layer2_outputs(4840)) and not (layer2_outputs(1868));
    outputs(2410) <= not(layer2_outputs(1543));
    outputs(2411) <= layer2_outputs(1483);
    outputs(2412) <= not(layer2_outputs(4334));
    outputs(2413) <= not(layer2_outputs(1834));
    outputs(2414) <= layer2_outputs(3732);
    outputs(2415) <= (layer2_outputs(3768)) and (layer2_outputs(2880));
    outputs(2416) <= layer2_outputs(1443);
    outputs(2417) <= not((layer2_outputs(5066)) and (layer2_outputs(3531)));
    outputs(2418) <= not((layer2_outputs(808)) or (layer2_outputs(4708)));
    outputs(2419) <= (layer2_outputs(4297)) and not (layer2_outputs(2759));
    outputs(2420) <= not(layer2_outputs(3453));
    outputs(2421) <= (layer2_outputs(3104)) and (layer2_outputs(3902));
    outputs(2422) <= layer2_outputs(2179);
    outputs(2423) <= not((layer2_outputs(1516)) or (layer2_outputs(3053)));
    outputs(2424) <= (layer2_outputs(1409)) and not (layer2_outputs(4084));
    outputs(2425) <= not((layer2_outputs(2246)) xor (layer2_outputs(5015)));
    outputs(2426) <= not(layer2_outputs(2387));
    outputs(2427) <= layer2_outputs(4423);
    outputs(2428) <= not(layer2_outputs(4342));
    outputs(2429) <= not(layer2_outputs(3376));
    outputs(2430) <= layer2_outputs(2267);
    outputs(2431) <= not(layer2_outputs(216));
    outputs(2432) <= (layer2_outputs(4966)) xor (layer2_outputs(352));
    outputs(2433) <= (layer2_outputs(4622)) xor (layer2_outputs(1801));
    outputs(2434) <= not(layer2_outputs(3329));
    outputs(2435) <= layer2_outputs(4095);
    outputs(2436) <= not(layer2_outputs(1813));
    outputs(2437) <= layer2_outputs(4578);
    outputs(2438) <= layer2_outputs(2228);
    outputs(2439) <= layer2_outputs(4881);
    outputs(2440) <= not((layer2_outputs(1833)) or (layer2_outputs(772)));
    outputs(2441) <= layer2_outputs(4466);
    outputs(2442) <= layer2_outputs(874);
    outputs(2443) <= not((layer2_outputs(4080)) or (layer2_outputs(3900)));
    outputs(2444) <= not(layer2_outputs(4756));
    outputs(2445) <= not(layer2_outputs(970));
    outputs(2446) <= layer2_outputs(4433);
    outputs(2447) <= layer2_outputs(1917);
    outputs(2448) <= layer2_outputs(775);
    outputs(2449) <= not(layer2_outputs(3420));
    outputs(2450) <= (layer2_outputs(686)) and not (layer2_outputs(4724));
    outputs(2451) <= (layer2_outputs(252)) and not (layer2_outputs(2117));
    outputs(2452) <= (layer2_outputs(4380)) and not (layer2_outputs(2868));
    outputs(2453) <= (layer2_outputs(4257)) and not (layer2_outputs(4791));
    outputs(2454) <= not((layer2_outputs(313)) and (layer2_outputs(68)));
    outputs(2455) <= (layer2_outputs(4750)) xor (layer2_outputs(4403));
    outputs(2456) <= not(layer2_outputs(5063));
    outputs(2457) <= layer2_outputs(3609);
    outputs(2458) <= not(layer2_outputs(1560));
    outputs(2459) <= layer2_outputs(2799);
    outputs(2460) <= (layer2_outputs(1187)) and not (layer2_outputs(1030));
    outputs(2461) <= layer2_outputs(3169);
    outputs(2462) <= layer2_outputs(2087);
    outputs(2463) <= layer2_outputs(4523);
    outputs(2464) <= not((layer2_outputs(2319)) xor (layer2_outputs(3503)));
    outputs(2465) <= not(layer2_outputs(1150));
    outputs(2466) <= not(layer2_outputs(2508));
    outputs(2467) <= not(layer2_outputs(137)) or (layer2_outputs(428));
    outputs(2468) <= not(layer2_outputs(1341));
    outputs(2469) <= not(layer2_outputs(4369));
    outputs(2470) <= not(layer2_outputs(2074));
    outputs(2471) <= (layer2_outputs(3198)) and (layer2_outputs(2453));
    outputs(2472) <= layer2_outputs(5112);
    outputs(2473) <= not(layer2_outputs(1289));
    outputs(2474) <= not((layer2_outputs(147)) or (layer2_outputs(3242)));
    outputs(2475) <= not(layer2_outputs(3044));
    outputs(2476) <= not(layer2_outputs(5050));
    outputs(2477) <= layer2_outputs(2773);
    outputs(2478) <= not((layer2_outputs(1126)) xor (layer2_outputs(3127)));
    outputs(2479) <= not(layer2_outputs(2166));
    outputs(2480) <= not(layer2_outputs(2511));
    outputs(2481) <= (layer2_outputs(1925)) and not (layer2_outputs(1004));
    outputs(2482) <= layer2_outputs(4157);
    outputs(2483) <= layer2_outputs(3248);
    outputs(2484) <= not(layer2_outputs(2093));
    outputs(2485) <= layer2_outputs(5085);
    outputs(2486) <= (layer2_outputs(3159)) and not (layer2_outputs(4054));
    outputs(2487) <= not(layer2_outputs(2467));
    outputs(2488) <= layer2_outputs(2023);
    outputs(2489) <= not(layer2_outputs(4165));
    outputs(2490) <= not(layer2_outputs(4532));
    outputs(2491) <= layer2_outputs(3214);
    outputs(2492) <= not(layer2_outputs(1119));
    outputs(2493) <= not(layer2_outputs(2330));
    outputs(2494) <= (layer2_outputs(584)) and not (layer2_outputs(2627));
    outputs(2495) <= layer2_outputs(3084);
    outputs(2496) <= not((layer2_outputs(1032)) xor (layer2_outputs(3908)));
    outputs(2497) <= not(layer2_outputs(4995));
    outputs(2498) <= not(layer2_outputs(3612));
    outputs(2499) <= layer2_outputs(3554);
    outputs(2500) <= (layer2_outputs(1185)) or (layer2_outputs(3089));
    outputs(2501) <= not(layer2_outputs(3819));
    outputs(2502) <= not(layer2_outputs(4631));
    outputs(2503) <= not(layer2_outputs(448));
    outputs(2504) <= (layer2_outputs(1679)) and not (layer2_outputs(2014));
    outputs(2505) <= layer2_outputs(99);
    outputs(2506) <= (layer2_outputs(1948)) and not (layer2_outputs(855));
    outputs(2507) <= not(layer2_outputs(2533));
    outputs(2508) <= not(layer2_outputs(2202));
    outputs(2509) <= (layer2_outputs(2830)) or (layer2_outputs(1320));
    outputs(2510) <= layer2_outputs(1949);
    outputs(2511) <= not(layer2_outputs(4432));
    outputs(2512) <= layer2_outputs(4993);
    outputs(2513) <= layer2_outputs(3088);
    outputs(2514) <= layer2_outputs(2695);
    outputs(2515) <= layer2_outputs(429);
    outputs(2516) <= layer2_outputs(4728);
    outputs(2517) <= layer2_outputs(3955);
    outputs(2518) <= not((layer2_outputs(3704)) or (layer2_outputs(1914)));
    outputs(2519) <= (layer2_outputs(4363)) or (layer2_outputs(2143));
    outputs(2520) <= not(layer2_outputs(3980));
    outputs(2521) <= layer2_outputs(2907);
    outputs(2522) <= layer2_outputs(2320);
    outputs(2523) <= (layer2_outputs(4426)) and not (layer2_outputs(1735));
    outputs(2524) <= layer2_outputs(4099);
    outputs(2525) <= layer2_outputs(1060);
    outputs(2526) <= not(layer2_outputs(4962));
    outputs(2527) <= not(layer2_outputs(4416));
    outputs(2528) <= (layer2_outputs(655)) and not (layer2_outputs(2338));
    outputs(2529) <= layer2_outputs(2037);
    outputs(2530) <= layer2_outputs(89);
    outputs(2531) <= layer2_outputs(1185);
    outputs(2532) <= (layer2_outputs(1783)) and (layer2_outputs(2851));
    outputs(2533) <= layer2_outputs(197);
    outputs(2534) <= not(layer2_outputs(1037));
    outputs(2535) <= not((layer2_outputs(4794)) xor (layer2_outputs(321)));
    outputs(2536) <= (layer2_outputs(4840)) and not (layer2_outputs(5));
    outputs(2537) <= (layer2_outputs(671)) and not (layer2_outputs(2671));
    outputs(2538) <= (layer2_outputs(2369)) and (layer2_outputs(2077));
    outputs(2539) <= layer2_outputs(529);
    outputs(2540) <= not(layer2_outputs(39));
    outputs(2541) <= (layer2_outputs(2135)) and not (layer2_outputs(611));
    outputs(2542) <= layer2_outputs(924);
    outputs(2543) <= layer2_outputs(2026);
    outputs(2544) <= layer2_outputs(910);
    outputs(2545) <= not(layer2_outputs(2874)) or (layer2_outputs(1205));
    outputs(2546) <= layer2_outputs(467);
    outputs(2547) <= (layer2_outputs(2109)) and not (layer2_outputs(1885));
    outputs(2548) <= not((layer2_outputs(459)) and (layer2_outputs(4019)));
    outputs(2549) <= not(layer2_outputs(2886));
    outputs(2550) <= (layer2_outputs(4047)) and (layer2_outputs(2428));
    outputs(2551) <= not(layer2_outputs(3718));
    outputs(2552) <= layer2_outputs(301);
    outputs(2553) <= not(layer2_outputs(1945));
    outputs(2554) <= layer2_outputs(3029);
    outputs(2555) <= layer2_outputs(1414);
    outputs(2556) <= not(layer2_outputs(2515));
    outputs(2557) <= (layer2_outputs(3907)) and not (layer2_outputs(3210));
    outputs(2558) <= not(layer2_outputs(1299));
    outputs(2559) <= (layer2_outputs(922)) and not (layer2_outputs(1826));
    outputs(2560) <= layer2_outputs(2120);
    outputs(2561) <= (layer2_outputs(4651)) xor (layer2_outputs(2124));
    outputs(2562) <= not(layer2_outputs(5018));
    outputs(2563) <= layer2_outputs(1774);
    outputs(2564) <= (layer2_outputs(3894)) xor (layer2_outputs(3514));
    outputs(2565) <= layer2_outputs(1715);
    outputs(2566) <= layer2_outputs(4645);
    outputs(2567) <= layer2_outputs(3391);
    outputs(2568) <= layer2_outputs(3964);
    outputs(2569) <= not((layer2_outputs(149)) and (layer2_outputs(4244)));
    outputs(2570) <= not((layer2_outputs(2714)) xor (layer2_outputs(439)));
    outputs(2571) <= not(layer2_outputs(2122));
    outputs(2572) <= not((layer2_outputs(5065)) or (layer2_outputs(647)));
    outputs(2573) <= not(layer2_outputs(578));
    outputs(2574) <= layer2_outputs(2541);
    outputs(2575) <= not(layer2_outputs(4133));
    outputs(2576) <= layer2_outputs(679);
    outputs(2577) <= not((layer2_outputs(1390)) and (layer2_outputs(2466)));
    outputs(2578) <= not((layer2_outputs(1896)) xor (layer2_outputs(1149)));
    outputs(2579) <= layer2_outputs(2472);
    outputs(2580) <= (layer2_outputs(4895)) xor (layer2_outputs(534));
    outputs(2581) <= not((layer2_outputs(2984)) and (layer2_outputs(1222)));
    outputs(2582) <= not((layer2_outputs(1130)) xor (layer2_outputs(2998)));
    outputs(2583) <= layer2_outputs(4021);
    outputs(2584) <= not((layer2_outputs(359)) or (layer2_outputs(87)));
    outputs(2585) <= layer2_outputs(1798);
    outputs(2586) <= not(layer2_outputs(2151));
    outputs(2587) <= (layer2_outputs(2700)) xor (layer2_outputs(3811));
    outputs(2588) <= not(layer2_outputs(3782));
    outputs(2589) <= not(layer2_outputs(1875));
    outputs(2590) <= (layer2_outputs(215)) and (layer2_outputs(3628));
    outputs(2591) <= (layer2_outputs(2071)) xor (layer2_outputs(3367));
    outputs(2592) <= (layer2_outputs(1154)) xor (layer2_outputs(1357));
    outputs(2593) <= not(layer2_outputs(729));
    outputs(2594) <= layer2_outputs(4676);
    outputs(2595) <= (layer2_outputs(2842)) xor (layer2_outputs(123));
    outputs(2596) <= not(layer2_outputs(2729));
    outputs(2597) <= not(layer2_outputs(918));
    outputs(2598) <= layer2_outputs(3517);
    outputs(2599) <= not(layer2_outputs(2963));
    outputs(2600) <= layer2_outputs(2379);
    outputs(2601) <= not(layer2_outputs(1650));
    outputs(2602) <= not(layer2_outputs(291));
    outputs(2603) <= not((layer2_outputs(536)) xor (layer2_outputs(3354)));
    outputs(2604) <= not((layer2_outputs(4573)) or (layer2_outputs(2203)));
    outputs(2605) <= (layer2_outputs(4507)) and not (layer2_outputs(2943));
    outputs(2606) <= not(layer2_outputs(1749));
    outputs(2607) <= layer2_outputs(1045);
    outputs(2608) <= (layer2_outputs(1466)) and not (layer2_outputs(1646));
    outputs(2609) <= not((layer2_outputs(354)) xor (layer2_outputs(4002)));
    outputs(2610) <= layer2_outputs(2715);
    outputs(2611) <= not(layer2_outputs(1851)) or (layer2_outputs(2183));
    outputs(2612) <= not(layer2_outputs(16));
    outputs(2613) <= not(layer2_outputs(815));
    outputs(2614) <= layer2_outputs(2367);
    outputs(2615) <= not(layer2_outputs(1942));
    outputs(2616) <= not(layer2_outputs(4914));
    outputs(2617) <= layer2_outputs(1225);
    outputs(2618) <= not(layer2_outputs(4));
    outputs(2619) <= layer2_outputs(2622);
    outputs(2620) <= (layer2_outputs(61)) and not (layer2_outputs(4839));
    outputs(2621) <= not((layer2_outputs(3677)) xor (layer2_outputs(799)));
    outputs(2622) <= (layer2_outputs(2688)) xor (layer2_outputs(4439));
    outputs(2623) <= layer2_outputs(2856);
    outputs(2624) <= layer2_outputs(2274);
    outputs(2625) <= not(layer2_outputs(3244));
    outputs(2626) <= not(layer2_outputs(1646));
    outputs(2627) <= (layer2_outputs(2504)) and (layer2_outputs(1277));
    outputs(2628) <= (layer2_outputs(4319)) and not (layer2_outputs(134));
    outputs(2629) <= not(layer2_outputs(4390));
    outputs(2630) <= not(layer2_outputs(3046));
    outputs(2631) <= layer2_outputs(5078);
    outputs(2632) <= not(layer2_outputs(4975));
    outputs(2633) <= (layer2_outputs(1380)) xor (layer2_outputs(2025));
    outputs(2634) <= layer2_outputs(2632);
    outputs(2635) <= not(layer2_outputs(2840));
    outputs(2636) <= not(layer2_outputs(4797));
    outputs(2637) <= layer2_outputs(4764);
    outputs(2638) <= not((layer2_outputs(2465)) xor (layer2_outputs(835)));
    outputs(2639) <= not(layer2_outputs(1863));
    outputs(2640) <= not((layer2_outputs(1734)) xor (layer2_outputs(4361)));
    outputs(2641) <= not(layer2_outputs(3522));
    outputs(2642) <= not((layer2_outputs(4174)) xor (layer2_outputs(4149)));
    outputs(2643) <= not(layer2_outputs(4693));
    outputs(2644) <= layer2_outputs(2541);
    outputs(2645) <= (layer2_outputs(2044)) and (layer2_outputs(2506));
    outputs(2646) <= layer2_outputs(3135);
    outputs(2647) <= layer2_outputs(4516);
    outputs(2648) <= not(layer2_outputs(4530)) or (layer2_outputs(789));
    outputs(2649) <= (layer2_outputs(36)) or (layer2_outputs(3164));
    outputs(2650) <= (layer2_outputs(2837)) and not (layer2_outputs(190));
    outputs(2651) <= layer2_outputs(1598);
    outputs(2652) <= not(layer2_outputs(2003));
    outputs(2653) <= not(layer2_outputs(3873)) or (layer2_outputs(4323));
    outputs(2654) <= (layer2_outputs(2961)) xor (layer2_outputs(3338));
    outputs(2655) <= (layer2_outputs(4407)) and (layer2_outputs(4387));
    outputs(2656) <= not((layer2_outputs(3947)) xor (layer2_outputs(1467)));
    outputs(2657) <= not((layer2_outputs(3781)) xor (layer2_outputs(2977)));
    outputs(2658) <= (layer2_outputs(2762)) xor (layer2_outputs(3411));
    outputs(2659) <= layer2_outputs(4981);
    outputs(2660) <= (layer2_outputs(639)) and not (layer2_outputs(1260));
    outputs(2661) <= (layer2_outputs(3823)) and not (layer2_outputs(4947));
    outputs(2662) <= not(layer2_outputs(4610));
    outputs(2663) <= not(layer2_outputs(919));
    outputs(2664) <= layer2_outputs(4652);
    outputs(2665) <= not(layer2_outputs(4252));
    outputs(2666) <= not((layer2_outputs(5097)) xor (layer2_outputs(1067)));
    outputs(2667) <= not(layer2_outputs(3096));
    outputs(2668) <= layer2_outputs(3006);
    outputs(2669) <= not((layer2_outputs(2898)) xor (layer2_outputs(1248)));
    outputs(2670) <= (layer2_outputs(2312)) and not (layer2_outputs(1282));
    outputs(2671) <= layer2_outputs(335);
    outputs(2672) <= layer2_outputs(2199);
    outputs(2673) <= not(layer2_outputs(963));
    outputs(2674) <= not(layer2_outputs(3114));
    outputs(2675) <= (layer2_outputs(1584)) xor (layer2_outputs(4579));
    outputs(2676) <= layer2_outputs(3814);
    outputs(2677) <= not(layer2_outputs(1847));
    outputs(2678) <= (layer2_outputs(1296)) and (layer2_outputs(1448));
    outputs(2679) <= layer2_outputs(3603);
    outputs(2680) <= layer2_outputs(1144);
    outputs(2681) <= layer2_outputs(2082);
    outputs(2682) <= (layer2_outputs(76)) xor (layer2_outputs(3979));
    outputs(2683) <= (layer2_outputs(1334)) and (layer2_outputs(2404));
    outputs(2684) <= not(layer2_outputs(3944));
    outputs(2685) <= not(layer2_outputs(773));
    outputs(2686) <= layer2_outputs(4185);
    outputs(2687) <= layer2_outputs(3315);
    outputs(2688) <= layer2_outputs(2988);
    outputs(2689) <= not(layer2_outputs(2392));
    outputs(2690) <= (layer2_outputs(5056)) and not (layer2_outputs(3610));
    outputs(2691) <= layer2_outputs(4971);
    outputs(2692) <= not((layer2_outputs(537)) or (layer2_outputs(3571)));
    outputs(2693) <= layer2_outputs(20);
    outputs(2694) <= not(layer2_outputs(5024));
    outputs(2695) <= not((layer2_outputs(4876)) or (layer2_outputs(2152)));
    outputs(2696) <= layer2_outputs(4276);
    outputs(2697) <= (layer2_outputs(3158)) and not (layer2_outputs(1041));
    outputs(2698) <= not(layer2_outputs(3818));
    outputs(2699) <= not(layer2_outputs(2954));
    outputs(2700) <= layer2_outputs(2163);
    outputs(2701) <= (layer2_outputs(2976)) and not (layer2_outputs(2539));
    outputs(2702) <= layer2_outputs(780);
    outputs(2703) <= not(layer2_outputs(241)) or (layer2_outputs(187));
    outputs(2704) <= not((layer2_outputs(915)) xor (layer2_outputs(950)));
    outputs(2705) <= layer2_outputs(2627);
    outputs(2706) <= (layer2_outputs(3839)) xor (layer2_outputs(46));
    outputs(2707) <= not((layer2_outputs(3327)) xor (layer2_outputs(3276)));
    outputs(2708) <= not(layer2_outputs(823));
    outputs(2709) <= layer2_outputs(3890);
    outputs(2710) <= (layer2_outputs(1549)) xor (layer2_outputs(792));
    outputs(2711) <= not((layer2_outputs(4453)) xor (layer2_outputs(4525)));
    outputs(2712) <= not((layer2_outputs(4605)) xor (layer2_outputs(714)));
    outputs(2713) <= not(layer2_outputs(2265)) or (layer2_outputs(2720));
    outputs(2714) <= layer2_outputs(4539);
    outputs(2715) <= not((layer2_outputs(2805)) xor (layer2_outputs(428)));
    outputs(2716) <= not((layer2_outputs(3079)) and (layer2_outputs(2950)));
    outputs(2717) <= not(layer2_outputs(2735));
    outputs(2718) <= not(layer2_outputs(1266));
    outputs(2719) <= layer2_outputs(3796);
    outputs(2720) <= layer2_outputs(92);
    outputs(2721) <= not((layer2_outputs(4358)) xor (layer2_outputs(897)));
    outputs(2722) <= (layer2_outputs(4351)) or (layer2_outputs(2503));
    outputs(2723) <= layer2_outputs(346);
    outputs(2724) <= layer2_outputs(615);
    outputs(2725) <= (layer2_outputs(1067)) xor (layer2_outputs(4485));
    outputs(2726) <= not((layer2_outputs(78)) and (layer2_outputs(3437)));
    outputs(2727) <= layer2_outputs(1806);
    outputs(2728) <= (layer2_outputs(2598)) and not (layer2_outputs(3835));
    outputs(2729) <= layer2_outputs(4055);
    outputs(2730) <= not((layer2_outputs(3832)) xor (layer2_outputs(3535)));
    outputs(2731) <= (layer2_outputs(4773)) xor (layer2_outputs(2294));
    outputs(2732) <= layer2_outputs(1627);
    outputs(2733) <= not(layer2_outputs(2846));
    outputs(2734) <= layer2_outputs(3526);
    outputs(2735) <= layer2_outputs(2914);
    outputs(2736) <= not((layer2_outputs(837)) or (layer2_outputs(4134)));
    outputs(2737) <= not((layer2_outputs(4891)) xor (layer2_outputs(4314)));
    outputs(2738) <= not((layer2_outputs(585)) and (layer2_outputs(632)));
    outputs(2739) <= layer2_outputs(2902);
    outputs(2740) <= layer2_outputs(796);
    outputs(2741) <= layer2_outputs(604);
    outputs(2742) <= (layer2_outputs(787)) and (layer2_outputs(4833));
    outputs(2743) <= (layer2_outputs(1916)) and not (layer2_outputs(2847));
    outputs(2744) <= (layer2_outputs(1313)) xor (layer2_outputs(4418));
    outputs(2745) <= layer2_outputs(1521);
    outputs(2746) <= layer2_outputs(3208);
    outputs(2747) <= not(layer2_outputs(929));
    outputs(2748) <= (layer2_outputs(507)) and not (layer2_outputs(5052));
    outputs(2749) <= not(layer2_outputs(2214));
    outputs(2750) <= not(layer2_outputs(2697));
    outputs(2751) <= (layer2_outputs(223)) xor (layer2_outputs(4856));
    outputs(2752) <= not(layer2_outputs(2463));
    outputs(2753) <= (layer2_outputs(2196)) xor (layer2_outputs(2624));
    outputs(2754) <= not((layer2_outputs(1396)) xor (layer2_outputs(2777)));
    outputs(2755) <= not(layer2_outputs(2601));
    outputs(2756) <= (layer2_outputs(781)) xor (layer2_outputs(4828));
    outputs(2757) <= layer2_outputs(1634);
    outputs(2758) <= (layer2_outputs(2723)) and (layer2_outputs(1500));
    outputs(2759) <= not((layer2_outputs(1404)) and (layer2_outputs(973)));
    outputs(2760) <= not((layer2_outputs(5005)) xor (layer2_outputs(4770)));
    outputs(2761) <= not((layer2_outputs(526)) and (layer2_outputs(3178)));
    outputs(2762) <= layer2_outputs(1943);
    outputs(2763) <= not((layer2_outputs(4902)) xor (layer2_outputs(461)));
    outputs(2764) <= not(layer2_outputs(3248));
    outputs(2765) <= not(layer2_outputs(4588));
    outputs(2766) <= layer2_outputs(1157);
    outputs(2767) <= (layer2_outputs(2310)) xor (layer2_outputs(1760));
    outputs(2768) <= not(layer2_outputs(309)) or (layer2_outputs(1073));
    outputs(2769) <= not(layer2_outputs(3431));
    outputs(2770) <= layer2_outputs(330);
    outputs(2771) <= (layer2_outputs(3031)) and not (layer2_outputs(2599));
    outputs(2772) <= layer2_outputs(4510);
    outputs(2773) <= (layer2_outputs(3957)) or (layer2_outputs(2808));
    outputs(2774) <= not((layer2_outputs(1729)) xor (layer2_outputs(343)));
    outputs(2775) <= not(layer2_outputs(2110));
    outputs(2776) <= not(layer2_outputs(3280));
    outputs(2777) <= (layer2_outputs(4039)) and not (layer2_outputs(4236));
    outputs(2778) <= not((layer2_outputs(2966)) xor (layer2_outputs(2380)));
    outputs(2779) <= layer2_outputs(948);
    outputs(2780) <= (layer2_outputs(3755)) and not (layer2_outputs(1854));
    outputs(2781) <= not(layer2_outputs(534)) or (layer2_outputs(555));
    outputs(2782) <= (layer2_outputs(3232)) xor (layer2_outputs(1880));
    outputs(2783) <= not(layer2_outputs(4183));
    outputs(2784) <= layer2_outputs(579);
    outputs(2785) <= layer2_outputs(1887);
    outputs(2786) <= layer2_outputs(4462);
    outputs(2787) <= not(layer2_outputs(3266));
    outputs(2788) <= not(layer2_outputs(3507));
    outputs(2789) <= (layer2_outputs(2299)) xor (layer2_outputs(3501));
    outputs(2790) <= layer2_outputs(618);
    outputs(2791) <= not(layer2_outputs(1241));
    outputs(2792) <= not((layer2_outputs(1632)) xor (layer2_outputs(3029)));
    outputs(2793) <= not(layer2_outputs(3174));
    outputs(2794) <= not(layer2_outputs(2690));
    outputs(2795) <= not((layer2_outputs(784)) xor (layer2_outputs(5076)));
    outputs(2796) <= (layer2_outputs(711)) and not (layer2_outputs(3641));
    outputs(2797) <= not(layer2_outputs(4358));
    outputs(2798) <= (layer2_outputs(472)) and not (layer2_outputs(2863));
    outputs(2799) <= not((layer2_outputs(180)) xor (layer2_outputs(377)));
    outputs(2800) <= layer2_outputs(2764);
    outputs(2801) <= not(layer2_outputs(4224));
    outputs(2802) <= (layer2_outputs(811)) and (layer2_outputs(732));
    outputs(2803) <= not((layer2_outputs(2709)) xor (layer2_outputs(3495)));
    outputs(2804) <= (layer2_outputs(4108)) and (layer2_outputs(698));
    outputs(2805) <= not((layer2_outputs(4326)) xor (layer2_outputs(4459)));
    outputs(2806) <= not(layer2_outputs(3856)) or (layer2_outputs(122));
    outputs(2807) <= not(layer2_outputs(4691));
    outputs(2808) <= not((layer2_outputs(4172)) or (layer2_outputs(4389)));
    outputs(2809) <= not(layer2_outputs(2388));
    outputs(2810) <= not(layer2_outputs(4426));
    outputs(2811) <= (layer2_outputs(3408)) xor (layer2_outputs(2144));
    outputs(2812) <= not(layer2_outputs(4384));
    outputs(2813) <= not(layer2_outputs(5085));
    outputs(2814) <= layer2_outputs(2657);
    outputs(2815) <= not(layer2_outputs(1078));
    outputs(2816) <= not(layer2_outputs(3555));
    outputs(2817) <= not(layer2_outputs(3913));
    outputs(2818) <= not((layer2_outputs(2741)) or (layer2_outputs(4910)));
    outputs(2819) <= not(layer2_outputs(3958));
    outputs(2820) <= layer2_outputs(2753);
    outputs(2821) <= not(layer2_outputs(1589));
    outputs(2822) <= not(layer2_outputs(4062)) or (layer2_outputs(3202));
    outputs(2823) <= not(layer2_outputs(3334));
    outputs(2824) <= (layer2_outputs(3395)) and not (layer2_outputs(4904));
    outputs(2825) <= not(layer2_outputs(5051));
    outputs(2826) <= not(layer2_outputs(3953));
    outputs(2827) <= (layer2_outputs(4489)) or (layer2_outputs(1724));
    outputs(2828) <= layer2_outputs(4052);
    outputs(2829) <= not(layer2_outputs(3855));
    outputs(2830) <= not(layer2_outputs(3566));
    outputs(2831) <= not(layer2_outputs(2876));
    outputs(2832) <= layer2_outputs(5041);
    outputs(2833) <= layer2_outputs(2490);
    outputs(2834) <= not(layer2_outputs(1295));
    outputs(2835) <= not(layer2_outputs(1755));
    outputs(2836) <= not((layer2_outputs(3673)) xor (layer2_outputs(3831)));
    outputs(2837) <= layer2_outputs(3382);
    outputs(2838) <= not((layer2_outputs(188)) xor (layer2_outputs(2631)));
    outputs(2839) <= not((layer2_outputs(940)) or (layer2_outputs(1999)));
    outputs(2840) <= not(layer2_outputs(186));
    outputs(2841) <= (layer2_outputs(1714)) and not (layer2_outputs(1110));
    outputs(2842) <= layer2_outputs(2823);
    outputs(2843) <= not((layer2_outputs(4160)) or (layer2_outputs(2932)));
    outputs(2844) <= layer2_outputs(262);
    outputs(2845) <= layer2_outputs(2290);
    outputs(2846) <= layer2_outputs(2946);
    outputs(2847) <= not(layer2_outputs(2363));
    outputs(2848) <= layer2_outputs(1865);
    outputs(2849) <= not(layer2_outputs(645)) or (layer2_outputs(110));
    outputs(2850) <= layer2_outputs(2351);
    outputs(2851) <= (layer2_outputs(4131)) and (layer2_outputs(1531));
    outputs(2852) <= not((layer2_outputs(514)) or (layer2_outputs(71)));
    outputs(2853) <= (layer2_outputs(178)) and not (layer2_outputs(2550));
    outputs(2854) <= not(layer2_outputs(1532));
    outputs(2855) <= layer2_outputs(1801);
    outputs(2856) <= not(layer2_outputs(4408));
    outputs(2857) <= not((layer2_outputs(1858)) or (layer2_outputs(4621)));
    outputs(2858) <= (layer2_outputs(3698)) and not (layer2_outputs(3016));
    outputs(2859) <= not(layer2_outputs(1018));
    outputs(2860) <= not(layer2_outputs(158));
    outputs(2861) <= layer2_outputs(3733);
    outputs(2862) <= not(layer2_outputs(740));
    outputs(2863) <= layer2_outputs(2915);
    outputs(2864) <= layer2_outputs(867);
    outputs(2865) <= (layer2_outputs(1013)) and (layer2_outputs(4271));
    outputs(2866) <= layer2_outputs(892);
    outputs(2867) <= layer2_outputs(1930);
    outputs(2868) <= not(layer2_outputs(4316)) or (layer2_outputs(1489));
    outputs(2869) <= (layer2_outputs(3273)) xor (layer2_outputs(4941));
    outputs(2870) <= not((layer2_outputs(1259)) or (layer2_outputs(748)));
    outputs(2871) <= not((layer2_outputs(3546)) and (layer2_outputs(5067)));
    outputs(2872) <= not(layer2_outputs(1135));
    outputs(2873) <= layer2_outputs(794);
    outputs(2874) <= not(layer2_outputs(4614));
    outputs(2875) <= layer2_outputs(3158);
    outputs(2876) <= not((layer2_outputs(3558)) and (layer2_outputs(4066)));
    outputs(2877) <= not((layer2_outputs(485)) or (layer2_outputs(2864)));
    outputs(2878) <= layer2_outputs(3284);
    outputs(2879) <= not(layer2_outputs(3344)) or (layer2_outputs(164));
    outputs(2880) <= layer2_outputs(1111);
    outputs(2881) <= layer2_outputs(3333);
    outputs(2882) <= not(layer2_outputs(1695));
    outputs(2883) <= not(layer2_outputs(902));
    outputs(2884) <= (layer2_outputs(1107)) and (layer2_outputs(1624));
    outputs(2885) <= not(layer2_outputs(4058));
    outputs(2886) <= not((layer2_outputs(1209)) and (layer2_outputs(4047)));
    outputs(2887) <= not((layer2_outputs(1156)) or (layer2_outputs(3392)));
    outputs(2888) <= not((layer2_outputs(1953)) and (layer2_outputs(1008)));
    outputs(2889) <= not((layer2_outputs(2476)) xor (layer2_outputs(4798)));
    outputs(2890) <= not(layer2_outputs(4854));
    outputs(2891) <= layer2_outputs(2923);
    outputs(2892) <= layer2_outputs(1173);
    outputs(2893) <= not(layer2_outputs(3215));
    outputs(2894) <= layer2_outputs(575);
    outputs(2895) <= layer2_outputs(680);
    outputs(2896) <= (layer2_outputs(4141)) xor (layer2_outputs(1819));
    outputs(2897) <= layer2_outputs(581);
    outputs(2898) <= not(layer2_outputs(4303));
    outputs(2899) <= layer2_outputs(480);
    outputs(2900) <= (layer2_outputs(3308)) xor (layer2_outputs(1123));
    outputs(2901) <= layer2_outputs(2828);
    outputs(2902) <= not((layer2_outputs(1696)) and (layer2_outputs(1988)));
    outputs(2903) <= layer2_outputs(4921);
    outputs(2904) <= not(layer2_outputs(1790)) or (layer2_outputs(583));
    outputs(2905) <= not(layer2_outputs(4010));
    outputs(2906) <= not(layer2_outputs(1215)) or (layer2_outputs(5046));
    outputs(2907) <= not(layer2_outputs(1709));
    outputs(2908) <= not((layer2_outputs(2666)) and (layer2_outputs(1307)));
    outputs(2909) <= (layer2_outputs(1533)) xor (layer2_outputs(4005));
    outputs(2910) <= not(layer2_outputs(1381));
    outputs(2911) <= layer2_outputs(174);
    outputs(2912) <= not(layer2_outputs(3274)) or (layer2_outputs(2556));
    outputs(2913) <= not(layer2_outputs(4686));
    outputs(2914) <= (layer2_outputs(1750)) and not (layer2_outputs(3893));
    outputs(2915) <= not(layer2_outputs(3115));
    outputs(2916) <= (layer2_outputs(4291)) and not (layer2_outputs(1234));
    outputs(2917) <= not(layer2_outputs(573));
    outputs(2918) <= not(layer2_outputs(4608));
    outputs(2919) <= layer2_outputs(376);
    outputs(2920) <= (layer2_outputs(1402)) xor (layer2_outputs(1731));
    outputs(2921) <= not((layer2_outputs(716)) xor (layer2_outputs(988)));
    outputs(2922) <= layer2_outputs(1440);
    outputs(2923) <= not(layer2_outputs(631));
    outputs(2924) <= layer2_outputs(214);
    outputs(2925) <= layer2_outputs(3373);
    outputs(2926) <= (layer2_outputs(781)) xor (layer2_outputs(1343));
    outputs(2927) <= layer2_outputs(580);
    outputs(2928) <= not(layer2_outputs(3985));
    outputs(2929) <= not(layer2_outputs(2867));
    outputs(2930) <= layer2_outputs(1774);
    outputs(2931) <= layer2_outputs(2596);
    outputs(2932) <= not(layer2_outputs(1403));
    outputs(2933) <= layer2_outputs(4559);
    outputs(2934) <= not((layer2_outputs(1319)) xor (layer2_outputs(273)));
    outputs(2935) <= (layer2_outputs(297)) and (layer2_outputs(2185));
    outputs(2936) <= layer2_outputs(4753);
    outputs(2937) <= layer2_outputs(4769);
    outputs(2938) <= layer2_outputs(271);
    outputs(2939) <= (layer2_outputs(374)) and not (layer2_outputs(3555));
    outputs(2940) <= not(layer2_outputs(2713));
    outputs(2941) <= (layer2_outputs(2093)) or (layer2_outputs(3579));
    outputs(2942) <= not(layer2_outputs(513));
    outputs(2943) <= layer2_outputs(4330);
    outputs(2944) <= (layer2_outputs(4310)) and not (layer2_outputs(1000));
    outputs(2945) <= (layer2_outputs(150)) and not (layer2_outputs(248));
    outputs(2946) <= not(layer2_outputs(2727));
    outputs(2947) <= (layer2_outputs(280)) or (layer2_outputs(1752));
    outputs(2948) <= not(layer2_outputs(2774));
    outputs(2949) <= layer2_outputs(984);
    outputs(2950) <= layer2_outputs(3928);
    outputs(2951) <= not((layer2_outputs(3925)) and (layer2_outputs(1097)));
    outputs(2952) <= layer2_outputs(5017);
    outputs(2953) <= not(layer2_outputs(903));
    outputs(2954) <= not(layer2_outputs(647));
    outputs(2955) <= layer2_outputs(3427);
    outputs(2956) <= not((layer2_outputs(1101)) xor (layer2_outputs(681)));
    outputs(2957) <= not(layer2_outputs(2774)) or (layer2_outputs(2406));
    outputs(2958) <= not(layer2_outputs(1080)) or (layer2_outputs(3767));
    outputs(2959) <= not((layer2_outputs(2864)) or (layer2_outputs(1789)));
    outputs(2960) <= not(layer2_outputs(2369));
    outputs(2961) <= layer2_outputs(644);
    outputs(2962) <= layer2_outputs(3848);
    outputs(2963) <= not((layer2_outputs(3520)) xor (layer2_outputs(3478)));
    outputs(2964) <= not((layer2_outputs(1367)) or (layer2_outputs(3841)));
    outputs(2965) <= not((layer2_outputs(3468)) or (layer2_outputs(167)));
    outputs(2966) <= (layer2_outputs(4006)) xor (layer2_outputs(4672));
    outputs(2967) <= not(layer2_outputs(4205));
    outputs(2968) <= not(layer2_outputs(1615));
    outputs(2969) <= not(layer2_outputs(1967));
    outputs(2970) <= layer2_outputs(4785);
    outputs(2971) <= not((layer2_outputs(4871)) or (layer2_outputs(2112)));
    outputs(2972) <= not(layer2_outputs(4434));
    outputs(2973) <= not(layer2_outputs(2153)) or (layer2_outputs(3448));
    outputs(2974) <= not((layer2_outputs(4927)) xor (layer2_outputs(2636)));
    outputs(2975) <= layer2_outputs(3592);
    outputs(2976) <= not(layer2_outputs(4192));
    outputs(2977) <= not(layer2_outputs(1665));
    outputs(2978) <= not(layer2_outputs(75));
    outputs(2979) <= not((layer2_outputs(3752)) and (layer2_outputs(1056)));
    outputs(2980) <= (layer2_outputs(2514)) xor (layer2_outputs(4607));
    outputs(2981) <= not(layer2_outputs(4087));
    outputs(2982) <= layer2_outputs(3061);
    outputs(2983) <= not(layer2_outputs(2838));
    outputs(2984) <= not((layer2_outputs(3297)) xor (layer2_outputs(3451)));
    outputs(2985) <= layer2_outputs(1799);
    outputs(2986) <= not(layer2_outputs(963));
    outputs(2987) <= not(layer2_outputs(3394));
    outputs(2988) <= (layer2_outputs(1036)) and (layer2_outputs(1955));
    outputs(2989) <= not((layer2_outputs(3994)) xor (layer2_outputs(1261)));
    outputs(2990) <= layer2_outputs(4790);
    outputs(2991) <= layer2_outputs(776);
    outputs(2992) <= not((layer2_outputs(4053)) and (layer2_outputs(4332)));
    outputs(2993) <= not(layer2_outputs(2997)) or (layer2_outputs(2566));
    outputs(2994) <= layer2_outputs(693);
    outputs(2995) <= not((layer2_outputs(2651)) xor (layer2_outputs(288)));
    outputs(2996) <= layer2_outputs(3192);
    outputs(2997) <= not(layer2_outputs(3650));
    outputs(2998) <= (layer2_outputs(1940)) and not (layer2_outputs(5098));
    outputs(2999) <= not(layer2_outputs(2184)) or (layer2_outputs(1396));
    outputs(3000) <= not(layer2_outputs(4917));
    outputs(3001) <= not(layer2_outputs(554));
    outputs(3002) <= (layer2_outputs(3373)) xor (layer2_outputs(3636));
    outputs(3003) <= layer2_outputs(2038);
    outputs(3004) <= not(layer2_outputs(1049));
    outputs(3005) <= not(layer2_outputs(3552));
    outputs(3006) <= not(layer2_outputs(3700));
    outputs(3007) <= (layer2_outputs(2729)) xor (layer2_outputs(4430));
    outputs(3008) <= not(layer2_outputs(3934));
    outputs(3009) <= (layer2_outputs(1609)) and not (layer2_outputs(3805));
    outputs(3010) <= not(layer2_outputs(1826));
    outputs(3011) <= not(layer2_outputs(4292)) or (layer2_outputs(906));
    outputs(3012) <= not((layer2_outputs(548)) or (layer2_outputs(1859)));
    outputs(3013) <= not((layer2_outputs(2217)) xor (layer2_outputs(5026)));
    outputs(3014) <= layer2_outputs(1555);
    outputs(3015) <= layer2_outputs(3066);
    outputs(3016) <= not((layer2_outputs(4171)) and (layer2_outputs(1696)));
    outputs(3017) <= layer2_outputs(4961);
    outputs(3018) <= not(layer2_outputs(758));
    outputs(3019) <= layer2_outputs(184);
    outputs(3020) <= not(layer2_outputs(1418));
    outputs(3021) <= (layer2_outputs(1991)) xor (layer2_outputs(657));
    outputs(3022) <= not(layer2_outputs(3620));
    outputs(3023) <= not(layer2_outputs(61));
    outputs(3024) <= layer2_outputs(2326);
    outputs(3025) <= not(layer2_outputs(4997));
    outputs(3026) <= (layer2_outputs(3776)) xor (layer2_outputs(3267));
    outputs(3027) <= not(layer2_outputs(3641));
    outputs(3028) <= layer2_outputs(4566);
    outputs(3029) <= not(layer2_outputs(1875));
    outputs(3030) <= layer2_outputs(2279);
    outputs(3031) <= (layer2_outputs(2385)) xor (layer2_outputs(4414));
    outputs(3032) <= layer2_outputs(1751);
    outputs(3033) <= not(layer2_outputs(1134));
    outputs(3034) <= layer2_outputs(4097);
    outputs(3035) <= layer2_outputs(1441);
    outputs(3036) <= layer2_outputs(182);
    outputs(3037) <= layer2_outputs(282);
    outputs(3038) <= (layer2_outputs(2299)) and (layer2_outputs(1576));
    outputs(3039) <= not(layer2_outputs(4816));
    outputs(3040) <= (layer2_outputs(1476)) and not (layer2_outputs(1234));
    outputs(3041) <= layer2_outputs(417);
    outputs(3042) <= not(layer2_outputs(5068));
    outputs(3043) <= (layer2_outputs(4890)) and (layer2_outputs(4823));
    outputs(3044) <= not(layer2_outputs(4014));
    outputs(3045) <= not(layer2_outputs(2821));
    outputs(3046) <= not(layer2_outputs(2460));
    outputs(3047) <= not((layer2_outputs(3440)) xor (layer2_outputs(4871)));
    outputs(3048) <= layer2_outputs(507);
    outputs(3049) <= not(layer2_outputs(219)) or (layer2_outputs(4537));
    outputs(3050) <= layer2_outputs(3966);
    outputs(3051) <= (layer2_outputs(1887)) and not (layer2_outputs(3976));
    outputs(3052) <= not(layer2_outputs(1733));
    outputs(3053) <= layer2_outputs(1409);
    outputs(3054) <= (layer2_outputs(720)) and (layer2_outputs(4185));
    outputs(3055) <= not(layer2_outputs(2512));
    outputs(3056) <= not(layer2_outputs(3317));
    outputs(3057) <= layer2_outputs(96);
    outputs(3058) <= not(layer2_outputs(3560));
    outputs(3059) <= not(layer2_outputs(2807));
    outputs(3060) <= not(layer2_outputs(3867));
    outputs(3061) <= not(layer2_outputs(3335));
    outputs(3062) <= layer2_outputs(4602);
    outputs(3063) <= not(layer2_outputs(3424));
    outputs(3064) <= layer2_outputs(4333);
    outputs(3065) <= layer2_outputs(811);
    outputs(3066) <= (layer2_outputs(5013)) and not (layer2_outputs(2749));
    outputs(3067) <= (layer2_outputs(3445)) and (layer2_outputs(1938));
    outputs(3068) <= layer2_outputs(4557);
    outputs(3069) <= (layer2_outputs(2986)) or (layer2_outputs(1111));
    outputs(3070) <= not(layer2_outputs(4284));
    outputs(3071) <= not(layer2_outputs(3290));
    outputs(3072) <= not(layer2_outputs(4778)) or (layer2_outputs(2221));
    outputs(3073) <= layer2_outputs(3226);
    outputs(3074) <= not(layer2_outputs(282));
    outputs(3075) <= not(layer2_outputs(4225));
    outputs(3076) <= layer2_outputs(1046);
    outputs(3077) <= not(layer2_outputs(1051));
    outputs(3078) <= not(layer2_outputs(4056));
    outputs(3079) <= layer2_outputs(2489);
    outputs(3080) <= not(layer2_outputs(234));
    outputs(3081) <= layer2_outputs(4389);
    outputs(3082) <= layer2_outputs(349);
    outputs(3083) <= (layer2_outputs(3557)) xor (layer2_outputs(3688));
    outputs(3084) <= layer2_outputs(2102);
    outputs(3085) <= layer2_outputs(450);
    outputs(3086) <= layer2_outputs(3955);
    outputs(3087) <= layer2_outputs(2926);
    outputs(3088) <= layer2_outputs(3951);
    outputs(3089) <= layer2_outputs(3712);
    outputs(3090) <= layer2_outputs(2752);
    outputs(3091) <= not(layer2_outputs(3572));
    outputs(3092) <= layer2_outputs(4861);
    outputs(3093) <= not((layer2_outputs(2684)) or (layer2_outputs(2885)));
    outputs(3094) <= not(layer2_outputs(2568));
    outputs(3095) <= (layer2_outputs(3085)) xor (layer2_outputs(3466));
    outputs(3096) <= layer2_outputs(3195);
    outputs(3097) <= layer2_outputs(540);
    outputs(3098) <= not(layer2_outputs(476));
    outputs(3099) <= not(layer2_outputs(4868));
    outputs(3100) <= layer2_outputs(2629);
    outputs(3101) <= layer2_outputs(1642);
    outputs(3102) <= layer2_outputs(1927);
    outputs(3103) <= (layer2_outputs(3002)) xor (layer2_outputs(3201));
    outputs(3104) <= (layer2_outputs(2138)) or (layer2_outputs(152));
    outputs(3105) <= not(layer2_outputs(3771));
    outputs(3106) <= layer2_outputs(670);
    outputs(3107) <= layer2_outputs(2118);
    outputs(3108) <= not(layer2_outputs(3043));
    outputs(3109) <= not(layer2_outputs(956));
    outputs(3110) <= not(layer2_outputs(140)) or (layer2_outputs(4238));
    outputs(3111) <= not(layer2_outputs(37));
    outputs(3112) <= not((layer2_outputs(2829)) and (layer2_outputs(4473)));
    outputs(3113) <= not(layer2_outputs(2563)) or (layer2_outputs(453));
    outputs(3114) <= layer2_outputs(1815);
    outputs(3115) <= layer2_outputs(136);
    outputs(3116) <= layer2_outputs(2358);
    outputs(3117) <= layer2_outputs(1246);
    outputs(3118) <= not((layer2_outputs(4217)) and (layer2_outputs(1090)));
    outputs(3119) <= not(layer2_outputs(2978));
    outputs(3120) <= not(layer2_outputs(813));
    outputs(3121) <= (layer2_outputs(319)) and (layer2_outputs(1485));
    outputs(3122) <= not(layer2_outputs(228));
    outputs(3123) <= layer2_outputs(5110);
    outputs(3124) <= not(layer2_outputs(4767));
    outputs(3125) <= not(layer2_outputs(4896));
    outputs(3126) <= layer2_outputs(152);
    outputs(3127) <= layer2_outputs(1105);
    outputs(3128) <= (layer2_outputs(1169)) or (layer2_outputs(2444));
    outputs(3129) <= layer2_outputs(3464);
    outputs(3130) <= layer2_outputs(4521);
    outputs(3131) <= not(layer2_outputs(3256)) or (layer2_outputs(1752));
    outputs(3132) <= layer2_outputs(1452);
    outputs(3133) <= layer2_outputs(3331);
    outputs(3134) <= (layer2_outputs(3425)) and not (layer2_outputs(564));
    outputs(3135) <= (layer2_outputs(3449)) and not (layer2_outputs(2357));
    outputs(3136) <= (layer2_outputs(4461)) or (layer2_outputs(4379));
    outputs(3137) <= not((layer2_outputs(1619)) xor (layer2_outputs(4320)));
    outputs(3138) <= not(layer2_outputs(1380));
    outputs(3139) <= not(layer2_outputs(1670));
    outputs(3140) <= not((layer2_outputs(2335)) or (layer2_outputs(2594)));
    outputs(3141) <= (layer2_outputs(2157)) and (layer2_outputs(404));
    outputs(3142) <= not(layer2_outputs(4580));
    outputs(3143) <= layer2_outputs(2801);
    outputs(3144) <= not(layer2_outputs(587));
    outputs(3145) <= layer2_outputs(105);
    outputs(3146) <= not(layer2_outputs(393));
    outputs(3147) <= (layer2_outputs(3975)) and not (layer2_outputs(3940));
    outputs(3148) <= not((layer2_outputs(3070)) xor (layer2_outputs(2426)));
    outputs(3149) <= not(layer2_outputs(598)) or (layer2_outputs(31));
    outputs(3150) <= layer2_outputs(4248);
    outputs(3151) <= layer2_outputs(4694);
    outputs(3152) <= layer2_outputs(4987);
    outputs(3153) <= layer2_outputs(2292);
    outputs(3154) <= not(layer2_outputs(3672));
    outputs(3155) <= not((layer2_outputs(2643)) xor (layer2_outputs(2835)));
    outputs(3156) <= layer2_outputs(4898);
    outputs(3157) <= layer2_outputs(5010);
    outputs(3158) <= not(layer2_outputs(756));
    outputs(3159) <= layer2_outputs(735);
    outputs(3160) <= not(layer2_outputs(3352));
    outputs(3161) <= layer2_outputs(1843);
    outputs(3162) <= not(layer2_outputs(2176));
    outputs(3163) <= not(layer2_outputs(4213));
    outputs(3164) <= not(layer2_outputs(1081));
    outputs(3165) <= not(layer2_outputs(4204));
    outputs(3166) <= not(layer2_outputs(921));
    outputs(3167) <= layer2_outputs(1407);
    outputs(3168) <= not(layer2_outputs(4385));
    outputs(3169) <= layer2_outputs(824);
    outputs(3170) <= not(layer2_outputs(2612)) or (layer2_outputs(2090));
    outputs(3171) <= layer2_outputs(4961);
    outputs(3172) <= layer2_outputs(3046);
    outputs(3173) <= layer2_outputs(1793);
    outputs(3174) <= layer2_outputs(4051);
    outputs(3175) <= layer2_outputs(1003);
    outputs(3176) <= not(layer2_outputs(4171));
    outputs(3177) <= not(layer2_outputs(1993));
    outputs(3178) <= not((layer2_outputs(1285)) xor (layer2_outputs(4722)));
    outputs(3179) <= layer2_outputs(4191);
    outputs(3180) <= layer2_outputs(641);
    outputs(3181) <= layer2_outputs(4096);
    outputs(3182) <= not(layer2_outputs(1854));
    outputs(3183) <= layer2_outputs(3323);
    outputs(3184) <= not(layer2_outputs(2377));
    outputs(3185) <= not(layer2_outputs(3330));
    outputs(3186) <= layer2_outputs(2047);
    outputs(3187) <= (layer2_outputs(1128)) and (layer2_outputs(3097));
    outputs(3188) <= (layer2_outputs(3748)) or (layer2_outputs(2053));
    outputs(3189) <= layer2_outputs(1832);
    outputs(3190) <= not(layer2_outputs(1022));
    outputs(3191) <= (layer2_outputs(1764)) and not (layer2_outputs(2481));
    outputs(3192) <= (layer2_outputs(3177)) and not (layer2_outputs(1891));
    outputs(3193) <= not(layer2_outputs(2594));
    outputs(3194) <= not(layer2_outputs(3852));
    outputs(3195) <= not(layer2_outputs(3873));
    outputs(3196) <= not(layer2_outputs(3988));
    outputs(3197) <= layer2_outputs(4021);
    outputs(3198) <= not(layer2_outputs(1232));
    outputs(3199) <= (layer2_outputs(2048)) xor (layer2_outputs(3299));
    outputs(3200) <= layer2_outputs(3498);
    outputs(3201) <= not(layer2_outputs(4452));
    outputs(3202) <= not(layer2_outputs(4958));
    outputs(3203) <= layer2_outputs(2020);
    outputs(3204) <= layer2_outputs(2047);
    outputs(3205) <= layer2_outputs(1217);
    outputs(3206) <= layer2_outputs(820);
    outputs(3207) <= layer2_outputs(1505);
    outputs(3208) <= layer2_outputs(2110);
    outputs(3209) <= not((layer2_outputs(1655)) xor (layer2_outputs(4912)));
    outputs(3210) <= not(layer2_outputs(3107));
    outputs(3211) <= not(layer2_outputs(3724));
    outputs(3212) <= not(layer2_outputs(3216));
    outputs(3213) <= not((layer2_outputs(1011)) or (layer2_outputs(3149)));
    outputs(3214) <= layer2_outputs(3127);
    outputs(3215) <= layer2_outputs(872);
    outputs(3216) <= not(layer2_outputs(192));
    outputs(3217) <= layer2_outputs(4233);
    outputs(3218) <= layer2_outputs(1800);
    outputs(3219) <= not(layer2_outputs(259));
    outputs(3220) <= not(layer2_outputs(909)) or (layer2_outputs(4937));
    outputs(3221) <= (layer2_outputs(1439)) and not (layer2_outputs(3833));
    outputs(3222) <= not(layer2_outputs(3311));
    outputs(3223) <= not(layer2_outputs(3532));
    outputs(3224) <= (layer2_outputs(3859)) and not (layer2_outputs(4478));
    outputs(3225) <= not(layer2_outputs(1325));
    outputs(3226) <= layer2_outputs(3524);
    outputs(3227) <= (layer2_outputs(1831)) and not (layer2_outputs(3284));
    outputs(3228) <= (layer2_outputs(296)) and (layer2_outputs(170));
    outputs(3229) <= not(layer2_outputs(3028));
    outputs(3230) <= layer2_outputs(977);
    outputs(3231) <= layer2_outputs(3059);
    outputs(3232) <= not(layer2_outputs(4382));
    outputs(3233) <= not(layer2_outputs(2866));
    outputs(3234) <= layer2_outputs(1239);
    outputs(3235) <= not(layer2_outputs(4690));
    outputs(3236) <= (layer2_outputs(3465)) and (layer2_outputs(531));
    outputs(3237) <= not(layer2_outputs(2298)) or (layer2_outputs(5087));
    outputs(3238) <= not(layer2_outputs(1809));
    outputs(3239) <= not(layer2_outputs(5055));
    outputs(3240) <= layer2_outputs(1333);
    outputs(3241) <= not(layer2_outputs(444));
    outputs(3242) <= not((layer2_outputs(1637)) xor (layer2_outputs(1619)));
    outputs(3243) <= not(layer2_outputs(2343));
    outputs(3244) <= not((layer2_outputs(3372)) or (layer2_outputs(1343)));
    outputs(3245) <= layer2_outputs(1190);
    outputs(3246) <= layer2_outputs(154);
    outputs(3247) <= not(layer2_outputs(1022));
    outputs(3248) <= layer2_outputs(4353);
    outputs(3249) <= layer2_outputs(1456);
    outputs(3250) <= layer2_outputs(3410);
    outputs(3251) <= not(layer2_outputs(5118));
    outputs(3252) <= not(layer2_outputs(5019)) or (layer2_outputs(4703));
    outputs(3253) <= not(layer2_outputs(2545));
    outputs(3254) <= not(layer2_outputs(3254));
    outputs(3255) <= layer2_outputs(3325);
    outputs(3256) <= not((layer2_outputs(1313)) or (layer2_outputs(3111)));
    outputs(3257) <= not(layer2_outputs(2377)) or (layer2_outputs(5110));
    outputs(3258) <= not(layer2_outputs(624));
    outputs(3259) <= layer2_outputs(1814);
    outputs(3260) <= not(layer2_outputs(3801));
    outputs(3261) <= not((layer2_outputs(1824)) xor (layer2_outputs(689)));
    outputs(3262) <= (layer2_outputs(295)) or (layer2_outputs(2574));
    outputs(3263) <= not(layer2_outputs(498));
    outputs(3264) <= layer2_outputs(3938);
    outputs(3265) <= not(layer2_outputs(3853));
    outputs(3266) <= not(layer2_outputs(3874));
    outputs(3267) <= not(layer2_outputs(4778));
    outputs(3268) <= (layer2_outputs(10)) xor (layer2_outputs(4998));
    outputs(3269) <= not(layer2_outputs(3259)) or (layer2_outputs(4582));
    outputs(3270) <= layer2_outputs(1271);
    outputs(3271) <= layer2_outputs(2678);
    outputs(3272) <= not(layer2_outputs(2417));
    outputs(3273) <= not(layer2_outputs(37));
    outputs(3274) <= not(layer2_outputs(2176));
    outputs(3275) <= not((layer2_outputs(1518)) or (layer2_outputs(2257)));
    outputs(3276) <= (layer2_outputs(2271)) and not (layer2_outputs(4348));
    outputs(3277) <= layer2_outputs(340);
    outputs(3278) <= layer2_outputs(2954);
    outputs(3279) <= layer2_outputs(1415);
    outputs(3280) <= not(layer2_outputs(1464));
    outputs(3281) <= layer2_outputs(4345);
    outputs(3282) <= layer2_outputs(4206);
    outputs(3283) <= layer2_outputs(989);
    outputs(3284) <= not(layer2_outputs(3034));
    outputs(3285) <= (layer2_outputs(2641)) and not (layer2_outputs(2407));
    outputs(3286) <= not(layer2_outputs(1345));
    outputs(3287) <= not((layer2_outputs(2810)) xor (layer2_outputs(5113)));
    outputs(3288) <= layer2_outputs(3318);
    outputs(3289) <= layer2_outputs(3747);
    outputs(3290) <= not(layer2_outputs(3929));
    outputs(3291) <= (layer2_outputs(3117)) xor (layer2_outputs(3970));
    outputs(3292) <= layer2_outputs(2412);
    outputs(3293) <= not(layer2_outputs(2483));
    outputs(3294) <= not(layer2_outputs(597));
    outputs(3295) <= layer2_outputs(4898);
    outputs(3296) <= layer2_outputs(151);
    outputs(3297) <= layer2_outputs(1458);
    outputs(3298) <= layer2_outputs(3770);
    outputs(3299) <= (layer2_outputs(2254)) and not (layer2_outputs(441));
    outputs(3300) <= (layer2_outputs(4106)) and (layer2_outputs(2427));
    outputs(3301) <= (layer2_outputs(1174)) and not (layer2_outputs(5088));
    outputs(3302) <= not(layer2_outputs(3249));
    outputs(3303) <= not(layer2_outputs(2724));
    outputs(3304) <= layer2_outputs(4096);
    outputs(3305) <= not(layer2_outputs(2917));
    outputs(3306) <= not(layer2_outputs(5039)) or (layer2_outputs(4283));
    outputs(3307) <= not(layer2_outputs(4979));
    outputs(3308) <= layer2_outputs(1603);
    outputs(3309) <= layer2_outputs(1456);
    outputs(3310) <= not(layer2_outputs(3825));
    outputs(3311) <= not(layer2_outputs(3259));
    outputs(3312) <= (layer2_outputs(4616)) and not (layer2_outputs(2687));
    outputs(3313) <= layer2_outputs(819);
    outputs(3314) <= layer2_outputs(3975);
    outputs(3315) <= not(layer2_outputs(144));
    outputs(3316) <= layer2_outputs(1573);
    outputs(3317) <= layer2_outputs(984);
    outputs(3318) <= (layer2_outputs(3480)) and not (layer2_outputs(3663));
    outputs(3319) <= (layer2_outputs(3978)) xor (layer2_outputs(3013));
    outputs(3320) <= not(layer2_outputs(1287));
    outputs(3321) <= (layer2_outputs(3512)) and not (layer2_outputs(2525));
    outputs(3322) <= not(layer2_outputs(2728));
    outputs(3323) <= (layer2_outputs(5065)) and not (layer2_outputs(2744));
    outputs(3324) <= not(layer2_outputs(2454));
    outputs(3325) <= layer2_outputs(177);
    outputs(3326) <= layer2_outputs(740);
    outputs(3327) <= layer2_outputs(169);
    outputs(3328) <= not(layer2_outputs(3905));
    outputs(3329) <= not(layer2_outputs(4477));
    outputs(3330) <= not((layer2_outputs(5060)) and (layer2_outputs(222)));
    outputs(3331) <= layer2_outputs(4184);
    outputs(3332) <= not(layer2_outputs(2984));
    outputs(3333) <= (layer2_outputs(3545)) and not (layer2_outputs(1348));
    outputs(3334) <= not((layer2_outputs(2602)) and (layer2_outputs(2382)));
    outputs(3335) <= layer2_outputs(2447);
    outputs(3336) <= not(layer2_outputs(4981));
    outputs(3337) <= not((layer2_outputs(368)) xor (layer2_outputs(3756)));
    outputs(3338) <= not(layer2_outputs(126));
    outputs(3339) <= not(layer2_outputs(1310));
    outputs(3340) <= not((layer2_outputs(1837)) or (layer2_outputs(3837)));
    outputs(3341) <= not(layer2_outputs(3882)) or (layer2_outputs(54));
    outputs(3342) <= (layer2_outputs(2455)) and (layer2_outputs(26));
    outputs(3343) <= not((layer2_outputs(1364)) xor (layer2_outputs(2556)));
    outputs(3344) <= layer2_outputs(3684);
    outputs(3345) <= layer2_outputs(4867);
    outputs(3346) <= layer2_outputs(1501);
    outputs(3347) <= not((layer2_outputs(3096)) xor (layer2_outputs(446)));
    outputs(3348) <= layer2_outputs(2368);
    outputs(3349) <= layer2_outputs(648);
    outputs(3350) <= not((layer2_outputs(5028)) or (layer2_outputs(1411)));
    outputs(3351) <= layer2_outputs(4265);
    outputs(3352) <= (layer2_outputs(1206)) xor (layer2_outputs(849));
    outputs(3353) <= (layer2_outputs(4702)) xor (layer2_outputs(2081));
    outputs(3354) <= not(layer2_outputs(3479));
    outputs(3355) <= not(layer2_outputs(16)) or (layer2_outputs(741));
    outputs(3356) <= not(layer2_outputs(2789));
    outputs(3357) <= layer2_outputs(2064);
    outputs(3358) <= not((layer2_outputs(778)) xor (layer2_outputs(1791)));
    outputs(3359) <= layer2_outputs(1983);
    outputs(3360) <= not(layer2_outputs(4359));
    outputs(3361) <= not((layer2_outputs(3226)) xor (layer2_outputs(404)));
    outputs(3362) <= layer2_outputs(218);
    outputs(3363) <= layer2_outputs(3086);
    outputs(3364) <= layer2_outputs(3927);
    outputs(3365) <= (layer2_outputs(3918)) and not (layer2_outputs(3603));
    outputs(3366) <= layer2_outputs(3082);
    outputs(3367) <= layer2_outputs(399);
    outputs(3368) <= layer2_outputs(4345);
    outputs(3369) <= layer2_outputs(2600);
    outputs(3370) <= not((layer2_outputs(3568)) or (layer2_outputs(2852)));
    outputs(3371) <= not((layer2_outputs(1841)) xor (layer2_outputs(313)));
    outputs(3372) <= not(layer2_outputs(673));
    outputs(3373) <= (layer2_outputs(4657)) and not (layer2_outputs(446));
    outputs(3374) <= not((layer2_outputs(4221)) xor (layer2_outputs(415)));
    outputs(3375) <= not(layer2_outputs(1042));
    outputs(3376) <= layer2_outputs(2913);
    outputs(3377) <= layer2_outputs(4073);
    outputs(3378) <= layer2_outputs(861);
    outputs(3379) <= layer2_outputs(4864);
    outputs(3380) <= not(layer2_outputs(2003));
    outputs(3381) <= not(layer2_outputs(3730));
    outputs(3382) <= (layer2_outputs(1096)) xor (layer2_outputs(139));
    outputs(3383) <= not(layer2_outputs(922));
    outputs(3384) <= layer2_outputs(3159);
    outputs(3385) <= not(layer2_outputs(2981));
    outputs(3386) <= not(layer2_outputs(4350));
    outputs(3387) <= (layer2_outputs(730)) and (layer2_outputs(3862));
    outputs(3388) <= not(layer2_outputs(4451));
    outputs(3389) <= layer2_outputs(3747);
    outputs(3390) <= not((layer2_outputs(204)) xor (layer2_outputs(2169)));
    outputs(3391) <= not(layer2_outputs(2995));
    outputs(3392) <= layer2_outputs(2513);
    outputs(3393) <= layer2_outputs(2362);
    outputs(3394) <= not(layer2_outputs(481));
    outputs(3395) <= not(layer2_outputs(1819));
    outputs(3396) <= not(layer2_outputs(492));
    outputs(3397) <= not(layer2_outputs(1689));
    outputs(3398) <= layer2_outputs(3393);
    outputs(3399) <= not(layer2_outputs(3864));
    outputs(3400) <= not(layer2_outputs(30));
    outputs(3401) <= layer2_outputs(4813);
    outputs(3402) <= (layer2_outputs(2933)) and not (layer2_outputs(2111));
    outputs(3403) <= not(layer2_outputs(797));
    outputs(3404) <= not(layer2_outputs(2265));
    outputs(3405) <= layer2_outputs(148);
    outputs(3406) <= not(layer2_outputs(5027));
    outputs(3407) <= (layer2_outputs(4137)) xor (layer2_outputs(3405));
    outputs(3408) <= not(layer2_outputs(4969));
    outputs(3409) <= not(layer2_outputs(324));
    outputs(3410) <= (layer2_outputs(1775)) xor (layer2_outputs(1031));
    outputs(3411) <= layer2_outputs(2472);
    outputs(3412) <= layer2_outputs(1699);
    outputs(3413) <= layer2_outputs(3389);
    outputs(3414) <= layer2_outputs(3422);
    outputs(3415) <= not(layer2_outputs(4611));
    outputs(3416) <= (layer2_outputs(1582)) and (layer2_outputs(2233));
    outputs(3417) <= layer2_outputs(3989);
    outputs(3418) <= not(layer2_outputs(456));
    outputs(3419) <= (layer2_outputs(1203)) xor (layer2_outputs(2473));
    outputs(3420) <= not(layer2_outputs(1211));
    outputs(3421) <= layer2_outputs(874);
    outputs(3422) <= layer2_outputs(2302);
    outputs(3423) <= layer2_outputs(2677);
    outputs(3424) <= not((layer2_outputs(3974)) and (layer2_outputs(1534)));
    outputs(3425) <= not(layer2_outputs(3941));
    outputs(3426) <= (layer2_outputs(2991)) and not (layer2_outputs(4637));
    outputs(3427) <= not(layer2_outputs(4307));
    outputs(3428) <= not((layer2_outputs(821)) and (layer2_outputs(2232)));
    outputs(3429) <= layer2_outputs(2832);
    outputs(3430) <= not(layer2_outputs(1902));
    outputs(3431) <= not(layer2_outputs(3663));
    outputs(3432) <= not(layer2_outputs(91));
    outputs(3433) <= not(layer2_outputs(1678));
    outputs(3434) <= not(layer2_outputs(3147));
    outputs(3435) <= not(layer2_outputs(196));
    outputs(3436) <= layer2_outputs(4315);
    outputs(3437) <= layer2_outputs(5115);
    outputs(3438) <= not(layer2_outputs(3241));
    outputs(3439) <= not(layer2_outputs(3774));
    outputs(3440) <= layer2_outputs(3696);
    outputs(3441) <= (layer2_outputs(2306)) and not (layer2_outputs(1024));
    outputs(3442) <= not(layer2_outputs(904));
    outputs(3443) <= not(layer2_outputs(2374));
    outputs(3444) <= (layer2_outputs(2035)) and not (layer2_outputs(559));
    outputs(3445) <= not(layer2_outputs(2052));
    outputs(3446) <= not(layer2_outputs(870));
    outputs(3447) <= layer2_outputs(695);
    outputs(3448) <= not((layer2_outputs(2983)) or (layer2_outputs(3772)));
    outputs(3449) <= (layer2_outputs(1946)) and (layer2_outputs(3289));
    outputs(3450) <= not(layer2_outputs(3553));
    outputs(3451) <= layer2_outputs(620);
    outputs(3452) <= layer2_outputs(895);
    outputs(3453) <= layer2_outputs(715);
    outputs(3454) <= (layer2_outputs(1172)) and not (layer2_outputs(4942));
    outputs(3455) <= not(layer2_outputs(3718));
    outputs(3456) <= not((layer2_outputs(3511)) or (layer2_outputs(1924)));
    outputs(3457) <= not(layer2_outputs(2308));
    outputs(3458) <= layer2_outputs(2286);
    outputs(3459) <= not(layer2_outputs(1779));
    outputs(3460) <= not(layer2_outputs(4119));
    outputs(3461) <= layer2_outputs(4877);
    outputs(3462) <= not(layer2_outputs(2998));
    outputs(3463) <= not(layer2_outputs(3679));
    outputs(3464) <= layer2_outputs(1117);
    outputs(3465) <= (layer2_outputs(2714)) and (layer2_outputs(4433));
    outputs(3466) <= not(layer2_outputs(674)) or (layer2_outputs(3535));
    outputs(3467) <= not(layer2_outputs(3537));
    outputs(3468) <= (layer2_outputs(584)) xor (layer2_outputs(1718));
    outputs(3469) <= (layer2_outputs(419)) xor (layer2_outputs(743));
    outputs(3470) <= layer2_outputs(1145);
    outputs(3471) <= not(layer2_outputs(3626));
    outputs(3472) <= layer2_outputs(1958);
    outputs(3473) <= not((layer2_outputs(4422)) xor (layer2_outputs(2786)));
    outputs(3474) <= layer2_outputs(2405);
    outputs(3475) <= not(layer2_outputs(2399));
    outputs(3476) <= not(layer2_outputs(1005));
    outputs(3477) <= layer2_outputs(4806);
    outputs(3478) <= not(layer2_outputs(657));
    outputs(3479) <= layer2_outputs(4747);
    outputs(3480) <= not(layer2_outputs(4025));
    outputs(3481) <= layer2_outputs(3389);
    outputs(3482) <= layer2_outputs(193);
    outputs(3483) <= (layer2_outputs(4339)) and not (layer2_outputs(1388));
    outputs(3484) <= not(layer2_outputs(655));
    outputs(3485) <= layer2_outputs(1853);
    outputs(3486) <= not(layer2_outputs(557));
    outputs(3487) <= layer2_outputs(327);
    outputs(3488) <= not(layer2_outputs(3868));
    outputs(3489) <= (layer2_outputs(837)) and not (layer2_outputs(3860));
    outputs(3490) <= (layer2_outputs(1866)) xor (layer2_outputs(2424));
    outputs(3491) <= not(layer2_outputs(1438));
    outputs(3492) <= layer2_outputs(2609);
    outputs(3493) <= layer2_outputs(1444);
    outputs(3494) <= (layer2_outputs(2064)) and not (layer2_outputs(791));
    outputs(3495) <= not(layer2_outputs(3390));
    outputs(3496) <= not(layer2_outputs(124));
    outputs(3497) <= (layer2_outputs(2139)) xor (layer2_outputs(375));
    outputs(3498) <= (layer2_outputs(2625)) xor (layer2_outputs(4974));
    outputs(3499) <= not(layer2_outputs(261));
    outputs(3500) <= layer2_outputs(5096);
    outputs(3501) <= not(layer2_outputs(4396));
    outputs(3502) <= not(layer2_outputs(23));
    outputs(3503) <= not(layer2_outputs(3847));
    outputs(3504) <= not(layer2_outputs(4280));
    outputs(3505) <= not(layer2_outputs(3980));
    outputs(3506) <= not(layer2_outputs(2177));
    outputs(3507) <= (layer2_outputs(2125)) or (layer2_outputs(1434));
    outputs(3508) <= (layer2_outputs(722)) xor (layer2_outputs(3243));
    outputs(3509) <= not(layer2_outputs(2730));
    outputs(3510) <= not(layer2_outputs(2766));
    outputs(3511) <= not(layer2_outputs(4906));
    outputs(3512) <= layer2_outputs(3328);
    outputs(3513) <= layer2_outputs(458);
    outputs(3514) <= not(layer2_outputs(3707));
    outputs(3515) <= not(layer2_outputs(1539));
    outputs(3516) <= not(layer2_outputs(4181));
    outputs(3517) <= not(layer2_outputs(589));
    outputs(3518) <= not(layer2_outputs(656));
    outputs(3519) <= not(layer2_outputs(2725));
    outputs(3520) <= layer2_outputs(3282);
    outputs(3521) <= not(layer2_outputs(3521));
    outputs(3522) <= layer2_outputs(4196);
    outputs(3523) <= layer2_outputs(3775);
    outputs(3524) <= (layer2_outputs(4784)) and not (layer2_outputs(2569));
    outputs(3525) <= (layer2_outputs(2644)) or (layer2_outputs(828));
    outputs(3526) <= not((layer2_outputs(2213)) xor (layer2_outputs(3804)));
    outputs(3527) <= not(layer2_outputs(3433));
    outputs(3528) <= (layer2_outputs(2008)) xor (layer2_outputs(1483));
    outputs(3529) <= (layer2_outputs(3275)) and not (layer2_outputs(1578));
    outputs(3530) <= layer2_outputs(1651);
    outputs(3531) <= not(layer2_outputs(972));
    outputs(3532) <= (layer2_outputs(4900)) and not (layer2_outputs(498));
    outputs(3533) <= layer2_outputs(4353);
    outputs(3534) <= not(layer2_outputs(1347));
    outputs(3535) <= not(layer2_outputs(2602));
    outputs(3536) <= layer2_outputs(1004);
    outputs(3537) <= not(layer2_outputs(4796));
    outputs(3538) <= layer2_outputs(1016);
    outputs(3539) <= not(layer2_outputs(2457));
    outputs(3540) <= layer2_outputs(1161);
    outputs(3541) <= layer2_outputs(582);
    outputs(3542) <= not(layer2_outputs(1847));
    outputs(3543) <= not(layer2_outputs(2200));
    outputs(3544) <= layer2_outputs(2600);
    outputs(3545) <= layer2_outputs(334);
    outputs(3546) <= not(layer2_outputs(4734));
    outputs(3547) <= (layer2_outputs(591)) and not (layer2_outputs(1554));
    outputs(3548) <= layer2_outputs(2676);
    outputs(3549) <= not(layer2_outputs(966));
    outputs(3550) <= layer2_outputs(1359);
    outputs(3551) <= not((layer2_outputs(83)) xor (layer2_outputs(2534)));
    outputs(3552) <= not(layer2_outputs(3424));
    outputs(3553) <= not(layer2_outputs(2171));
    outputs(3554) <= not(layer2_outputs(2177));
    outputs(3555) <= (layer2_outputs(3721)) and (layer2_outputs(3165));
    outputs(3556) <= layer2_outputs(4460);
    outputs(3557) <= layer2_outputs(1226);
    outputs(3558) <= (layer2_outputs(3045)) and (layer2_outputs(1147));
    outputs(3559) <= layer2_outputs(4199);
    outputs(3560) <= not(layer2_outputs(2605)) or (layer2_outputs(2574));
    outputs(3561) <= layer2_outputs(933);
    outputs(3562) <= (layer2_outputs(4493)) and (layer2_outputs(1623));
    outputs(3563) <= not((layer2_outputs(3656)) and (layer2_outputs(3300)));
    outputs(3564) <= not((layer2_outputs(1403)) xor (layer2_outputs(5023)));
    outputs(3565) <= layer2_outputs(1876);
    outputs(3566) <= not(layer2_outputs(2978));
    outputs(3567) <= not(layer2_outputs(1518));
    outputs(3568) <= not(layer2_outputs(4951));
    outputs(3569) <= not(layer2_outputs(1705));
    outputs(3570) <= not(layer2_outputs(4084));
    outputs(3571) <= not((layer2_outputs(4483)) and (layer2_outputs(2129)));
    outputs(3572) <= (layer2_outputs(4470)) and not (layer2_outputs(4214));
    outputs(3573) <= layer2_outputs(3923);
    outputs(3574) <= not(layer2_outputs(1743));
    outputs(3575) <= not(layer2_outputs(823));
    outputs(3576) <= layer2_outputs(641);
    outputs(3577) <= layer2_outputs(2734);
    outputs(3578) <= layer2_outputs(2504);
    outputs(3579) <= (layer2_outputs(709)) xor (layer2_outputs(4850));
    outputs(3580) <= layer2_outputs(3014);
    outputs(3581) <= not(layer2_outputs(444));
    outputs(3582) <= (layer2_outputs(1890)) and not (layer2_outputs(115));
    outputs(3583) <= (layer2_outputs(3292)) and not (layer2_outputs(2698));
    outputs(3584) <= layer2_outputs(1668);
    outputs(3585) <= (layer2_outputs(2595)) and not (layer2_outputs(1724));
    outputs(3586) <= (layer2_outputs(4109)) xor (layer2_outputs(4391));
    outputs(3587) <= not(layer2_outputs(1382));
    outputs(3588) <= (layer2_outputs(3412)) and not (layer2_outputs(2305));
    outputs(3589) <= layer2_outputs(1960);
    outputs(3590) <= (layer2_outputs(3650)) and (layer2_outputs(1182));
    outputs(3591) <= layer2_outputs(401);
    outputs(3592) <= layer2_outputs(1125);
    outputs(3593) <= not(layer2_outputs(351));
    outputs(3594) <= (layer2_outputs(1972)) or (layer2_outputs(2244));
    outputs(3595) <= layer2_outputs(1741);
    outputs(3596) <= not(layer2_outputs(3708));
    outputs(3597) <= layer2_outputs(2160);
    outputs(3598) <= (layer2_outputs(1525)) and not (layer2_outputs(3435));
    outputs(3599) <= layer2_outputs(2282);
    outputs(3600) <= (layer2_outputs(5036)) and (layer2_outputs(5043));
    outputs(3601) <= not(layer2_outputs(3184));
    outputs(3602) <= layer2_outputs(5043);
    outputs(3603) <= not((layer2_outputs(3270)) or (layer2_outputs(2188)));
    outputs(3604) <= not(layer2_outputs(4742));
    outputs(3605) <= (layer2_outputs(3071)) and not (layer2_outputs(1221));
    outputs(3606) <= (layer2_outputs(398)) and not (layer2_outputs(1138));
    outputs(3607) <= not(layer2_outputs(4643));
    outputs(3608) <= layer2_outputs(2932);
    outputs(3609) <= layer2_outputs(2846);
    outputs(3610) <= layer2_outputs(2066);
    outputs(3611) <= (layer2_outputs(2128)) and not (layer2_outputs(4287));
    outputs(3612) <= not(layer2_outputs(118));
    outputs(3613) <= not(layer2_outputs(279));
    outputs(3614) <= layer2_outputs(3240);
    outputs(3615) <= layer2_outputs(3335);
    outputs(3616) <= not(layer2_outputs(4100));
    outputs(3617) <= not(layer2_outputs(3239));
    outputs(3618) <= (layer2_outputs(758)) and not (layer2_outputs(4007));
    outputs(3619) <= (layer2_outputs(871)) xor (layer2_outputs(161));
    outputs(3620) <= not(layer2_outputs(2499));
    outputs(3621) <= (layer2_outputs(4436)) and not (layer2_outputs(3701));
    outputs(3622) <= (layer2_outputs(4031)) and (layer2_outputs(1647));
    outputs(3623) <= (layer2_outputs(4331)) and not (layer2_outputs(3));
    outputs(3624) <= layer2_outputs(1918);
    outputs(3625) <= layer2_outputs(2756);
    outputs(3626) <= layer2_outputs(721);
    outputs(3627) <= layer2_outputs(848);
    outputs(3628) <= layer2_outputs(3706);
    outputs(3629) <= not((layer2_outputs(2845)) or (layer2_outputs(4603)));
    outputs(3630) <= layer2_outputs(3122);
    outputs(3631) <= layer2_outputs(2001);
    outputs(3632) <= layer2_outputs(3021);
    outputs(3633) <= (layer2_outputs(1061)) xor (layer2_outputs(378));
    outputs(3634) <= not(layer2_outputs(304));
    outputs(3635) <= not((layer2_outputs(284)) or (layer2_outputs(2897)));
    outputs(3636) <= (layer2_outputs(4748)) and (layer2_outputs(1442));
    outputs(3637) <= not(layer2_outputs(4679));
    outputs(3638) <= layer2_outputs(1905);
    outputs(3639) <= layer2_outputs(1921);
    outputs(3640) <= layer2_outputs(2904);
    outputs(3641) <= (layer2_outputs(2531)) and (layer2_outputs(2100));
    outputs(3642) <= not(layer2_outputs(1657)) or (layer2_outputs(4668));
    outputs(3643) <= not(layer2_outputs(1109));
    outputs(3644) <= layer2_outputs(765);
    outputs(3645) <= not(layer2_outputs(2589));
    outputs(3646) <= layer2_outputs(3386);
    outputs(3647) <= layer2_outputs(1782);
    outputs(3648) <= layer2_outputs(3846);
    outputs(3649) <= not(layer2_outputs(1748));
    outputs(3650) <= not(layer2_outputs(4496));
    outputs(3651) <= (layer2_outputs(4765)) and not (layer2_outputs(1739));
    outputs(3652) <= not(layer2_outputs(4133));
    outputs(3653) <= not(layer2_outputs(3681));
    outputs(3654) <= layer2_outputs(1088);
    outputs(3655) <= (layer2_outputs(4631)) xor (layer2_outputs(385));
    outputs(3656) <= not(layer2_outputs(4973));
    outputs(3657) <= layer2_outputs(2196);
    outputs(3658) <= layer2_outputs(564);
    outputs(3659) <= not((layer2_outputs(4713)) and (layer2_outputs(4807)));
    outputs(3660) <= (layer2_outputs(4445)) and not (layer2_outputs(3673));
    outputs(3661) <= not(layer2_outputs(287));
    outputs(3662) <= (layer2_outputs(1114)) and not (layer2_outputs(4954));
    outputs(3663) <= (layer2_outputs(1978)) and not (layer2_outputs(1484));
    outputs(3664) <= not(layer2_outputs(902));
    outputs(3665) <= not((layer2_outputs(3879)) or (layer2_outputs(3494)));
    outputs(3666) <= not(layer2_outputs(1867));
    outputs(3667) <= layer2_outputs(4761);
    outputs(3668) <= layer2_outputs(1445);
    outputs(3669) <= not(layer2_outputs(666));
    outputs(3670) <= (layer2_outputs(3917)) xor (layer2_outputs(3711));
    outputs(3671) <= not((layer2_outputs(3228)) or (layer2_outputs(1103)));
    outputs(3672) <= layer2_outputs(151);
    outputs(3673) <= layer2_outputs(2448);
    outputs(3674) <= not(layer2_outputs(2845));
    outputs(3675) <= not((layer2_outputs(1815)) xor (layer2_outputs(582)));
    outputs(3676) <= (layer2_outputs(4397)) and not (layer2_outputs(432));
    outputs(3677) <= not(layer2_outputs(1959));
    outputs(3678) <= not(layer2_outputs(4228));
    outputs(3679) <= not(layer2_outputs(20));
    outputs(3680) <= not(layer2_outputs(4504));
    outputs(3681) <= not(layer2_outputs(1244));
    outputs(3682) <= not(layer2_outputs(987));
    outputs(3683) <= not(layer2_outputs(1925));
    outputs(3684) <= not((layer2_outputs(2636)) or (layer2_outputs(2980)));
    outputs(3685) <= layer2_outputs(2905);
    outputs(3686) <= layer2_outputs(3671);
    outputs(3687) <= (layer2_outputs(3998)) and not (layer2_outputs(95));
    outputs(3688) <= not(layer2_outputs(3473)) or (layer2_outputs(1942));
    outputs(3689) <= layer2_outputs(4809);
    outputs(3690) <= (layer2_outputs(1499)) and (layer2_outputs(3949));
    outputs(3691) <= layer2_outputs(4810);
    outputs(3692) <= not(layer2_outputs(3));
    outputs(3693) <= not(layer2_outputs(174));
    outputs(3694) <= (layer2_outputs(411)) and (layer2_outputs(3589));
    outputs(3695) <= layer2_outputs(3751);
    outputs(3696) <= not(layer2_outputs(2370));
    outputs(3697) <= not(layer2_outputs(3108));
    outputs(3698) <= (layer2_outputs(621)) and (layer2_outputs(5038));
    outputs(3699) <= not((layer2_outputs(3071)) xor (layer2_outputs(2587)));
    outputs(3700) <= layer2_outputs(4793);
    outputs(3701) <= layer2_outputs(4396);
    outputs(3702) <= not((layer2_outputs(4164)) xor (layer2_outputs(1938)));
    outputs(3703) <= not((layer2_outputs(697)) and (layer2_outputs(4612)));
    outputs(3704) <= layer2_outputs(827);
    outputs(3705) <= layer2_outputs(957);
    outputs(3706) <= not(layer2_outputs(1630));
    outputs(3707) <= layer2_outputs(1640);
    outputs(3708) <= layer2_outputs(1749);
    outputs(3709) <= not(layer2_outputs(715));
    outputs(3710) <= (layer2_outputs(2641)) and not (layer2_outputs(4855));
    outputs(3711) <= not(layer2_outputs(1996));
    outputs(3712) <= not(layer2_outputs(242));
    outputs(3713) <= not(layer2_outputs(4223));
    outputs(3714) <= not(layer2_outputs(2827));
    outputs(3715) <= not(layer2_outputs(610));
    outputs(3716) <= not(layer2_outputs(1558));
    outputs(3717) <= not(layer2_outputs(4599));
    outputs(3718) <= (layer2_outputs(4082)) and not (layer2_outputs(4678));
    outputs(3719) <= layer2_outputs(2630);
    outputs(3720) <= (layer2_outputs(3691)) and (layer2_outputs(420));
    outputs(3721) <= layer2_outputs(1647);
    outputs(3722) <= not(layer2_outputs(3627));
    outputs(3723) <= not(layer2_outputs(4324));
    outputs(3724) <= layer2_outputs(643);
    outputs(3725) <= (layer2_outputs(2896)) and not (layer2_outputs(1965));
    outputs(3726) <= not((layer2_outputs(4897)) xor (layer2_outputs(2766)));
    outputs(3727) <= layer2_outputs(1477);
    outputs(3728) <= not(layer2_outputs(2870));
    outputs(3729) <= layer2_outputs(1451);
    outputs(3730) <= not(layer2_outputs(1382));
    outputs(3731) <= layer2_outputs(159);
    outputs(3732) <= (layer2_outputs(4538)) or (layer2_outputs(3587));
    outputs(3733) <= layer2_outputs(4920);
    outputs(3734) <= (layer2_outputs(3504)) xor (layer2_outputs(3375));
    outputs(3735) <= not(layer2_outputs(4277));
    outputs(3736) <= (layer2_outputs(3238)) xor (layer2_outputs(4789));
    outputs(3737) <= (layer2_outputs(4598)) and (layer2_outputs(3511));
    outputs(3738) <= (layer2_outputs(2700)) and not (layer2_outputs(1723));
    outputs(3739) <= (layer2_outputs(231)) and not (layer2_outputs(2652));
    outputs(3740) <= (layer2_outputs(4893)) and not (layer2_outputs(3717));
    outputs(3741) <= not(layer2_outputs(2646));
    outputs(3742) <= not(layer2_outputs(2928));
    outputs(3743) <= (layer2_outputs(2437)) or (layer2_outputs(4721));
    outputs(3744) <= layer2_outputs(2596);
    outputs(3745) <= layer2_outputs(4800);
    outputs(3746) <= (layer2_outputs(3252)) and not (layer2_outputs(1892));
    outputs(3747) <= layer2_outputs(4935);
    outputs(3748) <= not(layer2_outputs(4274));
    outputs(3749) <= layer2_outputs(1270);
    outputs(3750) <= layer2_outputs(4706);
    outputs(3751) <= (layer2_outputs(3047)) and not (layer2_outputs(4844));
    outputs(3752) <= (layer2_outputs(3502)) and not (layer2_outputs(2297));
    outputs(3753) <= layer2_outputs(2697);
    outputs(3754) <= (layer2_outputs(1036)) xor (layer2_outputs(416));
    outputs(3755) <= not(layer2_outputs(1526));
    outputs(3756) <= not((layer2_outputs(2053)) or (layer2_outputs(3682)));
    outputs(3757) <= not(layer2_outputs(4625));
    outputs(3758) <= layer2_outputs(4059);
    outputs(3759) <= not(layer2_outputs(338));
    outputs(3760) <= not(layer2_outputs(4420)) or (layer2_outputs(2736));
    outputs(3761) <= not(layer2_outputs(4111)) or (layer2_outputs(205));
    outputs(3762) <= not(layer2_outputs(1487));
    outputs(3763) <= not(layer2_outputs(516));
    outputs(3764) <= (layer2_outputs(3934)) and not (layer2_outputs(2038));
    outputs(3765) <= not(layer2_outputs(4323));
    outputs(3766) <= not(layer2_outputs(2597));
    outputs(3767) <= not(layer2_outputs(2078));
    outputs(3768) <= (layer2_outputs(2639)) or (layer2_outputs(2878));
    outputs(3769) <= layer2_outputs(2659);
    outputs(3770) <= not(layer2_outputs(1274));
    outputs(3771) <= (layer2_outputs(4924)) and not (layer2_outputs(2809));
    outputs(3772) <= layer2_outputs(4574);
    outputs(3773) <= layer2_outputs(3835);
    outputs(3774) <= (layer2_outputs(4974)) and not (layer2_outputs(4309));
    outputs(3775) <= (layer2_outputs(2818)) xor (layer2_outputs(1430));
    outputs(3776) <= (layer2_outputs(3189)) and not (layer2_outputs(2027));
    outputs(3777) <= layer2_outputs(108);
    outputs(3778) <= not(layer2_outputs(3533));
    outputs(3779) <= layer2_outputs(2413);
    outputs(3780) <= layer2_outputs(4399);
    outputs(3781) <= layer2_outputs(1163);
    outputs(3782) <= layer2_outputs(3241);
    outputs(3783) <= layer2_outputs(1557);
    outputs(3784) <= not((layer2_outputs(5092)) xor (layer2_outputs(4759)));
    outputs(3785) <= layer2_outputs(3355);
    outputs(3786) <= not(layer2_outputs(3493));
    outputs(3787) <= (layer2_outputs(3819)) and not (layer2_outputs(3820));
    outputs(3788) <= layer2_outputs(1726);
    outputs(3789) <= not(layer2_outputs(341));
    outputs(3790) <= (layer2_outputs(3899)) and not (layer2_outputs(2782));
    outputs(3791) <= layer2_outputs(2507);
    outputs(3792) <= not((layer2_outputs(4179)) or (layer2_outputs(4153)));
    outputs(3793) <= not(layer2_outputs(3082));
    outputs(3794) <= not(layer2_outputs(2251));
    outputs(3795) <= layer2_outputs(1102);
    outputs(3796) <= layer2_outputs(5022);
    outputs(3797) <= layer2_outputs(1640);
    outputs(3798) <= not(layer2_outputs(4597));
    outputs(3799) <= layer2_outputs(1872);
    outputs(3800) <= not(layer2_outputs(358));
    outputs(3801) <= not((layer2_outputs(1899)) or (layer2_outputs(3633)));
    outputs(3802) <= layer2_outputs(3956);
    outputs(3803) <= (layer2_outputs(499)) xor (layer2_outputs(1979));
    outputs(3804) <= not(layer2_outputs(81));
    outputs(3805) <= (layer2_outputs(1252)) and (layer2_outputs(1335));
    outputs(3806) <= layer2_outputs(2612);
    outputs(3807) <= not(layer2_outputs(1886));
    outputs(3808) <= layer2_outputs(4988);
    outputs(3809) <= layer2_outputs(2197);
    outputs(3810) <= layer2_outputs(2548);
    outputs(3811) <= not(layer2_outputs(4277));
    outputs(3812) <= not((layer2_outputs(3774)) xor (layer2_outputs(4980)));
    outputs(3813) <= not((layer2_outputs(547)) and (layer2_outputs(1298)));
    outputs(3814) <= not((layer2_outputs(4357)) xor (layer2_outputs(219)));
    outputs(3815) <= not(layer2_outputs(4415));
    outputs(3816) <= layer2_outputs(3346);
    outputs(3817) <= not(layer2_outputs(4673)) or (layer2_outputs(739));
    outputs(3818) <= not(layer2_outputs(2144));
    outputs(3819) <= (layer2_outputs(899)) and not (layer2_outputs(4272));
    outputs(3820) <= (layer2_outputs(4440)) xor (layer2_outputs(2537));
    outputs(3821) <= not(layer2_outputs(3495));
    outputs(3822) <= layer2_outputs(4392);
    outputs(3823) <= (layer2_outputs(1241)) and not (layer2_outputs(2327));
    outputs(3824) <= (layer2_outputs(523)) xor (layer2_outputs(682));
    outputs(3825) <= layer2_outputs(2128);
    outputs(3826) <= not(layer2_outputs(4606));
    outputs(3827) <= not((layer2_outputs(4468)) and (layer2_outputs(4207)));
    outputs(3828) <= layer2_outputs(2786);
    outputs(3829) <= not((layer2_outputs(3749)) and (layer2_outputs(4848)));
    outputs(3830) <= (layer2_outputs(479)) xor (layer2_outputs(3619));
    outputs(3831) <= (layer2_outputs(1070)) or (layer2_outputs(3462));
    outputs(3832) <= (layer2_outputs(3910)) and not (layer2_outputs(1820));
    outputs(3833) <= not(layer2_outputs(630)) or (layer2_outputs(5073));
    outputs(3834) <= not(layer2_outputs(3305)) or (layer2_outputs(3170));
    outputs(3835) <= not((layer2_outputs(1912)) xor (layer2_outputs(1354)));
    outputs(3836) <= not(layer2_outputs(1602));
    outputs(3837) <= not(layer2_outputs(4115));
    outputs(3838) <= not(layer2_outputs(3078));
    outputs(3839) <= not(layer2_outputs(2293)) or (layer2_outputs(1034));
    outputs(3840) <= not(layer2_outputs(279));
    outputs(3841) <= not(layer2_outputs(1693));
    outputs(3842) <= layer2_outputs(3382);
    outputs(3843) <= not(layer2_outputs(3134));
    outputs(3844) <= (layer2_outputs(3882)) and not (layer2_outputs(3012));
    outputs(3845) <= not(layer2_outputs(3233));
    outputs(3846) <= not(layer2_outputs(148));
    outputs(3847) <= not(layer2_outputs(1018)) or (layer2_outputs(153));
    outputs(3848) <= not(layer2_outputs(2088));
    outputs(3849) <= not(layer2_outputs(3895));
    outputs(3850) <= (layer2_outputs(2194)) xor (layer2_outputs(3174));
    outputs(3851) <= layer2_outputs(2219);
    outputs(3852) <= (layer2_outputs(2554)) and (layer2_outputs(1074));
    outputs(3853) <= layer2_outputs(2381);
    outputs(3854) <= layer2_outputs(140);
    outputs(3855) <= (layer2_outputs(2347)) xor (layer2_outputs(945));
    outputs(3856) <= layer2_outputs(1740);
    outputs(3857) <= (layer2_outputs(1945)) and not (layer2_outputs(4318));
    outputs(3858) <= (layer2_outputs(4429)) and (layer2_outputs(4677));
    outputs(3859) <= layer2_outputs(601);
    outputs(3860) <= layer2_outputs(1469);
    outputs(3861) <= not((layer2_outputs(312)) or (layer2_outputs(2469)));
    outputs(3862) <= not(layer2_outputs(450));
    outputs(3863) <= (layer2_outputs(1062)) and (layer2_outputs(2193));
    outputs(3864) <= not(layer2_outputs(17));
    outputs(3865) <= not(layer2_outputs(4018));
    outputs(3866) <= layer2_outputs(3183);
    outputs(3867) <= not(layer2_outputs(552));
    outputs(3868) <= not((layer2_outputs(4835)) xor (layer2_outputs(991)));
    outputs(3869) <= not(layer2_outputs(184));
    outputs(3870) <= not((layer2_outputs(1235)) or (layer2_outputs(3234)));
    outputs(3871) <= layer2_outputs(141);
    outputs(3872) <= (layer2_outputs(3287)) and (layer2_outputs(880));
    outputs(3873) <= not(layer2_outputs(5092));
    outputs(3874) <= (layer2_outputs(3197)) xor (layer2_outputs(1572));
    outputs(3875) <= not(layer2_outputs(2055));
    outputs(3876) <= not(layer2_outputs(948));
    outputs(3877) <= layer2_outputs(2242);
    outputs(3878) <= layer2_outputs(2493);
    outputs(3879) <= not((layer2_outputs(2261)) or (layer2_outputs(1122)));
    outputs(3880) <= not((layer2_outputs(3261)) or (layer2_outputs(2558)));
    outputs(3881) <= (layer2_outputs(2539)) and not (layer2_outputs(4564));
    outputs(3882) <= layer2_outputs(1652);
    outputs(3883) <= layer2_outputs(885);
    outputs(3884) <= not(layer2_outputs(4509));
    outputs(3885) <= not(layer2_outputs(4797));
    outputs(3886) <= not(layer2_outputs(1306));
    outputs(3887) <= (layer2_outputs(1525)) and (layer2_outputs(1118));
    outputs(3888) <= not((layer2_outputs(873)) or (layer2_outputs(4757)));
    outputs(3889) <= not(layer2_outputs(309));
    outputs(3890) <= not(layer2_outputs(830));
    outputs(3891) <= not(layer2_outputs(3864));
    outputs(3892) <= (layer2_outputs(3833)) or (layer2_outputs(2615));
    outputs(3893) <= not(layer2_outputs(3776));
    outputs(3894) <= layer2_outputs(4003);
    outputs(3895) <= layer2_outputs(2592);
    outputs(3896) <= not(layer2_outputs(2731));
    outputs(3897) <= not((layer2_outputs(3685)) xor (layer2_outputs(4427)));
    outputs(3898) <= layer2_outputs(1586);
    outputs(3899) <= (layer2_outputs(2495)) and not (layer2_outputs(1909));
    outputs(3900) <= not(layer2_outputs(3268));
    outputs(3901) <= layer2_outputs(4795);
    outputs(3902) <= (layer2_outputs(1408)) xor (layer2_outputs(2066));
    outputs(3903) <= not(layer2_outputs(1758));
    outputs(3904) <= (layer2_outputs(2005)) and (layer2_outputs(4331));
    outputs(3905) <= layer2_outputs(905);
    outputs(3906) <= layer2_outputs(764);
    outputs(3907) <= layer2_outputs(2851);
    outputs(3908) <= layer2_outputs(4841);
    outputs(3909) <= layer2_outputs(3731);
    outputs(3910) <= not(layer2_outputs(4510));
    outputs(3911) <= not((layer2_outputs(3203)) or (layer2_outputs(5041)));
    outputs(3912) <= not((layer2_outputs(5114)) or (layer2_outputs(2734)));
    outputs(3913) <= layer2_outputs(2424);
    outputs(3914) <= not(layer2_outputs(857)) or (layer2_outputs(2655));
    outputs(3915) <= layer2_outputs(4704);
    outputs(3916) <= not(layer2_outputs(613));
    outputs(3917) <= (layer2_outputs(1535)) and not (layer2_outputs(5059));
    outputs(3918) <= (layer2_outputs(770)) and (layer2_outputs(2771));
    outputs(3919) <= (layer2_outputs(2488)) and (layer2_outputs(1508));
    outputs(3920) <= not((layer2_outputs(12)) or (layer2_outputs(3371)));
    outputs(3921) <= layer2_outputs(4014);
    outputs(3922) <= layer2_outputs(4304);
    outputs(3923) <= (layer2_outputs(5072)) and (layer2_outputs(734));
    outputs(3924) <= not(layer2_outputs(2758)) or (layer2_outputs(2426));
    outputs(3925) <= (layer2_outputs(2559)) and not (layer2_outputs(1979));
    outputs(3926) <= layer2_outputs(993);
    outputs(3927) <= (layer2_outputs(406)) and not (layer2_outputs(416));
    outputs(3928) <= not(layer2_outputs(4419));
    outputs(3929) <= not(layer2_outputs(900));
    outputs(3930) <= layer2_outputs(4454);
    outputs(3931) <= not(layer2_outputs(3760));
    outputs(3932) <= (layer2_outputs(5039)) and (layer2_outputs(726));
    outputs(3933) <= not(layer2_outputs(3467)) or (layer2_outputs(4548));
    outputs(3934) <= layer2_outputs(1613);
    outputs(3935) <= not(layer2_outputs(1137));
    outputs(3936) <= not((layer2_outputs(2336)) xor (layer2_outputs(1361)));
    outputs(3937) <= layer2_outputs(3484);
    outputs(3938) <= layer2_outputs(2834);
    outputs(3939) <= not((layer2_outputs(5057)) xor (layer2_outputs(1748)));
    outputs(3940) <= not(layer2_outputs(73));
    outputs(3941) <= layer2_outputs(1140);
    outputs(3942) <= not(layer2_outputs(2677));
    outputs(3943) <= (layer2_outputs(4040)) xor (layer2_outputs(1079));
    outputs(3944) <= layer2_outputs(998);
    outputs(3945) <= (layer2_outputs(3337)) and not (layer2_outputs(809));
    outputs(3946) <= not(layer2_outputs(3310));
    outputs(3947) <= not((layer2_outputs(1151)) or (layer2_outputs(915)));
    outputs(3948) <= (layer2_outputs(4320)) and not (layer2_outputs(3109));
    outputs(3949) <= layer2_outputs(4425);
    outputs(3950) <= layer2_outputs(834);
    outputs(3951) <= not(layer2_outputs(3403)) or (layer2_outputs(762));
    outputs(3952) <= (layer2_outputs(3340)) and not (layer2_outputs(3720));
    outputs(3953) <= layer2_outputs(4515);
    outputs(3954) <= layer2_outputs(1683);
    outputs(3955) <= layer2_outputs(2218);
    outputs(3956) <= not(layer2_outputs(2871));
    outputs(3957) <= (layer2_outputs(3383)) and not (layer2_outputs(3992));
    outputs(3958) <= not(layer2_outputs(3442));
    outputs(3959) <= layer2_outputs(2508);
    outputs(3960) <= (layer2_outputs(3972)) xor (layer2_outputs(4077));
    outputs(3961) <= not(layer2_outputs(4878));
    outputs(3962) <= not(layer2_outputs(531)) or (layer2_outputs(4555));
    outputs(3963) <= (layer2_outputs(5054)) xor (layer2_outputs(2344));
    outputs(3964) <= not(layer2_outputs(1415));
    outputs(3965) <= not(layer2_outputs(4970)) or (layer2_outputs(1194));
    outputs(3966) <= (layer2_outputs(294)) and not (layer2_outputs(2569));
    outputs(3967) <= layer2_outputs(4741);
    outputs(3968) <= layer2_outputs(3447);
    outputs(3969) <= (layer2_outputs(1566)) and (layer2_outputs(3865));
    outputs(3970) <= (layer2_outputs(4948)) and (layer2_outputs(69));
    outputs(3971) <= layer2_outputs(4942);
    outputs(3972) <= (layer2_outputs(2348)) or (layer2_outputs(1592));
    outputs(3973) <= not((layer2_outputs(455)) xor (layer2_outputs(530)));
    outputs(3974) <= not(layer2_outputs(4271));
    outputs(3975) <= (layer2_outputs(2540)) xor (layer2_outputs(267));
    outputs(3976) <= not(layer2_outputs(2695));
    outputs(3977) <= (layer2_outputs(1621)) xor (layer2_outputs(3563));
    outputs(3978) <= not(layer2_outputs(2938));
    outputs(3979) <= (layer2_outputs(4615)) and (layer2_outputs(4708));
    outputs(3980) <= not((layer2_outputs(642)) xor (layer2_outputs(4692)));
    outputs(3981) <= layer2_outputs(1789);
    outputs(3982) <= layer2_outputs(1075);
    outputs(3983) <= not(layer2_outputs(3347));
    outputs(3984) <= layer2_outputs(1348);
    outputs(3985) <= not(layer2_outputs(1296));
    outputs(3986) <= layer2_outputs(2812);
    outputs(3987) <= (layer2_outputs(2210)) and (layer2_outputs(3960));
    outputs(3988) <= (layer2_outputs(2300)) and not (layer2_outputs(3843));
    outputs(3989) <= not(layer2_outputs(2491));
    outputs(3990) <= not(layer2_outputs(825));
    outputs(3991) <= not(layer2_outputs(4486));
    outputs(3992) <= layer2_outputs(308);
    outputs(3993) <= (layer2_outputs(2014)) and not (layer2_outputs(1705));
    outputs(3994) <= not(layer2_outputs(4736));
    outputs(3995) <= not(layer2_outputs(4064)) or (layer2_outputs(1288));
    outputs(3996) <= layer2_outputs(2655);
    outputs(3997) <= (layer2_outputs(2990)) xor (layer2_outputs(3617));
    outputs(3998) <= (layer2_outputs(3842)) xor (layer2_outputs(4893));
    outputs(3999) <= (layer2_outputs(3451)) and (layer2_outputs(4926));
    outputs(4000) <= not(layer2_outputs(370));
    outputs(4001) <= not(layer2_outputs(85));
    outputs(4002) <= layer2_outputs(3470);
    outputs(4003) <= (layer2_outputs(247)) and not (layer2_outputs(1725));
    outputs(4004) <= not(layer2_outputs(1574));
    outputs(4005) <= not(layer2_outputs(665));
    outputs(4006) <= (layer2_outputs(1342)) and not (layer2_outputs(1853));
    outputs(4007) <= (layer2_outputs(3881)) xor (layer2_outputs(2151));
    outputs(4008) <= layer2_outputs(675);
    outputs(4009) <= (layer2_outputs(4407)) and not (layer2_outputs(2420));
    outputs(4010) <= (layer2_outputs(2433)) and not (layer2_outputs(3686));
    outputs(4011) <= not((layer2_outputs(4848)) and (layer2_outputs(80)));
    outputs(4012) <= not(layer2_outputs(3399));
    outputs(4013) <= layer2_outputs(2200);
    outputs(4014) <= (layer2_outputs(2089)) and not (layer2_outputs(3186));
    outputs(4015) <= (layer2_outputs(1342)) and not (layer2_outputs(2029));
    outputs(4016) <= not(layer2_outputs(4495));
    outputs(4017) <= (layer2_outputs(241)) and (layer2_outputs(2130));
    outputs(4018) <= not(layer2_outputs(1101));
    outputs(4019) <= not(layer2_outputs(4878));
    outputs(4020) <= layer2_outputs(2019);
    outputs(4021) <= not((layer2_outputs(474)) xor (layer2_outputs(1601)));
    outputs(4022) <= (layer2_outputs(4554)) or (layer2_outputs(4851));
    outputs(4023) <= layer2_outputs(46);
    outputs(4024) <= not((layer2_outputs(1256)) or (layer2_outputs(3209)));
    outputs(4025) <= not((layer2_outputs(935)) xor (layer2_outputs(4691)));
    outputs(4026) <= not(layer2_outputs(4356));
    outputs(4027) <= layer2_outputs(953);
    outputs(4028) <= layer2_outputs(3080);
    outputs(4029) <= not(layer2_outputs(112));
    outputs(4030) <= layer2_outputs(3286);
    outputs(4031) <= (layer2_outputs(3215)) and not (layer2_outputs(1697));
    outputs(4032) <= not((layer2_outputs(4550)) xor (layer2_outputs(4834)));
    outputs(4033) <= not(layer2_outputs(1599));
    outputs(4034) <= (layer2_outputs(3745)) and (layer2_outputs(3732));
    outputs(4035) <= not(layer2_outputs(4266));
    outputs(4036) <= not(layer2_outputs(221));
    outputs(4037) <= not(layer2_outputs(3576));
    outputs(4038) <= layer2_outputs(2962);
    outputs(4039) <= not(layer2_outputs(491));
    outputs(4040) <= not(layer2_outputs(4061)) or (layer2_outputs(12));
    outputs(4041) <= not((layer2_outputs(101)) xor (layer2_outputs(264)));
    outputs(4042) <= layer2_outputs(662);
    outputs(4043) <= (layer2_outputs(1661)) and (layer2_outputs(4162));
    outputs(4044) <= layer2_outputs(48);
    outputs(4045) <= not(layer2_outputs(2815));
    outputs(4046) <= layer2_outputs(1678);
    outputs(4047) <= (layer2_outputs(2415)) and not (layer2_outputs(890));
    outputs(4048) <= not((layer2_outputs(4779)) xor (layer2_outputs(3292)));
    outputs(4049) <= not(layer2_outputs(1688));
    outputs(4050) <= layer2_outputs(2262);
    outputs(4051) <= layer2_outputs(4321);
    outputs(4052) <= not(layer2_outputs(1032));
    outputs(4053) <= layer2_outputs(2855);
    outputs(4054) <= layer2_outputs(476);
    outputs(4055) <= (layer2_outputs(3076)) and not (layer2_outputs(4233));
    outputs(4056) <= not(layer2_outputs(4865)) or (layer2_outputs(3263));
    outputs(4057) <= layer2_outputs(13);
    outputs(4058) <= layer2_outputs(3044);
    outputs(4059) <= not(layer2_outputs(2049));
    outputs(4060) <= not((layer2_outputs(2572)) or (layer2_outputs(34)));
    outputs(4061) <= (layer2_outputs(2429)) and (layer2_outputs(2415));
    outputs(4062) <= not((layer2_outputs(1115)) or (layer2_outputs(4986)));
    outputs(4063) <= layer2_outputs(971);
    outputs(4064) <= not(layer2_outputs(1626));
    outputs(4065) <= not((layer2_outputs(1119)) and (layer2_outputs(3565)));
    outputs(4066) <= not(layer2_outputs(370));
    outputs(4067) <= not((layer2_outputs(798)) xor (layer2_outputs(339)));
    outputs(4068) <= layer2_outputs(4771);
    outputs(4069) <= not((layer2_outputs(4907)) or (layer2_outputs(1546)));
    outputs(4070) <= layer2_outputs(3949);
    outputs(4071) <= layer2_outputs(4201);
    outputs(4072) <= layer2_outputs(4936);
    outputs(4073) <= (layer2_outputs(3581)) and not (layer2_outputs(1244));
    outputs(4074) <= layer2_outputs(2174);
    outputs(4075) <= layer2_outputs(3558);
    outputs(4076) <= not(layer2_outputs(3079));
    outputs(4077) <= layer2_outputs(3179);
    outputs(4078) <= not((layer2_outputs(2253)) xor (layer2_outputs(4256)));
    outputs(4079) <= (layer2_outputs(2382)) and (layer2_outputs(785));
    outputs(4080) <= (layer2_outputs(1215)) and (layer2_outputs(2724));
    outputs(4081) <= not(layer2_outputs(3017));
    outputs(4082) <= (layer2_outputs(2959)) and (layer2_outputs(901));
    outputs(4083) <= layer2_outputs(1589);
    outputs(4084) <= not(layer2_outputs(3992));
    outputs(4085) <= not(layer2_outputs(2467));
    outputs(4086) <= not(layer2_outputs(3078));
    outputs(4087) <= not(layer2_outputs(4129)) or (layer2_outputs(4979));
    outputs(4088) <= (layer2_outputs(4552)) and not (layer2_outputs(2239));
    outputs(4089) <= layer2_outputs(1966);
    outputs(4090) <= not(layer2_outputs(3926));
    outputs(4091) <= layer2_outputs(2277);
    outputs(4092) <= not(layer2_outputs(239)) or (layer2_outputs(4918));
    outputs(4093) <= (layer2_outputs(4167)) and not (layer2_outputs(65));
    outputs(4094) <= not(layer2_outputs(1763));
    outputs(4095) <= (layer2_outputs(3810)) and not (layer2_outputs(2164));
    outputs(4096) <= not((layer2_outputs(4692)) xor (layer2_outputs(345)));
    outputs(4097) <= not(layer2_outputs(1419));
    outputs(4098) <= layer2_outputs(2340);
    outputs(4099) <= (layer2_outputs(1384)) or (layer2_outputs(5099));
    outputs(4100) <= not(layer2_outputs(3959));
    outputs(4101) <= not(layer2_outputs(1214));
    outputs(4102) <= layer2_outputs(4920);
    outputs(4103) <= not(layer2_outputs(4230));
    outputs(4104) <= layer2_outputs(4623);
    outputs(4105) <= not(layer2_outputs(965));
    outputs(4106) <= (layer2_outputs(3260)) xor (layer2_outputs(3302));
    outputs(4107) <= not(layer2_outputs(2336));
    outputs(4108) <= (layer2_outputs(1756)) xor (layer2_outputs(5001));
    outputs(4109) <= not(layer2_outputs(3708));
    outputs(4110) <= layer2_outputs(129);
    outputs(4111) <= (layer2_outputs(3454)) or (layer2_outputs(3859));
    outputs(4112) <= layer2_outputs(2958);
    outputs(4113) <= (layer2_outputs(4090)) and (layer2_outputs(4513));
    outputs(4114) <= layer2_outputs(1237);
    outputs(4115) <= not(layer2_outputs(3556));
    outputs(4116) <= layer2_outputs(3133);
    outputs(4117) <= layer2_outputs(1257);
    outputs(4118) <= not(layer2_outputs(4567));
    outputs(4119) <= layer2_outputs(3816);
    outputs(4120) <= not((layer2_outputs(60)) and (layer2_outputs(2123)));
    outputs(4121) <= not(layer2_outputs(1397));
    outputs(4122) <= not(layer2_outputs(1535));
    outputs(4123) <= (layer2_outputs(1989)) or (layer2_outputs(2325));
    outputs(4124) <= not((layer2_outputs(3596)) xor (layer2_outputs(2669)));
    outputs(4125) <= layer2_outputs(2652);
    outputs(4126) <= not((layer2_outputs(1834)) or (layer2_outputs(1340)));
    outputs(4127) <= (layer2_outputs(2105)) or (layer2_outputs(897));
    outputs(4128) <= (layer2_outputs(774)) and not (layer2_outputs(3585));
    outputs(4129) <= not(layer2_outputs(2439));
    outputs(4130) <= (layer2_outputs(526)) and (layer2_outputs(598));
    outputs(4131) <= layer2_outputs(3027);
    outputs(4132) <= layer2_outputs(4670);
    outputs(4133) <= not(layer2_outputs(7));
    outputs(4134) <= not(layer2_outputs(3161));
    outputs(4135) <= not((layer2_outputs(3386)) xor (layer2_outputs(1929)));
    outputs(4136) <= (layer2_outputs(4896)) and not (layer2_outputs(3795));
    outputs(4137) <= layer2_outputs(102);
    outputs(4138) <= layer2_outputs(4785);
    outputs(4139) <= layer2_outputs(2076);
    outputs(4140) <= not(layer2_outputs(143));
    outputs(4141) <= not((layer2_outputs(451)) xor (layer2_outputs(311)));
    outputs(4142) <= layer2_outputs(1310);
    outputs(4143) <= not(layer2_outputs(692));
    outputs(4144) <= layer2_outputs(2335);
    outputs(4145) <= layer2_outputs(4205);
    outputs(4146) <= not((layer2_outputs(1197)) xor (layer2_outputs(997)));
    outputs(4147) <= not(layer2_outputs(1719));
    outputs(4148) <= not(layer2_outputs(1358));
    outputs(4149) <= not(layer2_outputs(3891));
    outputs(4150) <= not(layer2_outputs(4129));
    outputs(4151) <= not(layer2_outputs(2580));
    outputs(4152) <= (layer2_outputs(3939)) or (layer2_outputs(24));
    outputs(4153) <= not((layer2_outputs(5014)) xor (layer2_outputs(3559)));
    outputs(4154) <= not((layer2_outputs(3179)) xor (layer2_outputs(1155)));
    outputs(4155) <= not(layer2_outputs(3854));
    outputs(4156) <= layer2_outputs(2941);
    outputs(4157) <= not(layer2_outputs(4079));
    outputs(4158) <= (layer2_outputs(2829)) xor (layer2_outputs(1157));
    outputs(4159) <= layer2_outputs(63);
    outputs(4160) <= not(layer2_outputs(2795));
    outputs(4161) <= not(layer2_outputs(3792));
    outputs(4162) <= not(layer2_outputs(1612));
    outputs(4163) <= (layer2_outputs(2383)) and not (layer2_outputs(1370));
    outputs(4164) <= layer2_outputs(2813);
    outputs(4165) <= not(layer2_outputs(4633));
    outputs(4166) <= (layer2_outputs(2498)) and (layer2_outputs(3397));
    outputs(4167) <= (layer2_outputs(2638)) and not (layer2_outputs(937));
    outputs(4168) <= not(layer2_outputs(981));
    outputs(4169) <= (layer2_outputs(1702)) xor (layer2_outputs(290));
    outputs(4170) <= not(layer2_outputs(3279));
    outputs(4171) <= not(layer2_outputs(168));
    outputs(4172) <= not((layer2_outputs(1846)) or (layer2_outputs(4695)));
    outputs(4173) <= not(layer2_outputs(3509)) or (layer2_outputs(2798));
    outputs(4174) <= layer2_outputs(1425);
    outputs(4175) <= (layer2_outputs(3522)) or (layer2_outputs(5055));
    outputs(4176) <= not(layer2_outputs(4837)) or (layer2_outputs(2735));
    outputs(4177) <= not((layer2_outputs(2148)) xor (layer2_outputs(3623)));
    outputs(4178) <= (layer2_outputs(3065)) xor (layer2_outputs(1765));
    outputs(4179) <= (layer2_outputs(3146)) xor (layer2_outputs(3465));
    outputs(4180) <= (layer2_outputs(1577)) xor (layer2_outputs(1785));
    outputs(4181) <= not(layer2_outputs(3703));
    outputs(4182) <= not(layer2_outputs(3761));
    outputs(4183) <= not(layer2_outputs(2746)) or (layer2_outputs(3904));
    outputs(4184) <= not((layer2_outputs(3507)) xor (layer2_outputs(3286)));
    outputs(4185) <= not(layer2_outputs(2826));
    outputs(4186) <= (layer2_outputs(2293)) and not (layer2_outputs(42));
    outputs(4187) <= layer2_outputs(4106);
    outputs(4188) <= not(layer2_outputs(2942)) or (layer2_outputs(2638));
    outputs(4189) <= not((layer2_outputs(1413)) xor (layer2_outputs(4083)));
    outputs(4190) <= not((layer2_outputs(72)) xor (layer2_outputs(597)));
    outputs(4191) <= not(layer2_outputs(1446));
    outputs(4192) <= (layer2_outputs(2562)) xor (layer2_outputs(2782));
    outputs(4193) <= layer2_outputs(911);
    outputs(4194) <= not(layer2_outputs(2189));
    outputs(4195) <= layer2_outputs(2402);
    outputs(4196) <= not(layer2_outputs(4960)) or (layer2_outputs(2440));
    outputs(4197) <= layer2_outputs(2206);
    outputs(4198) <= layer2_outputs(4955);
    outputs(4199) <= not((layer2_outputs(1414)) or (layer2_outputs(2330)));
    outputs(4200) <= not(layer2_outputs(4430));
    outputs(4201) <= not((layer2_outputs(2085)) xor (layer2_outputs(1262)));
    outputs(4202) <= layer2_outputs(3360);
    outputs(4203) <= (layer2_outputs(1871)) xor (layer2_outputs(1407));
    outputs(4204) <= layer2_outputs(2889);
    outputs(4205) <= layer2_outputs(550);
    outputs(4206) <= layer2_outputs(360);
    outputs(4207) <= not(layer2_outputs(2069));
    outputs(4208) <= not(layer2_outputs(4432));
    outputs(4209) <= layer2_outputs(2773);
    outputs(4210) <= not((layer2_outputs(505)) xor (layer2_outputs(1607)));
    outputs(4211) <= not(layer2_outputs(1144));
    outputs(4212) <= not(layer2_outputs(2082));
    outputs(4213) <= (layer2_outputs(3456)) xor (layer2_outputs(4751));
    outputs(4214) <= not(layer2_outputs(1604));
    outputs(4215) <= (layer2_outputs(1891)) and not (layer2_outputs(953));
    outputs(4216) <= not(layer2_outputs(2935)) or (layer2_outputs(2759));
    outputs(4217) <= not(layer2_outputs(2856));
    outputs(4218) <= (layer2_outputs(3221)) xor (layer2_outputs(108));
    outputs(4219) <= (layer2_outputs(38)) xor (layer2_outputs(1237));
    outputs(4220) <= layer2_outputs(3817);
    outputs(4221) <= not(layer2_outputs(3580));
    outputs(4222) <= layer2_outputs(1575);
    outputs(4223) <= not(layer2_outputs(3797)) or (layer2_outputs(2283));
    outputs(4224) <= layer2_outputs(1305);
    outputs(4225) <= not((layer2_outputs(817)) xor (layer2_outputs(1867)));
    outputs(4226) <= layer2_outputs(1245);
    outputs(4227) <= layer2_outputs(4857);
    outputs(4228) <= not(layer2_outputs(3968));
    outputs(4229) <= not(layer2_outputs(4404)) or (layer2_outputs(1606));
    outputs(4230) <= not(layer2_outputs(2342)) or (layer2_outputs(2278));
    outputs(4231) <= not(layer2_outputs(2620));
    outputs(4232) <= not(layer2_outputs(2888));
    outputs(4233) <= not(layer2_outputs(2568));
    outputs(4234) <= layer2_outputs(3812);
    outputs(4235) <= layer2_outputs(3943);
    outputs(4236) <= not(layer2_outputs(2254));
    outputs(4237) <= (layer2_outputs(3917)) or (layer2_outputs(1857));
    outputs(4238) <= layer2_outputs(761);
    outputs(4239) <= (layer2_outputs(4719)) xor (layer2_outputs(4033));
    outputs(4240) <= not((layer2_outputs(1995)) xor (layer2_outputs(195)));
    outputs(4241) <= not(layer2_outputs(4672));
    outputs(4242) <= not(layer2_outputs(3177)) or (layer2_outputs(1722));
    outputs(4243) <= not((layer2_outputs(2240)) xor (layer2_outputs(856)));
    outputs(4244) <= '1';
    outputs(4245) <= layer2_outputs(2229);
    outputs(4246) <= not((layer2_outputs(2286)) or (layer2_outputs(2059)));
    outputs(4247) <= (layer2_outputs(787)) and (layer2_outputs(1048));
    outputs(4248) <= layer2_outputs(1268);
    outputs(4249) <= not(layer2_outputs(1292));
    outputs(4250) <= not(layer2_outputs(3991));
    outputs(4251) <= not((layer2_outputs(821)) xor (layer2_outputs(4491)));
    outputs(4252) <= not((layer2_outputs(4732)) xor (layer2_outputs(2663)));
    outputs(4253) <= not(layer2_outputs(3913)) or (layer2_outputs(1044));
    outputs(4254) <= not(layer2_outputs(3320));
    outputs(4255) <= not((layer2_outputs(3358)) or (layer2_outputs(3069)));
    outputs(4256) <= not(layer2_outputs(1078));
    outputs(4257) <= not((layer2_outputs(4838)) xor (layer2_outputs(4264)));
    outputs(4258) <= not(layer2_outputs(4810));
    outputs(4259) <= (layer2_outputs(3309)) xor (layer2_outputs(348));
    outputs(4260) <= not(layer2_outputs(727));
    outputs(4261) <= layer2_outputs(4422);
    outputs(4262) <= not(layer2_outputs(1662)) or (layer2_outputs(4170));
    outputs(4263) <= layer2_outputs(943);
    outputs(4264) <= (layer2_outputs(3923)) and not (layer2_outputs(1513));
    outputs(4265) <= (layer2_outputs(4327)) xor (layer2_outputs(1893));
    outputs(4266) <= (layer2_outputs(1301)) and not (layer2_outputs(802));
    outputs(4267) <= layer2_outputs(2229);
    outputs(4268) <= layer2_outputs(1970);
    outputs(4269) <= layer2_outputs(2725);
    outputs(4270) <= not(layer2_outputs(3520));
    outputs(4271) <= not((layer2_outputs(73)) xor (layer2_outputs(2767)));
    outputs(4272) <= not(layer2_outputs(2855));
    outputs(4273) <= layer2_outputs(2964);
    outputs(4274) <= layer2_outputs(363);
    outputs(4275) <= (layer2_outputs(3437)) and not (layer2_outputs(4240));
    outputs(4276) <= not(layer2_outputs(1054));
    outputs(4277) <= (layer2_outputs(3289)) and not (layer2_outputs(3336));
    outputs(4278) <= layer2_outputs(907);
    outputs(4279) <= layer2_outputs(1981);
    outputs(4280) <= not((layer2_outputs(3670)) xor (layer2_outputs(2885)));
    outputs(4281) <= (layer2_outputs(4648)) and (layer2_outputs(2983));
    outputs(4282) <= (layer2_outputs(3488)) xor (layer2_outputs(2305));
    outputs(4283) <= not(layer2_outputs(121));
    outputs(4284) <= not(layer2_outputs(587));
    outputs(4285) <= layer2_outputs(4184);
    outputs(4286) <= layer2_outputs(3094);
    outputs(4287) <= not((layer2_outputs(3069)) xor (layer2_outputs(551)));
    outputs(4288) <= layer2_outputs(4745);
    outputs(4289) <= layer2_outputs(10);
    outputs(4290) <= not(layer2_outputs(477)) or (layer2_outputs(5105));
    outputs(4291) <= (layer2_outputs(2691)) and (layer2_outputs(825));
    outputs(4292) <= layer2_outputs(4062);
    outputs(4293) <= layer2_outputs(5008);
    outputs(4294) <= not((layer2_outputs(4037)) xor (layer2_outputs(2974)));
    outputs(4295) <= not((layer2_outputs(214)) or (layer2_outputs(504)));
    outputs(4296) <= (layer2_outputs(4735)) and not (layer2_outputs(1825));
    outputs(4297) <= (layer2_outputs(3921)) and not (layer2_outputs(3746));
    outputs(4298) <= (layer2_outputs(3322)) and not (layer2_outputs(1276));
    outputs(4299) <= layer2_outputs(4151);
    outputs(4300) <= layer2_outputs(703);
    outputs(4301) <= not(layer2_outputs(289));
    outputs(4302) <= not((layer2_outputs(3565)) and (layer2_outputs(2794)));
    outputs(4303) <= layer2_outputs(4231);
    outputs(4304) <= not(layer2_outputs(3783));
    outputs(4305) <= layer2_outputs(2022);
    outputs(4306) <= not(layer2_outputs(3738));
    outputs(4307) <= not(layer2_outputs(4254));
    outputs(4308) <= layer2_outputs(2332);
    outputs(4309) <= not((layer2_outputs(283)) xor (layer2_outputs(2667)));
    outputs(4310) <= (layer2_outputs(337)) xor (layer2_outputs(1558));
    outputs(4311) <= not((layer2_outputs(3621)) xor (layer2_outputs(1505)));
    outputs(4312) <= layer2_outputs(4463);
    outputs(4313) <= layer2_outputs(3234);
    outputs(4314) <= not((layer2_outputs(5044)) xor (layer2_outputs(4883)));
    outputs(4315) <= layer2_outputs(3889);
    outputs(4316) <= (layer2_outputs(2209)) xor (layer2_outputs(3596));
    outputs(4317) <= (layer2_outputs(4431)) xor (layer2_outputs(603));
    outputs(4318) <= layer2_outputs(3171);
    outputs(4319) <= not(layer2_outputs(1963));
    outputs(4320) <= not(layer2_outputs(3791));
    outputs(4321) <= (layer2_outputs(737)) or (layer2_outputs(405));
    outputs(4322) <= (layer2_outputs(1507)) or (layer2_outputs(3043));
    outputs(4323) <= layer2_outputs(4569);
    outputs(4324) <= (layer2_outputs(3869)) xor (layer2_outputs(2686));
    outputs(4325) <= layer2_outputs(985);
    outputs(4326) <= layer2_outputs(947);
    outputs(4327) <= layer2_outputs(4520);
    outputs(4328) <= not((layer2_outputs(342)) and (layer2_outputs(1227)));
    outputs(4329) <= not((layer2_outputs(4404)) xor (layer2_outputs(3844)));
    outputs(4330) <= not(layer2_outputs(2634)) or (layer2_outputs(3737));
    outputs(4331) <= layer2_outputs(1534);
    outputs(4332) <= layer2_outputs(4589);
    outputs(4333) <= layer2_outputs(4944);
    outputs(4334) <= layer2_outputs(3725);
    outputs(4335) <= (layer2_outputs(4794)) and not (layer2_outputs(1704));
    outputs(4336) <= not((layer2_outputs(4999)) and (layer2_outputs(1142)));
    outputs(4337) <= (layer2_outputs(2289)) xor (layer2_outputs(2663));
    outputs(4338) <= not((layer2_outputs(4435)) or (layer2_outputs(2398)));
    outputs(4339) <= not((layer2_outputs(1597)) xor (layer2_outputs(4580)));
    outputs(4340) <= (layer2_outputs(1428)) and not (layer2_outputs(2479));
    outputs(4341) <= layer2_outputs(3766);
    outputs(4342) <= layer2_outputs(447);
    outputs(4343) <= not(layer2_outputs(1762));
    outputs(4344) <= not((layer2_outputs(2634)) or (layer2_outputs(4464)));
    outputs(4345) <= (layer2_outputs(2421)) xor (layer2_outputs(2485));
    outputs(4346) <= (layer2_outputs(2256)) xor (layer2_outputs(2009));
    outputs(4347) <= layer2_outputs(3621);
    outputs(4348) <= (layer2_outputs(162)) and not (layer2_outputs(115));
    outputs(4349) <= (layer2_outputs(5104)) and (layer2_outputs(3342));
    outputs(4350) <= not(layer2_outputs(356));
    outputs(4351) <= layer2_outputs(659);
    outputs(4352) <= (layer2_outputs(3849)) and (layer2_outputs(345));
    outputs(4353) <= (layer2_outputs(1069)) xor (layer2_outputs(4093));
    outputs(4354) <= not(layer2_outputs(4413));
    outputs(4355) <= not((layer2_outputs(2688)) xor (layer2_outputs(962)));
    outputs(4356) <= not(layer2_outputs(4997));
    outputs(4357) <= not(layer2_outputs(258));
    outputs(4358) <= layer2_outputs(3571);
    outputs(4359) <= (layer2_outputs(2359)) xor (layer2_outputs(3253));
    outputs(4360) <= not((layer2_outputs(5081)) and (layer2_outputs(5006)));
    outputs(4361) <= not(layer2_outputs(1802)) or (layer2_outputs(595));
    outputs(4362) <= (layer2_outputs(3679)) xor (layer2_outputs(3965));
    outputs(4363) <= not(layer2_outputs(4782));
    outputs(4364) <= not(layer2_outputs(4292)) or (layer2_outputs(2943));
    outputs(4365) <= layer2_outputs(4599);
    outputs(4366) <= layer2_outputs(1778);
    outputs(4367) <= not(layer2_outputs(876)) or (layer2_outputs(3616));
    outputs(4368) <= not(layer2_outputs(1509)) or (layer2_outputs(4610));
    outputs(4369) <= layer2_outputs(1277);
    outputs(4370) <= layer2_outputs(4288);
    outputs(4371) <= not(layer2_outputs(2235));
    outputs(4372) <= not(layer2_outputs(4921));
    outputs(4373) <= layer2_outputs(5011);
    outputs(4374) <= layer2_outputs(3037);
    outputs(4375) <= not((layer2_outputs(2237)) xor (layer2_outputs(4310)));
    outputs(4376) <= layer2_outputs(4303);
    outputs(4377) <= not(layer2_outputs(1093));
    outputs(4378) <= layer2_outputs(1978);
    outputs(4379) <= not(layer2_outputs(403));
    outputs(4380) <= (layer2_outputs(1427)) xor (layer2_outputs(3674));
    outputs(4381) <= not(layer2_outputs(2322));
    outputs(4382) <= not(layer2_outputs(1129));
    outputs(4383) <= not((layer2_outputs(1405)) xor (layer2_outputs(4212)));
    outputs(4384) <= layer2_outputs(4463);
    outputs(4385) <= (layer2_outputs(1711)) xor (layer2_outputs(3108));
    outputs(4386) <= not(layer2_outputs(1800));
    outputs(4387) <= not((layer2_outputs(3911)) xor (layer2_outputs(2494)));
    outputs(4388) <= not(layer2_outputs(2193));
    outputs(4389) <= not((layer2_outputs(590)) and (layer2_outputs(2819)));
    outputs(4390) <= not(layer2_outputs(3590));
    outputs(4391) <= layer2_outputs(5104);
    outputs(4392) <= not(layer2_outputs(1373));
    outputs(4393) <= not(layer2_outputs(2679)) or (layer2_outputs(3606));
    outputs(4394) <= not(layer2_outputs(2020));
    outputs(4395) <= not(layer2_outputs(3787));
    outputs(4396) <= not(layer2_outputs(3863)) or (layer2_outputs(2739));
    outputs(4397) <= not(layer2_outputs(4379));
    outputs(4398) <= not((layer2_outputs(3385)) or (layer2_outputs(4626)));
    outputs(4399) <= layer2_outputs(2992);
    outputs(4400) <= not((layer2_outputs(1455)) or (layer2_outputs(4747)));
    outputs(4401) <= not((layer2_outputs(3390)) xor (layer2_outputs(3612)));
    outputs(4402) <= not(layer2_outputs(4827));
    outputs(4403) <= layer2_outputs(1229);
    outputs(4404) <= not(layer2_outputs(3973));
    outputs(4405) <= layer2_outputs(3155);
    outputs(4406) <= layer2_outputs(3409);
    outputs(4407) <= not(layer2_outputs(2318));
    outputs(4408) <= layer2_outputs(1146);
    outputs(4409) <= layer2_outputs(202);
    outputs(4410) <= not(layer2_outputs(4471)) or (layer2_outputs(105));
    outputs(4411) <= layer2_outputs(3360);
    outputs(4412) <= not(layer2_outputs(249));
    outputs(4413) <= (layer2_outputs(2606)) and (layer2_outputs(484));
    outputs(4414) <= not((layer2_outputs(2861)) xor (layer2_outputs(306)));
    outputs(4415) <= not(layer2_outputs(1493));
    outputs(4416) <= not(layer2_outputs(718)) or (layer2_outputs(2121));
    outputs(4417) <= (layer2_outputs(1983)) xor (layer2_outputs(1390));
    outputs(4418) <= (layer2_outputs(2814)) and (layer2_outputs(4900));
    outputs(4419) <= layer2_outputs(3928);
    outputs(4420) <= layer2_outputs(4995);
    outputs(4421) <= layer2_outputs(1338);
    outputs(4422) <= not(layer2_outputs(1605));
    outputs(4423) <= not(layer2_outputs(2459));
    outputs(4424) <= layer2_outputs(4370);
    outputs(4425) <= (layer2_outputs(2349)) or (layer2_outputs(2360));
    outputs(4426) <= layer2_outputs(1912);
    outputs(4427) <= (layer2_outputs(2772)) xor (layer2_outputs(2323));
    outputs(4428) <= (layer2_outputs(1860)) xor (layer2_outputs(1651));
    outputs(4429) <= not((layer2_outputs(3662)) xor (layer2_outputs(2423)));
    outputs(4430) <= not((layer2_outputs(636)) or (layer2_outputs(4089)));
    outputs(4431) <= (layer2_outputs(3930)) or (layer2_outputs(2120));
    outputs(4432) <= layer2_outputs(846);
    outputs(4433) <= not(layer2_outputs(3462));
    outputs(4434) <= layer2_outputs(4617);
    outputs(4435) <= (layer2_outputs(3586)) xor (layer2_outputs(367));
    outputs(4436) <= (layer2_outputs(4728)) and (layer2_outputs(1188));
    outputs(4437) <= layer2_outputs(623);
    outputs(4438) <= (layer2_outputs(3132)) xor (layer2_outputs(2328));
    outputs(4439) <= not(layer2_outputs(4400));
    outputs(4440) <= layer2_outputs(3611);
    outputs(4441) <= not(layer2_outputs(1764));
    outputs(4442) <= layer2_outputs(4162);
    outputs(4443) <= (layer2_outputs(3231)) xor (layer2_outputs(1368));
    outputs(4444) <= layer2_outputs(3281);
    outputs(4445) <= not(layer2_outputs(1135));
    outputs(4446) <= not(layer2_outputs(1708));
    outputs(4447) <= layer2_outputs(1820);
    outputs(4448) <= not((layer2_outputs(4544)) or (layer2_outputs(1803)));
    outputs(4449) <= (layer2_outputs(408)) or (layer2_outputs(4269));
    outputs(4450) <= layer2_outputs(4685);
    outputs(4451) <= not(layer2_outputs(2410));
    outputs(4452) <= layer2_outputs(536);
    outputs(4453) <= (layer2_outputs(2665)) and (layer2_outputs(70));
    outputs(4454) <= layer2_outputs(3472);
    outputs(4455) <= not(layer2_outputs(25));
    outputs(4456) <= layer2_outputs(1087);
    outputs(4457) <= not(layer2_outputs(1997)) or (layer2_outputs(4845));
    outputs(4458) <= layer2_outputs(4328);
    outputs(4459) <= not(layer2_outputs(1459));
    outputs(4460) <= layer2_outputs(4913);
    outputs(4461) <= layer2_outputs(2538);
    outputs(4462) <= not(layer2_outputs(3669));
    outputs(4463) <= layer2_outputs(2952);
    outputs(4464) <= not(layer2_outputs(3929));
    outputs(4465) <= layer2_outputs(232);
    outputs(4466) <= layer2_outputs(1183);
    outputs(4467) <= not((layer2_outputs(410)) and (layer2_outputs(2059)));
    outputs(4468) <= not((layer2_outputs(5002)) and (layer2_outputs(2994)));
    outputs(4469) <= not(layer2_outputs(4182));
    outputs(4470) <= layer2_outputs(3160);
    outputs(4471) <= (layer2_outputs(4830)) xor (layer2_outputs(583));
    outputs(4472) <= not(layer2_outputs(92)) or (layer2_outputs(325));
    outputs(4473) <= not((layer2_outputs(3173)) xor (layer2_outputs(5012)));
    outputs(4474) <= (layer2_outputs(1861)) and not (layer2_outputs(1053));
    outputs(4475) <= not(layer2_outputs(2874));
    outputs(4476) <= not(layer2_outputs(1743));
    outputs(4477) <= not(layer2_outputs(1542));
    outputs(4478) <= not(layer2_outputs(2134));
    outputs(4479) <= not(layer2_outputs(180));
    outputs(4480) <= (layer2_outputs(4410)) xor (layer2_outputs(635));
    outputs(4481) <= not(layer2_outputs(3551)) or (layer2_outputs(3476));
    outputs(4482) <= not(layer2_outputs(3684));
    outputs(4483) <= (layer2_outputs(2280)) xor (layer2_outputs(2770));
    outputs(4484) <= (layer2_outputs(3288)) xor (layer2_outputs(3109));
    outputs(4485) <= layer2_outputs(316);
    outputs(4486) <= not((layer2_outputs(3581)) xor (layer2_outputs(3995)));
    outputs(4487) <= not(layer2_outputs(3042)) or (layer2_outputs(4607));
    outputs(4488) <= (layer2_outputs(2389)) and not (layer2_outputs(3400));
    outputs(4489) <= (layer2_outputs(1019)) and not (layer2_outputs(2859));
    outputs(4490) <= layer2_outputs(1985);
    outputs(4491) <= layer2_outputs(566);
    outputs(4492) <= not((layer2_outputs(1454)) xor (layer2_outputs(4850)));
    outputs(4493) <= layer2_outputs(485);
    outputs(4494) <= layer2_outputs(1714);
    outputs(4495) <= layer2_outputs(4994);
    outputs(4496) <= not((layer2_outputs(1965)) or (layer2_outputs(3099)));
    outputs(4497) <= layer2_outputs(750);
    outputs(4498) <= not((layer2_outputs(4799)) xor (layer2_outputs(2241)));
    outputs(4499) <= layer2_outputs(3802);
    outputs(4500) <= not(layer2_outputs(4198));
    outputs(4501) <= (layer2_outputs(2593)) or (layer2_outputs(2698));
    outputs(4502) <= not(layer2_outputs(2523));
    outputs(4503) <= (layer2_outputs(571)) and not (layer2_outputs(801));
    outputs(4504) <= not(layer2_outputs(3173));
    outputs(4505) <= (layer2_outputs(4969)) xor (layer2_outputs(2622));
    outputs(4506) <= (layer2_outputs(4718)) and not (layer2_outputs(19));
    outputs(4507) <= not(layer2_outputs(1933));
    outputs(4508) <= not(layer2_outputs(3713));
    outputs(4509) <= layer2_outputs(304);
    outputs(4510) <= not(layer2_outputs(2016)) or (layer2_outputs(1725));
    outputs(4511) <= not(layer2_outputs(4340));
    outputs(4512) <= (layer2_outputs(3391)) xor (layer2_outputs(637));
    outputs(4513) <= not((layer2_outputs(765)) xor (layer2_outputs(3860)));
    outputs(4514) <= (layer2_outputs(2730)) and not (layer2_outputs(3081));
    outputs(4515) <= (layer2_outputs(4417)) and not (layer2_outputs(4657));
    outputs(4516) <= (layer2_outputs(974)) and (layer2_outputs(946));
    outputs(4517) <= (layer2_outputs(112)) or (layer2_outputs(4376));
    outputs(4518) <= not((layer2_outputs(100)) or (layer2_outputs(1573)));
    outputs(4519) <= layer2_outputs(202);
    outputs(4520) <= not(layer2_outputs(652));
    outputs(4521) <= layer2_outputs(1529);
    outputs(4522) <= layer2_outputs(1722);
    outputs(4523) <= not(layer2_outputs(3894));
    outputs(4524) <= not(layer2_outputs(4704));
    outputs(4525) <= layer2_outputs(4769);
    outputs(4526) <= not(layer2_outputs(2745));
    outputs(4527) <= layer2_outputs(1540);
    outputs(4528) <= not(layer2_outputs(2073));
    outputs(4529) <= (layer2_outputs(175)) xor (layer2_outputs(1276));
    outputs(4530) <= (layer2_outputs(4683)) or (layer2_outputs(5034));
    outputs(4531) <= (layer2_outputs(1585)) and (layer2_outputs(974));
    outputs(4532) <= not(layer2_outputs(3480));
    outputs(4533) <= not(layer2_outputs(709));
    outputs(4534) <= not(layer2_outputs(365));
    outputs(4535) <= not((layer2_outputs(681)) xor (layer2_outputs(203)));
    outputs(4536) <= layer2_outputs(2837);
    outputs(4537) <= not(layer2_outputs(3791));
    outputs(4538) <= layer2_outputs(1957);
    outputs(4539) <= not(layer2_outputs(2119));
    outputs(4540) <= layer2_outputs(155);
    outputs(4541) <= not(layer2_outputs(2826));
    outputs(4542) <= (layer2_outputs(2166)) and not (layer2_outputs(72));
    outputs(4543) <= not((layer2_outputs(3866)) xor (layer2_outputs(2391)));
    outputs(4544) <= not((layer2_outputs(188)) or (layer2_outputs(4286)));
    outputs(4545) <= layer2_outputs(4578);
    outputs(4546) <= not(layer2_outputs(2843));
    outputs(4547) <= not(layer2_outputs(1529)) or (layer2_outputs(4734));
    outputs(4548) <= layer2_outputs(4416);
    outputs(4549) <= not(layer2_outputs(3023));
    outputs(4550) <= layer2_outputs(4857);
    outputs(4551) <= not((layer2_outputs(420)) and (layer2_outputs(1828)));
    outputs(4552) <= (layer2_outputs(1795)) and (layer2_outputs(4661));
    outputs(4553) <= not((layer2_outputs(1998)) xor (layer2_outputs(2409)));
    outputs(4554) <= not(layer2_outputs(165));
    outputs(4555) <= (layer2_outputs(4350)) and not (layer2_outputs(1054));
    outputs(4556) <= (layer2_outputs(91)) and not (layer2_outputs(1236));
    outputs(4557) <= layer2_outputs(4348);
    outputs(4558) <= (layer2_outputs(3528)) and not (layer2_outputs(4447));
    outputs(4559) <= not((layer2_outputs(3735)) xor (layer2_outputs(550)));
    outputs(4560) <= layer2_outputs(5024);
    outputs(4561) <= layer2_outputs(437);
    outputs(4562) <= not((layer2_outputs(619)) xor (layer2_outputs(822)));
    outputs(4563) <= not(layer2_outputs(1410));
    outputs(4564) <= (layer2_outputs(2373)) and not (layer2_outputs(100));
    outputs(4565) <= layer2_outputs(750);
    outputs(4566) <= not(layer2_outputs(1303));
    outputs(4567) <= not((layer2_outputs(4245)) or (layer2_outputs(5053)));
    outputs(4568) <= layer2_outputs(2928);
    outputs(4569) <= not(layer2_outputs(1109));
    outputs(4570) <= layer2_outputs(1180);
    outputs(4571) <= not(layer2_outputs(880));
    outputs(4572) <= (layer2_outputs(4695)) xor (layer2_outputs(2790));
    outputs(4573) <= layer2_outputs(905);
    outputs(4574) <= layer2_outputs(2199);
    outputs(4575) <= not(layer2_outputs(2430));
    outputs(4576) <= not((layer2_outputs(1449)) xor (layer2_outputs(3706)));
    outputs(4577) <= layer2_outputs(3599);
    outputs(4578) <= (layer2_outputs(4811)) and not (layer2_outputs(2609));
    outputs(4579) <= not(layer2_outputs(1501));
    outputs(4580) <= layer2_outputs(1181);
    outputs(4581) <= not(layer2_outputs(4415));
    outputs(4582) <= not((layer2_outputs(1944)) xor (layer2_outputs(4032)));
    outputs(4583) <= not(layer2_outputs(2560));
    outputs(4584) <= layer2_outputs(2926);
    outputs(4585) <= layer2_outputs(4906);
    outputs(4586) <= layer2_outputs(3409);
    outputs(4587) <= not((layer2_outputs(4108)) xor (layer2_outputs(4803)));
    outputs(4588) <= layer2_outputs(487);
    outputs(4589) <= (layer2_outputs(1097)) xor (layer2_outputs(751));
    outputs(4590) <= not(layer2_outputs(3019));
    outputs(4591) <= layer2_outputs(1488);
    outputs(4592) <= (layer2_outputs(1671)) and (layer2_outputs(877));
    outputs(4593) <= layer2_outputs(4469);
    outputs(4594) <= layer2_outputs(4401);
    outputs(4595) <= (layer2_outputs(1426)) xor (layer2_outputs(4911));
    outputs(4596) <= not((layer2_outputs(4600)) xor (layer2_outputs(4584)));
    outputs(4597) <= (layer2_outputs(3353)) and not (layer2_outputs(3993));
    outputs(4598) <= not((layer2_outputs(2288)) and (layer2_outputs(5093)));
    outputs(4599) <= not(layer2_outputs(2633));
    outputs(4600) <= (layer2_outputs(2289)) xor (layer2_outputs(605));
    outputs(4601) <= not(layer2_outputs(3552)) or (layer2_outputs(2402));
    outputs(4602) <= not((layer2_outputs(2244)) or (layer2_outputs(1376)));
    outputs(4603) <= not(layer2_outputs(2256));
    outputs(4604) <= not(layer2_outputs(517)) or (layer2_outputs(3471));
    outputs(4605) <= not(layer2_outputs(2063)) or (layer2_outputs(302));
    outputs(4606) <= (layer2_outputs(276)) and not (layer2_outputs(3056));
    outputs(4607) <= not(layer2_outputs(569));
    outputs(4608) <= layer2_outputs(144);
    outputs(4609) <= (layer2_outputs(1975)) xor (layer2_outputs(3379));
    outputs(4610) <= (layer2_outputs(2515)) and not (layer2_outputs(3562));
    outputs(4611) <= not((layer2_outputs(1934)) or (layer2_outputs(3270)));
    outputs(4612) <= not((layer2_outputs(3773)) and (layer2_outputs(4886)));
    outputs(4613) <= layer2_outputs(3193);
    outputs(4614) <= (layer2_outputs(3489)) xor (layer2_outputs(2163));
    outputs(4615) <= not(layer2_outputs(3204));
    outputs(4616) <= not(layer2_outputs(1113));
    outputs(4617) <= layer2_outputs(5069);
    outputs(4618) <= not(layer2_outputs(1595));
    outputs(4619) <= not(layer2_outputs(1321));
    outputs(4620) <= not((layer2_outputs(497)) or (layer2_outputs(4740)));
    outputs(4621) <= layer2_outputs(111);
    outputs(4622) <= layer2_outputs(812);
    outputs(4623) <= (layer2_outputs(4341)) and (layer2_outputs(4666));
    outputs(4624) <= (layer2_outputs(2326)) and not (layer2_outputs(2878));
    outputs(4625) <= layer2_outputs(3912);
    outputs(4626) <= layer2_outputs(172);
    outputs(4627) <= (layer2_outputs(1042)) xor (layer2_outputs(786));
    outputs(4628) <= not(layer2_outputs(4176));
    outputs(4629) <= not(layer2_outputs(1129));
    outputs(4630) <= layer2_outputs(1425);
    outputs(4631) <= layer2_outputs(4447);
    outputs(4632) <= (layer2_outputs(562)) and not (layer2_outputs(4834));
    outputs(4633) <= not(layer2_outputs(3187));
    outputs(4634) <= not(layer2_outputs(1590));
    outputs(4635) <= (layer2_outputs(2012)) and not (layer2_outputs(592));
    outputs(4636) <= layer2_outputs(3380);
    outputs(4637) <= layer2_outputs(2797);
    outputs(4638) <= (layer2_outputs(639)) and (layer2_outputs(1865));
    outputs(4639) <= not(layer2_outputs(4207));
    outputs(4640) <= layer2_outputs(1009);
    outputs(4641) <= not((layer2_outputs(2156)) xor (layer2_outputs(2601)));
    outputs(4642) <= (layer2_outputs(2012)) and not (layer2_outputs(620));
    outputs(4643) <= not(layer2_outputs(2013));
    outputs(4644) <= layer2_outputs(2309);
    outputs(4645) <= not((layer2_outputs(1767)) xor (layer2_outputs(3255)));
    outputs(4646) <= not(layer2_outputs(3618));
    outputs(4647) <= layer2_outputs(4275);
    outputs(4648) <= (layer2_outputs(2866)) and not (layer2_outputs(1653));
    outputs(4649) <= not(layer2_outputs(2469));
    outputs(4650) <= not((layer2_outputs(1095)) and (layer2_outputs(215)));
    outputs(4651) <= layer2_outputs(387);
    outputs(4652) <= not(layer2_outputs(3866));
    outputs(4653) <= (layer2_outputs(1179)) and not (layer2_outputs(302));
    outputs(4654) <= layer2_outputs(528);
    outputs(4655) <= not((layer2_outputs(2039)) xor (layer2_outputs(2739)));
    outputs(4656) <= (layer2_outputs(1922)) and (layer2_outputs(3789));
    outputs(4657) <= not(layer2_outputs(882));
    outputs(4658) <= not(layer2_outputs(2516));
    outputs(4659) <= layer2_outputs(3374);
    outputs(4660) <= not((layer2_outputs(3251)) xor (layer2_outputs(3921)));
    outputs(4661) <= not(layer2_outputs(1563));
    outputs(4662) <= not((layer2_outputs(2260)) or (layer2_outputs(1110)));
    outputs(4663) <= layer2_outputs(779);
    outputs(4664) <= not(layer2_outputs(4032));
    outputs(4665) <= layer2_outputs(2682);
    outputs(4666) <= layer2_outputs(4029);
    outputs(4667) <= (layer2_outputs(4139)) and (layer2_outputs(1849));
    outputs(4668) <= not(layer2_outputs(2501));
    outputs(4669) <= not(layer2_outputs(5058));
    outputs(4670) <= (layer2_outputs(1809)) and not (layer2_outputs(2557));
    outputs(4671) <= (layer2_outputs(286)) and not (layer2_outputs(2238));
    outputs(4672) <= not((layer2_outputs(4929)) or (layer2_outputs(2334)));
    outputs(4673) <= not(layer2_outputs(4573));
    outputs(4674) <= layer2_outputs(562);
    outputs(4675) <= not(layer2_outputs(4189));
    outputs(4676) <= layer2_outputs(1674);
    outputs(4677) <= not(layer2_outputs(659));
    outputs(4678) <= (layer2_outputs(2186)) and (layer2_outputs(2418));
    outputs(4679) <= not((layer2_outputs(3180)) or (layer2_outputs(4262)));
    outputs(4680) <= (layer2_outputs(2514)) and (layer2_outputs(841));
    outputs(4681) <= (layer2_outputs(3765)) xor (layer2_outputs(1539));
    outputs(4682) <= (layer2_outputs(1031)) xor (layer2_outputs(4924));
    outputs(4683) <= not(layer2_outputs(4880));
    outputs(4684) <= not(layer2_outputs(4311));
    outputs(4685) <= not(layer2_outputs(44));
    outputs(4686) <= not(layer2_outputs(1582));
    outputs(4687) <= layer2_outputs(4317);
    outputs(4688) <= (layer2_outputs(164)) and not (layer2_outputs(2028));
    outputs(4689) <= not((layer2_outputs(4629)) or (layer2_outputs(4414)));
    outputs(4690) <= layer2_outputs(3482);
    outputs(4691) <= (layer2_outputs(4297)) and not (layer2_outputs(3441));
    outputs(4692) <= layer2_outputs(1278);
    outputs(4693) <= not(layer2_outputs(2078));
    outputs(4694) <= (layer2_outputs(3589)) and (layer2_outputs(3097));
    outputs(4695) <= layer2_outputs(3727);
    outputs(4696) <= layer2_outputs(658);
    outputs(4697) <= layer2_outputs(3630);
    outputs(4698) <= layer2_outputs(3836);
    outputs(4699) <= (layer2_outputs(4824)) and (layer2_outputs(595));
    outputs(4700) <= not(layer2_outputs(1208));
    outputs(4701) <= not((layer2_outputs(3255)) xor (layer2_outputs(1961)));
    outputs(4702) <= (layer2_outputs(4116)) and not (layer2_outputs(1934));
    outputs(4703) <= layer2_outputs(3553);
    outputs(4704) <= not((layer2_outputs(1698)) or (layer2_outputs(2857)));
    outputs(4705) <= not((layer2_outputs(2447)) or (layer2_outputs(2325)));
    outputs(4706) <= not((layer2_outputs(2675)) xor (layer2_outputs(3345)));
    outputs(4707) <= (layer2_outputs(2032)) xor (layer2_outputs(710));
    outputs(4708) <= (layer2_outputs(4267)) xor (layer2_outputs(1681));
    outputs(4709) <= not((layer2_outputs(142)) and (layer2_outputs(2375)));
    outputs(4710) <= not(layer2_outputs(4894));
    outputs(4711) <= not((layer2_outputs(2599)) xor (layer2_outputs(4384)));
    outputs(4712) <= layer2_outputs(3515);
    outputs(4713) <= layer2_outputs(2777);
    outputs(4714) <= not((layer2_outputs(3191)) xor (layer2_outputs(979)));
    outputs(4715) <= layer2_outputs(5081);
    outputs(4716) <= not(layer2_outputs(1436));
    outputs(4717) <= (layer2_outputs(3138)) and not (layer2_outputs(322));
    outputs(4718) <= not(layer2_outputs(3445));
    outputs(4719) <= not(layer2_outputs(3952));
    outputs(4720) <= (layer2_outputs(1544)) xor (layer2_outputs(3384));
    outputs(4721) <= layer2_outputs(3182);
    outputs(4722) <= layer2_outputs(711);
    outputs(4723) <= layer2_outputs(687);
    outputs(4724) <= layer2_outputs(2298);
    outputs(4725) <= not(layer2_outputs(640));
    outputs(4726) <= layer2_outputs(539);
    outputs(4727) <= layer2_outputs(4554);
    outputs(4728) <= (layer2_outputs(782)) and not (layer2_outputs(4929));
    outputs(4729) <= not(layer2_outputs(4179));
    outputs(4730) <= layer2_outputs(58);
    outputs(4731) <= (layer2_outputs(668)) and (layer2_outputs(2930));
    outputs(4732) <= (layer2_outputs(266)) and not (layer2_outputs(4545));
    outputs(4733) <= layer2_outputs(2206);
    outputs(4734) <= (layer2_outputs(4172)) or (layer2_outputs(1255));
    outputs(4735) <= not(layer2_outputs(5031)) or (layer2_outputs(2757));
    outputs(4736) <= layer2_outputs(4507);
    outputs(4737) <= (layer2_outputs(4013)) and not (layer2_outputs(2302));
    outputs(4738) <= (layer2_outputs(4156)) xor (layer2_outputs(138));
    outputs(4739) <= layer2_outputs(663);
    outputs(4740) <= not(layer2_outputs(2478));
    outputs(4741) <= (layer2_outputs(33)) and not (layer2_outputs(2384));
    outputs(4742) <= not(layer2_outputs(3458));
    outputs(4743) <= not((layer2_outputs(368)) and (layer2_outputs(3656)));
    outputs(4744) <= layer2_outputs(1289);
    outputs(4745) <= not(layer2_outputs(1581));
    outputs(4746) <= layer2_outputs(369);
    outputs(4747) <= not((layer2_outputs(4514)) xor (layer2_outputs(3587)));
    outputs(4748) <= not(layer2_outputs(4344));
    outputs(4749) <= not(layer2_outputs(4372)) or (layer2_outputs(2761));
    outputs(4750) <= layer2_outputs(4781);
    outputs(4751) <= (layer2_outputs(2751)) and (layer2_outputs(4690));
    outputs(4752) <= not(layer2_outputs(4194));
    outputs(4753) <= not(layer2_outputs(2181));
    outputs(4754) <= (layer2_outputs(47)) and not (layer2_outputs(862));
    outputs(4755) <= not(layer2_outputs(1280));
    outputs(4756) <= not(layer2_outputs(511));
    outputs(4757) <= not(layer2_outputs(1416));
    outputs(4758) <= (layer2_outputs(1421)) and (layer2_outputs(1323));
    outputs(4759) <= not(layer2_outputs(986));
    outputs(4760) <= not(layer2_outputs(4670));
    outputs(4761) <= (layer2_outputs(3857)) xor (layer2_outputs(2234));
    outputs(4762) <= not(layer2_outputs(592));
    outputs(4763) <= layer2_outputs(4525);
    outputs(4764) <= (layer2_outputs(1445)) xor (layer2_outputs(3539));
    outputs(4765) <= layer2_outputs(3990);
    outputs(4766) <= not((layer2_outputs(502)) or (layer2_outputs(2350)));
    outputs(4767) <= (layer2_outputs(2489)) xor (layer2_outputs(1841));
    outputs(4768) <= not(layer2_outputs(3203));
    outputs(4769) <= layer2_outputs(1928);
    outputs(4770) <= (layer2_outputs(2283)) and not (layer2_outputs(506));
    outputs(4771) <= layer2_outputs(4477);
    outputs(4772) <= layer2_outputs(435);
    outputs(4773) <= layer2_outputs(3076);
    outputs(4774) <= not(layer2_outputs(74)) or (layer2_outputs(2214));
    outputs(4775) <= not((layer2_outputs(4034)) xor (layer2_outputs(2339)));
    outputs(4776) <= (layer2_outputs(904)) and not (layer2_outputs(206));
    outputs(4777) <= not((layer2_outputs(3510)) xor (layer2_outputs(4812)));
    outputs(4778) <= layer2_outputs(1412);
    outputs(4779) <= (layer2_outputs(4473)) and not (layer2_outputs(690));
    outputs(4780) <= not((layer2_outputs(2158)) or (layer2_outputs(1016)));
    outputs(4781) <= not(layer2_outputs(3223));
    outputs(4782) <= not((layer2_outputs(1350)) xor (layer2_outputs(848)));
    outputs(4783) <= not(layer2_outputs(628));
    outputs(4784) <= (layer2_outputs(612)) and not (layer2_outputs(667));
    outputs(4785) <= not(layer2_outputs(1851)) or (layer2_outputs(4044));
    outputs(4786) <= not((layer2_outputs(3786)) xor (layer2_outputs(3090)));
    outputs(4787) <= (layer2_outputs(3367)) and not (layer2_outputs(4086));
    outputs(4788) <= (layer2_outputs(1506)) and not (layer2_outputs(3124));
    outputs(4789) <= not((layer2_outputs(2451)) or (layer2_outputs(4173)));
    outputs(4790) <= not(layer2_outputs(3666)) or (layer2_outputs(402));
    outputs(4791) <= layer2_outputs(3112);
    outputs(4792) <= not((layer2_outputs(4212)) xor (layer2_outputs(1753)));
    outputs(4793) <= (layer2_outputs(2311)) xor (layer2_outputs(3544));
    outputs(4794) <= layer2_outputs(3415);
    outputs(4795) <= (layer2_outputs(3946)) or (layer2_outputs(4642));
    outputs(4796) <= (layer2_outputs(4818)) or (layer2_outputs(2994));
    outputs(4797) <= (layer2_outputs(1701)) and not (layer2_outputs(3168));
    outputs(4798) <= not(layer2_outputs(570));
    outputs(4799) <= not((layer2_outputs(4533)) xor (layer2_outputs(1997)));
    outputs(4800) <= not(layer2_outputs(2054));
    outputs(4801) <= not(layer2_outputs(594)) or (layer2_outputs(5021));
    outputs(4802) <= not(layer2_outputs(79));
    outputs(4803) <= (layer2_outputs(3126)) and not (layer2_outputs(1817));
    outputs(4804) <= layer2_outputs(212);
    outputs(4805) <= (layer2_outputs(3875)) xor (layer2_outputs(132));
    outputs(4806) <= layer2_outputs(1432);
    outputs(4807) <= layer2_outputs(1372);
    outputs(4808) <= not(layer2_outputs(2315));
    outputs(4809) <= layer2_outputs(1526);
    outputs(4810) <= not(layer2_outputs(2857));
    outputs(4811) <= not(layer2_outputs(1069));
    outputs(4812) <= (layer2_outputs(55)) and not (layer2_outputs(2290));
    outputs(4813) <= layer2_outputs(978);
    outputs(4814) <= not((layer2_outputs(523)) xor (layer2_outputs(634)));
    outputs(4815) <= layer2_outputs(4434);
    outputs(4816) <= layer2_outputs(652);
    outputs(4817) <= not(layer2_outputs(347));
    outputs(4818) <= layer2_outputs(2434);
    outputs(4819) <= layer2_outputs(2089);
    outputs(4820) <= (layer2_outputs(379)) and not (layer2_outputs(2291));
    outputs(4821) <= (layer2_outputs(2099)) and not (layer2_outputs(2084));
    outputs(4822) <= layer2_outputs(323);
    outputs(4823) <= not(layer2_outputs(500)) or (layer2_outputs(5044));
    outputs(4824) <= layer2_outputs(4660);
    outputs(4825) <= not(layer2_outputs(1827)) or (layer2_outputs(688));
    outputs(4826) <= layer2_outputs(1090);
    outputs(4827) <= layer2_outputs(281);
    outputs(4828) <= not(layer2_outputs(719));
    outputs(4829) <= not(layer2_outputs(3217));
    outputs(4830) <= not(layer2_outputs(187));
    outputs(4831) <= not(layer2_outputs(2807)) or (layer2_outputs(1306));
    outputs(4832) <= layer2_outputs(4932);
    outputs(4833) <= not(layer2_outputs(2122));
    outputs(4834) <= not(layer2_outputs(1060));
    outputs(4835) <= not(layer2_outputs(1196));
    outputs(4836) <= layer2_outputs(760);
    outputs(4837) <= layer2_outputs(1964);
    outputs(4838) <= not(layer2_outputs(326));
    outputs(4839) <= not(layer2_outputs(177));
    outputs(4840) <= layer2_outputs(2760);
    outputs(4841) <= not(layer2_outputs(4973));
    outputs(4842) <= (layer2_outputs(405)) and not (layer2_outputs(5111));
    outputs(4843) <= layer2_outputs(2179);
    outputs(4844) <= (layer2_outputs(510)) and (layer2_outputs(2619));
    outputs(4845) <= (layer2_outputs(4163)) or (layer2_outputs(673));
    outputs(4846) <= not(layer2_outputs(4278));
    outputs(4847) <= not(layer2_outputs(1982));
    outputs(4848) <= not(layer2_outputs(3952));
    outputs(4849) <= (layer2_outputs(465)) and (layer2_outputs(3338));
    outputs(4850) <= layer2_outputs(742);
    outputs(4851) <= not((layer2_outputs(990)) xor (layer2_outputs(2883)));
    outputs(4852) <= (layer2_outputs(2391)) and not (layer2_outputs(1898));
    outputs(4853) <= layer2_outputs(2623);
    outputs(4854) <= not((layer2_outputs(4872)) and (layer2_outputs(4536)));
    outputs(4855) <= not((layer2_outputs(3351)) or (layer2_outputs(1176)));
    outputs(4856) <= not((layer2_outputs(887)) and (layer2_outputs(4915)));
    outputs(4857) <= layer2_outputs(4696);
    outputs(4858) <= not((layer2_outputs(4114)) or (layer2_outputs(4561)));
    outputs(4859) <= (layer2_outputs(617)) xor (layer2_outputs(908));
    outputs(4860) <= (layer2_outputs(3885)) and not (layer2_outputs(300));
    outputs(4861) <= layer2_outputs(816);
    outputs(4862) <= not(layer2_outputs(4802)) or (layer2_outputs(4889));
    outputs(4863) <= (layer2_outputs(67)) and (layer2_outputs(3112));
    outputs(4864) <= layer2_outputs(2017);
    outputs(4865) <= not(layer2_outputs(1312));
    outputs(4866) <= (layer2_outputs(2981)) and not (layer2_outputs(4754));
    outputs(4867) <= layer2_outputs(2317);
    outputs(4868) <= layer2_outputs(2007);
    outputs(4869) <= not(layer2_outputs(56));
    outputs(4870) <= (layer2_outputs(3693)) xor (layer2_outputs(2180));
    outputs(4871) <= layer2_outputs(2107);
    outputs(4872) <= layer2_outputs(2546);
    outputs(4873) <= layer2_outputs(1791);
    outputs(4874) <= layer2_outputs(4752);
    outputs(4875) <= not(layer2_outputs(1561));
    outputs(4876) <= not(layer2_outputs(3032));
    outputs(4877) <= not(layer2_outputs(1271));
    outputs(4878) <= not(layer2_outputs(1954));
    outputs(4879) <= not((layer2_outputs(994)) or (layer2_outputs(4264)));
    outputs(4880) <= layer2_outputs(4565);
    outputs(4881) <= (layer2_outputs(3311)) and (layer2_outputs(3787));
    outputs(4882) <= layer2_outputs(1233);
    outputs(4883) <= (layer2_outputs(4355)) and (layer2_outputs(4575));
    outputs(4884) <= not(layer2_outputs(4130));
    outputs(4885) <= layer2_outputs(1207);
    outputs(4886) <= not(layer2_outputs(3931));
    outputs(4887) <= not(layer2_outputs(2839));
    outputs(4888) <= not(layer2_outputs(4530));
    outputs(4889) <= not(layer2_outputs(165));
    outputs(4890) <= layer2_outputs(1143);
    outputs(4891) <= not(layer2_outputs(4342));
    outputs(4892) <= not(layer2_outputs(4503));
    outputs(4893) <= layer2_outputs(3728);
    outputs(4894) <= layer2_outputs(2880);
    outputs(4895) <= not(layer2_outputs(4671));
    outputs(4896) <= layer2_outputs(4558);
    outputs(4897) <= layer2_outputs(832);
    outputs(4898) <= not(layer2_outputs(4539));
    outputs(4899) <= not(layer2_outputs(3813));
    outputs(4900) <= not(layer2_outputs(1105));
    outputs(4901) <= (layer2_outputs(1302)) xor (layer2_outputs(2617));
    outputs(4902) <= layer2_outputs(1318);
    outputs(4903) <= layer2_outputs(2703);
    outputs(4904) <= not(layer2_outputs(3670));
    outputs(4905) <= layer2_outputs(726);
    outputs(4906) <= not(layer2_outputs(95));
    outputs(4907) <= layer2_outputs(4932);
    outputs(4908) <= layer2_outputs(3954);
    outputs(4909) <= (layer2_outputs(4023)) and not (layer2_outputs(640));
    outputs(4910) <= layer2_outputs(777);
    outputs(4911) <= (layer2_outputs(2955)) and not (layer2_outputs(4028));
    outputs(4912) <= layer2_outputs(2046);
    outputs(4913) <= not((layer2_outputs(4405)) or (layer2_outputs(541)));
    outputs(4914) <= (layer2_outputs(2252)) and not (layer2_outputs(4196));
    outputs(4915) <= layer2_outputs(1024);
    outputs(4916) <= layer2_outputs(4418);
    outputs(4917) <= (layer2_outputs(950)) and not (layer2_outputs(2863));
    outputs(4918) <= layer2_outputs(5012);
    outputs(4919) <= layer2_outputs(1437);
    outputs(4920) <= layer2_outputs(1290);
    outputs(4921) <= (layer2_outputs(5048)) and (layer2_outputs(4492));
    outputs(4922) <= not(layer2_outputs(2918));
    outputs(4923) <= layer2_outputs(1929);
    outputs(4924) <= layer2_outputs(408);
    outputs(4925) <= (layer2_outputs(269)) and (layer2_outputs(4472));
    outputs(4926) <= layer2_outputs(3739);
    outputs(4927) <= not((layer2_outputs(3418)) and (layer2_outputs(4688)));
    outputs(4928) <= not(layer2_outputs(4068));
    outputs(4929) <= not(layer2_outputs(4786));
    outputs(4930) <= not(layer2_outputs(3113));
    outputs(4931) <= (layer2_outputs(1684)) and not (layer2_outputs(4443));
    outputs(4932) <= layer2_outputs(4895);
    outputs(4933) <= not(layer2_outputs(3122)) or (layer2_outputs(2349));
    outputs(4934) <= (layer2_outputs(4934)) and (layer2_outputs(1973));
    outputs(4935) <= not((layer2_outputs(4474)) and (layer2_outputs(952)));
    outputs(4936) <= layer2_outputs(1301);
    outputs(4937) <= layer2_outputs(3491);
    outputs(4938) <= not(layer2_outputs(4075));
    outputs(4939) <= layer2_outputs(3547);
    outputs(4940) <= layer2_outputs(3973);
    outputs(4941) <= not(layer2_outputs(1498));
    outputs(4942) <= not((layer2_outputs(4627)) xor (layer2_outputs(421)));
    outputs(4943) <= layer2_outputs(2597);
    outputs(4944) <= layer2_outputs(4668);
    outputs(4945) <= layer2_outputs(3125);
    outputs(4946) <= layer2_outputs(69);
    outputs(4947) <= not(layer2_outputs(2027));
    outputs(4948) <= not(layer2_outputs(1567));
    outputs(4949) <= not(layer2_outputs(1599));
    outputs(4950) <= layer2_outputs(1219);
    outputs(4951) <= (layer2_outputs(1660)) and (layer2_outputs(367));
    outputs(4952) <= not(layer2_outputs(898));
    outputs(4953) <= layer2_outputs(1812);
    outputs(4954) <= not((layer2_outputs(3777)) or (layer2_outputs(1168)));
    outputs(4955) <= not(layer2_outputs(533));
    outputs(4956) <= (layer2_outputs(1924)) and not (layer2_outputs(2970));
    outputs(4957) <= not(layer2_outputs(788));
    outputs(4958) <= not(layer2_outputs(2370));
    outputs(4959) <= layer2_outputs(2852);
    outputs(4960) <= not(layer2_outputs(357));
    outputs(4961) <= (layer2_outputs(4956)) and not (layer2_outputs(784));
    outputs(4962) <= not((layer2_outputs(1624)) or (layer2_outputs(4446)));
    outputs(4963) <= not(layer2_outputs(1911));
    outputs(4964) <= (layer2_outputs(2893)) or (layer2_outputs(3523));
    outputs(4965) <= not(layer2_outputs(3785));
    outputs(4966) <= not(layer2_outputs(3442));
    outputs(4967) <= not((layer2_outputs(633)) and (layer2_outputs(320)));
    outputs(4968) <= not((layer2_outputs(4465)) and (layer2_outputs(4875)));
    outputs(4969) <= not((layer2_outputs(4811)) xor (layer2_outputs(2921)));
    outputs(4970) <= layer2_outputs(4148);
    outputs(4971) <= (layer2_outputs(4991)) and not (layer2_outputs(3398));
    outputs(4972) <= not((layer2_outputs(1007)) or (layer2_outputs(2872)));
    outputs(4973) <= not(layer2_outputs(4395));
    outputs(4974) <= layer2_outputs(1632);
    outputs(4975) <= (layer2_outputs(3823)) and (layer2_outputs(3688));
    outputs(4976) <= not(layer2_outputs(5026)) or (layer2_outputs(1538));
    outputs(4977) <= not((layer2_outputs(1332)) xor (layer2_outputs(1823)));
    outputs(4978) <= (layer2_outputs(3986)) and not (layer2_outputs(147));
    outputs(4979) <= layer2_outputs(2728);
    outputs(4980) <= not(layer2_outputs(4908));
    outputs(4981) <= layer2_outputs(3152);
    outputs(4982) <= not(layer2_outputs(2877)) or (layer2_outputs(1201));
    outputs(4983) <= not(layer2_outputs(2608));
    outputs(4984) <= layer2_outputs(3971);
    outputs(4985) <= layer2_outputs(1770);
    outputs(4986) <= not(layer2_outputs(2664));
    outputs(4987) <= layer2_outputs(3689);
    outputs(4988) <= (layer2_outputs(2980)) or (layer2_outputs(3624));
    outputs(4989) <= not((layer2_outputs(3551)) xor (layer2_outputs(3072)));
    outputs(4990) <= not(layer2_outputs(4050));
    outputs(4991) <= layer2_outputs(555);
    outputs(4992) <= not(layer2_outputs(4219));
    outputs(4993) <= layer2_outputs(2909);
    outputs(4994) <= not(layer2_outputs(1297));
    outputs(4995) <= layer2_outputs(224);
    outputs(4996) <= (layer2_outputs(4826)) or (layer2_outputs(433));
    outputs(4997) <= layer2_outputs(2995);
    outputs(4998) <= layer2_outputs(1915);
    outputs(4999) <= layer2_outputs(4367);
    outputs(5000) <= not(layer2_outputs(3770));
    outputs(5001) <= layer2_outputs(1071);
    outputs(5002) <= not(layer2_outputs(4570));
    outputs(5003) <= not(layer2_outputs(2394));
    outputs(5004) <= layer2_outputs(2249);
    outputs(5005) <= layer2_outputs(424);
    outputs(5006) <= not((layer2_outputs(4169)) or (layer2_outputs(545)));
    outputs(5007) <= not((layer2_outputs(3963)) xor (layer2_outputs(312)));
    outputs(5008) <= (layer2_outputs(1400)) and (layer2_outputs(3303));
    outputs(5009) <= not(layer2_outputs(468));
    outputs(5010) <= not(layer2_outputs(4273));
    outputs(5011) <= not(layer2_outputs(2419));
    outputs(5012) <= not(layer2_outputs(2084));
    outputs(5013) <= layer2_outputs(2392);
    outputs(5014) <= not(layer2_outputs(4671));
    outputs(5015) <= not(layer2_outputs(3145));
    outputs(5016) <= not(layer2_outputs(201));
    outputs(5017) <= layer2_outputs(2552);
    outputs(5018) <= not(layer2_outputs(2371));
    outputs(5019) <= layer2_outputs(13);
    outputs(5020) <= not(layer2_outputs(3900));
    outputs(5021) <= not(layer2_outputs(2013));
    outputs(5022) <= layer2_outputs(2094);
    outputs(5023) <= not((layer2_outputs(4273)) or (layer2_outputs(4938)));
    outputs(5024) <= not(layer2_outputs(4654));
    outputs(5025) <= layer2_outputs(3901);
    outputs(5026) <= not(layer2_outputs(1585));
    outputs(5027) <= layer2_outputs(1674);
    outputs(5028) <= (layer2_outputs(5047)) xor (layer2_outputs(3144));
    outputs(5029) <= layer2_outputs(4227);
    outputs(5030) <= not(layer2_outputs(4561));
    outputs(5031) <= not((layer2_outputs(4606)) xor (layer2_outputs(1884)));
    outputs(5032) <= not(layer2_outputs(330));
    outputs(5033) <= layer2_outputs(1692);
    outputs(5034) <= (layer2_outputs(3895)) and not (layer2_outputs(1401));
    outputs(5035) <= not(layer2_outputs(1131));
    outputs(5036) <= (layer2_outputs(3033)) xor (layer2_outputs(4059));
    outputs(5037) <= (layer2_outputs(1638)) xor (layer2_outputs(2740));
    outputs(5038) <= not(layer2_outputs(4839));
    outputs(5039) <= not(layer2_outputs(4195));
    outputs(5040) <= not(layer2_outputs(227));
    outputs(5041) <= (layer2_outputs(831)) and not (layer2_outputs(1730));
    outputs(5042) <= layer2_outputs(1998);
    outputs(5043) <= layer2_outputs(346);
    outputs(5044) <= layer2_outputs(2388);
    outputs(5045) <= layer2_outputs(199);
    outputs(5046) <= (layer2_outputs(395)) and not (layer2_outputs(3738));
    outputs(5047) <= not(layer2_outputs(850)) or (layer2_outputs(3716));
    outputs(5048) <= not((layer2_outputs(3876)) xor (layer2_outputs(208)));
    outputs(5049) <= not((layer2_outputs(2637)) or (layer2_outputs(4370)));
    outputs(5050) <= not(layer2_outputs(3282));
    outputs(5051) <= layer2_outputs(1835);
    outputs(5052) <= layer2_outputs(3249);
    outputs(5053) <= (layer2_outputs(4312)) xor (layer2_outputs(4779));
    outputs(5054) <= not(layer2_outputs(4085));
    outputs(5055) <= not(layer2_outputs(2031));
    outputs(5056) <= not(layer2_outputs(2716));
    outputs(5057) <= (layer2_outputs(5100)) and not (layer2_outputs(59));
    outputs(5058) <= layer2_outputs(4989);
    outputs(5059) <= (layer2_outputs(3807)) xor (layer2_outputs(696));
    outputs(5060) <= not(layer2_outputs(1156));
    outputs(5061) <= layer2_outputs(1431);
    outputs(5062) <= layer2_outputs(2481);
    outputs(5063) <= not((layer2_outputs(850)) and (layer2_outputs(4601)));
    outputs(5064) <= (layer2_outputs(746)) and (layer2_outputs(2564));
    outputs(5065) <= not((layer2_outputs(2015)) and (layer2_outputs(1935)));
    outputs(5066) <= (layer2_outputs(2936)) and not (layer2_outputs(496));
    outputs(5067) <= not(layer2_outputs(3639));
    outputs(5068) <= not(layer2_outputs(2512));
    outputs(5069) <= layer2_outputs(9);
    outputs(5070) <= not(layer2_outputs(683));
    outputs(5071) <= layer2_outputs(2853);
    outputs(5072) <= not(layer2_outputs(1273));
    outputs(5073) <= (layer2_outputs(4145)) and (layer2_outputs(4598));
    outputs(5074) <= not(layer2_outputs(3006));
    outputs(5075) <= (layer2_outputs(3085)) and (layer2_outputs(2719));
    outputs(5076) <= not(layer2_outputs(2664));
    outputs(5077) <= not(layer2_outputs(1560));
    outputs(5078) <= (layer2_outputs(3997)) and (layer2_outputs(1807));
    outputs(5079) <= layer2_outputs(4246);
    outputs(5080) <= not((layer2_outputs(1493)) and (layer2_outputs(4513)));
    outputs(5081) <= not(layer2_outputs(3889));
    outputs(5082) <= (layer2_outputs(5090)) and not (layer2_outputs(3593));
    outputs(5083) <= layer2_outputs(2575);
    outputs(5084) <= not(layer2_outputs(4189));
    outputs(5085) <= layer2_outputs(3037);
    outputs(5086) <= (layer2_outputs(1712)) and (layer2_outputs(4698));
    outputs(5087) <= (layer2_outputs(3626)) and (layer2_outputs(4965));
    outputs(5088) <= (layer2_outputs(664)) and not (layer2_outputs(2141));
    outputs(5089) <= (layer2_outputs(4633)) xor (layer2_outputs(4722));
    outputs(5090) <= layer2_outputs(2803);
    outputs(5091) <= layer2_outputs(2001);
    outputs(5092) <= layer2_outputs(3306);
    outputs(5093) <= not(layer2_outputs(4724));
    outputs(5094) <= layer2_outputs(4611);
    outputs(5095) <= not(layer2_outputs(4471));
    outputs(5096) <= layer2_outputs(2413);
    outputs(5097) <= not(layer2_outputs(1349));
    outputs(5098) <= not(layer2_outputs(883));
    outputs(5099) <= (layer2_outputs(1935)) xor (layer2_outputs(1392));
    outputs(5100) <= layer2_outputs(395);
    outputs(5101) <= layer2_outputs(260);
    outputs(5102) <= (layer2_outputs(4544)) xor (layer2_outputs(4088));
    outputs(5103) <= not(layer2_outputs(4356));
    outputs(5104) <= layer2_outputs(2689);
    outputs(5105) <= layer2_outputs(538);
    outputs(5106) <= (layer2_outputs(4104)) and (layer2_outputs(593));
    outputs(5107) <= not(layer2_outputs(1888));
    outputs(5108) <= layer2_outputs(3020);
    outputs(5109) <= layer2_outputs(1707);
    outputs(5110) <= not((layer2_outputs(3357)) xor (layer2_outputs(3397)));
    outputs(5111) <= not((layer2_outputs(4091)) xor (layer2_outputs(2945)));
    outputs(5112) <= layer2_outputs(634);
    outputs(5113) <= not((layer2_outputs(3387)) or (layer2_outputs(3524)));
    outputs(5114) <= (layer2_outputs(4738)) and not (layer2_outputs(225));
    outputs(5115) <= not((layer2_outputs(4571)) or (layer2_outputs(2646)));
    outputs(5116) <= not((layer2_outputs(4255)) xor (layer2_outputs(4321)));
    outputs(5117) <= (layer2_outputs(2787)) and not (layer2_outputs(3329));
    outputs(5118) <= not(layer2_outputs(2934)) or (layer2_outputs(1628));
    outputs(5119) <= layer2_outputs(3434);

end Behavioral;
