library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(10239 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(10239 downto 0);

begin

    layer0_outputs(0) <= inputs(130);
    layer0_outputs(1) <= not((inputs(222)) or (inputs(91)));
    layer0_outputs(2) <= not((inputs(255)) xor (inputs(69)));
    layer0_outputs(3) <= not((inputs(247)) or (inputs(93)));
    layer0_outputs(4) <= not(inputs(234));
    layer0_outputs(5) <= (inputs(8)) or (inputs(34));
    layer0_outputs(6) <= not((inputs(80)) xor (inputs(49)));
    layer0_outputs(7) <= inputs(109);
    layer0_outputs(8) <= (inputs(205)) xor (inputs(51));
    layer0_outputs(9) <= (inputs(185)) or (inputs(172));
    layer0_outputs(10) <= (inputs(211)) or (inputs(72));
    layer0_outputs(11) <= (inputs(124)) and (inputs(78));
    layer0_outputs(12) <= not(inputs(171)) or (inputs(106));
    layer0_outputs(13) <= (inputs(130)) xor (inputs(148));
    layer0_outputs(14) <= not(inputs(41));
    layer0_outputs(15) <= (inputs(196)) or (inputs(143));
    layer0_outputs(16) <= not(inputs(170));
    layer0_outputs(17) <= (inputs(58)) xor (inputs(250));
    layer0_outputs(18) <= (inputs(34)) and not (inputs(77));
    layer0_outputs(19) <= inputs(18);
    layer0_outputs(20) <= (inputs(181)) and not (inputs(137));
    layer0_outputs(21) <= (inputs(87)) and not (inputs(95));
    layer0_outputs(22) <= not((inputs(111)) or (inputs(254)));
    layer0_outputs(23) <= inputs(8);
    layer0_outputs(24) <= inputs(85);
    layer0_outputs(25) <= not((inputs(39)) and (inputs(119)));
    layer0_outputs(26) <= not((inputs(223)) or (inputs(91)));
    layer0_outputs(27) <= not(inputs(106));
    layer0_outputs(28) <= not(inputs(232)) or (inputs(32));
    layer0_outputs(29) <= inputs(8);
    layer0_outputs(30) <= not(inputs(168)) or (inputs(28));
    layer0_outputs(31) <= not(inputs(195));
    layer0_outputs(32) <= (inputs(226)) and not (inputs(67));
    layer0_outputs(33) <= not(inputs(236));
    layer0_outputs(34) <= not(inputs(25)) or (inputs(223));
    layer0_outputs(35) <= (inputs(50)) and not (inputs(160));
    layer0_outputs(36) <= not((inputs(156)) or (inputs(116)));
    layer0_outputs(37) <= not(inputs(87));
    layer0_outputs(38) <= (inputs(151)) or (inputs(162));
    layer0_outputs(39) <= (inputs(229)) and (inputs(164));
    layer0_outputs(40) <= not(inputs(26));
    layer0_outputs(41) <= not((inputs(59)) or (inputs(130)));
    layer0_outputs(42) <= inputs(201);
    layer0_outputs(43) <= not((inputs(3)) or (inputs(192)));
    layer0_outputs(44) <= (inputs(185)) and not (inputs(33));
    layer0_outputs(45) <= '1';
    layer0_outputs(46) <= not(inputs(37));
    layer0_outputs(47) <= (inputs(248)) and not (inputs(184));
    layer0_outputs(48) <= not(inputs(105)) or (inputs(144));
    layer0_outputs(49) <= (inputs(131)) xor (inputs(11));
    layer0_outputs(50) <= inputs(127);
    layer0_outputs(51) <= (inputs(85)) or (inputs(189));
    layer0_outputs(52) <= not(inputs(98)) or (inputs(239));
    layer0_outputs(53) <= (inputs(44)) and not (inputs(192));
    layer0_outputs(54) <= not((inputs(73)) xor (inputs(151)));
    layer0_outputs(55) <= not(inputs(147));
    layer0_outputs(56) <= (inputs(20)) and not (inputs(255));
    layer0_outputs(57) <= '0';
    layer0_outputs(58) <= not(inputs(105)) or (inputs(238));
    layer0_outputs(59) <= not((inputs(68)) or (inputs(2)));
    layer0_outputs(60) <= (inputs(22)) and not (inputs(138));
    layer0_outputs(61) <= (inputs(80)) or (inputs(143));
    layer0_outputs(62) <= (inputs(207)) xor (inputs(89));
    layer0_outputs(63) <= inputs(102);
    layer0_outputs(64) <= not(inputs(254));
    layer0_outputs(65) <= not(inputs(11)) or (inputs(102));
    layer0_outputs(66) <= not(inputs(106)) or (inputs(109));
    layer0_outputs(67) <= (inputs(244)) and not (inputs(98));
    layer0_outputs(68) <= inputs(113);
    layer0_outputs(69) <= not(inputs(166)) or (inputs(225));
    layer0_outputs(70) <= not(inputs(24));
    layer0_outputs(71) <= inputs(90);
    layer0_outputs(72) <= inputs(108);
    layer0_outputs(73) <= (inputs(97)) and not (inputs(243));
    layer0_outputs(74) <= not(inputs(100));
    layer0_outputs(75) <= (inputs(203)) or (inputs(9));
    layer0_outputs(76) <= (inputs(117)) and not (inputs(227));
    layer0_outputs(77) <= inputs(10);
    layer0_outputs(78) <= not((inputs(221)) or (inputs(82)));
    layer0_outputs(79) <= not(inputs(30));
    layer0_outputs(80) <= (inputs(107)) and (inputs(36));
    layer0_outputs(81) <= not((inputs(125)) xor (inputs(172)));
    layer0_outputs(82) <= not((inputs(218)) xor (inputs(163)));
    layer0_outputs(83) <= not(inputs(146));
    layer0_outputs(84) <= inputs(37);
    layer0_outputs(85) <= (inputs(138)) and (inputs(90));
    layer0_outputs(86) <= not((inputs(141)) xor (inputs(93)));
    layer0_outputs(87) <= not(inputs(236));
    layer0_outputs(88) <= (inputs(214)) and (inputs(73));
    layer0_outputs(89) <= (inputs(26)) or (inputs(205));
    layer0_outputs(90) <= not((inputs(116)) xor (inputs(44)));
    layer0_outputs(91) <= inputs(14);
    layer0_outputs(92) <= (inputs(196)) and not (inputs(129));
    layer0_outputs(93) <= not((inputs(195)) and (inputs(145)));
    layer0_outputs(94) <= '1';
    layer0_outputs(95) <= (inputs(154)) xor (inputs(114));
    layer0_outputs(96) <= (inputs(5)) xor (inputs(143));
    layer0_outputs(97) <= not(inputs(76));
    layer0_outputs(98) <= (inputs(119)) and (inputs(100));
    layer0_outputs(99) <= (inputs(249)) xor (inputs(145));
    layer0_outputs(100) <= not(inputs(248)) or (inputs(254));
    layer0_outputs(101) <= not(inputs(6));
    layer0_outputs(102) <= not((inputs(0)) or (inputs(221)));
    layer0_outputs(103) <= not(inputs(246)) or (inputs(64));
    layer0_outputs(104) <= inputs(181);
    layer0_outputs(105) <= inputs(72);
    layer0_outputs(106) <= not(inputs(228)) or (inputs(1));
    layer0_outputs(107) <= (inputs(43)) and (inputs(109));
    layer0_outputs(108) <= not((inputs(207)) or (inputs(93)));
    layer0_outputs(109) <= inputs(24);
    layer0_outputs(110) <= (inputs(127)) or (inputs(17));
    layer0_outputs(111) <= inputs(65);
    layer0_outputs(112) <= not(inputs(22));
    layer0_outputs(113) <= (inputs(149)) or (inputs(6));
    layer0_outputs(114) <= inputs(8);
    layer0_outputs(115) <= (inputs(63)) or (inputs(128));
    layer0_outputs(116) <= (inputs(254)) or (inputs(226));
    layer0_outputs(117) <= (inputs(22)) and not (inputs(251));
    layer0_outputs(118) <= not(inputs(216));
    layer0_outputs(119) <= not(inputs(79));
    layer0_outputs(120) <= not(inputs(187)) or (inputs(28));
    layer0_outputs(121) <= (inputs(216)) xor (inputs(217));
    layer0_outputs(122) <= (inputs(139)) or (inputs(245));
    layer0_outputs(123) <= not((inputs(4)) or (inputs(165)));
    layer0_outputs(124) <= (inputs(2)) and not (inputs(239));
    layer0_outputs(125) <= not(inputs(91));
    layer0_outputs(126) <= not((inputs(193)) or (inputs(159)));
    layer0_outputs(127) <= not(inputs(92));
    layer0_outputs(128) <= not((inputs(191)) or (inputs(190)));
    layer0_outputs(129) <= not((inputs(49)) xor (inputs(1)));
    layer0_outputs(130) <= inputs(131);
    layer0_outputs(131) <= not((inputs(28)) xor (inputs(22)));
    layer0_outputs(132) <= inputs(113);
    layer0_outputs(133) <= inputs(228);
    layer0_outputs(134) <= (inputs(183)) and not (inputs(61));
    layer0_outputs(135) <= (inputs(156)) xor (inputs(122));
    layer0_outputs(136) <= not(inputs(105));
    layer0_outputs(137) <= (inputs(173)) xor (inputs(12));
    layer0_outputs(138) <= inputs(11);
    layer0_outputs(139) <= inputs(137);
    layer0_outputs(140) <= not(inputs(39)) or (inputs(162));
    layer0_outputs(141) <= not((inputs(254)) or (inputs(153)));
    layer0_outputs(142) <= (inputs(247)) xor (inputs(130));
    layer0_outputs(143) <= (inputs(203)) or (inputs(227));
    layer0_outputs(144) <= (inputs(81)) or (inputs(247));
    layer0_outputs(145) <= not((inputs(198)) or (inputs(14)));
    layer0_outputs(146) <= not(inputs(197)) or (inputs(161));
    layer0_outputs(147) <= not((inputs(217)) and (inputs(198)));
    layer0_outputs(148) <= not(inputs(177));
    layer0_outputs(149) <= (inputs(2)) xor (inputs(84));
    layer0_outputs(150) <= (inputs(101)) xor (inputs(125));
    layer0_outputs(151) <= not((inputs(255)) or (inputs(14)));
    layer0_outputs(152) <= inputs(41);
    layer0_outputs(153) <= (inputs(57)) and not (inputs(109));
    layer0_outputs(154) <= (inputs(96)) or (inputs(124));
    layer0_outputs(155) <= inputs(11);
    layer0_outputs(156) <= inputs(215);
    layer0_outputs(157) <= not((inputs(154)) or (inputs(110)));
    layer0_outputs(158) <= not(inputs(87));
    layer0_outputs(159) <= not((inputs(172)) xor (inputs(176)));
    layer0_outputs(160) <= (inputs(163)) or (inputs(47));
    layer0_outputs(161) <= not(inputs(83));
    layer0_outputs(162) <= not(inputs(113));
    layer0_outputs(163) <= not(inputs(98)) or (inputs(56));
    layer0_outputs(164) <= not(inputs(62)) or (inputs(11));
    layer0_outputs(165) <= (inputs(202)) xor (inputs(104));
    layer0_outputs(166) <= (inputs(161)) or (inputs(255));
    layer0_outputs(167) <= inputs(230);
    layer0_outputs(168) <= (inputs(84)) or (inputs(157));
    layer0_outputs(169) <= not(inputs(152));
    layer0_outputs(170) <= (inputs(225)) xor (inputs(103));
    layer0_outputs(171) <= inputs(90);
    layer0_outputs(172) <= not((inputs(213)) or (inputs(56)));
    layer0_outputs(173) <= not((inputs(47)) or (inputs(37)));
    layer0_outputs(174) <= (inputs(156)) and (inputs(100));
    layer0_outputs(175) <= (inputs(249)) xor (inputs(111));
    layer0_outputs(176) <= not((inputs(146)) or (inputs(149)));
    layer0_outputs(177) <= (inputs(167)) or (inputs(185));
    layer0_outputs(178) <= (inputs(121)) or (inputs(128));
    layer0_outputs(179) <= (inputs(181)) and not (inputs(34));
    layer0_outputs(180) <= inputs(232);
    layer0_outputs(181) <= not((inputs(148)) xor (inputs(2)));
    layer0_outputs(182) <= inputs(107);
    layer0_outputs(183) <= not((inputs(111)) xor (inputs(165)));
    layer0_outputs(184) <= inputs(52);
    layer0_outputs(185) <= not((inputs(163)) or (inputs(2)));
    layer0_outputs(186) <= inputs(103);
    layer0_outputs(187) <= inputs(197);
    layer0_outputs(188) <= not((inputs(142)) or (inputs(190)));
    layer0_outputs(189) <= (inputs(19)) or (inputs(94));
    layer0_outputs(190) <= inputs(94);
    layer0_outputs(191) <= '1';
    layer0_outputs(192) <= not(inputs(215));
    layer0_outputs(193) <= not(inputs(214));
    layer0_outputs(194) <= (inputs(254)) xor (inputs(122));
    layer0_outputs(195) <= inputs(76);
    layer0_outputs(196) <= (inputs(124)) xor (inputs(170));
    layer0_outputs(197) <= (inputs(60)) and (inputs(125));
    layer0_outputs(198) <= not((inputs(142)) or (inputs(119)));
    layer0_outputs(199) <= not((inputs(86)) and (inputs(203)));
    layer0_outputs(200) <= (inputs(235)) and not (inputs(65));
    layer0_outputs(201) <= not((inputs(42)) or (inputs(208)));
    layer0_outputs(202) <= (inputs(105)) or (inputs(72));
    layer0_outputs(203) <= not(inputs(26)) or (inputs(233));
    layer0_outputs(204) <= inputs(102);
    layer0_outputs(205) <= (inputs(226)) xor (inputs(74));
    layer0_outputs(206) <= inputs(68);
    layer0_outputs(207) <= (inputs(251)) or (inputs(151));
    layer0_outputs(208) <= not(inputs(200));
    layer0_outputs(209) <= not(inputs(92)) or (inputs(191));
    layer0_outputs(210) <= inputs(161);
    layer0_outputs(211) <= (inputs(107)) or (inputs(246));
    layer0_outputs(212) <= (inputs(115)) or (inputs(70));
    layer0_outputs(213) <= (inputs(244)) or (inputs(190));
    layer0_outputs(214) <= inputs(75);
    layer0_outputs(215) <= not(inputs(154)) or (inputs(78));
    layer0_outputs(216) <= not((inputs(156)) or (inputs(35)));
    layer0_outputs(217) <= not((inputs(252)) and (inputs(174)));
    layer0_outputs(218) <= (inputs(106)) and not (inputs(129));
    layer0_outputs(219) <= not(inputs(69)) or (inputs(55));
    layer0_outputs(220) <= inputs(203);
    layer0_outputs(221) <= not((inputs(52)) and (inputs(33)));
    layer0_outputs(222) <= (inputs(166)) and not (inputs(7));
    layer0_outputs(223) <= inputs(229);
    layer0_outputs(224) <= not(inputs(58)) or (inputs(230));
    layer0_outputs(225) <= (inputs(153)) and not (inputs(36));
    layer0_outputs(226) <= not((inputs(106)) xor (inputs(193)));
    layer0_outputs(227) <= inputs(238);
    layer0_outputs(228) <= not((inputs(44)) xor (inputs(82)));
    layer0_outputs(229) <= inputs(176);
    layer0_outputs(230) <= not((inputs(170)) xor (inputs(140)));
    layer0_outputs(231) <= not(inputs(191)) or (inputs(187));
    layer0_outputs(232) <= inputs(185);
    layer0_outputs(233) <= (inputs(102)) xor (inputs(67));
    layer0_outputs(234) <= inputs(145);
    layer0_outputs(235) <= not(inputs(20)) or (inputs(166));
    layer0_outputs(236) <= not((inputs(80)) or (inputs(151)));
    layer0_outputs(237) <= not((inputs(200)) xor (inputs(149)));
    layer0_outputs(238) <= (inputs(232)) and not (inputs(60));
    layer0_outputs(239) <= inputs(209);
    layer0_outputs(240) <= (inputs(220)) and not (inputs(128));
    layer0_outputs(241) <= not(inputs(177));
    layer0_outputs(242) <= not((inputs(116)) or (inputs(174)));
    layer0_outputs(243) <= (inputs(107)) xor (inputs(227));
    layer0_outputs(244) <= inputs(9);
    layer0_outputs(245) <= not(inputs(42));
    layer0_outputs(246) <= inputs(232);
    layer0_outputs(247) <= inputs(67);
    layer0_outputs(248) <= not((inputs(77)) or (inputs(187)));
    layer0_outputs(249) <= not(inputs(149));
    layer0_outputs(250) <= (inputs(77)) and (inputs(210));
    layer0_outputs(251) <= not(inputs(117));
    layer0_outputs(252) <= not(inputs(88)) or (inputs(177));
    layer0_outputs(253) <= inputs(88);
    layer0_outputs(254) <= not((inputs(216)) and (inputs(106)));
    layer0_outputs(255) <= (inputs(117)) and not (inputs(64));
    layer0_outputs(256) <= inputs(215);
    layer0_outputs(257) <= inputs(234);
    layer0_outputs(258) <= (inputs(246)) and not (inputs(128));
    layer0_outputs(259) <= (inputs(38)) xor (inputs(14));
    layer0_outputs(260) <= not(inputs(232)) or (inputs(113));
    layer0_outputs(261) <= not((inputs(164)) xor (inputs(174)));
    layer0_outputs(262) <= (inputs(52)) and not (inputs(141));
    layer0_outputs(263) <= (inputs(139)) xor (inputs(167));
    layer0_outputs(264) <= (inputs(147)) and not (inputs(240));
    layer0_outputs(265) <= not(inputs(12)) or (inputs(24));
    layer0_outputs(266) <= (inputs(236)) xor (inputs(219));
    layer0_outputs(267) <= not(inputs(167)) or (inputs(117));
    layer0_outputs(268) <= (inputs(231)) and not (inputs(0));
    layer0_outputs(269) <= (inputs(198)) or (inputs(219));
    layer0_outputs(270) <= not((inputs(89)) or (inputs(129)));
    layer0_outputs(271) <= not(inputs(31));
    layer0_outputs(272) <= (inputs(103)) or (inputs(191));
    layer0_outputs(273) <= not(inputs(92)) or (inputs(47));
    layer0_outputs(274) <= not((inputs(102)) or (inputs(101)));
    layer0_outputs(275) <= not((inputs(117)) or (inputs(228)));
    layer0_outputs(276) <= inputs(241);
    layer0_outputs(277) <= not(inputs(30));
    layer0_outputs(278) <= not(inputs(131)) or (inputs(240));
    layer0_outputs(279) <= inputs(180);
    layer0_outputs(280) <= not(inputs(33));
    layer0_outputs(281) <= inputs(210);
    layer0_outputs(282) <= not((inputs(128)) or (inputs(31)));
    layer0_outputs(283) <= not((inputs(131)) or (inputs(100)));
    layer0_outputs(284) <= (inputs(114)) or (inputs(14));
    layer0_outputs(285) <= not(inputs(231));
    layer0_outputs(286) <= (inputs(141)) xor (inputs(189));
    layer0_outputs(287) <= not(inputs(191));
    layer0_outputs(288) <= (inputs(152)) and not (inputs(18));
    layer0_outputs(289) <= (inputs(169)) or (inputs(115));
    layer0_outputs(290) <= inputs(124);
    layer0_outputs(291) <= (inputs(0)) and not (inputs(9));
    layer0_outputs(292) <= not(inputs(103));
    layer0_outputs(293) <= not(inputs(101));
    layer0_outputs(294) <= not(inputs(238));
    layer0_outputs(295) <= not(inputs(31));
    layer0_outputs(296) <= not(inputs(170));
    layer0_outputs(297) <= (inputs(244)) or (inputs(148));
    layer0_outputs(298) <= (inputs(175)) or (inputs(217));
    layer0_outputs(299) <= not((inputs(63)) or (inputs(148)));
    layer0_outputs(300) <= (inputs(123)) and not (inputs(56));
    layer0_outputs(301) <= not(inputs(239));
    layer0_outputs(302) <= inputs(98);
    layer0_outputs(303) <= not(inputs(166)) or (inputs(36));
    layer0_outputs(304) <= (inputs(162)) xor (inputs(66));
    layer0_outputs(305) <= (inputs(138)) or (inputs(49));
    layer0_outputs(306) <= inputs(74);
    layer0_outputs(307) <= inputs(71);
    layer0_outputs(308) <= inputs(245);
    layer0_outputs(309) <= (inputs(20)) xor (inputs(69));
    layer0_outputs(310) <= (inputs(159)) xor (inputs(115));
    layer0_outputs(311) <= not(inputs(106)) or (inputs(216));
    layer0_outputs(312) <= not(inputs(179)) or (inputs(152));
    layer0_outputs(313) <= inputs(26);
    layer0_outputs(314) <= not(inputs(90));
    layer0_outputs(315) <= not((inputs(139)) and (inputs(107)));
    layer0_outputs(316) <= (inputs(120)) and (inputs(229));
    layer0_outputs(317) <= inputs(107);
    layer0_outputs(318) <= (inputs(87)) and not (inputs(35));
    layer0_outputs(319) <= not(inputs(179));
    layer0_outputs(320) <= not(inputs(46));
    layer0_outputs(321) <= not((inputs(153)) or (inputs(208)));
    layer0_outputs(322) <= not(inputs(220));
    layer0_outputs(323) <= (inputs(248)) xor (inputs(100));
    layer0_outputs(324) <= (inputs(76)) or (inputs(5));
    layer0_outputs(325) <= not((inputs(105)) or (inputs(135)));
    layer0_outputs(326) <= inputs(139);
    layer0_outputs(327) <= '0';
    layer0_outputs(328) <= not((inputs(4)) or (inputs(136)));
    layer0_outputs(329) <= (inputs(158)) xor (inputs(206));
    layer0_outputs(330) <= not((inputs(55)) or (inputs(158)));
    layer0_outputs(331) <= not((inputs(158)) xor (inputs(244)));
    layer0_outputs(332) <= not(inputs(222)) or (inputs(160));
    layer0_outputs(333) <= (inputs(221)) or (inputs(35));
    layer0_outputs(334) <= inputs(58);
    layer0_outputs(335) <= (inputs(107)) xor (inputs(172));
    layer0_outputs(336) <= not(inputs(18)) or (inputs(160));
    layer0_outputs(337) <= (inputs(199)) xor (inputs(181));
    layer0_outputs(338) <= not(inputs(205)) or (inputs(14));
    layer0_outputs(339) <= (inputs(103)) and not (inputs(2));
    layer0_outputs(340) <= inputs(198);
    layer0_outputs(341) <= (inputs(91)) or (inputs(13));
    layer0_outputs(342) <= inputs(44);
    layer0_outputs(343) <= (inputs(232)) and not (inputs(45));
    layer0_outputs(344) <= inputs(113);
    layer0_outputs(345) <= not(inputs(83));
    layer0_outputs(346) <= (inputs(22)) xor (inputs(192));
    layer0_outputs(347) <= not((inputs(219)) or (inputs(115)));
    layer0_outputs(348) <= inputs(61);
    layer0_outputs(349) <= not(inputs(133));
    layer0_outputs(350) <= not((inputs(246)) and (inputs(59)));
    layer0_outputs(351) <= not((inputs(143)) or (inputs(60)));
    layer0_outputs(352) <= not((inputs(66)) or (inputs(27)));
    layer0_outputs(353) <= not(inputs(181));
    layer0_outputs(354) <= inputs(187);
    layer0_outputs(355) <= not((inputs(93)) xor (inputs(177)));
    layer0_outputs(356) <= (inputs(73)) xor (inputs(36));
    layer0_outputs(357) <= inputs(128);
    layer0_outputs(358) <= not(inputs(56));
    layer0_outputs(359) <= not((inputs(239)) xor (inputs(190)));
    layer0_outputs(360) <= not(inputs(122)) or (inputs(217));
    layer0_outputs(361) <= (inputs(71)) xor (inputs(221));
    layer0_outputs(362) <= not(inputs(74)) or (inputs(172));
    layer0_outputs(363) <= inputs(93);
    layer0_outputs(364) <= not((inputs(180)) xor (inputs(254)));
    layer0_outputs(365) <= (inputs(112)) or (inputs(73));
    layer0_outputs(366) <= not((inputs(143)) xor (inputs(52)));
    layer0_outputs(367) <= not(inputs(192));
    layer0_outputs(368) <= (inputs(63)) or (inputs(214));
    layer0_outputs(369) <= not((inputs(196)) or (inputs(160)));
    layer0_outputs(370) <= (inputs(245)) xor (inputs(193));
    layer0_outputs(371) <= (inputs(7)) xor (inputs(37));
    layer0_outputs(372) <= (inputs(173)) or (inputs(141));
    layer0_outputs(373) <= inputs(129);
    layer0_outputs(374) <= not((inputs(221)) xor (inputs(93)));
    layer0_outputs(375) <= (inputs(150)) or (inputs(47));
    layer0_outputs(376) <= not((inputs(24)) xor (inputs(249)));
    layer0_outputs(377) <= (inputs(192)) or (inputs(171));
    layer0_outputs(378) <= (inputs(137)) and (inputs(23));
    layer0_outputs(379) <= not((inputs(100)) or (inputs(156)));
    layer0_outputs(380) <= (inputs(187)) and not (inputs(5));
    layer0_outputs(381) <= not(inputs(166));
    layer0_outputs(382) <= not(inputs(197));
    layer0_outputs(383) <= not((inputs(7)) or (inputs(24)));
    layer0_outputs(384) <= (inputs(187)) or (inputs(38));
    layer0_outputs(385) <= (inputs(24)) and not (inputs(3));
    layer0_outputs(386) <= (inputs(103)) xor (inputs(129));
    layer0_outputs(387) <= not((inputs(199)) or (inputs(222)));
    layer0_outputs(388) <= (inputs(157)) and not (inputs(159));
    layer0_outputs(389) <= inputs(16);
    layer0_outputs(390) <= (inputs(211)) or (inputs(141));
    layer0_outputs(391) <= not((inputs(37)) or (inputs(219)));
    layer0_outputs(392) <= (inputs(253)) or (inputs(179));
    layer0_outputs(393) <= (inputs(143)) or (inputs(209));
    layer0_outputs(394) <= not((inputs(219)) or (inputs(215)));
    layer0_outputs(395) <= not(inputs(222)) or (inputs(15));
    layer0_outputs(396) <= not(inputs(168));
    layer0_outputs(397) <= (inputs(164)) or (inputs(123));
    layer0_outputs(398) <= '0';
    layer0_outputs(399) <= not(inputs(115));
    layer0_outputs(400) <= inputs(57);
    layer0_outputs(401) <= inputs(198);
    layer0_outputs(402) <= not((inputs(39)) xor (inputs(105)));
    layer0_outputs(403) <= not((inputs(147)) and (inputs(51)));
    layer0_outputs(404) <= (inputs(171)) or (inputs(164));
    layer0_outputs(405) <= inputs(34);
    layer0_outputs(406) <= not(inputs(102));
    layer0_outputs(407) <= not(inputs(142)) or (inputs(141));
    layer0_outputs(408) <= inputs(85);
    layer0_outputs(409) <= (inputs(66)) or (inputs(185));
    layer0_outputs(410) <= not(inputs(214));
    layer0_outputs(411) <= not(inputs(57));
    layer0_outputs(412) <= not((inputs(115)) xor (inputs(101)));
    layer0_outputs(413) <= (inputs(245)) and not (inputs(80));
    layer0_outputs(414) <= not((inputs(109)) or (inputs(28)));
    layer0_outputs(415) <= not(inputs(93));
    layer0_outputs(416) <= inputs(111);
    layer0_outputs(417) <= not(inputs(219));
    layer0_outputs(418) <= (inputs(172)) xor (inputs(34));
    layer0_outputs(419) <= inputs(97);
    layer0_outputs(420) <= not(inputs(136));
    layer0_outputs(421) <= inputs(67);
    layer0_outputs(422) <= (inputs(73)) xor (inputs(74));
    layer0_outputs(423) <= not(inputs(43)) or (inputs(35));
    layer0_outputs(424) <= not(inputs(122));
    layer0_outputs(425) <= (inputs(233)) and not (inputs(80));
    layer0_outputs(426) <= (inputs(181)) and not (inputs(29));
    layer0_outputs(427) <= (inputs(212)) and not (inputs(92));
    layer0_outputs(428) <= not((inputs(194)) xor (inputs(135)));
    layer0_outputs(429) <= not(inputs(73));
    layer0_outputs(430) <= (inputs(32)) or (inputs(209));
    layer0_outputs(431) <= (inputs(161)) or (inputs(165));
    layer0_outputs(432) <= not((inputs(37)) and (inputs(77)));
    layer0_outputs(433) <= (inputs(161)) or (inputs(147));
    layer0_outputs(434) <= inputs(246);
    layer0_outputs(435) <= (inputs(12)) xor (inputs(253));
    layer0_outputs(436) <= (inputs(151)) or (inputs(233));
    layer0_outputs(437) <= inputs(165);
    layer0_outputs(438) <= (inputs(180)) and not (inputs(18));
    layer0_outputs(439) <= (inputs(188)) or (inputs(19));
    layer0_outputs(440) <= not(inputs(118));
    layer0_outputs(441) <= not((inputs(4)) or (inputs(216)));
    layer0_outputs(442) <= (inputs(125)) or (inputs(205));
    layer0_outputs(443) <= not(inputs(14));
    layer0_outputs(444) <= not(inputs(100));
    layer0_outputs(445) <= (inputs(200)) and (inputs(168));
    layer0_outputs(446) <= not((inputs(158)) xor (inputs(234)));
    layer0_outputs(447) <= not((inputs(99)) xor (inputs(24)));
    layer0_outputs(448) <= inputs(45);
    layer0_outputs(449) <= inputs(162);
    layer0_outputs(450) <= not(inputs(221)) or (inputs(30));
    layer0_outputs(451) <= not(inputs(59));
    layer0_outputs(452) <= (inputs(157)) and not (inputs(11));
    layer0_outputs(453) <= (inputs(80)) and not (inputs(126));
    layer0_outputs(454) <= inputs(117);
    layer0_outputs(455) <= not(inputs(164));
    layer0_outputs(456) <= (inputs(223)) xor (inputs(213));
    layer0_outputs(457) <= not(inputs(221));
    layer0_outputs(458) <= (inputs(128)) and (inputs(86));
    layer0_outputs(459) <= inputs(168);
    layer0_outputs(460) <= not(inputs(230));
    layer0_outputs(461) <= not((inputs(214)) and (inputs(187)));
    layer0_outputs(462) <= '1';
    layer0_outputs(463) <= inputs(216);
    layer0_outputs(464) <= (inputs(120)) and not (inputs(19));
    layer0_outputs(465) <= inputs(135);
    layer0_outputs(466) <= not(inputs(165));
    layer0_outputs(467) <= not(inputs(215)) or (inputs(255));
    layer0_outputs(468) <= inputs(181);
    layer0_outputs(469) <= '1';
    layer0_outputs(470) <= inputs(129);
    layer0_outputs(471) <= not(inputs(158));
    layer0_outputs(472) <= not((inputs(149)) xor (inputs(1)));
    layer0_outputs(473) <= not(inputs(244)) or (inputs(242));
    layer0_outputs(474) <= (inputs(199)) and (inputs(104));
    layer0_outputs(475) <= not(inputs(113));
    layer0_outputs(476) <= not((inputs(130)) or (inputs(207)));
    layer0_outputs(477) <= inputs(129);
    layer0_outputs(478) <= inputs(54);
    layer0_outputs(479) <= not(inputs(44)) or (inputs(229));
    layer0_outputs(480) <= (inputs(150)) and not (inputs(30));
    layer0_outputs(481) <= not(inputs(48)) or (inputs(97));
    layer0_outputs(482) <= (inputs(163)) and not (inputs(50));
    layer0_outputs(483) <= not((inputs(181)) xor (inputs(199)));
    layer0_outputs(484) <= (inputs(209)) or (inputs(130));
    layer0_outputs(485) <= (inputs(131)) xor (inputs(100));
    layer0_outputs(486) <= (inputs(39)) and not (inputs(202));
    layer0_outputs(487) <= inputs(222);
    layer0_outputs(488) <= (inputs(53)) and not (inputs(171));
    layer0_outputs(489) <= inputs(103);
    layer0_outputs(490) <= inputs(144);
    layer0_outputs(491) <= not(inputs(99));
    layer0_outputs(492) <= (inputs(144)) and (inputs(122));
    layer0_outputs(493) <= not(inputs(33));
    layer0_outputs(494) <= not((inputs(10)) xor (inputs(54)));
    layer0_outputs(495) <= (inputs(139)) and not (inputs(235));
    layer0_outputs(496) <= not(inputs(103)) or (inputs(112));
    layer0_outputs(497) <= inputs(193);
    layer0_outputs(498) <= (inputs(204)) and not (inputs(71));
    layer0_outputs(499) <= not(inputs(40)) or (inputs(183));
    layer0_outputs(500) <= not(inputs(103)) or (inputs(225));
    layer0_outputs(501) <= (inputs(239)) or (inputs(147));
    layer0_outputs(502) <= (inputs(20)) or (inputs(254));
    layer0_outputs(503) <= (inputs(219)) xor (inputs(241));
    layer0_outputs(504) <= not(inputs(172));
    layer0_outputs(505) <= not((inputs(236)) xor (inputs(195)));
    layer0_outputs(506) <= not((inputs(49)) xor (inputs(71)));
    layer0_outputs(507) <= not((inputs(162)) or (inputs(50)));
    layer0_outputs(508) <= (inputs(134)) and not (inputs(81));
    layer0_outputs(509) <= (inputs(170)) xor (inputs(219));
    layer0_outputs(510) <= not(inputs(31));
    layer0_outputs(511) <= not(inputs(228)) or (inputs(128));
    layer0_outputs(512) <= inputs(11);
    layer0_outputs(513) <= not((inputs(110)) and (inputs(204)));
    layer0_outputs(514) <= not(inputs(233));
    layer0_outputs(515) <= not((inputs(71)) xor (inputs(60)));
    layer0_outputs(516) <= not((inputs(208)) or (inputs(254)));
    layer0_outputs(517) <= (inputs(93)) and not (inputs(179));
    layer0_outputs(518) <= '0';
    layer0_outputs(519) <= not(inputs(67)) or (inputs(114));
    layer0_outputs(520) <= not(inputs(230)) or (inputs(0));
    layer0_outputs(521) <= not((inputs(4)) or (inputs(228)));
    layer0_outputs(522) <= not((inputs(189)) and (inputs(168)));
    layer0_outputs(523) <= not(inputs(216)) or (inputs(47));
    layer0_outputs(524) <= (inputs(177)) and not (inputs(251));
    layer0_outputs(525) <= inputs(56);
    layer0_outputs(526) <= not(inputs(70)) or (inputs(187));
    layer0_outputs(527) <= inputs(178);
    layer0_outputs(528) <= (inputs(121)) or (inputs(78));
    layer0_outputs(529) <= (inputs(180)) and not (inputs(114));
    layer0_outputs(530) <= (inputs(67)) or (inputs(120));
    layer0_outputs(531) <= not((inputs(207)) or (inputs(218)));
    layer0_outputs(532) <= not((inputs(202)) or (inputs(177)));
    layer0_outputs(533) <= (inputs(17)) or (inputs(235));
    layer0_outputs(534) <= not(inputs(43));
    layer0_outputs(535) <= (inputs(131)) or (inputs(15));
    layer0_outputs(536) <= not(inputs(70));
    layer0_outputs(537) <= inputs(99);
    layer0_outputs(538) <= not(inputs(124));
    layer0_outputs(539) <= inputs(194);
    layer0_outputs(540) <= not(inputs(10)) or (inputs(163));
    layer0_outputs(541) <= not(inputs(27));
    layer0_outputs(542) <= (inputs(193)) and not (inputs(48));
    layer0_outputs(543) <= not((inputs(118)) or (inputs(236)));
    layer0_outputs(544) <= inputs(125);
    layer0_outputs(545) <= not((inputs(125)) or (inputs(255)));
    layer0_outputs(546) <= not((inputs(170)) or (inputs(57)));
    layer0_outputs(547) <= not(inputs(204));
    layer0_outputs(548) <= (inputs(253)) or (inputs(81));
    layer0_outputs(549) <= not((inputs(0)) or (inputs(232)));
    layer0_outputs(550) <= not((inputs(27)) xor (inputs(145)));
    layer0_outputs(551) <= not(inputs(155));
    layer0_outputs(552) <= not((inputs(102)) xor (inputs(109)));
    layer0_outputs(553) <= not((inputs(28)) xor (inputs(135)));
    layer0_outputs(554) <= not(inputs(73));
    layer0_outputs(555) <= '0';
    layer0_outputs(556) <= not(inputs(114));
    layer0_outputs(557) <= not(inputs(215));
    layer0_outputs(558) <= not((inputs(252)) xor (inputs(238)));
    layer0_outputs(559) <= not(inputs(233)) or (inputs(13));
    layer0_outputs(560) <= (inputs(27)) and not (inputs(115));
    layer0_outputs(561) <= not((inputs(170)) or (inputs(187)));
    layer0_outputs(562) <= (inputs(88)) or (inputs(253));
    layer0_outputs(563) <= not(inputs(229));
    layer0_outputs(564) <= not(inputs(169)) or (inputs(80));
    layer0_outputs(565) <= (inputs(27)) xor (inputs(31));
    layer0_outputs(566) <= inputs(40);
    layer0_outputs(567) <= not((inputs(72)) xor (inputs(53)));
    layer0_outputs(568) <= not(inputs(92)) or (inputs(121));
    layer0_outputs(569) <= not(inputs(122));
    layer0_outputs(570) <= inputs(32);
    layer0_outputs(571) <= (inputs(205)) or (inputs(151));
    layer0_outputs(572) <= inputs(234);
    layer0_outputs(573) <= (inputs(253)) or (inputs(209));
    layer0_outputs(574) <= not((inputs(129)) xor (inputs(115)));
    layer0_outputs(575) <= not(inputs(152)) or (inputs(203));
    layer0_outputs(576) <= (inputs(178)) xor (inputs(188));
    layer0_outputs(577) <= (inputs(250)) or (inputs(248));
    layer0_outputs(578) <= inputs(228);
    layer0_outputs(579) <= not((inputs(14)) xor (inputs(253)));
    layer0_outputs(580) <= (inputs(223)) or (inputs(205));
    layer0_outputs(581) <= not(inputs(21)) or (inputs(206));
    layer0_outputs(582) <= (inputs(72)) xor (inputs(6));
    layer0_outputs(583) <= (inputs(34)) xor (inputs(64));
    layer0_outputs(584) <= not((inputs(185)) or (inputs(130)));
    layer0_outputs(585) <= not(inputs(151));
    layer0_outputs(586) <= not((inputs(61)) xor (inputs(88)));
    layer0_outputs(587) <= inputs(199);
    layer0_outputs(588) <= inputs(229);
    layer0_outputs(589) <= not(inputs(187));
    layer0_outputs(590) <= inputs(84);
    layer0_outputs(591) <= '0';
    layer0_outputs(592) <= not((inputs(30)) xor (inputs(144)));
    layer0_outputs(593) <= not(inputs(90));
    layer0_outputs(594) <= inputs(179);
    layer0_outputs(595) <= inputs(180);
    layer0_outputs(596) <= not((inputs(86)) xor (inputs(106)));
    layer0_outputs(597) <= not((inputs(93)) or (inputs(206)));
    layer0_outputs(598) <= inputs(59);
    layer0_outputs(599) <= not((inputs(102)) or (inputs(207)));
    layer0_outputs(600) <= not(inputs(134));
    layer0_outputs(601) <= not((inputs(22)) xor (inputs(9)));
    layer0_outputs(602) <= (inputs(83)) or (inputs(95));
    layer0_outputs(603) <= not(inputs(133)) or (inputs(15));
    layer0_outputs(604) <= not(inputs(159));
    layer0_outputs(605) <= not(inputs(23)) or (inputs(129));
    layer0_outputs(606) <= '0';
    layer0_outputs(607) <= (inputs(101)) and (inputs(91));
    layer0_outputs(608) <= (inputs(195)) and (inputs(147));
    layer0_outputs(609) <= (inputs(25)) and (inputs(190));
    layer0_outputs(610) <= not((inputs(109)) or (inputs(4)));
    layer0_outputs(611) <= (inputs(16)) or (inputs(74));
    layer0_outputs(612) <= not((inputs(52)) and (inputs(170)));
    layer0_outputs(613) <= (inputs(60)) xor (inputs(22));
    layer0_outputs(614) <= (inputs(2)) or (inputs(191));
    layer0_outputs(615) <= not(inputs(100));
    layer0_outputs(616) <= inputs(86);
    layer0_outputs(617) <= (inputs(155)) or (inputs(130));
    layer0_outputs(618) <= inputs(99);
    layer0_outputs(619) <= (inputs(215)) and not (inputs(206));
    layer0_outputs(620) <= not(inputs(169)) or (inputs(94));
    layer0_outputs(621) <= inputs(114);
    layer0_outputs(622) <= not(inputs(161));
    layer0_outputs(623) <= inputs(194);
    layer0_outputs(624) <= inputs(129);
    layer0_outputs(625) <= (inputs(27)) or (inputs(48));
    layer0_outputs(626) <= inputs(218);
    layer0_outputs(627) <= not((inputs(37)) xor (inputs(183)));
    layer0_outputs(628) <= inputs(245);
    layer0_outputs(629) <= not(inputs(24));
    layer0_outputs(630) <= inputs(128);
    layer0_outputs(631) <= (inputs(38)) xor (inputs(73));
    layer0_outputs(632) <= not(inputs(166));
    layer0_outputs(633) <= inputs(120);
    layer0_outputs(634) <= not((inputs(10)) xor (inputs(94)));
    layer0_outputs(635) <= '0';
    layer0_outputs(636) <= inputs(14);
    layer0_outputs(637) <= not(inputs(228)) or (inputs(18));
    layer0_outputs(638) <= not(inputs(82));
    layer0_outputs(639) <= (inputs(54)) xor (inputs(243));
    layer0_outputs(640) <= inputs(27);
    layer0_outputs(641) <= (inputs(112)) xor (inputs(181));
    layer0_outputs(642) <= (inputs(97)) xor (inputs(146));
    layer0_outputs(643) <= (inputs(169)) or (inputs(45));
    layer0_outputs(644) <= not(inputs(67));
    layer0_outputs(645) <= (inputs(141)) and (inputs(174));
    layer0_outputs(646) <= not(inputs(199));
    layer0_outputs(647) <= (inputs(125)) or (inputs(160));
    layer0_outputs(648) <= not(inputs(176));
    layer0_outputs(649) <= inputs(212);
    layer0_outputs(650) <= (inputs(7)) and (inputs(25));
    layer0_outputs(651) <= (inputs(84)) xor (inputs(170));
    layer0_outputs(652) <= (inputs(101)) or (inputs(80));
    layer0_outputs(653) <= not((inputs(7)) xor (inputs(207)));
    layer0_outputs(654) <= not((inputs(165)) xor (inputs(167)));
    layer0_outputs(655) <= not((inputs(29)) xor (inputs(149)));
    layer0_outputs(656) <= inputs(77);
    layer0_outputs(657) <= (inputs(143)) xor (inputs(83));
    layer0_outputs(658) <= not(inputs(150));
    layer0_outputs(659) <= (inputs(142)) and not (inputs(121));
    layer0_outputs(660) <= not(inputs(104));
    layer0_outputs(661) <= (inputs(173)) or (inputs(78));
    layer0_outputs(662) <= (inputs(104)) and not (inputs(0));
    layer0_outputs(663) <= (inputs(92)) or (inputs(203));
    layer0_outputs(664) <= not((inputs(191)) and (inputs(221)));
    layer0_outputs(665) <= not((inputs(183)) or (inputs(128)));
    layer0_outputs(666) <= (inputs(218)) and not (inputs(78));
    layer0_outputs(667) <= not(inputs(103));
    layer0_outputs(668) <= inputs(193);
    layer0_outputs(669) <= (inputs(225)) xor (inputs(235));
    layer0_outputs(670) <= (inputs(43)) and not (inputs(237));
    layer0_outputs(671) <= not(inputs(75));
    layer0_outputs(672) <= not((inputs(44)) or (inputs(89)));
    layer0_outputs(673) <= not(inputs(122)) or (inputs(249));
    layer0_outputs(674) <= inputs(124);
    layer0_outputs(675) <= (inputs(49)) or (inputs(199));
    layer0_outputs(676) <= (inputs(88)) xor (inputs(13));
    layer0_outputs(677) <= '0';
    layer0_outputs(678) <= (inputs(99)) xor (inputs(246));
    layer0_outputs(679) <= (inputs(66)) or (inputs(252));
    layer0_outputs(680) <= inputs(9);
    layer0_outputs(681) <= not((inputs(15)) or (inputs(43)));
    layer0_outputs(682) <= not((inputs(175)) or (inputs(88)));
    layer0_outputs(683) <= inputs(209);
    layer0_outputs(684) <= not((inputs(174)) or (inputs(148)));
    layer0_outputs(685) <= (inputs(136)) and not (inputs(147));
    layer0_outputs(686) <= (inputs(240)) and not (inputs(35));
    layer0_outputs(687) <= not(inputs(126));
    layer0_outputs(688) <= not(inputs(80)) or (inputs(38));
    layer0_outputs(689) <= inputs(98);
    layer0_outputs(690) <= inputs(91);
    layer0_outputs(691) <= (inputs(21)) or (inputs(194));
    layer0_outputs(692) <= inputs(104);
    layer0_outputs(693) <= inputs(99);
    layer0_outputs(694) <= not(inputs(234));
    layer0_outputs(695) <= not(inputs(90)) or (inputs(217));
    layer0_outputs(696) <= (inputs(34)) or (inputs(79));
    layer0_outputs(697) <= (inputs(59)) and (inputs(233));
    layer0_outputs(698) <= inputs(109);
    layer0_outputs(699) <= (inputs(89)) and not (inputs(252));
    layer0_outputs(700) <= not((inputs(27)) and (inputs(21)));
    layer0_outputs(701) <= inputs(107);
    layer0_outputs(702) <= inputs(213);
    layer0_outputs(703) <= not((inputs(193)) xor (inputs(251)));
    layer0_outputs(704) <= not((inputs(197)) xor (inputs(192)));
    layer0_outputs(705) <= (inputs(14)) or (inputs(116));
    layer0_outputs(706) <= (inputs(41)) or (inputs(173));
    layer0_outputs(707) <= not(inputs(129));
    layer0_outputs(708) <= not(inputs(36)) or (inputs(203));
    layer0_outputs(709) <= not((inputs(121)) or (inputs(30)));
    layer0_outputs(710) <= not((inputs(48)) or (inputs(144)));
    layer0_outputs(711) <= (inputs(231)) and not (inputs(238));
    layer0_outputs(712) <= (inputs(146)) or (inputs(76));
    layer0_outputs(713) <= (inputs(255)) and not (inputs(15));
    layer0_outputs(714) <= not((inputs(0)) or (inputs(172)));
    layer0_outputs(715) <= (inputs(173)) and (inputs(139));
    layer0_outputs(716) <= inputs(88);
    layer0_outputs(717) <= '1';
    layer0_outputs(718) <= (inputs(5)) and not (inputs(113));
    layer0_outputs(719) <= (inputs(227)) and not (inputs(89));
    layer0_outputs(720) <= not(inputs(242));
    layer0_outputs(721) <= inputs(228);
    layer0_outputs(722) <= not((inputs(144)) or (inputs(174)));
    layer0_outputs(723) <= (inputs(24)) and not (inputs(129));
    layer0_outputs(724) <= not((inputs(209)) or (inputs(1)));
    layer0_outputs(725) <= (inputs(86)) xor (inputs(176));
    layer0_outputs(726) <= (inputs(74)) xor (inputs(42));
    layer0_outputs(727) <= (inputs(165)) and not (inputs(2));
    layer0_outputs(728) <= inputs(25);
    layer0_outputs(729) <= inputs(52);
    layer0_outputs(730) <= not(inputs(188)) or (inputs(109));
    layer0_outputs(731) <= (inputs(72)) and not (inputs(19));
    layer0_outputs(732) <= not((inputs(98)) or (inputs(244)));
    layer0_outputs(733) <= not(inputs(7));
    layer0_outputs(734) <= not(inputs(254));
    layer0_outputs(735) <= (inputs(85)) and not (inputs(78));
    layer0_outputs(736) <= (inputs(194)) and not (inputs(97));
    layer0_outputs(737) <= inputs(105);
    layer0_outputs(738) <= not(inputs(65)) or (inputs(6));
    layer0_outputs(739) <= (inputs(4)) and (inputs(232));
    layer0_outputs(740) <= not(inputs(236));
    layer0_outputs(741) <= (inputs(202)) and not (inputs(34));
    layer0_outputs(742) <= (inputs(172)) and not (inputs(37));
    layer0_outputs(743) <= (inputs(69)) or (inputs(127));
    layer0_outputs(744) <= not((inputs(23)) xor (inputs(211)));
    layer0_outputs(745) <= not(inputs(104));
    layer0_outputs(746) <= not(inputs(147));
    layer0_outputs(747) <= (inputs(173)) or (inputs(96));
    layer0_outputs(748) <= (inputs(115)) or (inputs(8));
    layer0_outputs(749) <= not((inputs(51)) or (inputs(117)));
    layer0_outputs(750) <= not(inputs(120)) or (inputs(31));
    layer0_outputs(751) <= (inputs(167)) xor (inputs(164));
    layer0_outputs(752) <= inputs(226);
    layer0_outputs(753) <= (inputs(8)) and not (inputs(182));
    layer0_outputs(754) <= (inputs(171)) and not (inputs(81));
    layer0_outputs(755) <= not(inputs(77));
    layer0_outputs(756) <= (inputs(198)) and not (inputs(250));
    layer0_outputs(757) <= (inputs(204)) or (inputs(244));
    layer0_outputs(758) <= not(inputs(91));
    layer0_outputs(759) <= (inputs(25)) and not (inputs(164));
    layer0_outputs(760) <= (inputs(148)) and not (inputs(12));
    layer0_outputs(761) <= not((inputs(142)) xor (inputs(79)));
    layer0_outputs(762) <= inputs(197);
    layer0_outputs(763) <= not(inputs(136));
    layer0_outputs(764) <= (inputs(74)) and not (inputs(23));
    layer0_outputs(765) <= inputs(49);
    layer0_outputs(766) <= not((inputs(171)) xor (inputs(233)));
    layer0_outputs(767) <= not(inputs(170)) or (inputs(146));
    layer0_outputs(768) <= inputs(153);
    layer0_outputs(769) <= not(inputs(143));
    layer0_outputs(770) <= (inputs(169)) xor (inputs(246));
    layer0_outputs(771) <= not(inputs(66));
    layer0_outputs(772) <= not(inputs(9)) or (inputs(192));
    layer0_outputs(773) <= not(inputs(54));
    layer0_outputs(774) <= not((inputs(51)) xor (inputs(10)));
    layer0_outputs(775) <= inputs(226);
    layer0_outputs(776) <= not(inputs(82));
    layer0_outputs(777) <= (inputs(113)) and (inputs(41));
    layer0_outputs(778) <= not(inputs(76)) or (inputs(223));
    layer0_outputs(779) <= not(inputs(230));
    layer0_outputs(780) <= inputs(1);
    layer0_outputs(781) <= (inputs(137)) or (inputs(158));
    layer0_outputs(782) <= (inputs(160)) or (inputs(48));
    layer0_outputs(783) <= not((inputs(124)) xor (inputs(106)));
    layer0_outputs(784) <= inputs(10);
    layer0_outputs(785) <= not(inputs(36));
    layer0_outputs(786) <= inputs(92);
    layer0_outputs(787) <= not(inputs(247));
    layer0_outputs(788) <= (inputs(223)) or (inputs(218));
    layer0_outputs(789) <= (inputs(14)) and not (inputs(28));
    layer0_outputs(790) <= not(inputs(183)) or (inputs(111));
    layer0_outputs(791) <= (inputs(140)) xor (inputs(206));
    layer0_outputs(792) <= (inputs(116)) xor (inputs(140));
    layer0_outputs(793) <= not((inputs(177)) and (inputs(245)));
    layer0_outputs(794) <= (inputs(89)) or (inputs(224));
    layer0_outputs(795) <= not(inputs(232)) or (inputs(140));
    layer0_outputs(796) <= not(inputs(46)) or (inputs(80));
    layer0_outputs(797) <= not((inputs(51)) or (inputs(111)));
    layer0_outputs(798) <= (inputs(52)) or (inputs(127));
    layer0_outputs(799) <= inputs(54);
    layer0_outputs(800) <= not((inputs(15)) or (inputs(226)));
    layer0_outputs(801) <= (inputs(218)) and (inputs(232));
    layer0_outputs(802) <= (inputs(253)) or (inputs(238));
    layer0_outputs(803) <= (inputs(57)) or (inputs(92));
    layer0_outputs(804) <= not(inputs(68)) or (inputs(233));
    layer0_outputs(805) <= not((inputs(187)) xor (inputs(74)));
    layer0_outputs(806) <= inputs(106);
    layer0_outputs(807) <= inputs(82);
    layer0_outputs(808) <= '0';
    layer0_outputs(809) <= not(inputs(84));
    layer0_outputs(810) <= (inputs(56)) and not (inputs(250));
    layer0_outputs(811) <= not(inputs(173));
    layer0_outputs(812) <= (inputs(215)) and (inputs(120));
    layer0_outputs(813) <= not((inputs(202)) xor (inputs(116)));
    layer0_outputs(814) <= not((inputs(70)) xor (inputs(85)));
    layer0_outputs(815) <= not(inputs(174)) or (inputs(145));
    layer0_outputs(816) <= (inputs(0)) xor (inputs(156));
    layer0_outputs(817) <= inputs(124);
    layer0_outputs(818) <= '1';
    layer0_outputs(819) <= (inputs(35)) and (inputs(139));
    layer0_outputs(820) <= not((inputs(190)) xor (inputs(2)));
    layer0_outputs(821) <= (inputs(220)) or (inputs(127));
    layer0_outputs(822) <= not((inputs(120)) or (inputs(76)));
    layer0_outputs(823) <= not(inputs(203));
    layer0_outputs(824) <= not((inputs(216)) xor (inputs(243)));
    layer0_outputs(825) <= (inputs(146)) or (inputs(145));
    layer0_outputs(826) <= not(inputs(152)) or (inputs(15));
    layer0_outputs(827) <= not((inputs(138)) or (inputs(65)));
    layer0_outputs(828) <= not((inputs(204)) xor (inputs(105)));
    layer0_outputs(829) <= (inputs(42)) or (inputs(62));
    layer0_outputs(830) <= (inputs(135)) and not (inputs(65));
    layer0_outputs(831) <= (inputs(43)) and not (inputs(230));
    layer0_outputs(832) <= inputs(40);
    layer0_outputs(833) <= inputs(139);
    layer0_outputs(834) <= not(inputs(232));
    layer0_outputs(835) <= (inputs(228)) or (inputs(0));
    layer0_outputs(836) <= not(inputs(53));
    layer0_outputs(837) <= (inputs(245)) and not (inputs(2));
    layer0_outputs(838) <= not(inputs(94)) or (inputs(90));
    layer0_outputs(839) <= inputs(145);
    layer0_outputs(840) <= inputs(93);
    layer0_outputs(841) <= (inputs(159)) and not (inputs(14));
    layer0_outputs(842) <= not((inputs(196)) and (inputs(22)));
    layer0_outputs(843) <= not((inputs(135)) or (inputs(232)));
    layer0_outputs(844) <= not(inputs(192));
    layer0_outputs(845) <= (inputs(171)) and not (inputs(70));
    layer0_outputs(846) <= (inputs(32)) or (inputs(121));
    layer0_outputs(847) <= (inputs(205)) and not (inputs(35));
    layer0_outputs(848) <= not((inputs(17)) or (inputs(148)));
    layer0_outputs(849) <= inputs(220);
    layer0_outputs(850) <= (inputs(14)) or (inputs(156));
    layer0_outputs(851) <= not((inputs(33)) or (inputs(137)));
    layer0_outputs(852) <= not((inputs(205)) xor (inputs(128)));
    layer0_outputs(853) <= (inputs(248)) xor (inputs(30));
    layer0_outputs(854) <= (inputs(41)) xor (inputs(29));
    layer0_outputs(855) <= not(inputs(103)) or (inputs(176));
    layer0_outputs(856) <= (inputs(28)) or (inputs(34));
    layer0_outputs(857) <= not((inputs(177)) or (inputs(127)));
    layer0_outputs(858) <= inputs(224);
    layer0_outputs(859) <= inputs(23);
    layer0_outputs(860) <= (inputs(73)) xor (inputs(23));
    layer0_outputs(861) <= (inputs(123)) xor (inputs(154));
    layer0_outputs(862) <= (inputs(143)) or (inputs(132));
    layer0_outputs(863) <= not((inputs(150)) xor (inputs(156)));
    layer0_outputs(864) <= not(inputs(10));
    layer0_outputs(865) <= not(inputs(221)) or (inputs(230));
    layer0_outputs(866) <= (inputs(124)) and not (inputs(71));
    layer0_outputs(867) <= (inputs(66)) xor (inputs(176));
    layer0_outputs(868) <= (inputs(58)) or (inputs(44));
    layer0_outputs(869) <= not((inputs(104)) or (inputs(47)));
    layer0_outputs(870) <= not(inputs(227));
    layer0_outputs(871) <= (inputs(177)) and not (inputs(63));
    layer0_outputs(872) <= inputs(80);
    layer0_outputs(873) <= (inputs(77)) or (inputs(113));
    layer0_outputs(874) <= not(inputs(210));
    layer0_outputs(875) <= (inputs(238)) or (inputs(39));
    layer0_outputs(876) <= not((inputs(236)) or (inputs(131)));
    layer0_outputs(877) <= inputs(133);
    layer0_outputs(878) <= inputs(144);
    layer0_outputs(879) <= (inputs(17)) or (inputs(241));
    layer0_outputs(880) <= (inputs(217)) xor (inputs(80));
    layer0_outputs(881) <= not(inputs(227)) or (inputs(159));
    layer0_outputs(882) <= (inputs(95)) xor (inputs(167));
    layer0_outputs(883) <= inputs(26);
    layer0_outputs(884) <= not((inputs(20)) or (inputs(192)));
    layer0_outputs(885) <= (inputs(62)) or (inputs(62));
    layer0_outputs(886) <= not(inputs(225));
    layer0_outputs(887) <= not((inputs(102)) or (inputs(235)));
    layer0_outputs(888) <= (inputs(111)) and (inputs(193));
    layer0_outputs(889) <= inputs(123);
    layer0_outputs(890) <= not((inputs(211)) xor (inputs(209)));
    layer0_outputs(891) <= not(inputs(171));
    layer0_outputs(892) <= inputs(36);
    layer0_outputs(893) <= inputs(176);
    layer0_outputs(894) <= not(inputs(122));
    layer0_outputs(895) <= (inputs(208)) xor (inputs(249));
    layer0_outputs(896) <= (inputs(6)) or (inputs(47));
    layer0_outputs(897) <= not((inputs(139)) xor (inputs(188)));
    layer0_outputs(898) <= not((inputs(216)) or (inputs(207)));
    layer0_outputs(899) <= not((inputs(34)) xor (inputs(176)));
    layer0_outputs(900) <= (inputs(139)) and not (inputs(243));
    layer0_outputs(901) <= inputs(169);
    layer0_outputs(902) <= (inputs(199)) and not (inputs(62));
    layer0_outputs(903) <= not(inputs(102));
    layer0_outputs(904) <= (inputs(28)) and (inputs(76));
    layer0_outputs(905) <= not((inputs(132)) xor (inputs(50)));
    layer0_outputs(906) <= not((inputs(216)) xor (inputs(168)));
    layer0_outputs(907) <= (inputs(248)) and not (inputs(125));
    layer0_outputs(908) <= (inputs(66)) or (inputs(241));
    layer0_outputs(909) <= not((inputs(3)) or (inputs(220)));
    layer0_outputs(910) <= (inputs(235)) and not (inputs(157));
    layer0_outputs(911) <= inputs(23);
    layer0_outputs(912) <= inputs(251);
    layer0_outputs(913) <= not(inputs(74));
    layer0_outputs(914) <= not(inputs(45));
    layer0_outputs(915) <= not(inputs(24));
    layer0_outputs(916) <= not(inputs(29));
    layer0_outputs(917) <= (inputs(148)) or (inputs(172));
    layer0_outputs(918) <= inputs(8);
    layer0_outputs(919) <= not((inputs(52)) xor (inputs(3)));
    layer0_outputs(920) <= not((inputs(88)) and (inputs(121)));
    layer0_outputs(921) <= inputs(121);
    layer0_outputs(922) <= not(inputs(163)) or (inputs(150));
    layer0_outputs(923) <= not((inputs(12)) or (inputs(47)));
    layer0_outputs(924) <= inputs(206);
    layer0_outputs(925) <= not((inputs(217)) xor (inputs(193)));
    layer0_outputs(926) <= not((inputs(121)) or (inputs(116)));
    layer0_outputs(927) <= not(inputs(44)) or (inputs(164));
    layer0_outputs(928) <= (inputs(194)) or (inputs(28));
    layer0_outputs(929) <= not(inputs(169));
    layer0_outputs(930) <= (inputs(251)) xor (inputs(9));
    layer0_outputs(931) <= (inputs(239)) xor (inputs(45));
    layer0_outputs(932) <= inputs(114);
    layer0_outputs(933) <= not(inputs(101)) or (inputs(140));
    layer0_outputs(934) <= (inputs(165)) xor (inputs(46));
    layer0_outputs(935) <= not(inputs(114));
    layer0_outputs(936) <= not((inputs(132)) or (inputs(241)));
    layer0_outputs(937) <= (inputs(33)) and (inputs(71));
    layer0_outputs(938) <= (inputs(130)) or (inputs(36));
    layer0_outputs(939) <= not(inputs(249)) or (inputs(172));
    layer0_outputs(940) <= not((inputs(119)) and (inputs(8)));
    layer0_outputs(941) <= inputs(7);
    layer0_outputs(942) <= (inputs(0)) and (inputs(136));
    layer0_outputs(943) <= inputs(226);
    layer0_outputs(944) <= not(inputs(166)) or (inputs(16));
    layer0_outputs(945) <= not(inputs(249));
    layer0_outputs(946) <= (inputs(17)) xor (inputs(192));
    layer0_outputs(947) <= not(inputs(157)) or (inputs(87));
    layer0_outputs(948) <= inputs(142);
    layer0_outputs(949) <= not(inputs(83));
    layer0_outputs(950) <= not((inputs(209)) or (inputs(92)));
    layer0_outputs(951) <= inputs(57);
    layer0_outputs(952) <= not(inputs(71)) or (inputs(251));
    layer0_outputs(953) <= (inputs(4)) or (inputs(183));
    layer0_outputs(954) <= (inputs(94)) and not (inputs(106));
    layer0_outputs(955) <= not(inputs(224)) or (inputs(16));
    layer0_outputs(956) <= (inputs(65)) or (inputs(203));
    layer0_outputs(957) <= (inputs(254)) or (inputs(245));
    layer0_outputs(958) <= not((inputs(8)) and (inputs(5)));
    layer0_outputs(959) <= (inputs(140)) or (inputs(142));
    layer0_outputs(960) <= '1';
    layer0_outputs(961) <= (inputs(46)) xor (inputs(243));
    layer0_outputs(962) <= (inputs(111)) or (inputs(17));
    layer0_outputs(963) <= (inputs(20)) or (inputs(157));
    layer0_outputs(964) <= (inputs(77)) and (inputs(192));
    layer0_outputs(965) <= (inputs(47)) and (inputs(55));
    layer0_outputs(966) <= (inputs(62)) and not (inputs(193));
    layer0_outputs(967) <= (inputs(0)) xor (inputs(171));
    layer0_outputs(968) <= not(inputs(50)) or (inputs(214));
    layer0_outputs(969) <= inputs(9);
    layer0_outputs(970) <= not((inputs(60)) xor (inputs(51)));
    layer0_outputs(971) <= (inputs(100)) or (inputs(205));
    layer0_outputs(972) <= not(inputs(126));
    layer0_outputs(973) <= inputs(29);
    layer0_outputs(974) <= (inputs(237)) or (inputs(155));
    layer0_outputs(975) <= not((inputs(245)) xor (inputs(162)));
    layer0_outputs(976) <= inputs(135);
    layer0_outputs(977) <= not(inputs(216));
    layer0_outputs(978) <= (inputs(215)) and not (inputs(238));
    layer0_outputs(979) <= inputs(177);
    layer0_outputs(980) <= not(inputs(119));
    layer0_outputs(981) <= not((inputs(25)) xor (inputs(83)));
    layer0_outputs(982) <= not((inputs(87)) xor (inputs(102)));
    layer0_outputs(983) <= not(inputs(106));
    layer0_outputs(984) <= not(inputs(68));
    layer0_outputs(985) <= not(inputs(179));
    layer0_outputs(986) <= not(inputs(105));
    layer0_outputs(987) <= not(inputs(72)) or (inputs(17));
    layer0_outputs(988) <= not(inputs(135)) or (inputs(239));
    layer0_outputs(989) <= inputs(91);
    layer0_outputs(990) <= (inputs(127)) and not (inputs(49));
    layer0_outputs(991) <= not((inputs(235)) xor (inputs(192)));
    layer0_outputs(992) <= not(inputs(170));
    layer0_outputs(993) <= not(inputs(196));
    layer0_outputs(994) <= not(inputs(250));
    layer0_outputs(995) <= (inputs(209)) or (inputs(97));
    layer0_outputs(996) <= not((inputs(129)) xor (inputs(100)));
    layer0_outputs(997) <= not(inputs(253));
    layer0_outputs(998) <= not((inputs(150)) or (inputs(64)));
    layer0_outputs(999) <= not((inputs(117)) or (inputs(244)));
    layer0_outputs(1000) <= not(inputs(85)) or (inputs(193));
    layer0_outputs(1001) <= inputs(87);
    layer0_outputs(1002) <= (inputs(243)) or (inputs(14));
    layer0_outputs(1003) <= not((inputs(155)) xor (inputs(137)));
    layer0_outputs(1004) <= not(inputs(30)) or (inputs(135));
    layer0_outputs(1005) <= (inputs(15)) and not (inputs(97));
    layer0_outputs(1006) <= (inputs(105)) or (inputs(223));
    layer0_outputs(1007) <= (inputs(25)) or (inputs(48));
    layer0_outputs(1008) <= (inputs(0)) xor (inputs(183));
    layer0_outputs(1009) <= (inputs(73)) and not (inputs(81));
    layer0_outputs(1010) <= inputs(35);
    layer0_outputs(1011) <= not((inputs(82)) or (inputs(68)));
    layer0_outputs(1012) <= (inputs(45)) and not (inputs(227));
    layer0_outputs(1013) <= (inputs(18)) and not (inputs(81));
    layer0_outputs(1014) <= not(inputs(185)) or (inputs(163));
    layer0_outputs(1015) <= not(inputs(53)) or (inputs(62));
    layer0_outputs(1016) <= not(inputs(234));
    layer0_outputs(1017) <= not((inputs(223)) or (inputs(201)));
    layer0_outputs(1018) <= not(inputs(247)) or (inputs(57));
    layer0_outputs(1019) <= not(inputs(79));
    layer0_outputs(1020) <= not((inputs(247)) and (inputs(219)));
    layer0_outputs(1021) <= not((inputs(185)) and (inputs(206)));
    layer0_outputs(1022) <= (inputs(104)) and not (inputs(141));
    layer0_outputs(1023) <= inputs(245);
    layer0_outputs(1024) <= not((inputs(143)) or (inputs(63)));
    layer0_outputs(1025) <= (inputs(8)) and not (inputs(29));
    layer0_outputs(1026) <= (inputs(96)) and not (inputs(57));
    layer0_outputs(1027) <= inputs(36);
    layer0_outputs(1028) <= not((inputs(124)) and (inputs(48)));
    layer0_outputs(1029) <= not((inputs(237)) or (inputs(198)));
    layer0_outputs(1030) <= not(inputs(181));
    layer0_outputs(1031) <= not(inputs(229)) or (inputs(121));
    layer0_outputs(1032) <= not(inputs(158));
    layer0_outputs(1033) <= (inputs(91)) or (inputs(92));
    layer0_outputs(1034) <= inputs(166);
    layer0_outputs(1035) <= not(inputs(28));
    layer0_outputs(1036) <= not((inputs(32)) or (inputs(27)));
    layer0_outputs(1037) <= not((inputs(202)) or (inputs(239)));
    layer0_outputs(1038) <= inputs(164);
    layer0_outputs(1039) <= (inputs(25)) and not (inputs(177));
    layer0_outputs(1040) <= not(inputs(118)) or (inputs(137));
    layer0_outputs(1041) <= not(inputs(170)) or (inputs(30));
    layer0_outputs(1042) <= not(inputs(30));
    layer0_outputs(1043) <= (inputs(99)) and not (inputs(5));
    layer0_outputs(1044) <= (inputs(85)) or (inputs(22));
    layer0_outputs(1045) <= (inputs(124)) and not (inputs(46));
    layer0_outputs(1046) <= not(inputs(125)) or (inputs(109));
    layer0_outputs(1047) <= not(inputs(63));
    layer0_outputs(1048) <= not((inputs(177)) or (inputs(178)));
    layer0_outputs(1049) <= (inputs(233)) and not (inputs(111));
    layer0_outputs(1050) <= (inputs(190)) and not (inputs(42));
    layer0_outputs(1051) <= not(inputs(7)) or (inputs(172));
    layer0_outputs(1052) <= not(inputs(224));
    layer0_outputs(1053) <= not(inputs(10));
    layer0_outputs(1054) <= inputs(8);
    layer0_outputs(1055) <= not((inputs(219)) xor (inputs(202)));
    layer0_outputs(1056) <= not(inputs(91));
    layer0_outputs(1057) <= inputs(121);
    layer0_outputs(1058) <= not(inputs(239)) or (inputs(180));
    layer0_outputs(1059) <= not((inputs(157)) xor (inputs(102)));
    layer0_outputs(1060) <= (inputs(137)) and not (inputs(160));
    layer0_outputs(1061) <= not((inputs(72)) xor (inputs(42)));
    layer0_outputs(1062) <= (inputs(116)) xor (inputs(231));
    layer0_outputs(1063) <= not((inputs(199)) xor (inputs(147)));
    layer0_outputs(1064) <= (inputs(107)) and not (inputs(3));
    layer0_outputs(1065) <= not((inputs(77)) or (inputs(6)));
    layer0_outputs(1066) <= not((inputs(126)) xor (inputs(248)));
    layer0_outputs(1067) <= (inputs(29)) xor (inputs(196));
    layer0_outputs(1068) <= (inputs(125)) and not (inputs(220));
    layer0_outputs(1069) <= not((inputs(50)) and (inputs(240)));
    layer0_outputs(1070) <= not(inputs(58));
    layer0_outputs(1071) <= not(inputs(146)) or (inputs(94));
    layer0_outputs(1072) <= not(inputs(89));
    layer0_outputs(1073) <= inputs(199);
    layer0_outputs(1074) <= not((inputs(181)) and (inputs(0)));
    layer0_outputs(1075) <= not(inputs(93));
    layer0_outputs(1076) <= inputs(239);
    layer0_outputs(1077) <= not((inputs(139)) xor (inputs(62)));
    layer0_outputs(1078) <= (inputs(8)) or (inputs(161));
    layer0_outputs(1079) <= not(inputs(234));
    layer0_outputs(1080) <= not((inputs(219)) xor (inputs(49)));
    layer0_outputs(1081) <= (inputs(140)) xor (inputs(250));
    layer0_outputs(1082) <= inputs(135);
    layer0_outputs(1083) <= not(inputs(57));
    layer0_outputs(1084) <= not(inputs(193));
    layer0_outputs(1085) <= (inputs(176)) xor (inputs(180));
    layer0_outputs(1086) <= not((inputs(240)) or (inputs(75)));
    layer0_outputs(1087) <= (inputs(30)) and not (inputs(178));
    layer0_outputs(1088) <= not(inputs(214));
    layer0_outputs(1089) <= not((inputs(200)) or (inputs(37)));
    layer0_outputs(1090) <= not((inputs(254)) or (inputs(208)));
    layer0_outputs(1091) <= inputs(9);
    layer0_outputs(1092) <= not(inputs(82));
    layer0_outputs(1093) <= inputs(193);
    layer0_outputs(1094) <= not(inputs(245)) or (inputs(92));
    layer0_outputs(1095) <= not(inputs(37)) or (inputs(113));
    layer0_outputs(1096) <= (inputs(4)) or (inputs(8));
    layer0_outputs(1097) <= not((inputs(44)) xor (inputs(47)));
    layer0_outputs(1098) <= inputs(163);
    layer0_outputs(1099) <= (inputs(203)) and not (inputs(9));
    layer0_outputs(1100) <= not((inputs(81)) and (inputs(55)));
    layer0_outputs(1101) <= not((inputs(78)) or (inputs(127)));
    layer0_outputs(1102) <= not(inputs(60));
    layer0_outputs(1103) <= not(inputs(137)) or (inputs(158));
    layer0_outputs(1104) <= (inputs(118)) xor (inputs(222));
    layer0_outputs(1105) <= not(inputs(77)) or (inputs(204));
    layer0_outputs(1106) <= not(inputs(216)) or (inputs(10));
    layer0_outputs(1107) <= not(inputs(232)) or (inputs(88));
    layer0_outputs(1108) <= not((inputs(254)) or (inputs(214)));
    layer0_outputs(1109) <= not(inputs(199));
    layer0_outputs(1110) <= (inputs(50)) and not (inputs(113));
    layer0_outputs(1111) <= not((inputs(14)) or (inputs(155)));
    layer0_outputs(1112) <= inputs(253);
    layer0_outputs(1113) <= not(inputs(232));
    layer0_outputs(1114) <= not((inputs(205)) xor (inputs(193)));
    layer0_outputs(1115) <= '1';
    layer0_outputs(1116) <= (inputs(12)) and not (inputs(222));
    layer0_outputs(1117) <= not((inputs(168)) xor (inputs(136)));
    layer0_outputs(1118) <= (inputs(65)) or (inputs(20));
    layer0_outputs(1119) <= not((inputs(147)) or (inputs(50)));
    layer0_outputs(1120) <= (inputs(92)) or (inputs(83));
    layer0_outputs(1121) <= not((inputs(0)) or (inputs(106)));
    layer0_outputs(1122) <= inputs(94);
    layer0_outputs(1123) <= (inputs(58)) and not (inputs(162));
    layer0_outputs(1124) <= '0';
    layer0_outputs(1125) <= (inputs(247)) xor (inputs(213));
    layer0_outputs(1126) <= inputs(102);
    layer0_outputs(1127) <= not(inputs(38));
    layer0_outputs(1128) <= not(inputs(174));
    layer0_outputs(1129) <= not(inputs(208));
    layer0_outputs(1130) <= not(inputs(25));
    layer0_outputs(1131) <= not((inputs(92)) or (inputs(197)));
    layer0_outputs(1132) <= (inputs(73)) xor (inputs(0));
    layer0_outputs(1133) <= (inputs(157)) or (inputs(165));
    layer0_outputs(1134) <= (inputs(137)) and not (inputs(207));
    layer0_outputs(1135) <= not((inputs(157)) or (inputs(5)));
    layer0_outputs(1136) <= not((inputs(11)) xor (inputs(110)));
    layer0_outputs(1137) <= inputs(212);
    layer0_outputs(1138) <= not((inputs(160)) xor (inputs(243)));
    layer0_outputs(1139) <= (inputs(238)) xor (inputs(223));
    layer0_outputs(1140) <= inputs(165);
    layer0_outputs(1141) <= not(inputs(103));
    layer0_outputs(1142) <= not(inputs(62)) or (inputs(2));
    layer0_outputs(1143) <= inputs(163);
    layer0_outputs(1144) <= not((inputs(61)) and (inputs(241)));
    layer0_outputs(1145) <= not((inputs(169)) xor (inputs(108)));
    layer0_outputs(1146) <= not(inputs(16)) or (inputs(228));
    layer0_outputs(1147) <= not((inputs(4)) or (inputs(90)));
    layer0_outputs(1148) <= not(inputs(106)) or (inputs(250));
    layer0_outputs(1149) <= (inputs(32)) or (inputs(248));
    layer0_outputs(1150) <= (inputs(159)) or (inputs(8));
    layer0_outputs(1151) <= '0';
    layer0_outputs(1152) <= not((inputs(244)) or (inputs(49)));
    layer0_outputs(1153) <= inputs(177);
    layer0_outputs(1154) <= inputs(146);
    layer0_outputs(1155) <= not(inputs(138));
    layer0_outputs(1156) <= not(inputs(98));
    layer0_outputs(1157) <= (inputs(159)) or (inputs(115));
    layer0_outputs(1158) <= inputs(135);
    layer0_outputs(1159) <= not((inputs(227)) or (inputs(174)));
    layer0_outputs(1160) <= not(inputs(255)) or (inputs(138));
    layer0_outputs(1161) <= (inputs(220)) and not (inputs(161));
    layer0_outputs(1162) <= (inputs(64)) and not (inputs(157));
    layer0_outputs(1163) <= (inputs(136)) xor (inputs(84));
    layer0_outputs(1164) <= not(inputs(131));
    layer0_outputs(1165) <= inputs(91);
    layer0_outputs(1166) <= (inputs(23)) xor (inputs(207));
    layer0_outputs(1167) <= not(inputs(82));
    layer0_outputs(1168) <= not((inputs(12)) or (inputs(152)));
    layer0_outputs(1169) <= (inputs(212)) and not (inputs(93));
    layer0_outputs(1170) <= not(inputs(197)) or (inputs(55));
    layer0_outputs(1171) <= (inputs(55)) xor (inputs(68));
    layer0_outputs(1172) <= (inputs(142)) xor (inputs(4));
    layer0_outputs(1173) <= (inputs(146)) xor (inputs(220));
    layer0_outputs(1174) <= (inputs(1)) or (inputs(237));
    layer0_outputs(1175) <= (inputs(131)) xor (inputs(151));
    layer0_outputs(1176) <= inputs(129);
    layer0_outputs(1177) <= not(inputs(125));
    layer0_outputs(1178) <= not(inputs(152)) or (inputs(224));
    layer0_outputs(1179) <= (inputs(80)) xor (inputs(60));
    layer0_outputs(1180) <= not((inputs(147)) or (inputs(143)));
    layer0_outputs(1181) <= (inputs(6)) or (inputs(94));
    layer0_outputs(1182) <= inputs(69);
    layer0_outputs(1183) <= (inputs(14)) or (inputs(95));
    layer0_outputs(1184) <= (inputs(96)) xor (inputs(102));
    layer0_outputs(1185) <= '0';
    layer0_outputs(1186) <= (inputs(40)) xor (inputs(0));
    layer0_outputs(1187) <= (inputs(160)) or (inputs(22));
    layer0_outputs(1188) <= '1';
    layer0_outputs(1189) <= not(inputs(38));
    layer0_outputs(1190) <= (inputs(234)) or (inputs(16));
    layer0_outputs(1191) <= inputs(137);
    layer0_outputs(1192) <= inputs(38);
    layer0_outputs(1193) <= (inputs(73)) or (inputs(130));
    layer0_outputs(1194) <= (inputs(23)) and not (inputs(209));
    layer0_outputs(1195) <= inputs(226);
    layer0_outputs(1196) <= (inputs(171)) and (inputs(8));
    layer0_outputs(1197) <= not(inputs(23));
    layer0_outputs(1198) <= inputs(132);
    layer0_outputs(1199) <= not(inputs(26)) or (inputs(133));
    layer0_outputs(1200) <= '0';
    layer0_outputs(1201) <= not(inputs(182)) or (inputs(248));
    layer0_outputs(1202) <= (inputs(118)) and not (inputs(167));
    layer0_outputs(1203) <= (inputs(116)) and not (inputs(81));
    layer0_outputs(1204) <= (inputs(130)) xor (inputs(0));
    layer0_outputs(1205) <= not(inputs(59)) or (inputs(223));
    layer0_outputs(1206) <= not((inputs(104)) xor (inputs(180)));
    layer0_outputs(1207) <= (inputs(179)) or (inputs(126));
    layer0_outputs(1208) <= (inputs(212)) or (inputs(143));
    layer0_outputs(1209) <= not(inputs(25));
    layer0_outputs(1210) <= (inputs(69)) xor (inputs(104));
    layer0_outputs(1211) <= not(inputs(255)) or (inputs(238));
    layer0_outputs(1212) <= not(inputs(81));
    layer0_outputs(1213) <= not((inputs(166)) xor (inputs(164)));
    layer0_outputs(1214) <= (inputs(174)) xor (inputs(161));
    layer0_outputs(1215) <= inputs(63);
    layer0_outputs(1216) <= not(inputs(38)) or (inputs(49));
    layer0_outputs(1217) <= '1';
    layer0_outputs(1218) <= (inputs(249)) and not (inputs(211));
    layer0_outputs(1219) <= inputs(248);
    layer0_outputs(1220) <= not(inputs(70));
    layer0_outputs(1221) <= (inputs(44)) xor (inputs(105));
    layer0_outputs(1222) <= not((inputs(40)) and (inputs(38)));
    layer0_outputs(1223) <= not(inputs(222));
    layer0_outputs(1224) <= (inputs(254)) and (inputs(15));
    layer0_outputs(1225) <= not(inputs(60));
    layer0_outputs(1226) <= (inputs(186)) or (inputs(170));
    layer0_outputs(1227) <= (inputs(46)) xor (inputs(13));
    layer0_outputs(1228) <= not((inputs(206)) xor (inputs(42)));
    layer0_outputs(1229) <= (inputs(91)) and not (inputs(140));
    layer0_outputs(1230) <= not(inputs(176));
    layer0_outputs(1231) <= (inputs(57)) or (inputs(106));
    layer0_outputs(1232) <= not((inputs(55)) xor (inputs(4)));
    layer0_outputs(1233) <= not((inputs(197)) xor (inputs(161)));
    layer0_outputs(1234) <= not(inputs(217));
    layer0_outputs(1235) <= inputs(217);
    layer0_outputs(1236) <= inputs(102);
    layer0_outputs(1237) <= not(inputs(104)) or (inputs(204));
    layer0_outputs(1238) <= not(inputs(132));
    layer0_outputs(1239) <= (inputs(0)) and not (inputs(28));
    layer0_outputs(1240) <= not((inputs(103)) or (inputs(152)));
    layer0_outputs(1241) <= (inputs(226)) xor (inputs(71));
    layer0_outputs(1242) <= not((inputs(87)) or (inputs(224)));
    layer0_outputs(1243) <= (inputs(189)) and not (inputs(237));
    layer0_outputs(1244) <= not(inputs(136));
    layer0_outputs(1245) <= inputs(19);
    layer0_outputs(1246) <= not(inputs(117)) or (inputs(237));
    layer0_outputs(1247) <= (inputs(63)) xor (inputs(250));
    layer0_outputs(1248) <= not((inputs(175)) or (inputs(253)));
    layer0_outputs(1249) <= inputs(186);
    layer0_outputs(1250) <= inputs(38);
    layer0_outputs(1251) <= not(inputs(133)) or (inputs(253));
    layer0_outputs(1252) <= inputs(19);
    layer0_outputs(1253) <= (inputs(236)) or (inputs(120));
    layer0_outputs(1254) <= not((inputs(194)) or (inputs(176)));
    layer0_outputs(1255) <= (inputs(180)) xor (inputs(226));
    layer0_outputs(1256) <= not(inputs(142));
    layer0_outputs(1257) <= (inputs(100)) and not (inputs(239));
    layer0_outputs(1258) <= inputs(117);
    layer0_outputs(1259) <= (inputs(100)) and not (inputs(10));
    layer0_outputs(1260) <= not(inputs(170)) or (inputs(96));
    layer0_outputs(1261) <= inputs(212);
    layer0_outputs(1262) <= not(inputs(93)) or (inputs(154));
    layer0_outputs(1263) <= not((inputs(206)) or (inputs(21)));
    layer0_outputs(1264) <= not((inputs(165)) xor (inputs(88)));
    layer0_outputs(1265) <= not((inputs(231)) xor (inputs(183)));
    layer0_outputs(1266) <= (inputs(211)) and not (inputs(248));
    layer0_outputs(1267) <= (inputs(187)) xor (inputs(93));
    layer0_outputs(1268) <= (inputs(203)) and (inputs(182));
    layer0_outputs(1269) <= not((inputs(222)) or (inputs(2)));
    layer0_outputs(1270) <= not(inputs(75)) or (inputs(224));
    layer0_outputs(1271) <= inputs(30);
    layer0_outputs(1272) <= not(inputs(121));
    layer0_outputs(1273) <= inputs(24);
    layer0_outputs(1274) <= not((inputs(95)) or (inputs(93)));
    layer0_outputs(1275) <= (inputs(214)) or (inputs(207));
    layer0_outputs(1276) <= not(inputs(217)) or (inputs(18));
    layer0_outputs(1277) <= inputs(131);
    layer0_outputs(1278) <= inputs(84);
    layer0_outputs(1279) <= (inputs(101)) and not (inputs(65));
    layer0_outputs(1280) <= not((inputs(177)) xor (inputs(235)));
    layer0_outputs(1281) <= not(inputs(72)) or (inputs(204));
    layer0_outputs(1282) <= (inputs(45)) xor (inputs(169));
    layer0_outputs(1283) <= inputs(68);
    layer0_outputs(1284) <= not(inputs(192));
    layer0_outputs(1285) <= inputs(89);
    layer0_outputs(1286) <= not((inputs(14)) xor (inputs(230)));
    layer0_outputs(1287) <= not(inputs(28));
    layer0_outputs(1288) <= not((inputs(13)) or (inputs(16)));
    layer0_outputs(1289) <= (inputs(52)) xor (inputs(132));
    layer0_outputs(1290) <= not(inputs(71)) or (inputs(180));
    layer0_outputs(1291) <= (inputs(146)) xor (inputs(121));
    layer0_outputs(1292) <= (inputs(45)) or (inputs(115));
    layer0_outputs(1293) <= not(inputs(138)) or (inputs(253));
    layer0_outputs(1294) <= (inputs(20)) or (inputs(0));
    layer0_outputs(1295) <= (inputs(71)) xor (inputs(68));
    layer0_outputs(1296) <= not(inputs(160));
    layer0_outputs(1297) <= not((inputs(122)) xor (inputs(150)));
    layer0_outputs(1298) <= (inputs(118)) xor (inputs(132));
    layer0_outputs(1299) <= not(inputs(89));
    layer0_outputs(1300) <= not(inputs(91));
    layer0_outputs(1301) <= not(inputs(123));
    layer0_outputs(1302) <= not((inputs(245)) or (inputs(172)));
    layer0_outputs(1303) <= not(inputs(85));
    layer0_outputs(1304) <= not((inputs(244)) and (inputs(231)));
    layer0_outputs(1305) <= '0';
    layer0_outputs(1306) <= inputs(248);
    layer0_outputs(1307) <= not(inputs(171)) or (inputs(199));
    layer0_outputs(1308) <= not(inputs(62));
    layer0_outputs(1309) <= not(inputs(145));
    layer0_outputs(1310) <= inputs(54);
    layer0_outputs(1311) <= not(inputs(9));
    layer0_outputs(1312) <= (inputs(201)) or (inputs(212));
    layer0_outputs(1313) <= not(inputs(119));
    layer0_outputs(1314) <= (inputs(18)) or (inputs(224));
    layer0_outputs(1315) <= (inputs(144)) and (inputs(230));
    layer0_outputs(1316) <= not(inputs(211));
    layer0_outputs(1317) <= (inputs(223)) and not (inputs(35));
    layer0_outputs(1318) <= not((inputs(133)) xor (inputs(239)));
    layer0_outputs(1319) <= (inputs(134)) and not (inputs(214));
    layer0_outputs(1320) <= not(inputs(11));
    layer0_outputs(1321) <= (inputs(31)) xor (inputs(204));
    layer0_outputs(1322) <= '0';
    layer0_outputs(1323) <= (inputs(168)) and not (inputs(65));
    layer0_outputs(1324) <= (inputs(125)) and not (inputs(75));
    layer0_outputs(1325) <= not(inputs(173)) or (inputs(98));
    layer0_outputs(1326) <= inputs(62);
    layer0_outputs(1327) <= inputs(222);
    layer0_outputs(1328) <= not((inputs(2)) xor (inputs(176)));
    layer0_outputs(1329) <= not(inputs(120));
    layer0_outputs(1330) <= inputs(38);
    layer0_outputs(1331) <= inputs(79);
    layer0_outputs(1332) <= (inputs(168)) xor (inputs(150));
    layer0_outputs(1333) <= not(inputs(220));
    layer0_outputs(1334) <= (inputs(61)) xor (inputs(207));
    layer0_outputs(1335) <= inputs(230);
    layer0_outputs(1336) <= not((inputs(164)) and (inputs(228)));
    layer0_outputs(1337) <= inputs(216);
    layer0_outputs(1338) <= inputs(22);
    layer0_outputs(1339) <= inputs(85);
    layer0_outputs(1340) <= (inputs(79)) and not (inputs(253));
    layer0_outputs(1341) <= (inputs(220)) and not (inputs(158));
    layer0_outputs(1342) <= not((inputs(207)) xor (inputs(107)));
    layer0_outputs(1343) <= not((inputs(44)) or (inputs(58)));
    layer0_outputs(1344) <= not(inputs(100));
    layer0_outputs(1345) <= not((inputs(35)) and (inputs(144)));
    layer0_outputs(1346) <= not(inputs(115));
    layer0_outputs(1347) <= inputs(116);
    layer0_outputs(1348) <= not(inputs(148)) or (inputs(46));
    layer0_outputs(1349) <= inputs(167);
    layer0_outputs(1350) <= (inputs(151)) xor (inputs(212));
    layer0_outputs(1351) <= (inputs(104)) or (inputs(237));
    layer0_outputs(1352) <= (inputs(221)) xor (inputs(210));
    layer0_outputs(1353) <= (inputs(246)) xor (inputs(12));
    layer0_outputs(1354) <= not(inputs(75));
    layer0_outputs(1355) <= '1';
    layer0_outputs(1356) <= not((inputs(220)) xor (inputs(29)));
    layer0_outputs(1357) <= not(inputs(15));
    layer0_outputs(1358) <= (inputs(201)) and not (inputs(42));
    layer0_outputs(1359) <= not((inputs(66)) xor (inputs(79)));
    layer0_outputs(1360) <= not(inputs(5)) or (inputs(82));
    layer0_outputs(1361) <= not((inputs(57)) xor (inputs(21)));
    layer0_outputs(1362) <= (inputs(124)) or (inputs(244));
    layer0_outputs(1363) <= not(inputs(63));
    layer0_outputs(1364) <= (inputs(229)) and (inputs(208));
    layer0_outputs(1365) <= (inputs(203)) xor (inputs(84));
    layer0_outputs(1366) <= (inputs(53)) and not (inputs(109));
    layer0_outputs(1367) <= not(inputs(180));
    layer0_outputs(1368) <= (inputs(24)) xor (inputs(210));
    layer0_outputs(1369) <= inputs(160);
    layer0_outputs(1370) <= not(inputs(38)) or (inputs(209));
    layer0_outputs(1371) <= not((inputs(24)) xor (inputs(109)));
    layer0_outputs(1372) <= not(inputs(0));
    layer0_outputs(1373) <= not(inputs(158)) or (inputs(186));
    layer0_outputs(1374) <= (inputs(153)) and (inputs(203));
    layer0_outputs(1375) <= inputs(42);
    layer0_outputs(1376) <= (inputs(249)) or (inputs(42));
    layer0_outputs(1377) <= not((inputs(33)) xor (inputs(93)));
    layer0_outputs(1378) <= (inputs(154)) and not (inputs(41));
    layer0_outputs(1379) <= (inputs(130)) and not (inputs(36));
    layer0_outputs(1380) <= not(inputs(54)) or (inputs(63));
    layer0_outputs(1381) <= inputs(15);
    layer0_outputs(1382) <= not(inputs(159));
    layer0_outputs(1383) <= (inputs(116)) xor (inputs(48));
    layer0_outputs(1384) <= not((inputs(157)) xor (inputs(205)));
    layer0_outputs(1385) <= (inputs(179)) xor (inputs(192));
    layer0_outputs(1386) <= not(inputs(152));
    layer0_outputs(1387) <= not(inputs(99));
    layer0_outputs(1388) <= not(inputs(185));
    layer0_outputs(1389) <= not(inputs(197)) or (inputs(241));
    layer0_outputs(1390) <= not((inputs(18)) or (inputs(142)));
    layer0_outputs(1391) <= (inputs(21)) xor (inputs(98));
    layer0_outputs(1392) <= not(inputs(70)) or (inputs(206));
    layer0_outputs(1393) <= (inputs(127)) xor (inputs(180));
    layer0_outputs(1394) <= inputs(118);
    layer0_outputs(1395) <= (inputs(221)) and not (inputs(15));
    layer0_outputs(1396) <= not(inputs(149));
    layer0_outputs(1397) <= not(inputs(220));
    layer0_outputs(1398) <= not((inputs(187)) xor (inputs(98)));
    layer0_outputs(1399) <= (inputs(66)) and (inputs(237));
    layer0_outputs(1400) <= inputs(140);
    layer0_outputs(1401) <= (inputs(152)) xor (inputs(137));
    layer0_outputs(1402) <= not(inputs(89));
    layer0_outputs(1403) <= (inputs(87)) xor (inputs(134));
    layer0_outputs(1404) <= (inputs(216)) and not (inputs(96));
    layer0_outputs(1405) <= (inputs(243)) and (inputs(122));
    layer0_outputs(1406) <= (inputs(1)) and not (inputs(151));
    layer0_outputs(1407) <= not(inputs(117));
    layer0_outputs(1408) <= not((inputs(251)) or (inputs(235)));
    layer0_outputs(1409) <= (inputs(230)) or (inputs(234));
    layer0_outputs(1410) <= not(inputs(244)) or (inputs(253));
    layer0_outputs(1411) <= inputs(88);
    layer0_outputs(1412) <= (inputs(39)) or (inputs(79));
    layer0_outputs(1413) <= not((inputs(193)) or (inputs(230)));
    layer0_outputs(1414) <= (inputs(45)) or (inputs(255));
    layer0_outputs(1415) <= inputs(130);
    layer0_outputs(1416) <= inputs(132);
    layer0_outputs(1417) <= inputs(150);
    layer0_outputs(1418) <= not((inputs(253)) or (inputs(227)));
    layer0_outputs(1419) <= not((inputs(162)) xor (inputs(145)));
    layer0_outputs(1420) <= not(inputs(71));
    layer0_outputs(1421) <= inputs(61);
    layer0_outputs(1422) <= not((inputs(77)) or (inputs(160)));
    layer0_outputs(1423) <= inputs(126);
    layer0_outputs(1424) <= not((inputs(101)) or (inputs(40)));
    layer0_outputs(1425) <= not(inputs(5)) or (inputs(129));
    layer0_outputs(1426) <= not(inputs(244)) or (inputs(159));
    layer0_outputs(1427) <= '0';
    layer0_outputs(1428) <= not((inputs(98)) or (inputs(203)));
    layer0_outputs(1429) <= inputs(107);
    layer0_outputs(1430) <= (inputs(95)) xor (inputs(251));
    layer0_outputs(1431) <= (inputs(179)) and not (inputs(1));
    layer0_outputs(1432) <= inputs(129);
    layer0_outputs(1433) <= not(inputs(121));
    layer0_outputs(1434) <= inputs(201);
    layer0_outputs(1435) <= inputs(116);
    layer0_outputs(1436) <= not(inputs(41));
    layer0_outputs(1437) <= not((inputs(14)) or (inputs(113)));
    layer0_outputs(1438) <= (inputs(122)) xor (inputs(105));
    layer0_outputs(1439) <= (inputs(193)) or (inputs(49));
    layer0_outputs(1440) <= inputs(61);
    layer0_outputs(1441) <= (inputs(141)) or (inputs(67));
    layer0_outputs(1442) <= inputs(165);
    layer0_outputs(1443) <= inputs(144);
    layer0_outputs(1444) <= not((inputs(68)) and (inputs(152)));
    layer0_outputs(1445) <= not(inputs(168));
    layer0_outputs(1446) <= not(inputs(4));
    layer0_outputs(1447) <= inputs(219);
    layer0_outputs(1448) <= inputs(149);
    layer0_outputs(1449) <= not((inputs(224)) xor (inputs(248)));
    layer0_outputs(1450) <= not(inputs(192));
    layer0_outputs(1451) <= (inputs(129)) or (inputs(245));
    layer0_outputs(1452) <= not(inputs(8));
    layer0_outputs(1453) <= (inputs(108)) or (inputs(48));
    layer0_outputs(1454) <= (inputs(187)) xor (inputs(111));
    layer0_outputs(1455) <= not((inputs(166)) or (inputs(65)));
    layer0_outputs(1456) <= not((inputs(172)) or (inputs(116)));
    layer0_outputs(1457) <= (inputs(41)) and not (inputs(161));
    layer0_outputs(1458) <= (inputs(250)) xor (inputs(47));
    layer0_outputs(1459) <= inputs(79);
    layer0_outputs(1460) <= (inputs(163)) and not (inputs(78));
    layer0_outputs(1461) <= not(inputs(225));
    layer0_outputs(1462) <= inputs(244);
    layer0_outputs(1463) <= (inputs(39)) and not (inputs(130));
    layer0_outputs(1464) <= not(inputs(214));
    layer0_outputs(1465) <= inputs(67);
    layer0_outputs(1466) <= (inputs(238)) or (inputs(165));
    layer0_outputs(1467) <= (inputs(155)) and not (inputs(82));
    layer0_outputs(1468) <= inputs(106);
    layer0_outputs(1469) <= (inputs(214)) and (inputs(35));
    layer0_outputs(1470) <= not(inputs(95));
    layer0_outputs(1471) <= not((inputs(10)) xor (inputs(21)));
    layer0_outputs(1472) <= not(inputs(202));
    layer0_outputs(1473) <= not(inputs(122)) or (inputs(133));
    layer0_outputs(1474) <= (inputs(82)) or (inputs(212));
    layer0_outputs(1475) <= not(inputs(103)) or (inputs(157));
    layer0_outputs(1476) <= (inputs(179)) and not (inputs(139));
    layer0_outputs(1477) <= inputs(162);
    layer0_outputs(1478) <= (inputs(217)) and not (inputs(62));
    layer0_outputs(1479) <= not(inputs(199));
    layer0_outputs(1480) <= not((inputs(24)) xor (inputs(71)));
    layer0_outputs(1481) <= not(inputs(227));
    layer0_outputs(1482) <= not((inputs(131)) xor (inputs(148)));
    layer0_outputs(1483) <= not(inputs(244)) or (inputs(16));
    layer0_outputs(1484) <= inputs(37);
    layer0_outputs(1485) <= not(inputs(120));
    layer0_outputs(1486) <= (inputs(168)) xor (inputs(217));
    layer0_outputs(1487) <= not(inputs(215));
    layer0_outputs(1488) <= (inputs(91)) and not (inputs(189));
    layer0_outputs(1489) <= not((inputs(213)) or (inputs(197)));
    layer0_outputs(1490) <= not(inputs(199)) or (inputs(249));
    layer0_outputs(1491) <= not(inputs(151));
    layer0_outputs(1492) <= (inputs(214)) or (inputs(139));
    layer0_outputs(1493) <= (inputs(240)) or (inputs(244));
    layer0_outputs(1494) <= inputs(25);
    layer0_outputs(1495) <= not((inputs(20)) xor (inputs(50)));
    layer0_outputs(1496) <= (inputs(169)) or (inputs(150));
    layer0_outputs(1497) <= (inputs(169)) and not (inputs(126));
    layer0_outputs(1498) <= '0';
    layer0_outputs(1499) <= inputs(82);
    layer0_outputs(1500) <= (inputs(166)) and not (inputs(70));
    layer0_outputs(1501) <= (inputs(217)) or (inputs(31));
    layer0_outputs(1502) <= inputs(105);
    layer0_outputs(1503) <= (inputs(61)) and (inputs(51));
    layer0_outputs(1504) <= not(inputs(37));
    layer0_outputs(1505) <= inputs(148);
    layer0_outputs(1506) <= not((inputs(174)) or (inputs(185)));
    layer0_outputs(1507) <= inputs(249);
    layer0_outputs(1508) <= not(inputs(53)) or (inputs(132));
    layer0_outputs(1509) <= inputs(96);
    layer0_outputs(1510) <= (inputs(172)) or (inputs(243));
    layer0_outputs(1511) <= not((inputs(54)) xor (inputs(147)));
    layer0_outputs(1512) <= (inputs(86)) xor (inputs(253));
    layer0_outputs(1513) <= not(inputs(234));
    layer0_outputs(1514) <= (inputs(98)) or (inputs(211));
    layer0_outputs(1515) <= not((inputs(215)) or (inputs(4)));
    layer0_outputs(1516) <= (inputs(89)) and not (inputs(147));
    layer0_outputs(1517) <= not(inputs(131));
    layer0_outputs(1518) <= not((inputs(156)) and (inputs(157)));
    layer0_outputs(1519) <= not((inputs(150)) xor (inputs(6)));
    layer0_outputs(1520) <= not(inputs(76));
    layer0_outputs(1521) <= inputs(225);
    layer0_outputs(1522) <= inputs(157);
    layer0_outputs(1523) <= not((inputs(172)) xor (inputs(253)));
    layer0_outputs(1524) <= (inputs(228)) and not (inputs(112));
    layer0_outputs(1525) <= (inputs(209)) or (inputs(20));
    layer0_outputs(1526) <= not(inputs(203));
    layer0_outputs(1527) <= (inputs(133)) and not (inputs(125));
    layer0_outputs(1528) <= not(inputs(147));
    layer0_outputs(1529) <= not((inputs(61)) or (inputs(43)));
    layer0_outputs(1530) <= not(inputs(35)) or (inputs(113));
    layer0_outputs(1531) <= not((inputs(149)) xor (inputs(112)));
    layer0_outputs(1532) <= not(inputs(180)) or (inputs(187));
    layer0_outputs(1533) <= not((inputs(20)) or (inputs(75)));
    layer0_outputs(1534) <= (inputs(203)) or (inputs(60));
    layer0_outputs(1535) <= not(inputs(52)) or (inputs(162));
    layer0_outputs(1536) <= (inputs(254)) or (inputs(235));
    layer0_outputs(1537) <= not((inputs(155)) or (inputs(78)));
    layer0_outputs(1538) <= (inputs(159)) xor (inputs(163));
    layer0_outputs(1539) <= (inputs(233)) xor (inputs(54));
    layer0_outputs(1540) <= not((inputs(145)) xor (inputs(132)));
    layer0_outputs(1541) <= (inputs(250)) xor (inputs(237));
    layer0_outputs(1542) <= inputs(56);
    layer0_outputs(1543) <= (inputs(246)) or (inputs(235));
    layer0_outputs(1544) <= inputs(19);
    layer0_outputs(1545) <= not((inputs(125)) or (inputs(38)));
    layer0_outputs(1546) <= (inputs(147)) and not (inputs(66));
    layer0_outputs(1547) <= not((inputs(210)) and (inputs(246)));
    layer0_outputs(1548) <= not(inputs(182)) or (inputs(131));
    layer0_outputs(1549) <= not(inputs(156));
    layer0_outputs(1550) <= not((inputs(106)) and (inputs(221)));
    layer0_outputs(1551) <= (inputs(96)) and not (inputs(214));
    layer0_outputs(1552) <= inputs(160);
    layer0_outputs(1553) <= not((inputs(6)) xor (inputs(144)));
    layer0_outputs(1554) <= not(inputs(154)) or (inputs(200));
    layer0_outputs(1555) <= inputs(189);
    layer0_outputs(1556) <= inputs(98);
    layer0_outputs(1557) <= (inputs(160)) xor (inputs(100));
    layer0_outputs(1558) <= (inputs(181)) and not (inputs(191));
    layer0_outputs(1559) <= not((inputs(57)) or (inputs(225)));
    layer0_outputs(1560) <= (inputs(192)) or (inputs(111));
    layer0_outputs(1561) <= not(inputs(53)) or (inputs(13));
    layer0_outputs(1562) <= inputs(128);
    layer0_outputs(1563) <= not((inputs(46)) and (inputs(240)));
    layer0_outputs(1564) <= inputs(161);
    layer0_outputs(1565) <= (inputs(3)) and not (inputs(110));
    layer0_outputs(1566) <= not((inputs(233)) xor (inputs(72)));
    layer0_outputs(1567) <= (inputs(31)) or (inputs(224));
    layer0_outputs(1568) <= not(inputs(127));
    layer0_outputs(1569) <= not((inputs(81)) or (inputs(63)));
    layer0_outputs(1570) <= not(inputs(90)) or (inputs(67));
    layer0_outputs(1571) <= not(inputs(149)) or (inputs(139));
    layer0_outputs(1572) <= not(inputs(121)) or (inputs(165));
    layer0_outputs(1573) <= not(inputs(172));
    layer0_outputs(1574) <= not(inputs(229));
    layer0_outputs(1575) <= (inputs(19)) and not (inputs(239));
    layer0_outputs(1576) <= (inputs(240)) and not (inputs(255));
    layer0_outputs(1577) <= not((inputs(127)) xor (inputs(133)));
    layer0_outputs(1578) <= not((inputs(56)) or (inputs(230)));
    layer0_outputs(1579) <= inputs(57);
    layer0_outputs(1580) <= not(inputs(20)) or (inputs(31));
    layer0_outputs(1581) <= inputs(88);
    layer0_outputs(1582) <= (inputs(182)) and not (inputs(28));
    layer0_outputs(1583) <= (inputs(251)) xor (inputs(209));
    layer0_outputs(1584) <= (inputs(129)) or (inputs(183));
    layer0_outputs(1585) <= not((inputs(191)) xor (inputs(227)));
    layer0_outputs(1586) <= '0';
    layer0_outputs(1587) <= not((inputs(62)) and (inputs(242)));
    layer0_outputs(1588) <= (inputs(250)) and not (inputs(99));
    layer0_outputs(1589) <= not(inputs(27));
    layer0_outputs(1590) <= (inputs(215)) and (inputs(106));
    layer0_outputs(1591) <= not(inputs(89)) or (inputs(148));
    layer0_outputs(1592) <= (inputs(105)) and not (inputs(198));
    layer0_outputs(1593) <= inputs(61);
    layer0_outputs(1594) <= not(inputs(58));
    layer0_outputs(1595) <= not((inputs(142)) xor (inputs(160)));
    layer0_outputs(1596) <= not(inputs(21)) or (inputs(101));
    layer0_outputs(1597) <= (inputs(122)) and not (inputs(212));
    layer0_outputs(1598) <= not(inputs(182)) or (inputs(201));
    layer0_outputs(1599) <= not((inputs(180)) or (inputs(131)));
    layer0_outputs(1600) <= (inputs(215)) and (inputs(213));
    layer0_outputs(1601) <= not((inputs(50)) xor (inputs(46)));
    layer0_outputs(1602) <= (inputs(155)) and not (inputs(235));
    layer0_outputs(1603) <= '0';
    layer0_outputs(1604) <= inputs(101);
    layer0_outputs(1605) <= not(inputs(85));
    layer0_outputs(1606) <= not(inputs(81));
    layer0_outputs(1607) <= inputs(14);
    layer0_outputs(1608) <= not((inputs(217)) or (inputs(76)));
    layer0_outputs(1609) <= (inputs(1)) and not (inputs(98));
    layer0_outputs(1610) <= (inputs(172)) and not (inputs(2));
    layer0_outputs(1611) <= not(inputs(184));
    layer0_outputs(1612) <= (inputs(246)) and not (inputs(182));
    layer0_outputs(1613) <= not((inputs(3)) or (inputs(158)));
    layer0_outputs(1614) <= (inputs(213)) or (inputs(233));
    layer0_outputs(1615) <= not((inputs(33)) xor (inputs(27)));
    layer0_outputs(1616) <= not((inputs(117)) and (inputs(161)));
    layer0_outputs(1617) <= (inputs(41)) and not (inputs(127));
    layer0_outputs(1618) <= (inputs(106)) and not (inputs(99));
    layer0_outputs(1619) <= not(inputs(55));
    layer0_outputs(1620) <= not(inputs(165));
    layer0_outputs(1621) <= not((inputs(194)) and (inputs(231)));
    layer0_outputs(1622) <= (inputs(89)) xor (inputs(242));
    layer0_outputs(1623) <= not((inputs(2)) or (inputs(246)));
    layer0_outputs(1624) <= not(inputs(235));
    layer0_outputs(1625) <= not((inputs(9)) xor (inputs(43)));
    layer0_outputs(1626) <= (inputs(91)) or (inputs(112));
    layer0_outputs(1627) <= not(inputs(18)) or (inputs(65));
    layer0_outputs(1628) <= (inputs(27)) xor (inputs(74));
    layer0_outputs(1629) <= inputs(31);
    layer0_outputs(1630) <= not(inputs(88));
    layer0_outputs(1631) <= not((inputs(255)) xor (inputs(58)));
    layer0_outputs(1632) <= not(inputs(85));
    layer0_outputs(1633) <= not((inputs(88)) or (inputs(136)));
    layer0_outputs(1634) <= inputs(118);
    layer0_outputs(1635) <= (inputs(247)) and not (inputs(110));
    layer0_outputs(1636) <= not(inputs(21)) or (inputs(144));
    layer0_outputs(1637) <= inputs(210);
    layer0_outputs(1638) <= not((inputs(160)) or (inputs(213)));
    layer0_outputs(1639) <= not(inputs(65)) or (inputs(12));
    layer0_outputs(1640) <= not(inputs(210));
    layer0_outputs(1641) <= not(inputs(227));
    layer0_outputs(1642) <= not(inputs(43)) or (inputs(225));
    layer0_outputs(1643) <= not((inputs(77)) or (inputs(95)));
    layer0_outputs(1644) <= (inputs(219)) and not (inputs(115));
    layer0_outputs(1645) <= inputs(227);
    layer0_outputs(1646) <= not(inputs(74));
    layer0_outputs(1647) <= (inputs(165)) and not (inputs(114));
    layer0_outputs(1648) <= (inputs(45)) xor (inputs(75));
    layer0_outputs(1649) <= not(inputs(8));
    layer0_outputs(1650) <= (inputs(131)) and not (inputs(229));
    layer0_outputs(1651) <= not(inputs(198));
    layer0_outputs(1652) <= (inputs(234)) xor (inputs(86));
    layer0_outputs(1653) <= not(inputs(123)) or (inputs(71));
    layer0_outputs(1654) <= not((inputs(59)) xor (inputs(13)));
    layer0_outputs(1655) <= inputs(44);
    layer0_outputs(1656) <= not(inputs(25));
    layer0_outputs(1657) <= not((inputs(85)) or (inputs(205)));
    layer0_outputs(1658) <= not((inputs(169)) or (inputs(188)));
    layer0_outputs(1659) <= (inputs(232)) or (inputs(158));
    layer0_outputs(1660) <= not(inputs(80)) or (inputs(0));
    layer0_outputs(1661) <= not((inputs(90)) and (inputs(38)));
    layer0_outputs(1662) <= not((inputs(94)) or (inputs(108)));
    layer0_outputs(1663) <= not(inputs(223));
    layer0_outputs(1664) <= inputs(151);
    layer0_outputs(1665) <= not(inputs(221)) or (inputs(109));
    layer0_outputs(1666) <= not((inputs(214)) or (inputs(101)));
    layer0_outputs(1667) <= not(inputs(127));
    layer0_outputs(1668) <= inputs(189);
    layer0_outputs(1669) <= '0';
    layer0_outputs(1670) <= (inputs(25)) xor (inputs(56));
    layer0_outputs(1671) <= (inputs(166)) and not (inputs(102));
    layer0_outputs(1672) <= (inputs(161)) or (inputs(188));
    layer0_outputs(1673) <= not(inputs(230));
    layer0_outputs(1674) <= (inputs(13)) and (inputs(207));
    layer0_outputs(1675) <= inputs(246);
    layer0_outputs(1676) <= inputs(64);
    layer0_outputs(1677) <= (inputs(217)) xor (inputs(202));
    layer0_outputs(1678) <= not((inputs(112)) or (inputs(213)));
    layer0_outputs(1679) <= inputs(120);
    layer0_outputs(1680) <= not((inputs(112)) xor (inputs(69)));
    layer0_outputs(1681) <= inputs(27);
    layer0_outputs(1682) <= not(inputs(219)) or (inputs(77));
    layer0_outputs(1683) <= not((inputs(249)) or (inputs(195)));
    layer0_outputs(1684) <= (inputs(153)) and not (inputs(45));
    layer0_outputs(1685) <= not((inputs(231)) or (inputs(193)));
    layer0_outputs(1686) <= (inputs(172)) and not (inputs(17));
    layer0_outputs(1687) <= not((inputs(130)) or (inputs(131)));
    layer0_outputs(1688) <= (inputs(40)) and not (inputs(46));
    layer0_outputs(1689) <= not((inputs(98)) xor (inputs(210)));
    layer0_outputs(1690) <= (inputs(235)) or (inputs(89));
    layer0_outputs(1691) <= not(inputs(143));
    layer0_outputs(1692) <= not(inputs(231));
    layer0_outputs(1693) <= (inputs(121)) xor (inputs(114));
    layer0_outputs(1694) <= not(inputs(6)) or (inputs(195));
    layer0_outputs(1695) <= not((inputs(90)) or (inputs(65)));
    layer0_outputs(1696) <= not(inputs(229));
    layer0_outputs(1697) <= not((inputs(186)) or (inputs(182)));
    layer0_outputs(1698) <= not(inputs(183)) or (inputs(91));
    layer0_outputs(1699) <= not((inputs(199)) and (inputs(156)));
    layer0_outputs(1700) <= (inputs(58)) or (inputs(144));
    layer0_outputs(1701) <= not((inputs(98)) or (inputs(123)));
    layer0_outputs(1702) <= (inputs(31)) and not (inputs(76));
    layer0_outputs(1703) <= (inputs(172)) and not (inputs(236));
    layer0_outputs(1704) <= not(inputs(145));
    layer0_outputs(1705) <= not(inputs(190)) or (inputs(4));
    layer0_outputs(1706) <= inputs(19);
    layer0_outputs(1707) <= (inputs(188)) or (inputs(215));
    layer0_outputs(1708) <= inputs(17);
    layer0_outputs(1709) <= not(inputs(150)) or (inputs(2));
    layer0_outputs(1710) <= not((inputs(132)) xor (inputs(207)));
    layer0_outputs(1711) <= not((inputs(18)) or (inputs(46)));
    layer0_outputs(1712) <= not(inputs(197));
    layer0_outputs(1713) <= not(inputs(83)) or (inputs(205));
    layer0_outputs(1714) <= not(inputs(228));
    layer0_outputs(1715) <= (inputs(1)) or (inputs(138));
    layer0_outputs(1716) <= not(inputs(238)) or (inputs(211));
    layer0_outputs(1717) <= (inputs(64)) or (inputs(136));
    layer0_outputs(1718) <= not(inputs(222));
    layer0_outputs(1719) <= not((inputs(128)) or (inputs(123)));
    layer0_outputs(1720) <= inputs(65);
    layer0_outputs(1721) <= not(inputs(71)) or (inputs(170));
    layer0_outputs(1722) <= not((inputs(136)) or (inputs(238)));
    layer0_outputs(1723) <= inputs(166);
    layer0_outputs(1724) <= (inputs(180)) and not (inputs(11));
    layer0_outputs(1725) <= (inputs(169)) and not (inputs(212));
    layer0_outputs(1726) <= not((inputs(198)) or (inputs(119)));
    layer0_outputs(1727) <= not(inputs(56));
    layer0_outputs(1728) <= not(inputs(127));
    layer0_outputs(1729) <= not((inputs(59)) or (inputs(65)));
    layer0_outputs(1730) <= inputs(149);
    layer0_outputs(1731) <= not(inputs(29)) or (inputs(198));
    layer0_outputs(1732) <= not((inputs(35)) xor (inputs(42)));
    layer0_outputs(1733) <= (inputs(78)) xor (inputs(76));
    layer0_outputs(1734) <= not((inputs(9)) or (inputs(61)));
    layer0_outputs(1735) <= not((inputs(51)) or (inputs(193)));
    layer0_outputs(1736) <= (inputs(122)) and not (inputs(65));
    layer0_outputs(1737) <= inputs(191);
    layer0_outputs(1738) <= (inputs(231)) and not (inputs(34));
    layer0_outputs(1739) <= (inputs(191)) or (inputs(125));
    layer0_outputs(1740) <= not((inputs(176)) or (inputs(235)));
    layer0_outputs(1741) <= not((inputs(231)) and (inputs(7)));
    layer0_outputs(1742) <= (inputs(120)) and not (inputs(26));
    layer0_outputs(1743) <= inputs(37);
    layer0_outputs(1744) <= not((inputs(16)) or (inputs(194)));
    layer0_outputs(1745) <= not(inputs(31));
    layer0_outputs(1746) <= (inputs(70)) and not (inputs(17));
    layer0_outputs(1747) <= not(inputs(141)) or (inputs(227));
    layer0_outputs(1748) <= not((inputs(191)) and (inputs(200)));
    layer0_outputs(1749) <= not((inputs(82)) or (inputs(84)));
    layer0_outputs(1750) <= not(inputs(87));
    layer0_outputs(1751) <= '0';
    layer0_outputs(1752) <= (inputs(106)) and (inputs(28));
    layer0_outputs(1753) <= inputs(89);
    layer0_outputs(1754) <= (inputs(164)) xor (inputs(173));
    layer0_outputs(1755) <= inputs(110);
    layer0_outputs(1756) <= (inputs(24)) and not (inputs(183));
    layer0_outputs(1757) <= not(inputs(106)) or (inputs(50));
    layer0_outputs(1758) <= inputs(220);
    layer0_outputs(1759) <= not((inputs(205)) and (inputs(169)));
    layer0_outputs(1760) <= not((inputs(145)) or (inputs(242)));
    layer0_outputs(1761) <= (inputs(55)) xor (inputs(215));
    layer0_outputs(1762) <= not(inputs(120)) or (inputs(165));
    layer0_outputs(1763) <= inputs(146);
    layer0_outputs(1764) <= not(inputs(188)) or (inputs(59));
    layer0_outputs(1765) <= inputs(246);
    layer0_outputs(1766) <= not((inputs(157)) and (inputs(212)));
    layer0_outputs(1767) <= not(inputs(56));
    layer0_outputs(1768) <= not(inputs(108)) or (inputs(198));
    layer0_outputs(1769) <= not((inputs(132)) xor (inputs(160)));
    layer0_outputs(1770) <= inputs(165);
    layer0_outputs(1771) <= not((inputs(179)) or (inputs(225)));
    layer0_outputs(1772) <= not((inputs(97)) or (inputs(142)));
    layer0_outputs(1773) <= (inputs(171)) and (inputs(202));
    layer0_outputs(1774) <= inputs(21);
    layer0_outputs(1775) <= (inputs(187)) or (inputs(211));
    layer0_outputs(1776) <= inputs(22);
    layer0_outputs(1777) <= not((inputs(170)) and (inputs(197)));
    layer0_outputs(1778) <= not(inputs(198));
    layer0_outputs(1779) <= not((inputs(76)) or (inputs(97)));
    layer0_outputs(1780) <= inputs(116);
    layer0_outputs(1781) <= not(inputs(202)) or (inputs(238));
    layer0_outputs(1782) <= not(inputs(180));
    layer0_outputs(1783) <= inputs(209);
    layer0_outputs(1784) <= not(inputs(214));
    layer0_outputs(1785) <= '0';
    layer0_outputs(1786) <= inputs(221);
    layer0_outputs(1787) <= not(inputs(193));
    layer0_outputs(1788) <= (inputs(57)) or (inputs(255));
    layer0_outputs(1789) <= (inputs(58)) and not (inputs(252));
    layer0_outputs(1790) <= not((inputs(64)) or (inputs(208)));
    layer0_outputs(1791) <= not(inputs(225)) or (inputs(127));
    layer0_outputs(1792) <= (inputs(151)) or (inputs(230));
    layer0_outputs(1793) <= not((inputs(208)) xor (inputs(68)));
    layer0_outputs(1794) <= inputs(25);
    layer0_outputs(1795) <= (inputs(160)) or (inputs(206));
    layer0_outputs(1796) <= (inputs(129)) or (inputs(176));
    layer0_outputs(1797) <= not(inputs(157));
    layer0_outputs(1798) <= inputs(135);
    layer0_outputs(1799) <= inputs(43);
    layer0_outputs(1800) <= not(inputs(129)) or (inputs(34));
    layer0_outputs(1801) <= not((inputs(91)) xor (inputs(142)));
    layer0_outputs(1802) <= not((inputs(18)) xor (inputs(207)));
    layer0_outputs(1803) <= (inputs(146)) or (inputs(66));
    layer0_outputs(1804) <= not(inputs(197));
    layer0_outputs(1805) <= (inputs(88)) or (inputs(173));
    layer0_outputs(1806) <= not(inputs(135)) or (inputs(97));
    layer0_outputs(1807) <= not(inputs(137));
    layer0_outputs(1808) <= inputs(4);
    layer0_outputs(1809) <= not(inputs(122));
    layer0_outputs(1810) <= not(inputs(137));
    layer0_outputs(1811) <= (inputs(72)) xor (inputs(27));
    layer0_outputs(1812) <= (inputs(233)) and (inputs(182));
    layer0_outputs(1813) <= (inputs(46)) or (inputs(46));
    layer0_outputs(1814) <= (inputs(220)) and not (inputs(66));
    layer0_outputs(1815) <= not((inputs(35)) xor (inputs(13)));
    layer0_outputs(1816) <= not(inputs(168)) or (inputs(45));
    layer0_outputs(1817) <= (inputs(115)) and not (inputs(235));
    layer0_outputs(1818) <= not((inputs(58)) or (inputs(101)));
    layer0_outputs(1819) <= not((inputs(173)) and (inputs(244)));
    layer0_outputs(1820) <= (inputs(234)) xor (inputs(249));
    layer0_outputs(1821) <= not((inputs(16)) or (inputs(48)));
    layer0_outputs(1822) <= not((inputs(47)) or (inputs(36)));
    layer0_outputs(1823) <= not(inputs(214)) or (inputs(138));
    layer0_outputs(1824) <= not((inputs(16)) xor (inputs(123)));
    layer0_outputs(1825) <= not(inputs(147));
    layer0_outputs(1826) <= (inputs(246)) and not (inputs(192));
    layer0_outputs(1827) <= '0';
    layer0_outputs(1828) <= not((inputs(136)) xor (inputs(145)));
    layer0_outputs(1829) <= (inputs(201)) or (inputs(63));
    layer0_outputs(1830) <= not(inputs(66));
    layer0_outputs(1831) <= not((inputs(233)) xor (inputs(153)));
    layer0_outputs(1832) <= (inputs(213)) and (inputs(183));
    layer0_outputs(1833) <= inputs(170);
    layer0_outputs(1834) <= inputs(202);
    layer0_outputs(1835) <= inputs(232);
    layer0_outputs(1836) <= (inputs(6)) or (inputs(21));
    layer0_outputs(1837) <= inputs(98);
    layer0_outputs(1838) <= (inputs(179)) or (inputs(235));
    layer0_outputs(1839) <= '1';
    layer0_outputs(1840) <= not(inputs(38));
    layer0_outputs(1841) <= not(inputs(245)) or (inputs(64));
    layer0_outputs(1842) <= inputs(147);
    layer0_outputs(1843) <= (inputs(215)) and not (inputs(143));
    layer0_outputs(1844) <= not((inputs(102)) xor (inputs(63)));
    layer0_outputs(1845) <= not(inputs(113));
    layer0_outputs(1846) <= inputs(23);
    layer0_outputs(1847) <= (inputs(117)) and not (inputs(181));
    layer0_outputs(1848) <= not(inputs(93)) or (inputs(225));
    layer0_outputs(1849) <= (inputs(99)) and not (inputs(255));
    layer0_outputs(1850) <= not(inputs(50));
    layer0_outputs(1851) <= not((inputs(78)) xor (inputs(213)));
    layer0_outputs(1852) <= (inputs(82)) xor (inputs(116));
    layer0_outputs(1853) <= (inputs(122)) xor (inputs(156));
    layer0_outputs(1854) <= (inputs(230)) or (inputs(63));
    layer0_outputs(1855) <= inputs(170);
    layer0_outputs(1856) <= (inputs(106)) or (inputs(138));
    layer0_outputs(1857) <= inputs(218);
    layer0_outputs(1858) <= '1';
    layer0_outputs(1859) <= (inputs(119)) and (inputs(74));
    layer0_outputs(1860) <= not(inputs(89)) or (inputs(49));
    layer0_outputs(1861) <= (inputs(70)) and not (inputs(239));
    layer0_outputs(1862) <= not((inputs(200)) xor (inputs(18)));
    layer0_outputs(1863) <= inputs(107);
    layer0_outputs(1864) <= not(inputs(164));
    layer0_outputs(1865) <= not(inputs(141));
    layer0_outputs(1866) <= '0';
    layer0_outputs(1867) <= inputs(150);
    layer0_outputs(1868) <= not(inputs(30));
    layer0_outputs(1869) <= (inputs(49)) xor (inputs(3));
    layer0_outputs(1870) <= (inputs(185)) and not (inputs(111));
    layer0_outputs(1871) <= not(inputs(21));
    layer0_outputs(1872) <= not(inputs(104));
    layer0_outputs(1873) <= inputs(114);
    layer0_outputs(1874) <= not(inputs(159)) or (inputs(80));
    layer0_outputs(1875) <= not((inputs(214)) xor (inputs(247)));
    layer0_outputs(1876) <= not(inputs(175));
    layer0_outputs(1877) <= (inputs(142)) xor (inputs(12));
    layer0_outputs(1878) <= not(inputs(213));
    layer0_outputs(1879) <= (inputs(57)) and not (inputs(219));
    layer0_outputs(1880) <= (inputs(217)) and not (inputs(179));
    layer0_outputs(1881) <= (inputs(152)) xor (inputs(193));
    layer0_outputs(1882) <= (inputs(223)) or (inputs(30));
    layer0_outputs(1883) <= (inputs(107)) or (inputs(60));
    layer0_outputs(1884) <= not((inputs(187)) and (inputs(154)));
    layer0_outputs(1885) <= not((inputs(32)) and (inputs(30)));
    layer0_outputs(1886) <= not((inputs(164)) xor (inputs(46)));
    layer0_outputs(1887) <= inputs(249);
    layer0_outputs(1888) <= not(inputs(26)) or (inputs(226));
    layer0_outputs(1889) <= (inputs(18)) or (inputs(252));
    layer0_outputs(1890) <= (inputs(154)) xor (inputs(21));
    layer0_outputs(1891) <= inputs(94);
    layer0_outputs(1892) <= not(inputs(86));
    layer0_outputs(1893) <= not((inputs(73)) xor (inputs(104)));
    layer0_outputs(1894) <= not(inputs(73));
    layer0_outputs(1895) <= (inputs(166)) and not (inputs(47));
    layer0_outputs(1896) <= (inputs(251)) xor (inputs(180));
    layer0_outputs(1897) <= not(inputs(53));
    layer0_outputs(1898) <= not((inputs(42)) and (inputs(118)));
    layer0_outputs(1899) <= not(inputs(168));
    layer0_outputs(1900) <= (inputs(214)) and not (inputs(153));
    layer0_outputs(1901) <= (inputs(53)) or (inputs(63));
    layer0_outputs(1902) <= (inputs(30)) xor (inputs(19));
    layer0_outputs(1903) <= not(inputs(23));
    layer0_outputs(1904) <= not(inputs(58));
    layer0_outputs(1905) <= not(inputs(77));
    layer0_outputs(1906) <= not(inputs(109)) or (inputs(254));
    layer0_outputs(1907) <= inputs(173);
    layer0_outputs(1908) <= not(inputs(236));
    layer0_outputs(1909) <= not(inputs(17)) or (inputs(14));
    layer0_outputs(1910) <= (inputs(60)) xor (inputs(19));
    layer0_outputs(1911) <= inputs(48);
    layer0_outputs(1912) <= inputs(136);
    layer0_outputs(1913) <= (inputs(156)) or (inputs(60));
    layer0_outputs(1914) <= not((inputs(75)) or (inputs(187)));
    layer0_outputs(1915) <= not(inputs(73)) or (inputs(239));
    layer0_outputs(1916) <= not(inputs(135)) or (inputs(62));
    layer0_outputs(1917) <= (inputs(198)) and not (inputs(14));
    layer0_outputs(1918) <= (inputs(217)) and (inputs(182));
    layer0_outputs(1919) <= inputs(208);
    layer0_outputs(1920) <= (inputs(209)) or (inputs(158));
    layer0_outputs(1921) <= inputs(164);
    layer0_outputs(1922) <= inputs(182);
    layer0_outputs(1923) <= (inputs(10)) and not (inputs(252));
    layer0_outputs(1924) <= inputs(110);
    layer0_outputs(1925) <= not((inputs(129)) or (inputs(139)));
    layer0_outputs(1926) <= (inputs(153)) or (inputs(157));
    layer0_outputs(1927) <= inputs(145);
    layer0_outputs(1928) <= (inputs(202)) and not (inputs(238));
    layer0_outputs(1929) <= (inputs(8)) xor (inputs(78));
    layer0_outputs(1930) <= not((inputs(65)) or (inputs(68)));
    layer0_outputs(1931) <= inputs(247);
    layer0_outputs(1932) <= (inputs(0)) and not (inputs(161));
    layer0_outputs(1933) <= not((inputs(230)) or (inputs(229)));
    layer0_outputs(1934) <= (inputs(48)) or (inputs(235));
    layer0_outputs(1935) <= (inputs(36)) and not (inputs(157));
    layer0_outputs(1936) <= (inputs(167)) and not (inputs(222));
    layer0_outputs(1937) <= (inputs(112)) xor (inputs(146));
    layer0_outputs(1938) <= not(inputs(209));
    layer0_outputs(1939) <= (inputs(150)) and not (inputs(108));
    layer0_outputs(1940) <= inputs(222);
    layer0_outputs(1941) <= not((inputs(131)) xor (inputs(102)));
    layer0_outputs(1942) <= (inputs(170)) xor (inputs(186));
    layer0_outputs(1943) <= (inputs(87)) xor (inputs(243));
    layer0_outputs(1944) <= (inputs(158)) or (inputs(175));
    layer0_outputs(1945) <= inputs(147);
    layer0_outputs(1946) <= (inputs(247)) and not (inputs(110));
    layer0_outputs(1947) <= not(inputs(136)) or (inputs(210));
    layer0_outputs(1948) <= (inputs(82)) or (inputs(152));
    layer0_outputs(1949) <= (inputs(217)) xor (inputs(169));
    layer0_outputs(1950) <= (inputs(43)) or (inputs(96));
    layer0_outputs(1951) <= not((inputs(242)) xor (inputs(150)));
    layer0_outputs(1952) <= not((inputs(228)) or (inputs(22)));
    layer0_outputs(1953) <= not(inputs(246));
    layer0_outputs(1954) <= not((inputs(33)) or (inputs(24)));
    layer0_outputs(1955) <= not((inputs(89)) xor (inputs(175)));
    layer0_outputs(1956) <= not((inputs(132)) or (inputs(254)));
    layer0_outputs(1957) <= not(inputs(32)) or (inputs(65));
    layer0_outputs(1958) <= inputs(68);
    layer0_outputs(1959) <= (inputs(156)) and not (inputs(41));
    layer0_outputs(1960) <= not((inputs(10)) and (inputs(39)));
    layer0_outputs(1961) <= inputs(231);
    layer0_outputs(1962) <= inputs(63);
    layer0_outputs(1963) <= (inputs(35)) xor (inputs(82));
    layer0_outputs(1964) <= inputs(250);
    layer0_outputs(1965) <= (inputs(106)) and not (inputs(237));
    layer0_outputs(1966) <= not(inputs(168));
    layer0_outputs(1967) <= inputs(22);
    layer0_outputs(1968) <= (inputs(194)) or (inputs(237));
    layer0_outputs(1969) <= (inputs(108)) or (inputs(92));
    layer0_outputs(1970) <= (inputs(180)) or (inputs(113));
    layer0_outputs(1971) <= not(inputs(218)) or (inputs(29));
    layer0_outputs(1972) <= not(inputs(120)) or (inputs(171));
    layer0_outputs(1973) <= not(inputs(71)) or (inputs(151));
    layer0_outputs(1974) <= inputs(140);
    layer0_outputs(1975) <= (inputs(28)) xor (inputs(91));
    layer0_outputs(1976) <= not((inputs(127)) xor (inputs(181)));
    layer0_outputs(1977) <= not((inputs(229)) or (inputs(249)));
    layer0_outputs(1978) <= not((inputs(164)) or (inputs(234)));
    layer0_outputs(1979) <= not((inputs(130)) xor (inputs(18)));
    layer0_outputs(1980) <= (inputs(2)) xor (inputs(84));
    layer0_outputs(1981) <= inputs(70);
    layer0_outputs(1982) <= not(inputs(101));
    layer0_outputs(1983) <= not(inputs(179)) or (inputs(36));
    layer0_outputs(1984) <= (inputs(100)) and not (inputs(92));
    layer0_outputs(1985) <= not(inputs(132));
    layer0_outputs(1986) <= inputs(228);
    layer0_outputs(1987) <= (inputs(153)) and not (inputs(223));
    layer0_outputs(1988) <= inputs(158);
    layer0_outputs(1989) <= not((inputs(254)) or (inputs(218)));
    layer0_outputs(1990) <= (inputs(66)) and not (inputs(214));
    layer0_outputs(1991) <= (inputs(56)) and (inputs(59));
    layer0_outputs(1992) <= (inputs(235)) and not (inputs(117));
    layer0_outputs(1993) <= (inputs(8)) or (inputs(214));
    layer0_outputs(1994) <= not(inputs(121));
    layer0_outputs(1995) <= (inputs(43)) and not (inputs(193));
    layer0_outputs(1996) <= not(inputs(62));
    layer0_outputs(1997) <= (inputs(168)) xor (inputs(24));
    layer0_outputs(1998) <= not((inputs(223)) or (inputs(7)));
    layer0_outputs(1999) <= inputs(158);
    layer0_outputs(2000) <= (inputs(122)) and (inputs(217));
    layer0_outputs(2001) <= not(inputs(249)) or (inputs(91));
    layer0_outputs(2002) <= (inputs(242)) or (inputs(177));
    layer0_outputs(2003) <= (inputs(163)) or (inputs(223));
    layer0_outputs(2004) <= (inputs(243)) and (inputs(218));
    layer0_outputs(2005) <= not((inputs(13)) or (inputs(239)));
    layer0_outputs(2006) <= not((inputs(198)) or (inputs(186)));
    layer0_outputs(2007) <= inputs(226);
    layer0_outputs(2008) <= not((inputs(81)) xor (inputs(84)));
    layer0_outputs(2009) <= not(inputs(212)) or (inputs(222));
    layer0_outputs(2010) <= (inputs(180)) xor (inputs(179));
    layer0_outputs(2011) <= (inputs(207)) and (inputs(175));
    layer0_outputs(2012) <= (inputs(31)) and not (inputs(18));
    layer0_outputs(2013) <= inputs(153);
    layer0_outputs(2014) <= inputs(96);
    layer0_outputs(2015) <= (inputs(41)) xor (inputs(8));
    layer0_outputs(2016) <= not(inputs(83)) or (inputs(210));
    layer0_outputs(2017) <= not(inputs(87));
    layer0_outputs(2018) <= not(inputs(166));
    layer0_outputs(2019) <= (inputs(236)) and not (inputs(0));
    layer0_outputs(2020) <= inputs(174);
    layer0_outputs(2021) <= not(inputs(196));
    layer0_outputs(2022) <= inputs(108);
    layer0_outputs(2023) <= (inputs(168)) xor (inputs(138));
    layer0_outputs(2024) <= not((inputs(71)) or (inputs(195)));
    layer0_outputs(2025) <= not((inputs(36)) or (inputs(242)));
    layer0_outputs(2026) <= (inputs(14)) or (inputs(86));
    layer0_outputs(2027) <= (inputs(88)) xor (inputs(186));
    layer0_outputs(2028) <= (inputs(213)) or (inputs(242));
    layer0_outputs(2029) <= not(inputs(231)) or (inputs(220));
    layer0_outputs(2030) <= not(inputs(25));
    layer0_outputs(2031) <= (inputs(11)) and (inputs(17));
    layer0_outputs(2032) <= (inputs(14)) and not (inputs(155));
    layer0_outputs(2033) <= not(inputs(204)) or (inputs(95));
    layer0_outputs(2034) <= not(inputs(126));
    layer0_outputs(2035) <= inputs(108);
    layer0_outputs(2036) <= (inputs(212)) and not (inputs(14));
    layer0_outputs(2037) <= (inputs(161)) xor (inputs(104));
    layer0_outputs(2038) <= (inputs(74)) and not (inputs(23));
    layer0_outputs(2039) <= inputs(146);
    layer0_outputs(2040) <= (inputs(202)) or (inputs(0));
    layer0_outputs(2041) <= not(inputs(215));
    layer0_outputs(2042) <= not((inputs(184)) or (inputs(173)));
    layer0_outputs(2043) <= inputs(43);
    layer0_outputs(2044) <= not((inputs(172)) or (inputs(160)));
    layer0_outputs(2045) <= not(inputs(99)) or (inputs(245));
    layer0_outputs(2046) <= not((inputs(138)) xor (inputs(164)));
    layer0_outputs(2047) <= inputs(183);
    layer0_outputs(2048) <= not((inputs(250)) xor (inputs(201)));
    layer0_outputs(2049) <= not(inputs(164));
    layer0_outputs(2050) <= not(inputs(67)) or (inputs(19));
    layer0_outputs(2051) <= not(inputs(249));
    layer0_outputs(2052) <= not(inputs(210));
    layer0_outputs(2053) <= (inputs(115)) or (inputs(105));
    layer0_outputs(2054) <= (inputs(219)) or (inputs(173));
    layer0_outputs(2055) <= not((inputs(114)) or (inputs(104)));
    layer0_outputs(2056) <= inputs(189);
    layer0_outputs(2057) <= (inputs(210)) xor (inputs(26));
    layer0_outputs(2058) <= not((inputs(10)) xor (inputs(54)));
    layer0_outputs(2059) <= (inputs(136)) xor (inputs(168));
    layer0_outputs(2060) <= not(inputs(246)) or (inputs(114));
    layer0_outputs(2061) <= (inputs(138)) and (inputs(121));
    layer0_outputs(2062) <= not(inputs(79));
    layer0_outputs(2063) <= (inputs(15)) or (inputs(249));
    layer0_outputs(2064) <= not((inputs(56)) xor (inputs(20)));
    layer0_outputs(2065) <= (inputs(14)) xor (inputs(223));
    layer0_outputs(2066) <= inputs(91);
    layer0_outputs(2067) <= not((inputs(154)) or (inputs(105)));
    layer0_outputs(2068) <= not(inputs(135));
    layer0_outputs(2069) <= inputs(191);
    layer0_outputs(2070) <= (inputs(231)) and not (inputs(214));
    layer0_outputs(2071) <= (inputs(69)) xor (inputs(99));
    layer0_outputs(2072) <= not(inputs(60));
    layer0_outputs(2073) <= not((inputs(80)) or (inputs(23)));
    layer0_outputs(2074) <= not(inputs(47));
    layer0_outputs(2075) <= inputs(220);
    layer0_outputs(2076) <= not((inputs(204)) xor (inputs(218)));
    layer0_outputs(2077) <= (inputs(144)) or (inputs(49));
    layer0_outputs(2078) <= (inputs(16)) xor (inputs(117));
    layer0_outputs(2079) <= (inputs(47)) or (inputs(246));
    layer0_outputs(2080) <= inputs(26);
    layer0_outputs(2081) <= (inputs(127)) xor (inputs(177));
    layer0_outputs(2082) <= (inputs(110)) or (inputs(236));
    layer0_outputs(2083) <= (inputs(59)) xor (inputs(33));
    layer0_outputs(2084) <= not(inputs(92));
    layer0_outputs(2085) <= (inputs(101)) or (inputs(30));
    layer0_outputs(2086) <= not((inputs(18)) or (inputs(244)));
    layer0_outputs(2087) <= not(inputs(162));
    layer0_outputs(2088) <= inputs(130);
    layer0_outputs(2089) <= not(inputs(97)) or (inputs(46));
    layer0_outputs(2090) <= (inputs(110)) or (inputs(27));
    layer0_outputs(2091) <= (inputs(85)) or (inputs(106));
    layer0_outputs(2092) <= not(inputs(182));
    layer0_outputs(2093) <= not(inputs(72)) or (inputs(54));
    layer0_outputs(2094) <= not((inputs(221)) xor (inputs(28)));
    layer0_outputs(2095) <= (inputs(141)) or (inputs(70));
    layer0_outputs(2096) <= (inputs(255)) and (inputs(222));
    layer0_outputs(2097) <= inputs(21);
    layer0_outputs(2098) <= not(inputs(132));
    layer0_outputs(2099) <= not(inputs(89)) or (inputs(1));
    layer0_outputs(2100) <= (inputs(12)) xor (inputs(232));
    layer0_outputs(2101) <= not(inputs(13)) or (inputs(255));
    layer0_outputs(2102) <= (inputs(118)) or (inputs(32));
    layer0_outputs(2103) <= not(inputs(177)) or (inputs(48));
    layer0_outputs(2104) <= not((inputs(79)) xor (inputs(252)));
    layer0_outputs(2105) <= (inputs(152)) and not (inputs(41));
    layer0_outputs(2106) <= inputs(21);
    layer0_outputs(2107) <= (inputs(66)) xor (inputs(8));
    layer0_outputs(2108) <= (inputs(116)) xor (inputs(130));
    layer0_outputs(2109) <= (inputs(83)) or (inputs(110));
    layer0_outputs(2110) <= not(inputs(107)) or (inputs(180));
    layer0_outputs(2111) <= not((inputs(80)) or (inputs(190)));
    layer0_outputs(2112) <= not((inputs(243)) or (inputs(209)));
    layer0_outputs(2113) <= (inputs(26)) and (inputs(23));
    layer0_outputs(2114) <= (inputs(248)) and (inputs(247));
    layer0_outputs(2115) <= not(inputs(50)) or (inputs(33));
    layer0_outputs(2116) <= not(inputs(109));
    layer0_outputs(2117) <= (inputs(44)) or (inputs(153));
    layer0_outputs(2118) <= (inputs(32)) or (inputs(15));
    layer0_outputs(2119) <= (inputs(85)) and not (inputs(212));
    layer0_outputs(2120) <= inputs(245);
    layer0_outputs(2121) <= not(inputs(220));
    layer0_outputs(2122) <= not((inputs(127)) xor (inputs(189)));
    layer0_outputs(2123) <= (inputs(51)) and (inputs(13));
    layer0_outputs(2124) <= (inputs(53)) and not (inputs(79));
    layer0_outputs(2125) <= (inputs(241)) or (inputs(172));
    layer0_outputs(2126) <= not((inputs(103)) or (inputs(72)));
    layer0_outputs(2127) <= not(inputs(188));
    layer0_outputs(2128) <= not((inputs(92)) and (inputs(226)));
    layer0_outputs(2129) <= not((inputs(112)) or (inputs(144)));
    layer0_outputs(2130) <= not((inputs(241)) xor (inputs(210)));
    layer0_outputs(2131) <= inputs(91);
    layer0_outputs(2132) <= (inputs(119)) and not (inputs(155));
    layer0_outputs(2133) <= inputs(130);
    layer0_outputs(2134) <= not((inputs(141)) xor (inputs(74)));
    layer0_outputs(2135) <= not(inputs(25));
    layer0_outputs(2136) <= not((inputs(161)) xor (inputs(176)));
    layer0_outputs(2137) <= not((inputs(53)) and (inputs(24)));
    layer0_outputs(2138) <= inputs(177);
    layer0_outputs(2139) <= inputs(52);
    layer0_outputs(2140) <= (inputs(91)) and not (inputs(149));
    layer0_outputs(2141) <= (inputs(170)) xor (inputs(203));
    layer0_outputs(2142) <= not(inputs(119));
    layer0_outputs(2143) <= not(inputs(49)) or (inputs(11));
    layer0_outputs(2144) <= not(inputs(138)) or (inputs(94));
    layer0_outputs(2145) <= (inputs(162)) or (inputs(213));
    layer0_outputs(2146) <= not((inputs(8)) or (inputs(28)));
    layer0_outputs(2147) <= (inputs(85)) xor (inputs(54));
    layer0_outputs(2148) <= (inputs(65)) xor (inputs(86));
    layer0_outputs(2149) <= not((inputs(208)) and (inputs(43)));
    layer0_outputs(2150) <= not(inputs(4));
    layer0_outputs(2151) <= (inputs(220)) and not (inputs(47));
    layer0_outputs(2152) <= not(inputs(89)) or (inputs(47));
    layer0_outputs(2153) <= not(inputs(158));
    layer0_outputs(2154) <= (inputs(211)) and not (inputs(105));
    layer0_outputs(2155) <= (inputs(32)) and not (inputs(105));
    layer0_outputs(2156) <= not(inputs(206));
    layer0_outputs(2157) <= not((inputs(156)) xor (inputs(109)));
    layer0_outputs(2158) <= inputs(70);
    layer0_outputs(2159) <= inputs(179);
    layer0_outputs(2160) <= (inputs(106)) and not (inputs(11));
    layer0_outputs(2161) <= inputs(55);
    layer0_outputs(2162) <= not(inputs(210)) or (inputs(32));
    layer0_outputs(2163) <= inputs(118);
    layer0_outputs(2164) <= (inputs(105)) and not (inputs(148));
    layer0_outputs(2165) <= inputs(130);
    layer0_outputs(2166) <= (inputs(230)) and not (inputs(90));
    layer0_outputs(2167) <= inputs(44);
    layer0_outputs(2168) <= (inputs(14)) or (inputs(218));
    layer0_outputs(2169) <= not((inputs(165)) xor (inputs(240)));
    layer0_outputs(2170) <= not((inputs(146)) or (inputs(162)));
    layer0_outputs(2171) <= not((inputs(41)) or (inputs(31)));
    layer0_outputs(2172) <= inputs(146);
    layer0_outputs(2173) <= not(inputs(119));
    layer0_outputs(2174) <= (inputs(84)) and not (inputs(197));
    layer0_outputs(2175) <= inputs(138);
    layer0_outputs(2176) <= (inputs(252)) and not (inputs(191));
    layer0_outputs(2177) <= (inputs(227)) and not (inputs(64));
    layer0_outputs(2178) <= not(inputs(108));
    layer0_outputs(2179) <= (inputs(42)) and not (inputs(54));
    layer0_outputs(2180) <= inputs(101);
    layer0_outputs(2181) <= not((inputs(99)) xor (inputs(1)));
    layer0_outputs(2182) <= inputs(75);
    layer0_outputs(2183) <= (inputs(150)) or (inputs(164));
    layer0_outputs(2184) <= inputs(91);
    layer0_outputs(2185) <= (inputs(193)) or (inputs(49));
    layer0_outputs(2186) <= (inputs(83)) xor (inputs(178));
    layer0_outputs(2187) <= not(inputs(23));
    layer0_outputs(2188) <= not(inputs(157)) or (inputs(32));
    layer0_outputs(2189) <= (inputs(33)) and not (inputs(131));
    layer0_outputs(2190) <= not((inputs(205)) xor (inputs(224)));
    layer0_outputs(2191) <= (inputs(238)) xor (inputs(157));
    layer0_outputs(2192) <= not((inputs(24)) xor (inputs(196)));
    layer0_outputs(2193) <= inputs(230);
    layer0_outputs(2194) <= (inputs(144)) or (inputs(200));
    layer0_outputs(2195) <= not((inputs(4)) or (inputs(166)));
    layer0_outputs(2196) <= not((inputs(149)) xor (inputs(194)));
    layer0_outputs(2197) <= inputs(135);
    layer0_outputs(2198) <= not(inputs(233)) or (inputs(105));
    layer0_outputs(2199) <= not(inputs(246));
    layer0_outputs(2200) <= (inputs(23)) and not (inputs(180));
    layer0_outputs(2201) <= not((inputs(183)) xor (inputs(209)));
    layer0_outputs(2202) <= (inputs(205)) xor (inputs(115));
    layer0_outputs(2203) <= (inputs(73)) or (inputs(118));
    layer0_outputs(2204) <= inputs(120);
    layer0_outputs(2205) <= not((inputs(149)) or (inputs(240)));
    layer0_outputs(2206) <= not((inputs(134)) or (inputs(227)));
    layer0_outputs(2207) <= inputs(230);
    layer0_outputs(2208) <= (inputs(215)) and not (inputs(6));
    layer0_outputs(2209) <= not((inputs(36)) xor (inputs(255)));
    layer0_outputs(2210) <= not(inputs(115)) or (inputs(95));
    layer0_outputs(2211) <= inputs(42);
    layer0_outputs(2212) <= not((inputs(168)) xor (inputs(234)));
    layer0_outputs(2213) <= (inputs(156)) xor (inputs(188));
    layer0_outputs(2214) <= not(inputs(251)) or (inputs(171));
    layer0_outputs(2215) <= not((inputs(206)) or (inputs(60)));
    layer0_outputs(2216) <= not(inputs(222));
    layer0_outputs(2217) <= inputs(103);
    layer0_outputs(2218) <= inputs(232);
    layer0_outputs(2219) <= not((inputs(128)) or (inputs(230)));
    layer0_outputs(2220) <= not((inputs(208)) or (inputs(204)));
    layer0_outputs(2221) <= (inputs(5)) or (inputs(79));
    layer0_outputs(2222) <= inputs(149);
    layer0_outputs(2223) <= inputs(39);
    layer0_outputs(2224) <= (inputs(188)) and not (inputs(131));
    layer0_outputs(2225) <= not(inputs(116)) or (inputs(234));
    layer0_outputs(2226) <= not((inputs(16)) xor (inputs(210)));
    layer0_outputs(2227) <= not(inputs(146));
    layer0_outputs(2228) <= not((inputs(254)) or (inputs(88)));
    layer0_outputs(2229) <= (inputs(138)) or (inputs(57));
    layer0_outputs(2230) <= not((inputs(168)) xor (inputs(138)));
    layer0_outputs(2231) <= not((inputs(99)) or (inputs(15)));
    layer0_outputs(2232) <= inputs(142);
    layer0_outputs(2233) <= inputs(233);
    layer0_outputs(2234) <= not((inputs(41)) or (inputs(127)));
    layer0_outputs(2235) <= not(inputs(43)) or (inputs(191));
    layer0_outputs(2236) <= not(inputs(179));
    layer0_outputs(2237) <= (inputs(81)) xor (inputs(117));
    layer0_outputs(2238) <= (inputs(123)) and not (inputs(129));
    layer0_outputs(2239) <= not(inputs(177));
    layer0_outputs(2240) <= inputs(236);
    layer0_outputs(2241) <= inputs(165);
    layer0_outputs(2242) <= not(inputs(183));
    layer0_outputs(2243) <= not(inputs(164)) or (inputs(61));
    layer0_outputs(2244) <= not(inputs(106));
    layer0_outputs(2245) <= not(inputs(234));
    layer0_outputs(2246) <= (inputs(159)) or (inputs(124));
    layer0_outputs(2247) <= (inputs(99)) and not (inputs(214));
    layer0_outputs(2248) <= not((inputs(148)) or (inputs(100)));
    layer0_outputs(2249) <= inputs(130);
    layer0_outputs(2250) <= (inputs(202)) xor (inputs(93));
    layer0_outputs(2251) <= inputs(53);
    layer0_outputs(2252) <= (inputs(156)) xor (inputs(253));
    layer0_outputs(2253) <= (inputs(21)) or (inputs(61));
    layer0_outputs(2254) <= not(inputs(60)) or (inputs(254));
    layer0_outputs(2255) <= (inputs(156)) or (inputs(23));
    layer0_outputs(2256) <= (inputs(133)) or (inputs(35));
    layer0_outputs(2257) <= inputs(164);
    layer0_outputs(2258) <= inputs(163);
    layer0_outputs(2259) <= (inputs(254)) or (inputs(93));
    layer0_outputs(2260) <= not((inputs(234)) or (inputs(110)));
    layer0_outputs(2261) <= not(inputs(162)) or (inputs(45));
    layer0_outputs(2262) <= inputs(56);
    layer0_outputs(2263) <= (inputs(27)) or (inputs(45));
    layer0_outputs(2264) <= (inputs(233)) and (inputs(119));
    layer0_outputs(2265) <= not(inputs(35)) or (inputs(214));
    layer0_outputs(2266) <= inputs(120);
    layer0_outputs(2267) <= not((inputs(161)) xor (inputs(32)));
    layer0_outputs(2268) <= (inputs(151)) and not (inputs(41));
    layer0_outputs(2269) <= (inputs(190)) xor (inputs(64));
    layer0_outputs(2270) <= not(inputs(37)) or (inputs(224));
    layer0_outputs(2271) <= inputs(100);
    layer0_outputs(2272) <= (inputs(175)) xor (inputs(62));
    layer0_outputs(2273) <= (inputs(171)) and (inputs(210));
    layer0_outputs(2274) <= not((inputs(241)) or (inputs(245)));
    layer0_outputs(2275) <= not((inputs(161)) or (inputs(255)));
    layer0_outputs(2276) <= not((inputs(45)) xor (inputs(220)));
    layer0_outputs(2277) <= (inputs(221)) xor (inputs(50));
    layer0_outputs(2278) <= (inputs(132)) or (inputs(17));
    layer0_outputs(2279) <= not((inputs(69)) xor (inputs(144)));
    layer0_outputs(2280) <= not((inputs(254)) or (inputs(237)));
    layer0_outputs(2281) <= (inputs(181)) xor (inputs(162));
    layer0_outputs(2282) <= not((inputs(233)) xor (inputs(160)));
    layer0_outputs(2283) <= inputs(60);
    layer0_outputs(2284) <= inputs(73);
    layer0_outputs(2285) <= not(inputs(196)) or (inputs(79));
    layer0_outputs(2286) <= not((inputs(111)) xor (inputs(70)));
    layer0_outputs(2287) <= inputs(98);
    layer0_outputs(2288) <= not(inputs(13));
    layer0_outputs(2289) <= (inputs(237)) and (inputs(237));
    layer0_outputs(2290) <= inputs(122);
    layer0_outputs(2291) <= (inputs(242)) xor (inputs(113));
    layer0_outputs(2292) <= inputs(125);
    layer0_outputs(2293) <= not(inputs(217));
    layer0_outputs(2294) <= (inputs(241)) or (inputs(65));
    layer0_outputs(2295) <= '1';
    layer0_outputs(2296) <= inputs(215);
    layer0_outputs(2297) <= not((inputs(80)) or (inputs(31)));
    layer0_outputs(2298) <= inputs(39);
    layer0_outputs(2299) <= not((inputs(15)) xor (inputs(97)));
    layer0_outputs(2300) <= not((inputs(220)) xor (inputs(105)));
    layer0_outputs(2301) <= (inputs(158)) and not (inputs(101));
    layer0_outputs(2302) <= (inputs(90)) and not (inputs(39));
    layer0_outputs(2303) <= not(inputs(0)) or (inputs(188));
    layer0_outputs(2304) <= not((inputs(53)) or (inputs(21)));
    layer0_outputs(2305) <= not(inputs(133));
    layer0_outputs(2306) <= (inputs(141)) xor (inputs(241));
    layer0_outputs(2307) <= not((inputs(159)) or (inputs(145)));
    layer0_outputs(2308) <= not((inputs(250)) xor (inputs(161)));
    layer0_outputs(2309) <= not((inputs(196)) and (inputs(183)));
    layer0_outputs(2310) <= (inputs(160)) or (inputs(143));
    layer0_outputs(2311) <= not(inputs(55));
    layer0_outputs(2312) <= '0';
    layer0_outputs(2313) <= not((inputs(222)) xor (inputs(226)));
    layer0_outputs(2314) <= not(inputs(161));
    layer0_outputs(2315) <= inputs(111);
    layer0_outputs(2316) <= (inputs(179)) or (inputs(20));
    layer0_outputs(2317) <= (inputs(66)) xor (inputs(107));
    layer0_outputs(2318) <= (inputs(137)) and not (inputs(128));
    layer0_outputs(2319) <= not(inputs(84));
    layer0_outputs(2320) <= inputs(177);
    layer0_outputs(2321) <= (inputs(121)) and not (inputs(161));
    layer0_outputs(2322) <= not((inputs(96)) xor (inputs(98)));
    layer0_outputs(2323) <= inputs(69);
    layer0_outputs(2324) <= not(inputs(244));
    layer0_outputs(2325) <= not(inputs(214));
    layer0_outputs(2326) <= not(inputs(245));
    layer0_outputs(2327) <= not(inputs(104)) or (inputs(174));
    layer0_outputs(2328) <= (inputs(194)) xor (inputs(244));
    layer0_outputs(2329) <= inputs(231);
    layer0_outputs(2330) <= (inputs(99)) xor (inputs(82));
    layer0_outputs(2331) <= not(inputs(232)) or (inputs(30));
    layer0_outputs(2332) <= not(inputs(107));
    layer0_outputs(2333) <= not(inputs(5));
    layer0_outputs(2334) <= not(inputs(192)) or (inputs(31));
    layer0_outputs(2335) <= (inputs(71)) and not (inputs(137));
    layer0_outputs(2336) <= (inputs(91)) xor (inputs(45));
    layer0_outputs(2337) <= inputs(125);
    layer0_outputs(2338) <= '0';
    layer0_outputs(2339) <= not(inputs(133));
    layer0_outputs(2340) <= (inputs(167)) xor (inputs(195));
    layer0_outputs(2341) <= not((inputs(0)) and (inputs(87)));
    layer0_outputs(2342) <= not((inputs(188)) or (inputs(8)));
    layer0_outputs(2343) <= not((inputs(189)) or (inputs(135)));
    layer0_outputs(2344) <= (inputs(43)) or (inputs(33));
    layer0_outputs(2345) <= not(inputs(7)) or (inputs(160));
    layer0_outputs(2346) <= inputs(81);
    layer0_outputs(2347) <= (inputs(188)) and not (inputs(75));
    layer0_outputs(2348) <= inputs(135);
    layer0_outputs(2349) <= inputs(152);
    layer0_outputs(2350) <= inputs(37);
    layer0_outputs(2351) <= inputs(88);
    layer0_outputs(2352) <= not((inputs(5)) or (inputs(21)));
    layer0_outputs(2353) <= (inputs(173)) or (inputs(243));
    layer0_outputs(2354) <= not(inputs(117)) or (inputs(7));
    layer0_outputs(2355) <= not((inputs(40)) xor (inputs(64)));
    layer0_outputs(2356) <= not((inputs(178)) or (inputs(31)));
    layer0_outputs(2357) <= not((inputs(29)) or (inputs(35)));
    layer0_outputs(2358) <= not((inputs(2)) or (inputs(59)));
    layer0_outputs(2359) <= inputs(80);
    layer0_outputs(2360) <= (inputs(60)) or (inputs(108));
    layer0_outputs(2361) <= not((inputs(172)) or (inputs(42)));
    layer0_outputs(2362) <= not(inputs(101));
    layer0_outputs(2363) <= not((inputs(151)) xor (inputs(212)));
    layer0_outputs(2364) <= not(inputs(39)) or (inputs(131));
    layer0_outputs(2365) <= not(inputs(9));
    layer0_outputs(2366) <= not(inputs(132));
    layer0_outputs(2367) <= '0';
    layer0_outputs(2368) <= not((inputs(255)) or (inputs(251)));
    layer0_outputs(2369) <= (inputs(249)) xor (inputs(0));
    layer0_outputs(2370) <= not(inputs(243));
    layer0_outputs(2371) <= (inputs(25)) and (inputs(24));
    layer0_outputs(2372) <= not(inputs(165));
    layer0_outputs(2373) <= (inputs(197)) and not (inputs(207));
    layer0_outputs(2374) <= not(inputs(239));
    layer0_outputs(2375) <= not((inputs(160)) xor (inputs(196)));
    layer0_outputs(2376) <= not(inputs(248));
    layer0_outputs(2377) <= inputs(155);
    layer0_outputs(2378) <= (inputs(111)) and not (inputs(64));
    layer0_outputs(2379) <= (inputs(191)) and not (inputs(167));
    layer0_outputs(2380) <= not(inputs(8));
    layer0_outputs(2381) <= (inputs(233)) and not (inputs(73));
    layer0_outputs(2382) <= not((inputs(40)) xor (inputs(212)));
    layer0_outputs(2383) <= not(inputs(216)) or (inputs(146));
    layer0_outputs(2384) <= (inputs(224)) or (inputs(51));
    layer0_outputs(2385) <= (inputs(125)) and (inputs(43));
    layer0_outputs(2386) <= (inputs(187)) xor (inputs(2));
    layer0_outputs(2387) <= not(inputs(213)) or (inputs(58));
    layer0_outputs(2388) <= not(inputs(19));
    layer0_outputs(2389) <= not((inputs(68)) or (inputs(111)));
    layer0_outputs(2390) <= not((inputs(33)) or (inputs(143)));
    layer0_outputs(2391) <= inputs(117);
    layer0_outputs(2392) <= (inputs(26)) and not (inputs(69));
    layer0_outputs(2393) <= not((inputs(129)) and (inputs(145)));
    layer0_outputs(2394) <= inputs(60);
    layer0_outputs(2395) <= (inputs(154)) xor (inputs(13));
    layer0_outputs(2396) <= inputs(163);
    layer0_outputs(2397) <= not(inputs(230));
    layer0_outputs(2398) <= not((inputs(222)) or (inputs(50)));
    layer0_outputs(2399) <= not((inputs(6)) or (inputs(242)));
    layer0_outputs(2400) <= not((inputs(100)) and (inputs(254)));
    layer0_outputs(2401) <= (inputs(142)) and (inputs(166));
    layer0_outputs(2402) <= (inputs(136)) xor (inputs(124));
    layer0_outputs(2403) <= (inputs(194)) or (inputs(221));
    layer0_outputs(2404) <= inputs(38);
    layer0_outputs(2405) <= (inputs(146)) or (inputs(127));
    layer0_outputs(2406) <= (inputs(245)) and not (inputs(126));
    layer0_outputs(2407) <= (inputs(189)) or (inputs(223));
    layer0_outputs(2408) <= inputs(147);
    layer0_outputs(2409) <= not((inputs(125)) or (inputs(147)));
    layer0_outputs(2410) <= (inputs(18)) or (inputs(220));
    layer0_outputs(2411) <= inputs(97);
    layer0_outputs(2412) <= (inputs(16)) xor (inputs(175));
    layer0_outputs(2413) <= inputs(252);
    layer0_outputs(2414) <= not((inputs(96)) xor (inputs(101)));
    layer0_outputs(2415) <= (inputs(40)) and not (inputs(97));
    layer0_outputs(2416) <= (inputs(26)) and (inputs(67));
    layer0_outputs(2417) <= not(inputs(203)) or (inputs(70));
    layer0_outputs(2418) <= not((inputs(185)) xor (inputs(218)));
    layer0_outputs(2419) <= not((inputs(94)) or (inputs(58)));
    layer0_outputs(2420) <= not(inputs(133)) or (inputs(214));
    layer0_outputs(2421) <= inputs(17);
    layer0_outputs(2422) <= inputs(221);
    layer0_outputs(2423) <= not((inputs(166)) or (inputs(173)));
    layer0_outputs(2424) <= (inputs(92)) or (inputs(61));
    layer0_outputs(2425) <= (inputs(182)) and not (inputs(221));
    layer0_outputs(2426) <= (inputs(144)) xor (inputs(37));
    layer0_outputs(2427) <= inputs(227);
    layer0_outputs(2428) <= not((inputs(230)) or (inputs(81)));
    layer0_outputs(2429) <= not((inputs(9)) or (inputs(207)));
    layer0_outputs(2430) <= not(inputs(214));
    layer0_outputs(2431) <= not(inputs(35));
    layer0_outputs(2432) <= not(inputs(133));
    layer0_outputs(2433) <= not((inputs(4)) or (inputs(180)));
    layer0_outputs(2434) <= not(inputs(152)) or (inputs(11));
    layer0_outputs(2435) <= not(inputs(134)) or (inputs(252));
    layer0_outputs(2436) <= not((inputs(22)) or (inputs(44)));
    layer0_outputs(2437) <= not(inputs(105)) or (inputs(144));
    layer0_outputs(2438) <= not(inputs(172)) or (inputs(151));
    layer0_outputs(2439) <= not(inputs(221));
    layer0_outputs(2440) <= inputs(64);
    layer0_outputs(2441) <= (inputs(144)) and not (inputs(254));
    layer0_outputs(2442) <= not(inputs(24)) or (inputs(98));
    layer0_outputs(2443) <= not((inputs(232)) xor (inputs(27)));
    layer0_outputs(2444) <= not((inputs(163)) or (inputs(157)));
    layer0_outputs(2445) <= not(inputs(208)) or (inputs(99));
    layer0_outputs(2446) <= not((inputs(127)) or (inputs(174)));
    layer0_outputs(2447) <= inputs(165);
    layer0_outputs(2448) <= (inputs(206)) or (inputs(8));
    layer0_outputs(2449) <= inputs(166);
    layer0_outputs(2450) <= not(inputs(219)) or (inputs(40));
    layer0_outputs(2451) <= inputs(195);
    layer0_outputs(2452) <= not(inputs(183));
    layer0_outputs(2453) <= (inputs(52)) and not (inputs(176));
    layer0_outputs(2454) <= inputs(86);
    layer0_outputs(2455) <= inputs(234);
    layer0_outputs(2456) <= not(inputs(170)) or (inputs(219));
    layer0_outputs(2457) <= not((inputs(156)) xor (inputs(113)));
    layer0_outputs(2458) <= (inputs(173)) or (inputs(50));
    layer0_outputs(2459) <= not((inputs(36)) and (inputs(168)));
    layer0_outputs(2460) <= inputs(195);
    layer0_outputs(2461) <= (inputs(203)) and not (inputs(127));
    layer0_outputs(2462) <= (inputs(55)) or (inputs(0));
    layer0_outputs(2463) <= inputs(146);
    layer0_outputs(2464) <= not((inputs(32)) and (inputs(139)));
    layer0_outputs(2465) <= not(inputs(5));
    layer0_outputs(2466) <= not((inputs(214)) and (inputs(7)));
    layer0_outputs(2467) <= (inputs(122)) or (inputs(29));
    layer0_outputs(2468) <= not(inputs(237));
    layer0_outputs(2469) <= not(inputs(118)) or (inputs(32));
    layer0_outputs(2470) <= (inputs(31)) or (inputs(106));
    layer0_outputs(2471) <= (inputs(38)) xor (inputs(134));
    layer0_outputs(2472) <= not(inputs(2));
    layer0_outputs(2473) <= inputs(55);
    layer0_outputs(2474) <= inputs(25);
    layer0_outputs(2475) <= not(inputs(26));
    layer0_outputs(2476) <= inputs(147);
    layer0_outputs(2477) <= not(inputs(78));
    layer0_outputs(2478) <= not((inputs(182)) or (inputs(132)));
    layer0_outputs(2479) <= not(inputs(39)) or (inputs(248));
    layer0_outputs(2480) <= not((inputs(87)) or (inputs(118)));
    layer0_outputs(2481) <= not((inputs(227)) or (inputs(217)));
    layer0_outputs(2482) <= (inputs(221)) xor (inputs(219));
    layer0_outputs(2483) <= (inputs(232)) xor (inputs(3));
    layer0_outputs(2484) <= not(inputs(116));
    layer0_outputs(2485) <= inputs(237);
    layer0_outputs(2486) <= inputs(88);
    layer0_outputs(2487) <= inputs(81);
    layer0_outputs(2488) <= not((inputs(114)) or (inputs(112)));
    layer0_outputs(2489) <= (inputs(60)) xor (inputs(103));
    layer0_outputs(2490) <= not(inputs(86));
    layer0_outputs(2491) <= inputs(89);
    layer0_outputs(2492) <= not((inputs(195)) xor (inputs(178)));
    layer0_outputs(2493) <= not((inputs(250)) or (inputs(174)));
    layer0_outputs(2494) <= not((inputs(6)) xor (inputs(37)));
    layer0_outputs(2495) <= not((inputs(85)) or (inputs(160)));
    layer0_outputs(2496) <= (inputs(204)) xor (inputs(235));
    layer0_outputs(2497) <= not((inputs(248)) xor (inputs(20)));
    layer0_outputs(2498) <= not(inputs(236));
    layer0_outputs(2499) <= inputs(201);
    layer0_outputs(2500) <= inputs(75);
    layer0_outputs(2501) <= (inputs(176)) or (inputs(196));
    layer0_outputs(2502) <= not((inputs(179)) or (inputs(217)));
    layer0_outputs(2503) <= not(inputs(175)) or (inputs(25));
    layer0_outputs(2504) <= not(inputs(90)) or (inputs(235));
    layer0_outputs(2505) <= not(inputs(67));
    layer0_outputs(2506) <= not((inputs(46)) xor (inputs(136)));
    layer0_outputs(2507) <= (inputs(72)) and not (inputs(51));
    layer0_outputs(2508) <= inputs(167);
    layer0_outputs(2509) <= (inputs(108)) or (inputs(97));
    layer0_outputs(2510) <= not((inputs(143)) or (inputs(132)));
    layer0_outputs(2511) <= not(inputs(90));
    layer0_outputs(2512) <= not(inputs(117));
    layer0_outputs(2513) <= (inputs(124)) or (inputs(129));
    layer0_outputs(2514) <= (inputs(20)) and not (inputs(67));
    layer0_outputs(2515) <= not(inputs(159)) or (inputs(106));
    layer0_outputs(2516) <= inputs(120);
    layer0_outputs(2517) <= not(inputs(130));
    layer0_outputs(2518) <= inputs(219);
    layer0_outputs(2519) <= inputs(93);
    layer0_outputs(2520) <= not((inputs(182)) or (inputs(184)));
    layer0_outputs(2521) <= '1';
    layer0_outputs(2522) <= not(inputs(230));
    layer0_outputs(2523) <= not((inputs(131)) or (inputs(239)));
    layer0_outputs(2524) <= not(inputs(192)) or (inputs(210));
    layer0_outputs(2525) <= not((inputs(83)) xor (inputs(54)));
    layer0_outputs(2526) <= inputs(150);
    layer0_outputs(2527) <= not(inputs(185));
    layer0_outputs(2528) <= (inputs(211)) and (inputs(112));
    layer0_outputs(2529) <= (inputs(192)) xor (inputs(164));
    layer0_outputs(2530) <= (inputs(51)) or (inputs(181));
    layer0_outputs(2531) <= inputs(88);
    layer0_outputs(2532) <= inputs(245);
    layer0_outputs(2533) <= not((inputs(85)) xor (inputs(80)));
    layer0_outputs(2534) <= '1';
    layer0_outputs(2535) <= (inputs(21)) and not (inputs(116));
    layer0_outputs(2536) <= (inputs(195)) xor (inputs(201));
    layer0_outputs(2537) <= (inputs(73)) or (inputs(255));
    layer0_outputs(2538) <= not(inputs(181)) or (inputs(222));
    layer0_outputs(2539) <= not((inputs(180)) or (inputs(57)));
    layer0_outputs(2540) <= inputs(88);
    layer0_outputs(2541) <= inputs(101);
    layer0_outputs(2542) <= not((inputs(237)) or (inputs(220)));
    layer0_outputs(2543) <= inputs(19);
    layer0_outputs(2544) <= not((inputs(29)) or (inputs(4)));
    layer0_outputs(2545) <= not((inputs(247)) xor (inputs(19)));
    layer0_outputs(2546) <= inputs(60);
    layer0_outputs(2547) <= (inputs(14)) or (inputs(235));
    layer0_outputs(2548) <= not(inputs(63)) or (inputs(161));
    layer0_outputs(2549) <= (inputs(49)) xor (inputs(96));
    layer0_outputs(2550) <= not((inputs(88)) xor (inputs(226)));
    layer0_outputs(2551) <= not(inputs(148));
    layer0_outputs(2552) <= (inputs(240)) and not (inputs(113));
    layer0_outputs(2553) <= not(inputs(178));
    layer0_outputs(2554) <= not(inputs(24)) or (inputs(240));
    layer0_outputs(2555) <= inputs(114);
    layer0_outputs(2556) <= not(inputs(61));
    layer0_outputs(2557) <= not(inputs(169)) or (inputs(85));
    layer0_outputs(2558) <= not((inputs(29)) or (inputs(156)));
    layer0_outputs(2559) <= not(inputs(23));
    layer0_outputs(2560) <= not(inputs(235)) or (inputs(132));
    layer0_outputs(2561) <= (inputs(123)) and not (inputs(180));
    layer0_outputs(2562) <= (inputs(41)) or (inputs(4));
    layer0_outputs(2563) <= not((inputs(195)) xor (inputs(151)));
    layer0_outputs(2564) <= not(inputs(178)) or (inputs(153));
    layer0_outputs(2565) <= (inputs(181)) and not (inputs(253));
    layer0_outputs(2566) <= inputs(56);
    layer0_outputs(2567) <= inputs(6);
    layer0_outputs(2568) <= inputs(108);
    layer0_outputs(2569) <= (inputs(210)) or (inputs(78));
    layer0_outputs(2570) <= not((inputs(102)) or (inputs(219)));
    layer0_outputs(2571) <= (inputs(99)) and not (inputs(174));
    layer0_outputs(2572) <= inputs(38);
    layer0_outputs(2573) <= (inputs(158)) and not (inputs(11));
    layer0_outputs(2574) <= (inputs(37)) xor (inputs(45));
    layer0_outputs(2575) <= not(inputs(177)) or (inputs(14));
    layer0_outputs(2576) <= not(inputs(116)) or (inputs(38));
    layer0_outputs(2577) <= (inputs(126)) xor (inputs(210));
    layer0_outputs(2578) <= not((inputs(19)) or (inputs(42)));
    layer0_outputs(2579) <= not((inputs(97)) or (inputs(70)));
    layer0_outputs(2580) <= not(inputs(18));
    layer0_outputs(2581) <= (inputs(115)) and not (inputs(93));
    layer0_outputs(2582) <= not(inputs(165));
    layer0_outputs(2583) <= inputs(128);
    layer0_outputs(2584) <= not((inputs(247)) or (inputs(98)));
    layer0_outputs(2585) <= inputs(112);
    layer0_outputs(2586) <= not((inputs(173)) xor (inputs(160)));
    layer0_outputs(2587) <= (inputs(120)) and (inputs(106));
    layer0_outputs(2588) <= not((inputs(95)) or (inputs(113)));
    layer0_outputs(2589) <= not((inputs(28)) or (inputs(214)));
    layer0_outputs(2590) <= (inputs(125)) xor (inputs(44));
    layer0_outputs(2591) <= (inputs(156)) or (inputs(245));
    layer0_outputs(2592) <= not(inputs(103));
    layer0_outputs(2593) <= (inputs(180)) and not (inputs(124));
    layer0_outputs(2594) <= not(inputs(115)) or (inputs(55));
    layer0_outputs(2595) <= (inputs(5)) and not (inputs(0));
    layer0_outputs(2596) <= inputs(129);
    layer0_outputs(2597) <= not(inputs(85));
    layer0_outputs(2598) <= (inputs(223)) and not (inputs(160));
    layer0_outputs(2599) <= inputs(94);
    layer0_outputs(2600) <= not((inputs(164)) or (inputs(216)));
    layer0_outputs(2601) <= not((inputs(178)) or (inputs(124)));
    layer0_outputs(2602) <= (inputs(29)) and not (inputs(241));
    layer0_outputs(2603) <= inputs(118);
    layer0_outputs(2604) <= not(inputs(13)) or (inputs(126));
    layer0_outputs(2605) <= inputs(236);
    layer0_outputs(2606) <= (inputs(183)) xor (inputs(118));
    layer0_outputs(2607) <= not(inputs(33)) or (inputs(109));
    layer0_outputs(2608) <= (inputs(178)) and not (inputs(190));
    layer0_outputs(2609) <= inputs(109);
    layer0_outputs(2610) <= inputs(17);
    layer0_outputs(2611) <= not((inputs(112)) or (inputs(228)));
    layer0_outputs(2612) <= (inputs(78)) xor (inputs(6));
    layer0_outputs(2613) <= not((inputs(161)) or (inputs(229)));
    layer0_outputs(2614) <= not(inputs(68));
    layer0_outputs(2615) <= not((inputs(139)) xor (inputs(16)));
    layer0_outputs(2616) <= (inputs(172)) and (inputs(49));
    layer0_outputs(2617) <= (inputs(247)) xor (inputs(155));
    layer0_outputs(2618) <= not(inputs(211));
    layer0_outputs(2619) <= not(inputs(6)) or (inputs(251));
    layer0_outputs(2620) <= not((inputs(170)) xor (inputs(173)));
    layer0_outputs(2621) <= not(inputs(59));
    layer0_outputs(2622) <= (inputs(72)) and not (inputs(2));
    layer0_outputs(2623) <= (inputs(168)) and not (inputs(44));
    layer0_outputs(2624) <= not(inputs(98));
    layer0_outputs(2625) <= (inputs(217)) or (inputs(106));
    layer0_outputs(2626) <= inputs(237);
    layer0_outputs(2627) <= not((inputs(95)) or (inputs(6)));
    layer0_outputs(2628) <= (inputs(139)) and not (inputs(133));
    layer0_outputs(2629) <= (inputs(61)) xor (inputs(141));
    layer0_outputs(2630) <= (inputs(222)) or (inputs(189));
    layer0_outputs(2631) <= (inputs(201)) and (inputs(42));
    layer0_outputs(2632) <= not((inputs(84)) or (inputs(183)));
    layer0_outputs(2633) <= not(inputs(86));
    layer0_outputs(2634) <= not((inputs(230)) or (inputs(179)));
    layer0_outputs(2635) <= (inputs(174)) and not (inputs(94));
    layer0_outputs(2636) <= not((inputs(77)) xor (inputs(3)));
    layer0_outputs(2637) <= (inputs(53)) or (inputs(137));
    layer0_outputs(2638) <= (inputs(134)) and not (inputs(250));
    layer0_outputs(2639) <= not((inputs(121)) xor (inputs(251)));
    layer0_outputs(2640) <= not((inputs(5)) or (inputs(2)));
    layer0_outputs(2641) <= (inputs(1)) xor (inputs(70));
    layer0_outputs(2642) <= (inputs(128)) or (inputs(202));
    layer0_outputs(2643) <= inputs(131);
    layer0_outputs(2644) <= not(inputs(184));
    layer0_outputs(2645) <= not((inputs(176)) or (inputs(4)));
    layer0_outputs(2646) <= (inputs(59)) or (inputs(55));
    layer0_outputs(2647) <= inputs(115);
    layer0_outputs(2648) <= not(inputs(121)) or (inputs(164));
    layer0_outputs(2649) <= not(inputs(27));
    layer0_outputs(2650) <= not(inputs(22));
    layer0_outputs(2651) <= '1';
    layer0_outputs(2652) <= not(inputs(97));
    layer0_outputs(2653) <= (inputs(236)) or (inputs(55));
    layer0_outputs(2654) <= not((inputs(169)) xor (inputs(11)));
    layer0_outputs(2655) <= (inputs(96)) and not (inputs(28));
    layer0_outputs(2656) <= '0';
    layer0_outputs(2657) <= not((inputs(134)) and (inputs(163)));
    layer0_outputs(2658) <= (inputs(85)) xor (inputs(73));
    layer0_outputs(2659) <= (inputs(169)) xor (inputs(148));
    layer0_outputs(2660) <= (inputs(188)) or (inputs(93));
    layer0_outputs(2661) <= (inputs(176)) xor (inputs(27));
    layer0_outputs(2662) <= not(inputs(235)) or (inputs(127));
    layer0_outputs(2663) <= inputs(21);
    layer0_outputs(2664) <= not(inputs(209));
    layer0_outputs(2665) <= (inputs(126)) xor (inputs(5));
    layer0_outputs(2666) <= not(inputs(84));
    layer0_outputs(2667) <= not((inputs(76)) or (inputs(57)));
    layer0_outputs(2668) <= not(inputs(70)) or (inputs(221));
    layer0_outputs(2669) <= (inputs(175)) or (inputs(221));
    layer0_outputs(2670) <= not((inputs(92)) and (inputs(76)));
    layer0_outputs(2671) <= (inputs(45)) or (inputs(223));
    layer0_outputs(2672) <= not(inputs(197));
    layer0_outputs(2673) <= not(inputs(42));
    layer0_outputs(2674) <= (inputs(249)) or (inputs(245));
    layer0_outputs(2675) <= (inputs(137)) and not (inputs(146));
    layer0_outputs(2676) <= (inputs(15)) and not (inputs(185));
    layer0_outputs(2677) <= not((inputs(181)) xor (inputs(119)));
    layer0_outputs(2678) <= (inputs(233)) and not (inputs(166));
    layer0_outputs(2679) <= (inputs(80)) or (inputs(81));
    layer0_outputs(2680) <= not(inputs(82));
    layer0_outputs(2681) <= (inputs(21)) and not (inputs(183));
    layer0_outputs(2682) <= not((inputs(177)) or (inputs(111)));
    layer0_outputs(2683) <= not((inputs(246)) or (inputs(173)));
    layer0_outputs(2684) <= not((inputs(235)) xor (inputs(204)));
    layer0_outputs(2685) <= (inputs(70)) xor (inputs(18));
    layer0_outputs(2686) <= not((inputs(35)) xor (inputs(140)));
    layer0_outputs(2687) <= (inputs(100)) and not (inputs(173));
    layer0_outputs(2688) <= (inputs(22)) and not (inputs(253));
    layer0_outputs(2689) <= inputs(114);
    layer0_outputs(2690) <= inputs(177);
    layer0_outputs(2691) <= not((inputs(85)) or (inputs(68)));
    layer0_outputs(2692) <= not(inputs(230)) or (inputs(182));
    layer0_outputs(2693) <= not(inputs(241));
    layer0_outputs(2694) <= (inputs(84)) or (inputs(138));
    layer0_outputs(2695) <= inputs(73);
    layer0_outputs(2696) <= not(inputs(103));
    layer0_outputs(2697) <= inputs(192);
    layer0_outputs(2698) <= not((inputs(154)) or (inputs(14)));
    layer0_outputs(2699) <= (inputs(105)) or (inputs(243));
    layer0_outputs(2700) <= not(inputs(170)) or (inputs(127));
    layer0_outputs(2701) <= not(inputs(57)) or (inputs(107));
    layer0_outputs(2702) <= not(inputs(154));
    layer0_outputs(2703) <= inputs(20);
    layer0_outputs(2704) <= not((inputs(250)) xor (inputs(155)));
    layer0_outputs(2705) <= (inputs(173)) and (inputs(173));
    layer0_outputs(2706) <= (inputs(3)) or (inputs(158));
    layer0_outputs(2707) <= inputs(15);
    layer0_outputs(2708) <= (inputs(221)) and (inputs(198));
    layer0_outputs(2709) <= not((inputs(133)) or (inputs(149)));
    layer0_outputs(2710) <= not((inputs(21)) xor (inputs(170)));
    layer0_outputs(2711) <= inputs(103);
    layer0_outputs(2712) <= not((inputs(35)) xor (inputs(54)));
    layer0_outputs(2713) <= not(inputs(244));
    layer0_outputs(2714) <= (inputs(240)) and not (inputs(1));
    layer0_outputs(2715) <= not((inputs(106)) xor (inputs(43)));
    layer0_outputs(2716) <= not((inputs(5)) or (inputs(161)));
    layer0_outputs(2717) <= inputs(250);
    layer0_outputs(2718) <= (inputs(153)) or (inputs(16));
    layer0_outputs(2719) <= (inputs(131)) or (inputs(132));
    layer0_outputs(2720) <= '0';
    layer0_outputs(2721) <= (inputs(44)) xor (inputs(133));
    layer0_outputs(2722) <= (inputs(4)) xor (inputs(240));
    layer0_outputs(2723) <= not(inputs(30)) or (inputs(192));
    layer0_outputs(2724) <= not(inputs(238)) or (inputs(130));
    layer0_outputs(2725) <= (inputs(4)) and (inputs(185));
    layer0_outputs(2726) <= inputs(57);
    layer0_outputs(2727) <= not((inputs(39)) and (inputs(10)));
    layer0_outputs(2728) <= (inputs(73)) or (inputs(96));
    layer0_outputs(2729) <= inputs(231);
    layer0_outputs(2730) <= not(inputs(128));
    layer0_outputs(2731) <= (inputs(118)) and not (inputs(196));
    layer0_outputs(2732) <= (inputs(91)) xor (inputs(157));
    layer0_outputs(2733) <= not(inputs(165)) or (inputs(64));
    layer0_outputs(2734) <= not((inputs(28)) xor (inputs(30)));
    layer0_outputs(2735) <= inputs(133);
    layer0_outputs(2736) <= (inputs(162)) or (inputs(196));
    layer0_outputs(2737) <= not(inputs(236)) or (inputs(235));
    layer0_outputs(2738) <= not(inputs(150)) or (inputs(52));
    layer0_outputs(2739) <= (inputs(42)) and (inputs(68));
    layer0_outputs(2740) <= not((inputs(201)) or (inputs(6)));
    layer0_outputs(2741) <= not((inputs(116)) xor (inputs(248)));
    layer0_outputs(2742) <= (inputs(233)) and not (inputs(202));
    layer0_outputs(2743) <= not(inputs(167)) or (inputs(62));
    layer0_outputs(2744) <= inputs(243);
    layer0_outputs(2745) <= inputs(180);
    layer0_outputs(2746) <= (inputs(25)) and (inputs(11));
    layer0_outputs(2747) <= (inputs(224)) or (inputs(192));
    layer0_outputs(2748) <= not((inputs(53)) and (inputs(52)));
    layer0_outputs(2749) <= not((inputs(177)) or (inputs(210)));
    layer0_outputs(2750) <= (inputs(98)) and not (inputs(143));
    layer0_outputs(2751) <= not(inputs(30));
    layer0_outputs(2752) <= (inputs(243)) xor (inputs(248));
    layer0_outputs(2753) <= not((inputs(202)) xor (inputs(48)));
    layer0_outputs(2754) <= inputs(135);
    layer0_outputs(2755) <= (inputs(3)) and not (inputs(28));
    layer0_outputs(2756) <= not((inputs(28)) or (inputs(189)));
    layer0_outputs(2757) <= not((inputs(128)) or (inputs(69)));
    layer0_outputs(2758) <= not(inputs(113));
    layer0_outputs(2759) <= (inputs(236)) xor (inputs(246));
    layer0_outputs(2760) <= inputs(139);
    layer0_outputs(2761) <= (inputs(2)) or (inputs(159));
    layer0_outputs(2762) <= inputs(105);
    layer0_outputs(2763) <= not((inputs(135)) xor (inputs(89)));
    layer0_outputs(2764) <= not((inputs(124)) xor (inputs(160)));
    layer0_outputs(2765) <= (inputs(101)) and not (inputs(55));
    layer0_outputs(2766) <= not((inputs(122)) or (inputs(39)));
    layer0_outputs(2767) <= not((inputs(14)) or (inputs(15)));
    layer0_outputs(2768) <= not(inputs(136));
    layer0_outputs(2769) <= inputs(228);
    layer0_outputs(2770) <= not((inputs(211)) or (inputs(4)));
    layer0_outputs(2771) <= (inputs(54)) or (inputs(245));
    layer0_outputs(2772) <= not((inputs(124)) or (inputs(50)));
    layer0_outputs(2773) <= not((inputs(172)) xor (inputs(245)));
    layer0_outputs(2774) <= inputs(99);
    layer0_outputs(2775) <= not((inputs(40)) or (inputs(55)));
    layer0_outputs(2776) <= not(inputs(45));
    layer0_outputs(2777) <= not((inputs(177)) or (inputs(76)));
    layer0_outputs(2778) <= (inputs(158)) or (inputs(151));
    layer0_outputs(2779) <= not((inputs(162)) or (inputs(186)));
    layer0_outputs(2780) <= inputs(217);
    layer0_outputs(2781) <= not(inputs(21));
    layer0_outputs(2782) <= not((inputs(80)) or (inputs(67)));
    layer0_outputs(2783) <= (inputs(246)) xor (inputs(171));
    layer0_outputs(2784) <= (inputs(13)) or (inputs(252));
    layer0_outputs(2785) <= inputs(167);
    layer0_outputs(2786) <= (inputs(38)) xor (inputs(192));
    layer0_outputs(2787) <= (inputs(182)) and not (inputs(31));
    layer0_outputs(2788) <= '0';
    layer0_outputs(2789) <= not((inputs(230)) xor (inputs(24)));
    layer0_outputs(2790) <= (inputs(0)) xor (inputs(95));
    layer0_outputs(2791) <= not(inputs(126));
    layer0_outputs(2792) <= not(inputs(51)) or (inputs(31));
    layer0_outputs(2793) <= inputs(53);
    layer0_outputs(2794) <= not((inputs(74)) or (inputs(50)));
    layer0_outputs(2795) <= (inputs(169)) and not (inputs(195));
    layer0_outputs(2796) <= not(inputs(22));
    layer0_outputs(2797) <= (inputs(196)) and not (inputs(51));
    layer0_outputs(2798) <= inputs(114);
    layer0_outputs(2799) <= not((inputs(166)) and (inputs(215)));
    layer0_outputs(2800) <= not(inputs(146));
    layer0_outputs(2801) <= not(inputs(202));
    layer0_outputs(2802) <= inputs(192);
    layer0_outputs(2803) <= not(inputs(191)) or (inputs(216));
    layer0_outputs(2804) <= not((inputs(253)) xor (inputs(62)));
    layer0_outputs(2805) <= inputs(45);
    layer0_outputs(2806) <= (inputs(109)) xor (inputs(14));
    layer0_outputs(2807) <= '0';
    layer0_outputs(2808) <= not(inputs(41));
    layer0_outputs(2809) <= inputs(78);
    layer0_outputs(2810) <= (inputs(26)) and not (inputs(209));
    layer0_outputs(2811) <= (inputs(250)) or (inputs(210));
    layer0_outputs(2812) <= not((inputs(125)) and (inputs(58)));
    layer0_outputs(2813) <= not((inputs(36)) xor (inputs(211)));
    layer0_outputs(2814) <= not(inputs(59));
    layer0_outputs(2815) <= inputs(117);
    layer0_outputs(2816) <= not((inputs(209)) or (inputs(235)));
    layer0_outputs(2817) <= not(inputs(245));
    layer0_outputs(2818) <= not((inputs(54)) or (inputs(230)));
    layer0_outputs(2819) <= not((inputs(219)) xor (inputs(123)));
    layer0_outputs(2820) <= not(inputs(120));
    layer0_outputs(2821) <= not((inputs(106)) or (inputs(89)));
    layer0_outputs(2822) <= not((inputs(130)) or (inputs(129)));
    layer0_outputs(2823) <= not(inputs(110));
    layer0_outputs(2824) <= not(inputs(184));
    layer0_outputs(2825) <= inputs(136);
    layer0_outputs(2826) <= not(inputs(168)) or (inputs(175));
    layer0_outputs(2827) <= '1';
    layer0_outputs(2828) <= inputs(21);
    layer0_outputs(2829) <= (inputs(221)) or (inputs(138));
    layer0_outputs(2830) <= not((inputs(215)) and (inputs(183)));
    layer0_outputs(2831) <= not(inputs(63));
    layer0_outputs(2832) <= not((inputs(12)) or (inputs(65)));
    layer0_outputs(2833) <= not((inputs(99)) xor (inputs(239)));
    layer0_outputs(2834) <= (inputs(204)) or (inputs(233));
    layer0_outputs(2835) <= inputs(162);
    layer0_outputs(2836) <= not(inputs(39));
    layer0_outputs(2837) <= (inputs(233)) xor (inputs(41));
    layer0_outputs(2838) <= not(inputs(24)) or (inputs(147));
    layer0_outputs(2839) <= not(inputs(101));
    layer0_outputs(2840) <= not((inputs(65)) xor (inputs(149)));
    layer0_outputs(2841) <= not(inputs(70));
    layer0_outputs(2842) <= not((inputs(75)) xor (inputs(142)));
    layer0_outputs(2843) <= (inputs(123)) or (inputs(34));
    layer0_outputs(2844) <= inputs(40);
    layer0_outputs(2845) <= inputs(212);
    layer0_outputs(2846) <= not(inputs(6)) or (inputs(63));
    layer0_outputs(2847) <= not((inputs(205)) xor (inputs(25)));
    layer0_outputs(2848) <= not((inputs(10)) or (inputs(214)));
    layer0_outputs(2849) <= not(inputs(177)) or (inputs(68));
    layer0_outputs(2850) <= not(inputs(240));
    layer0_outputs(2851) <= not((inputs(230)) or (inputs(190)));
    layer0_outputs(2852) <= (inputs(242)) xor (inputs(12));
    layer0_outputs(2853) <= not((inputs(117)) xor (inputs(67)));
    layer0_outputs(2854) <= inputs(136);
    layer0_outputs(2855) <= not(inputs(172));
    layer0_outputs(2856) <= (inputs(230)) xor (inputs(90));
    layer0_outputs(2857) <= (inputs(26)) or (inputs(205));
    layer0_outputs(2858) <= (inputs(189)) xor (inputs(118));
    layer0_outputs(2859) <= (inputs(91)) or (inputs(144));
    layer0_outputs(2860) <= (inputs(231)) xor (inputs(53));
    layer0_outputs(2861) <= inputs(172);
    layer0_outputs(2862) <= inputs(146);
    layer0_outputs(2863) <= not(inputs(60));
    layer0_outputs(2864) <= not((inputs(71)) xor (inputs(202)));
    layer0_outputs(2865) <= inputs(236);
    layer0_outputs(2866) <= not(inputs(233)) or (inputs(124));
    layer0_outputs(2867) <= not(inputs(225));
    layer0_outputs(2868) <= (inputs(80)) xor (inputs(84));
    layer0_outputs(2869) <= (inputs(17)) or (inputs(44));
    layer0_outputs(2870) <= not((inputs(69)) or (inputs(228)));
    layer0_outputs(2871) <= inputs(164);
    layer0_outputs(2872) <= not(inputs(13)) or (inputs(12));
    layer0_outputs(2873) <= (inputs(48)) and not (inputs(148));
    layer0_outputs(2874) <= (inputs(171)) xor (inputs(3));
    layer0_outputs(2875) <= (inputs(201)) or (inputs(191));
    layer0_outputs(2876) <= not((inputs(38)) xor (inputs(88)));
    layer0_outputs(2877) <= not((inputs(162)) or (inputs(49)));
    layer0_outputs(2878) <= inputs(144);
    layer0_outputs(2879) <= (inputs(17)) or (inputs(201));
    layer0_outputs(2880) <= not((inputs(2)) or (inputs(128)));
    layer0_outputs(2881) <= not(inputs(221));
    layer0_outputs(2882) <= not((inputs(10)) xor (inputs(65)));
    layer0_outputs(2883) <= not(inputs(24));
    layer0_outputs(2884) <= not((inputs(29)) xor (inputs(123)));
    layer0_outputs(2885) <= inputs(26);
    layer0_outputs(2886) <= not(inputs(92));
    layer0_outputs(2887) <= (inputs(123)) xor (inputs(148));
    layer0_outputs(2888) <= (inputs(69)) and not (inputs(3));
    layer0_outputs(2889) <= (inputs(116)) xor (inputs(172));
    layer0_outputs(2890) <= not(inputs(102)) or (inputs(5));
    layer0_outputs(2891) <= not((inputs(143)) or (inputs(155)));
    layer0_outputs(2892) <= not((inputs(146)) or (inputs(10)));
    layer0_outputs(2893) <= (inputs(93)) or (inputs(59));
    layer0_outputs(2894) <= not((inputs(102)) xor (inputs(76)));
    layer0_outputs(2895) <= (inputs(94)) and not (inputs(57));
    layer0_outputs(2896) <= not(inputs(178));
    layer0_outputs(2897) <= not(inputs(176)) or (inputs(252));
    layer0_outputs(2898) <= inputs(151);
    layer0_outputs(2899) <= not(inputs(242)) or (inputs(102));
    layer0_outputs(2900) <= not(inputs(110));
    layer0_outputs(2901) <= (inputs(121)) and not (inputs(185));
    layer0_outputs(2902) <= (inputs(4)) xor (inputs(76));
    layer0_outputs(2903) <= not((inputs(80)) or (inputs(100)));
    layer0_outputs(2904) <= (inputs(29)) or (inputs(154));
    layer0_outputs(2905) <= not((inputs(114)) or (inputs(15)));
    layer0_outputs(2906) <= not((inputs(89)) and (inputs(7)));
    layer0_outputs(2907) <= (inputs(253)) or (inputs(40));
    layer0_outputs(2908) <= inputs(216);
    layer0_outputs(2909) <= not((inputs(251)) xor (inputs(48)));
    layer0_outputs(2910) <= not(inputs(236));
    layer0_outputs(2911) <= not((inputs(142)) or (inputs(187)));
    layer0_outputs(2912) <= not((inputs(229)) or (inputs(190)));
    layer0_outputs(2913) <= (inputs(57)) and not (inputs(112));
    layer0_outputs(2914) <= inputs(9);
    layer0_outputs(2915) <= not(inputs(237));
    layer0_outputs(2916) <= not(inputs(42));
    layer0_outputs(2917) <= not(inputs(69)) or (inputs(62));
    layer0_outputs(2918) <= (inputs(42)) and (inputs(121));
    layer0_outputs(2919) <= (inputs(33)) or (inputs(232));
    layer0_outputs(2920) <= (inputs(110)) or (inputs(156));
    layer0_outputs(2921) <= not((inputs(58)) and (inputs(139)));
    layer0_outputs(2922) <= not((inputs(10)) or (inputs(231)));
    layer0_outputs(2923) <= not(inputs(39)) or (inputs(203));
    layer0_outputs(2924) <= not(inputs(6)) or (inputs(143));
    layer0_outputs(2925) <= (inputs(244)) or (inputs(131));
    layer0_outputs(2926) <= not((inputs(111)) xor (inputs(244)));
    layer0_outputs(2927) <= (inputs(221)) xor (inputs(145));
    layer0_outputs(2928) <= not((inputs(239)) or (inputs(222)));
    layer0_outputs(2929) <= inputs(101);
    layer0_outputs(2930) <= not((inputs(149)) xor (inputs(73)));
    layer0_outputs(2931) <= not(inputs(149));
    layer0_outputs(2932) <= inputs(229);
    layer0_outputs(2933) <= not(inputs(27)) or (inputs(241));
    layer0_outputs(2934) <= not(inputs(130)) or (inputs(190));
    layer0_outputs(2935) <= not((inputs(22)) xor (inputs(109)));
    layer0_outputs(2936) <= (inputs(199)) xor (inputs(69));
    layer0_outputs(2937) <= not(inputs(152)) or (inputs(64));
    layer0_outputs(2938) <= inputs(27);
    layer0_outputs(2939) <= (inputs(86)) and not (inputs(3));
    layer0_outputs(2940) <= not(inputs(78)) or (inputs(222));
    layer0_outputs(2941) <= (inputs(98)) xor (inputs(252));
    layer0_outputs(2942) <= not((inputs(63)) xor (inputs(232)));
    layer0_outputs(2943) <= not(inputs(131));
    layer0_outputs(2944) <= not((inputs(226)) or (inputs(191)));
    layer0_outputs(2945) <= (inputs(139)) xor (inputs(169));
    layer0_outputs(2946) <= not(inputs(122));
    layer0_outputs(2947) <= (inputs(125)) and (inputs(161));
    layer0_outputs(2948) <= not(inputs(19));
    layer0_outputs(2949) <= (inputs(65)) or (inputs(223));
    layer0_outputs(2950) <= (inputs(164)) xor (inputs(135));
    layer0_outputs(2951) <= inputs(30);
    layer0_outputs(2952) <= not(inputs(9));
    layer0_outputs(2953) <= not(inputs(78));
    layer0_outputs(2954) <= not(inputs(44)) or (inputs(1));
    layer0_outputs(2955) <= inputs(100);
    layer0_outputs(2956) <= not((inputs(172)) and (inputs(247)));
    layer0_outputs(2957) <= (inputs(255)) and not (inputs(51));
    layer0_outputs(2958) <= inputs(61);
    layer0_outputs(2959) <= inputs(27);
    layer0_outputs(2960) <= (inputs(178)) and not (inputs(175));
    layer0_outputs(2961) <= inputs(106);
    layer0_outputs(2962) <= not((inputs(18)) or (inputs(180)));
    layer0_outputs(2963) <= not((inputs(162)) and (inputs(223)));
    layer0_outputs(2964) <= not(inputs(1));
    layer0_outputs(2965) <= not((inputs(199)) or (inputs(32)));
    layer0_outputs(2966) <= not((inputs(192)) or (inputs(195)));
    layer0_outputs(2967) <= (inputs(168)) and (inputs(69));
    layer0_outputs(2968) <= not((inputs(170)) or (inputs(113)));
    layer0_outputs(2969) <= inputs(210);
    layer0_outputs(2970) <= not(inputs(142));
    layer0_outputs(2971) <= (inputs(116)) and not (inputs(11));
    layer0_outputs(2972) <= inputs(231);
    layer0_outputs(2973) <= (inputs(189)) or (inputs(100));
    layer0_outputs(2974) <= (inputs(128)) xor (inputs(86));
    layer0_outputs(2975) <= not(inputs(152));
    layer0_outputs(2976) <= (inputs(48)) or (inputs(233));
    layer0_outputs(2977) <= not(inputs(82));
    layer0_outputs(2978) <= not(inputs(115));
    layer0_outputs(2979) <= inputs(84);
    layer0_outputs(2980) <= not((inputs(184)) or (inputs(104)));
    layer0_outputs(2981) <= (inputs(18)) and not (inputs(173));
    layer0_outputs(2982) <= not((inputs(78)) xor (inputs(45)));
    layer0_outputs(2983) <= (inputs(86)) xor (inputs(38));
    layer0_outputs(2984) <= (inputs(199)) and not (inputs(202));
    layer0_outputs(2985) <= not(inputs(242)) or (inputs(80));
    layer0_outputs(2986) <= (inputs(239)) xor (inputs(164));
    layer0_outputs(2987) <= not(inputs(157)) or (inputs(250));
    layer0_outputs(2988) <= (inputs(60)) xor (inputs(208));
    layer0_outputs(2989) <= not((inputs(76)) xor (inputs(255)));
    layer0_outputs(2990) <= (inputs(240)) xor (inputs(10));
    layer0_outputs(2991) <= not((inputs(2)) or (inputs(136)));
    layer0_outputs(2992) <= not(inputs(148));
    layer0_outputs(2993) <= (inputs(156)) and not (inputs(156));
    layer0_outputs(2994) <= not(inputs(163)) or (inputs(248));
    layer0_outputs(2995) <= (inputs(159)) or (inputs(246));
    layer0_outputs(2996) <= not((inputs(149)) or (inputs(20)));
    layer0_outputs(2997) <= inputs(86);
    layer0_outputs(2998) <= not((inputs(53)) and (inputs(138)));
    layer0_outputs(2999) <= inputs(24);
    layer0_outputs(3000) <= not(inputs(129));
    layer0_outputs(3001) <= not((inputs(25)) xor (inputs(203)));
    layer0_outputs(3002) <= (inputs(116)) and not (inputs(64));
    layer0_outputs(3003) <= (inputs(103)) or (inputs(238));
    layer0_outputs(3004) <= inputs(87);
    layer0_outputs(3005) <= '1';
    layer0_outputs(3006) <= not((inputs(155)) xor (inputs(74)));
    layer0_outputs(3007) <= '1';
    layer0_outputs(3008) <= '0';
    layer0_outputs(3009) <= (inputs(164)) xor (inputs(184));
    layer0_outputs(3010) <= inputs(89);
    layer0_outputs(3011) <= inputs(145);
    layer0_outputs(3012) <= inputs(161);
    layer0_outputs(3013) <= not(inputs(165));
    layer0_outputs(3014) <= inputs(110);
    layer0_outputs(3015) <= inputs(252);
    layer0_outputs(3016) <= not(inputs(82)) or (inputs(175));
    layer0_outputs(3017) <= not(inputs(196));
    layer0_outputs(3018) <= inputs(231);
    layer0_outputs(3019) <= (inputs(82)) or (inputs(81));
    layer0_outputs(3020) <= (inputs(101)) or (inputs(230));
    layer0_outputs(3021) <= inputs(2);
    layer0_outputs(3022) <= not(inputs(169));
    layer0_outputs(3023) <= (inputs(212)) and not (inputs(255));
    layer0_outputs(3024) <= (inputs(112)) or (inputs(117));
    layer0_outputs(3025) <= (inputs(176)) and not (inputs(151));
    layer0_outputs(3026) <= (inputs(109)) and not (inputs(221));
    layer0_outputs(3027) <= not(inputs(199)) or (inputs(63));
    layer0_outputs(3028) <= not(inputs(60));
    layer0_outputs(3029) <= (inputs(190)) or (inputs(62));
    layer0_outputs(3030) <= inputs(223);
    layer0_outputs(3031) <= (inputs(58)) and not (inputs(253));
    layer0_outputs(3032) <= not((inputs(245)) or (inputs(128)));
    layer0_outputs(3033) <= not((inputs(214)) or (inputs(64)));
    layer0_outputs(3034) <= (inputs(169)) and (inputs(228));
    layer0_outputs(3035) <= inputs(162);
    layer0_outputs(3036) <= not(inputs(96));
    layer0_outputs(3037) <= not(inputs(72)) or (inputs(147));
    layer0_outputs(3038) <= inputs(246);
    layer0_outputs(3039) <= not(inputs(188));
    layer0_outputs(3040) <= not((inputs(17)) and (inputs(34)));
    layer0_outputs(3041) <= (inputs(45)) or (inputs(58));
    layer0_outputs(3042) <= inputs(40);
    layer0_outputs(3043) <= not((inputs(130)) or (inputs(66)));
    layer0_outputs(3044) <= not(inputs(251)) or (inputs(144));
    layer0_outputs(3045) <= (inputs(239)) or (inputs(150));
    layer0_outputs(3046) <= (inputs(134)) and not (inputs(253));
    layer0_outputs(3047) <= inputs(239);
    layer0_outputs(3048) <= (inputs(120)) and not (inputs(182));
    layer0_outputs(3049) <= (inputs(205)) xor (inputs(56));
    layer0_outputs(3050) <= (inputs(29)) xor (inputs(40));
    layer0_outputs(3051) <= not((inputs(185)) and (inputs(45)));
    layer0_outputs(3052) <= not(inputs(178));
    layer0_outputs(3053) <= (inputs(60)) or (inputs(214));
    layer0_outputs(3054) <= not((inputs(210)) xor (inputs(218)));
    layer0_outputs(3055) <= not(inputs(230));
    layer0_outputs(3056) <= not((inputs(70)) xor (inputs(85)));
    layer0_outputs(3057) <= not(inputs(196));
    layer0_outputs(3058) <= inputs(4);
    layer0_outputs(3059) <= not((inputs(117)) xor (inputs(51)));
    layer0_outputs(3060) <= inputs(61);
    layer0_outputs(3061) <= (inputs(89)) or (inputs(105));
    layer0_outputs(3062) <= not((inputs(226)) xor (inputs(133)));
    layer0_outputs(3063) <= not(inputs(248)) or (inputs(90));
    layer0_outputs(3064) <= (inputs(248)) and not (inputs(4));
    layer0_outputs(3065) <= not((inputs(174)) xor (inputs(228)));
    layer0_outputs(3066) <= '1';
    layer0_outputs(3067) <= inputs(120);
    layer0_outputs(3068) <= not(inputs(142));
    layer0_outputs(3069) <= not((inputs(133)) or (inputs(128)));
    layer0_outputs(3070) <= (inputs(248)) and not (inputs(98));
    layer0_outputs(3071) <= not((inputs(164)) xor (inputs(98)));
    layer0_outputs(3072) <= (inputs(218)) or (inputs(239));
    layer0_outputs(3073) <= not(inputs(19));
    layer0_outputs(3074) <= (inputs(167)) and not (inputs(176));
    layer0_outputs(3075) <= (inputs(201)) and not (inputs(111));
    layer0_outputs(3076) <= not(inputs(29));
    layer0_outputs(3077) <= not(inputs(108)) or (inputs(144));
    layer0_outputs(3078) <= (inputs(57)) or (inputs(229));
    layer0_outputs(3079) <= not(inputs(92));
    layer0_outputs(3080) <= not((inputs(183)) or (inputs(125)));
    layer0_outputs(3081) <= not((inputs(87)) xor (inputs(26)));
    layer0_outputs(3082) <= not(inputs(231)) or (inputs(110));
    layer0_outputs(3083) <= not((inputs(227)) xor (inputs(199)));
    layer0_outputs(3084) <= not((inputs(222)) or (inputs(47)));
    layer0_outputs(3085) <= (inputs(224)) or (inputs(1));
    layer0_outputs(3086) <= (inputs(80)) xor (inputs(103));
    layer0_outputs(3087) <= not((inputs(166)) or (inputs(241)));
    layer0_outputs(3088) <= (inputs(168)) and (inputs(140));
    layer0_outputs(3089) <= (inputs(152)) and not (inputs(95));
    layer0_outputs(3090) <= inputs(182);
    layer0_outputs(3091) <= not(inputs(75));
    layer0_outputs(3092) <= not(inputs(52)) or (inputs(185));
    layer0_outputs(3093) <= not(inputs(126));
    layer0_outputs(3094) <= not((inputs(122)) or (inputs(154)));
    layer0_outputs(3095) <= not(inputs(85));
    layer0_outputs(3096) <= not(inputs(158));
    layer0_outputs(3097) <= not(inputs(163));
    layer0_outputs(3098) <= not(inputs(164));
    layer0_outputs(3099) <= not(inputs(51));
    layer0_outputs(3100) <= not((inputs(216)) xor (inputs(27)));
    layer0_outputs(3101) <= not(inputs(107));
    layer0_outputs(3102) <= not(inputs(168));
    layer0_outputs(3103) <= inputs(7);
    layer0_outputs(3104) <= not(inputs(5)) or (inputs(127));
    layer0_outputs(3105) <= inputs(110);
    layer0_outputs(3106) <= not(inputs(214)) or (inputs(153));
    layer0_outputs(3107) <= (inputs(86)) and not (inputs(54));
    layer0_outputs(3108) <= not((inputs(222)) or (inputs(204)));
    layer0_outputs(3109) <= (inputs(172)) xor (inputs(156));
    layer0_outputs(3110) <= (inputs(244)) or (inputs(190));
    layer0_outputs(3111) <= (inputs(163)) xor (inputs(167));
    layer0_outputs(3112) <= (inputs(159)) or (inputs(96));
    layer0_outputs(3113) <= inputs(231);
    layer0_outputs(3114) <= not((inputs(50)) xor (inputs(78)));
    layer0_outputs(3115) <= inputs(200);
    layer0_outputs(3116) <= '0';
    layer0_outputs(3117) <= inputs(113);
    layer0_outputs(3118) <= inputs(83);
    layer0_outputs(3119) <= inputs(234);
    layer0_outputs(3120) <= not((inputs(144)) and (inputs(255)));
    layer0_outputs(3121) <= not((inputs(39)) xor (inputs(52)));
    layer0_outputs(3122) <= (inputs(182)) and not (inputs(108));
    layer0_outputs(3123) <= inputs(234);
    layer0_outputs(3124) <= not((inputs(251)) or (inputs(171)));
    layer0_outputs(3125) <= not((inputs(24)) xor (inputs(72)));
    layer0_outputs(3126) <= inputs(124);
    layer0_outputs(3127) <= (inputs(45)) xor (inputs(190));
    layer0_outputs(3128) <= '1';
    layer0_outputs(3129) <= (inputs(52)) or (inputs(205));
    layer0_outputs(3130) <= not((inputs(247)) xor (inputs(75)));
    layer0_outputs(3131) <= inputs(107);
    layer0_outputs(3132) <= not((inputs(210)) xor (inputs(134)));
    layer0_outputs(3133) <= (inputs(64)) xor (inputs(63));
    layer0_outputs(3134) <= (inputs(15)) and not (inputs(11));
    layer0_outputs(3135) <= not((inputs(236)) or (inputs(223)));
    layer0_outputs(3136) <= not(inputs(236)) or (inputs(249));
    layer0_outputs(3137) <= not(inputs(14));
    layer0_outputs(3138) <= (inputs(26)) and not (inputs(133));
    layer0_outputs(3139) <= not(inputs(78));
    layer0_outputs(3140) <= (inputs(173)) xor (inputs(139));
    layer0_outputs(3141) <= not(inputs(131));
    layer0_outputs(3142) <= inputs(7);
    layer0_outputs(3143) <= not(inputs(140)) or (inputs(98));
    layer0_outputs(3144) <= not((inputs(91)) xor (inputs(248)));
    layer0_outputs(3145) <= not(inputs(98)) or (inputs(49));
    layer0_outputs(3146) <= not(inputs(197)) or (inputs(31));
    layer0_outputs(3147) <= not(inputs(157));
    layer0_outputs(3148) <= not(inputs(234));
    layer0_outputs(3149) <= (inputs(103)) or (inputs(219));
    layer0_outputs(3150) <= not((inputs(239)) or (inputs(16)));
    layer0_outputs(3151) <= not(inputs(198));
    layer0_outputs(3152) <= (inputs(138)) and not (inputs(96));
    layer0_outputs(3153) <= inputs(151);
    layer0_outputs(3154) <= not((inputs(189)) xor (inputs(185)));
    layer0_outputs(3155) <= not((inputs(116)) and (inputs(216)));
    layer0_outputs(3156) <= not((inputs(255)) or (inputs(186)));
    layer0_outputs(3157) <= not(inputs(50));
    layer0_outputs(3158) <= not(inputs(99));
    layer0_outputs(3159) <= not((inputs(95)) xor (inputs(203)));
    layer0_outputs(3160) <= (inputs(200)) and (inputs(147));
    layer0_outputs(3161) <= (inputs(108)) xor (inputs(17));
    layer0_outputs(3162) <= (inputs(135)) and not (inputs(191));
    layer0_outputs(3163) <= not(inputs(122));
    layer0_outputs(3164) <= (inputs(86)) xor (inputs(179));
    layer0_outputs(3165) <= not((inputs(204)) xor (inputs(37)));
    layer0_outputs(3166) <= (inputs(213)) and not (inputs(87));
    layer0_outputs(3167) <= not(inputs(205)) or (inputs(30));
    layer0_outputs(3168) <= not(inputs(14)) or (inputs(1));
    layer0_outputs(3169) <= not((inputs(134)) xor (inputs(55)));
    layer0_outputs(3170) <= not(inputs(112));
    layer0_outputs(3171) <= not((inputs(124)) or (inputs(10)));
    layer0_outputs(3172) <= not(inputs(75)) or (inputs(181));
    layer0_outputs(3173) <= not(inputs(180));
    layer0_outputs(3174) <= (inputs(195)) or (inputs(218));
    layer0_outputs(3175) <= inputs(140);
    layer0_outputs(3176) <= inputs(228);
    layer0_outputs(3177) <= not(inputs(119));
    layer0_outputs(3178) <= (inputs(195)) xor (inputs(31));
    layer0_outputs(3179) <= not((inputs(52)) xor (inputs(95)));
    layer0_outputs(3180) <= not((inputs(147)) xor (inputs(212)));
    layer0_outputs(3181) <= (inputs(246)) and not (inputs(1));
    layer0_outputs(3182) <= not(inputs(150)) or (inputs(8));
    layer0_outputs(3183) <= inputs(87);
    layer0_outputs(3184) <= not(inputs(41));
    layer0_outputs(3185) <= (inputs(1)) xor (inputs(25));
    layer0_outputs(3186) <= not((inputs(194)) or (inputs(160)));
    layer0_outputs(3187) <= not((inputs(91)) and (inputs(229)));
    layer0_outputs(3188) <= not((inputs(48)) or (inputs(227)));
    layer0_outputs(3189) <= (inputs(173)) and not (inputs(63));
    layer0_outputs(3190) <= not((inputs(36)) or (inputs(249)));
    layer0_outputs(3191) <= not(inputs(56)) or (inputs(137));
    layer0_outputs(3192) <= inputs(78);
    layer0_outputs(3193) <= (inputs(106)) and not (inputs(128));
    layer0_outputs(3194) <= not(inputs(16));
    layer0_outputs(3195) <= inputs(227);
    layer0_outputs(3196) <= inputs(226);
    layer0_outputs(3197) <= not(inputs(131));
    layer0_outputs(3198) <= inputs(210);
    layer0_outputs(3199) <= '1';
    layer0_outputs(3200) <= not(inputs(44)) or (inputs(171));
    layer0_outputs(3201) <= inputs(29);
    layer0_outputs(3202) <= not(inputs(253)) or (inputs(137));
    layer0_outputs(3203) <= not((inputs(77)) or (inputs(35)));
    layer0_outputs(3204) <= '0';
    layer0_outputs(3205) <= inputs(192);
    layer0_outputs(3206) <= inputs(237);
    layer0_outputs(3207) <= (inputs(29)) or (inputs(129));
    layer0_outputs(3208) <= (inputs(49)) and not (inputs(144));
    layer0_outputs(3209) <= inputs(117);
    layer0_outputs(3210) <= not(inputs(248));
    layer0_outputs(3211) <= not(inputs(173)) or (inputs(51));
    layer0_outputs(3212) <= not((inputs(79)) or (inputs(118)));
    layer0_outputs(3213) <= (inputs(217)) and not (inputs(54));
    layer0_outputs(3214) <= (inputs(231)) and not (inputs(17));
    layer0_outputs(3215) <= (inputs(41)) xor (inputs(10));
    layer0_outputs(3216) <= (inputs(255)) or (inputs(220));
    layer0_outputs(3217) <= not(inputs(88));
    layer0_outputs(3218) <= inputs(212);
    layer0_outputs(3219) <= not(inputs(25)) or (inputs(211));
    layer0_outputs(3220) <= inputs(83);
    layer0_outputs(3221) <= (inputs(146)) xor (inputs(104));
    layer0_outputs(3222) <= (inputs(66)) or (inputs(229));
    layer0_outputs(3223) <= not((inputs(175)) or (inputs(63)));
    layer0_outputs(3224) <= not(inputs(182)) or (inputs(51));
    layer0_outputs(3225) <= not(inputs(58));
    layer0_outputs(3226) <= not(inputs(84));
    layer0_outputs(3227) <= (inputs(23)) or (inputs(10));
    layer0_outputs(3228) <= (inputs(88)) or (inputs(137));
    layer0_outputs(3229) <= not(inputs(155));
    layer0_outputs(3230) <= (inputs(95)) or (inputs(26));
    layer0_outputs(3231) <= (inputs(56)) and not (inputs(200));
    layer0_outputs(3232) <= (inputs(141)) or (inputs(5));
    layer0_outputs(3233) <= inputs(122);
    layer0_outputs(3234) <= not(inputs(247)) or (inputs(59));
    layer0_outputs(3235) <= not((inputs(64)) or (inputs(118)));
    layer0_outputs(3236) <= (inputs(106)) xor (inputs(168));
    layer0_outputs(3237) <= not((inputs(37)) xor (inputs(31)));
    layer0_outputs(3238) <= (inputs(248)) xor (inputs(216));
    layer0_outputs(3239) <= not(inputs(54)) or (inputs(234));
    layer0_outputs(3240) <= not((inputs(240)) or (inputs(186)));
    layer0_outputs(3241) <= not((inputs(103)) xor (inputs(36)));
    layer0_outputs(3242) <= not((inputs(133)) xor (inputs(121)));
    layer0_outputs(3243) <= (inputs(229)) or (inputs(173));
    layer0_outputs(3244) <= inputs(86);
    layer0_outputs(3245) <= inputs(83);
    layer0_outputs(3246) <= (inputs(225)) and not (inputs(14));
    layer0_outputs(3247) <= inputs(189);
    layer0_outputs(3248) <= not(inputs(90)) or (inputs(194));
    layer0_outputs(3249) <= (inputs(221)) or (inputs(14));
    layer0_outputs(3250) <= '0';
    layer0_outputs(3251) <= (inputs(108)) or (inputs(12));
    layer0_outputs(3252) <= (inputs(68)) xor (inputs(25));
    layer0_outputs(3253) <= inputs(91);
    layer0_outputs(3254) <= inputs(42);
    layer0_outputs(3255) <= (inputs(161)) or (inputs(96));
    layer0_outputs(3256) <= (inputs(66)) or (inputs(205));
    layer0_outputs(3257) <= (inputs(24)) and not (inputs(197));
    layer0_outputs(3258) <= not(inputs(44)) or (inputs(156));
    layer0_outputs(3259) <= inputs(14);
    layer0_outputs(3260) <= not((inputs(228)) xor (inputs(248)));
    layer0_outputs(3261) <= (inputs(131)) and not (inputs(207));
    layer0_outputs(3262) <= not(inputs(194)) or (inputs(28));
    layer0_outputs(3263) <= not((inputs(0)) xor (inputs(65)));
    layer0_outputs(3264) <= not((inputs(169)) xor (inputs(182)));
    layer0_outputs(3265) <= (inputs(105)) and (inputs(15));
    layer0_outputs(3266) <= (inputs(70)) or (inputs(82));
    layer0_outputs(3267) <= not(inputs(3)) or (inputs(236));
    layer0_outputs(3268) <= (inputs(184)) or (inputs(169));
    layer0_outputs(3269) <= inputs(148);
    layer0_outputs(3270) <= inputs(179);
    layer0_outputs(3271) <= not(inputs(70));
    layer0_outputs(3272) <= not((inputs(225)) or (inputs(133)));
    layer0_outputs(3273) <= (inputs(113)) or (inputs(211));
    layer0_outputs(3274) <= not((inputs(133)) xor (inputs(205)));
    layer0_outputs(3275) <= not((inputs(254)) or (inputs(105)));
    layer0_outputs(3276) <= not(inputs(214));
    layer0_outputs(3277) <= not((inputs(93)) xor (inputs(112)));
    layer0_outputs(3278) <= not(inputs(61));
    layer0_outputs(3279) <= not(inputs(227)) or (inputs(255));
    layer0_outputs(3280) <= not(inputs(205)) or (inputs(162));
    layer0_outputs(3281) <= not(inputs(66)) or (inputs(144));
    layer0_outputs(3282) <= not((inputs(109)) xor (inputs(250)));
    layer0_outputs(3283) <= inputs(173);
    layer0_outputs(3284) <= not(inputs(148)) or (inputs(6));
    layer0_outputs(3285) <= not((inputs(210)) or (inputs(110)));
    layer0_outputs(3286) <= inputs(162);
    layer0_outputs(3287) <= not(inputs(255));
    layer0_outputs(3288) <= not(inputs(132));
    layer0_outputs(3289) <= not(inputs(224));
    layer0_outputs(3290) <= not((inputs(140)) or (inputs(111)));
    layer0_outputs(3291) <= not(inputs(219)) or (inputs(87));
    layer0_outputs(3292) <= (inputs(32)) or (inputs(75));
    layer0_outputs(3293) <= not(inputs(25)) or (inputs(147));
    layer0_outputs(3294) <= not(inputs(114));
    layer0_outputs(3295) <= not(inputs(126));
    layer0_outputs(3296) <= (inputs(68)) or (inputs(106));
    layer0_outputs(3297) <= (inputs(177)) or (inputs(96));
    layer0_outputs(3298) <= (inputs(229)) and not (inputs(76));
    layer0_outputs(3299) <= (inputs(124)) or (inputs(14));
    layer0_outputs(3300) <= inputs(109);
    layer0_outputs(3301) <= (inputs(201)) and not (inputs(151));
    layer0_outputs(3302) <= not((inputs(107)) or (inputs(247)));
    layer0_outputs(3303) <= not((inputs(88)) xor (inputs(104)));
    layer0_outputs(3304) <= inputs(112);
    layer0_outputs(3305) <= not(inputs(88));
    layer0_outputs(3306) <= not(inputs(73)) or (inputs(184));
    layer0_outputs(3307) <= (inputs(247)) and not (inputs(253));
    layer0_outputs(3308) <= inputs(190);
    layer0_outputs(3309) <= not(inputs(248)) or (inputs(2));
    layer0_outputs(3310) <= not(inputs(197)) or (inputs(232));
    layer0_outputs(3311) <= inputs(202);
    layer0_outputs(3312) <= not((inputs(7)) or (inputs(91)));
    layer0_outputs(3313) <= (inputs(43)) or (inputs(34));
    layer0_outputs(3314) <= (inputs(126)) xor (inputs(154));
    layer0_outputs(3315) <= (inputs(106)) and not (inputs(38));
    layer0_outputs(3316) <= not(inputs(87));
    layer0_outputs(3317) <= inputs(107);
    layer0_outputs(3318) <= inputs(149);
    layer0_outputs(3319) <= not(inputs(115));
    layer0_outputs(3320) <= (inputs(180)) or (inputs(96));
    layer0_outputs(3321) <= (inputs(55)) and not (inputs(95));
    layer0_outputs(3322) <= not(inputs(151));
    layer0_outputs(3323) <= (inputs(130)) xor (inputs(155));
    layer0_outputs(3324) <= (inputs(65)) or (inputs(188));
    layer0_outputs(3325) <= not((inputs(211)) or (inputs(160)));
    layer0_outputs(3326) <= (inputs(19)) or (inputs(47));
    layer0_outputs(3327) <= not(inputs(142));
    layer0_outputs(3328) <= not(inputs(215)) or (inputs(91));
    layer0_outputs(3329) <= not(inputs(22)) or (inputs(231));
    layer0_outputs(3330) <= not((inputs(11)) and (inputs(10)));
    layer0_outputs(3331) <= not((inputs(145)) or (inputs(159)));
    layer0_outputs(3332) <= not(inputs(237));
    layer0_outputs(3333) <= not(inputs(174));
    layer0_outputs(3334) <= (inputs(221)) and not (inputs(14));
    layer0_outputs(3335) <= not((inputs(250)) xor (inputs(51)));
    layer0_outputs(3336) <= inputs(55);
    layer0_outputs(3337) <= not((inputs(210)) or (inputs(190)));
    layer0_outputs(3338) <= (inputs(213)) xor (inputs(199));
    layer0_outputs(3339) <= (inputs(199)) or (inputs(141));
    layer0_outputs(3340) <= (inputs(185)) or (inputs(170));
    layer0_outputs(3341) <= inputs(51);
    layer0_outputs(3342) <= not(inputs(11)) or (inputs(188));
    layer0_outputs(3343) <= not((inputs(134)) and (inputs(28)));
    layer0_outputs(3344) <= (inputs(46)) and not (inputs(79));
    layer0_outputs(3345) <= (inputs(181)) and not (inputs(202));
    layer0_outputs(3346) <= (inputs(238)) or (inputs(8));
    layer0_outputs(3347) <= inputs(141);
    layer0_outputs(3348) <= '0';
    layer0_outputs(3349) <= (inputs(244)) or (inputs(28));
    layer0_outputs(3350) <= (inputs(112)) and not (inputs(47));
    layer0_outputs(3351) <= not(inputs(241)) or (inputs(46));
    layer0_outputs(3352) <= (inputs(183)) and (inputs(234));
    layer0_outputs(3353) <= not(inputs(178)) or (inputs(198));
    layer0_outputs(3354) <= not(inputs(180)) or (inputs(223));
    layer0_outputs(3355) <= not(inputs(153)) or (inputs(26));
    layer0_outputs(3356) <= not((inputs(16)) or (inputs(238)));
    layer0_outputs(3357) <= not(inputs(53));
    layer0_outputs(3358) <= inputs(70);
    layer0_outputs(3359) <= not((inputs(86)) xor (inputs(198)));
    layer0_outputs(3360) <= (inputs(208)) and (inputs(4));
    layer0_outputs(3361) <= (inputs(13)) and not (inputs(88));
    layer0_outputs(3362) <= (inputs(48)) xor (inputs(122));
    layer0_outputs(3363) <= not(inputs(148));
    layer0_outputs(3364) <= inputs(70);
    layer0_outputs(3365) <= not(inputs(9)) or (inputs(69));
    layer0_outputs(3366) <= inputs(61);
    layer0_outputs(3367) <= inputs(217);
    layer0_outputs(3368) <= not(inputs(104)) or (inputs(3));
    layer0_outputs(3369) <= not((inputs(253)) or (inputs(249)));
    layer0_outputs(3370) <= not((inputs(202)) and (inputs(215)));
    layer0_outputs(3371) <= (inputs(93)) or (inputs(111));
    layer0_outputs(3372) <= not((inputs(166)) or (inputs(21)));
    layer0_outputs(3373) <= not((inputs(71)) xor (inputs(6)));
    layer0_outputs(3374) <= (inputs(215)) or (inputs(171));
    layer0_outputs(3375) <= not(inputs(185));
    layer0_outputs(3376) <= '1';
    layer0_outputs(3377) <= not(inputs(170)) or (inputs(33));
    layer0_outputs(3378) <= not(inputs(75));
    layer0_outputs(3379) <= not((inputs(186)) or (inputs(175)));
    layer0_outputs(3380) <= (inputs(72)) and not (inputs(123));
    layer0_outputs(3381) <= (inputs(228)) xor (inputs(32));
    layer0_outputs(3382) <= not((inputs(196)) xor (inputs(167)));
    layer0_outputs(3383) <= (inputs(186)) xor (inputs(20));
    layer0_outputs(3384) <= inputs(58);
    layer0_outputs(3385) <= (inputs(23)) and not (inputs(15));
    layer0_outputs(3386) <= inputs(157);
    layer0_outputs(3387) <= not((inputs(205)) xor (inputs(211)));
    layer0_outputs(3388) <= not(inputs(28));
    layer0_outputs(3389) <= not(inputs(228)) or (inputs(68));
    layer0_outputs(3390) <= inputs(129);
    layer0_outputs(3391) <= (inputs(136)) xor (inputs(104));
    layer0_outputs(3392) <= not(inputs(27));
    layer0_outputs(3393) <= (inputs(196)) and (inputs(93));
    layer0_outputs(3394) <= (inputs(6)) or (inputs(179));
    layer0_outputs(3395) <= not(inputs(74));
    layer0_outputs(3396) <= (inputs(74)) and (inputs(221));
    layer0_outputs(3397) <= (inputs(61)) xor (inputs(62));
    layer0_outputs(3398) <= not(inputs(64));
    layer0_outputs(3399) <= (inputs(189)) or (inputs(45));
    layer0_outputs(3400) <= not(inputs(108));
    layer0_outputs(3401) <= not(inputs(217)) or (inputs(109));
    layer0_outputs(3402) <= inputs(226);
    layer0_outputs(3403) <= (inputs(44)) and (inputs(87));
    layer0_outputs(3404) <= (inputs(81)) or (inputs(178));
    layer0_outputs(3405) <= (inputs(247)) xor (inputs(36));
    layer0_outputs(3406) <= (inputs(29)) xor (inputs(62));
    layer0_outputs(3407) <= inputs(91);
    layer0_outputs(3408) <= inputs(204);
    layer0_outputs(3409) <= (inputs(142)) and (inputs(97));
    layer0_outputs(3410) <= inputs(50);
    layer0_outputs(3411) <= (inputs(176)) or (inputs(21));
    layer0_outputs(3412) <= not((inputs(68)) or (inputs(29)));
    layer0_outputs(3413) <= not(inputs(93));
    layer0_outputs(3414) <= (inputs(171)) and not (inputs(128));
    layer0_outputs(3415) <= inputs(46);
    layer0_outputs(3416) <= (inputs(168)) or (inputs(200));
    layer0_outputs(3417) <= not(inputs(200));
    layer0_outputs(3418) <= not((inputs(210)) xor (inputs(148)));
    layer0_outputs(3419) <= (inputs(178)) xor (inputs(228));
    layer0_outputs(3420) <= not((inputs(129)) or (inputs(13)));
    layer0_outputs(3421) <= not(inputs(27));
    layer0_outputs(3422) <= (inputs(153)) and not (inputs(48));
    layer0_outputs(3423) <= inputs(246);
    layer0_outputs(3424) <= not((inputs(180)) and (inputs(218)));
    layer0_outputs(3425) <= (inputs(142)) and not (inputs(43));
    layer0_outputs(3426) <= (inputs(197)) and not (inputs(32));
    layer0_outputs(3427) <= inputs(68);
    layer0_outputs(3428) <= not((inputs(72)) or (inputs(154)));
    layer0_outputs(3429) <= inputs(189);
    layer0_outputs(3430) <= inputs(230);
    layer0_outputs(3431) <= (inputs(110)) xor (inputs(33));
    layer0_outputs(3432) <= not((inputs(13)) and (inputs(74)));
    layer0_outputs(3433) <= not(inputs(4)) or (inputs(222));
    layer0_outputs(3434) <= not((inputs(229)) and (inputs(18)));
    layer0_outputs(3435) <= inputs(232);
    layer0_outputs(3436) <= (inputs(23)) or (inputs(46));
    layer0_outputs(3437) <= (inputs(93)) or (inputs(52));
    layer0_outputs(3438) <= not((inputs(110)) xor (inputs(191)));
    layer0_outputs(3439) <= not((inputs(140)) xor (inputs(248)));
    layer0_outputs(3440) <= not(inputs(104));
    layer0_outputs(3441) <= (inputs(92)) or (inputs(80));
    layer0_outputs(3442) <= not((inputs(173)) xor (inputs(203)));
    layer0_outputs(3443) <= not(inputs(107));
    layer0_outputs(3444) <= not(inputs(194));
    layer0_outputs(3445) <= not((inputs(160)) xor (inputs(232)));
    layer0_outputs(3446) <= inputs(119);
    layer0_outputs(3447) <= (inputs(46)) and not (inputs(161));
    layer0_outputs(3448) <= not(inputs(149));
    layer0_outputs(3449) <= not(inputs(243)) or (inputs(138));
    layer0_outputs(3450) <= not((inputs(115)) or (inputs(140)));
    layer0_outputs(3451) <= (inputs(51)) and not (inputs(217));
    layer0_outputs(3452) <= (inputs(194)) or (inputs(183));
    layer0_outputs(3453) <= not(inputs(211)) or (inputs(44));
    layer0_outputs(3454) <= (inputs(81)) xor (inputs(83));
    layer0_outputs(3455) <= not((inputs(8)) xor (inputs(5)));
    layer0_outputs(3456) <= inputs(190);
    layer0_outputs(3457) <= (inputs(237)) or (inputs(14));
    layer0_outputs(3458) <= not(inputs(229)) or (inputs(119));
    layer0_outputs(3459) <= inputs(245);
    layer0_outputs(3460) <= (inputs(134)) xor (inputs(102));
    layer0_outputs(3461) <= (inputs(41)) or (inputs(221));
    layer0_outputs(3462) <= inputs(56);
    layer0_outputs(3463) <= (inputs(67)) and not (inputs(72));
    layer0_outputs(3464) <= (inputs(188)) xor (inputs(83));
    layer0_outputs(3465) <= (inputs(191)) and not (inputs(145));
    layer0_outputs(3466) <= not(inputs(59));
    layer0_outputs(3467) <= not((inputs(234)) xor (inputs(154)));
    layer0_outputs(3468) <= (inputs(150)) and not (inputs(64));
    layer0_outputs(3469) <= (inputs(149)) and not (inputs(55));
    layer0_outputs(3470) <= not(inputs(126));
    layer0_outputs(3471) <= (inputs(11)) or (inputs(7));
    layer0_outputs(3472) <= not((inputs(68)) xor (inputs(51)));
    layer0_outputs(3473) <= not(inputs(162)) or (inputs(51));
    layer0_outputs(3474) <= not((inputs(250)) or (inputs(208)));
    layer0_outputs(3475) <= not((inputs(203)) or (inputs(242)));
    layer0_outputs(3476) <= not(inputs(197));
    layer0_outputs(3477) <= (inputs(155)) xor (inputs(181));
    layer0_outputs(3478) <= inputs(73);
    layer0_outputs(3479) <= inputs(21);
    layer0_outputs(3480) <= (inputs(58)) xor (inputs(38));
    layer0_outputs(3481) <= not(inputs(121));
    layer0_outputs(3482) <= not(inputs(210));
    layer0_outputs(3483) <= not((inputs(95)) or (inputs(109)));
    layer0_outputs(3484) <= not((inputs(111)) or (inputs(176)));
    layer0_outputs(3485) <= inputs(114);
    layer0_outputs(3486) <= inputs(245);
    layer0_outputs(3487) <= (inputs(214)) xor (inputs(7));
    layer0_outputs(3488) <= not(inputs(83));
    layer0_outputs(3489) <= not((inputs(237)) or (inputs(170)));
    layer0_outputs(3490) <= (inputs(73)) and (inputs(151));
    layer0_outputs(3491) <= not((inputs(169)) xor (inputs(0)));
    layer0_outputs(3492) <= (inputs(108)) xor (inputs(111));
    layer0_outputs(3493) <= (inputs(230)) or (inputs(159));
    layer0_outputs(3494) <= (inputs(190)) or (inputs(246));
    layer0_outputs(3495) <= (inputs(14)) or (inputs(200));
    layer0_outputs(3496) <= (inputs(77)) and not (inputs(252));
    layer0_outputs(3497) <= (inputs(103)) xor (inputs(116));
    layer0_outputs(3498) <= not((inputs(135)) or (inputs(87)));
    layer0_outputs(3499) <= not((inputs(105)) or (inputs(80)));
    layer0_outputs(3500) <= (inputs(52)) xor (inputs(178));
    layer0_outputs(3501) <= inputs(192);
    layer0_outputs(3502) <= not(inputs(228)) or (inputs(208));
    layer0_outputs(3503) <= not((inputs(10)) or (inputs(250)));
    layer0_outputs(3504) <= not(inputs(51));
    layer0_outputs(3505) <= (inputs(149)) and not (inputs(231));
    layer0_outputs(3506) <= not((inputs(48)) or (inputs(234)));
    layer0_outputs(3507) <= not(inputs(121));
    layer0_outputs(3508) <= not(inputs(120)) or (inputs(219));
    layer0_outputs(3509) <= not(inputs(54));
    layer0_outputs(3510) <= inputs(134);
    layer0_outputs(3511) <= inputs(158);
    layer0_outputs(3512) <= '0';
    layer0_outputs(3513) <= not(inputs(155));
    layer0_outputs(3514) <= not(inputs(230));
    layer0_outputs(3515) <= not(inputs(190));
    layer0_outputs(3516) <= not(inputs(165));
    layer0_outputs(3517) <= inputs(174);
    layer0_outputs(3518) <= not((inputs(103)) xor (inputs(13)));
    layer0_outputs(3519) <= (inputs(8)) xor (inputs(68));
    layer0_outputs(3520) <= not((inputs(157)) or (inputs(55)));
    layer0_outputs(3521) <= inputs(231);
    layer0_outputs(3522) <= not(inputs(161)) or (inputs(1));
    layer0_outputs(3523) <= not(inputs(196)) or (inputs(46));
    layer0_outputs(3524) <= (inputs(40)) and not (inputs(224));
    layer0_outputs(3525) <= not(inputs(207));
    layer0_outputs(3526) <= (inputs(131)) xor (inputs(251));
    layer0_outputs(3527) <= inputs(98);
    layer0_outputs(3528) <= not((inputs(198)) or (inputs(94)));
    layer0_outputs(3529) <= inputs(71);
    layer0_outputs(3530) <= not(inputs(208));
    layer0_outputs(3531) <= inputs(61);
    layer0_outputs(3532) <= (inputs(49)) or (inputs(86));
    layer0_outputs(3533) <= inputs(136);
    layer0_outputs(3534) <= not((inputs(78)) xor (inputs(203)));
    layer0_outputs(3535) <= not(inputs(84));
    layer0_outputs(3536) <= (inputs(121)) and not (inputs(178));
    layer0_outputs(3537) <= not(inputs(131));
    layer0_outputs(3538) <= inputs(98);
    layer0_outputs(3539) <= not(inputs(115));
    layer0_outputs(3540) <= (inputs(8)) and not (inputs(66));
    layer0_outputs(3541) <= (inputs(104)) and not (inputs(233));
    layer0_outputs(3542) <= not(inputs(57));
    layer0_outputs(3543) <= not(inputs(126));
    layer0_outputs(3544) <= inputs(79);
    layer0_outputs(3545) <= not(inputs(44)) or (inputs(252));
    layer0_outputs(3546) <= (inputs(5)) and not (inputs(202));
    layer0_outputs(3547) <= not((inputs(138)) or (inputs(63)));
    layer0_outputs(3548) <= (inputs(139)) xor (inputs(53));
    layer0_outputs(3549) <= (inputs(13)) xor (inputs(128));
    layer0_outputs(3550) <= not((inputs(47)) or (inputs(192)));
    layer0_outputs(3551) <= inputs(104);
    layer0_outputs(3552) <= (inputs(104)) and not (inputs(15));
    layer0_outputs(3553) <= (inputs(68)) and not (inputs(9));
    layer0_outputs(3554) <= not((inputs(25)) xor (inputs(234)));
    layer0_outputs(3555) <= inputs(46);
    layer0_outputs(3556) <= inputs(240);
    layer0_outputs(3557) <= inputs(106);
    layer0_outputs(3558) <= (inputs(133)) xor (inputs(136));
    layer0_outputs(3559) <= (inputs(191)) or (inputs(222));
    layer0_outputs(3560) <= (inputs(86)) and not (inputs(156));
    layer0_outputs(3561) <= (inputs(160)) and not (inputs(60));
    layer0_outputs(3562) <= '1';
    layer0_outputs(3563) <= (inputs(108)) or (inputs(168));
    layer0_outputs(3564) <= not((inputs(98)) or (inputs(129)));
    layer0_outputs(3565) <= '0';
    layer0_outputs(3566) <= inputs(125);
    layer0_outputs(3567) <= inputs(82);
    layer0_outputs(3568) <= (inputs(244)) and not (inputs(16));
    layer0_outputs(3569) <= inputs(67);
    layer0_outputs(3570) <= not(inputs(110)) or (inputs(223));
    layer0_outputs(3571) <= not((inputs(12)) and (inputs(131)));
    layer0_outputs(3572) <= not(inputs(253));
    layer0_outputs(3573) <= (inputs(205)) or (inputs(80));
    layer0_outputs(3574) <= (inputs(101)) and not (inputs(193));
    layer0_outputs(3575) <= (inputs(180)) xor (inputs(226));
    layer0_outputs(3576) <= not(inputs(213));
    layer0_outputs(3577) <= not(inputs(186)) or (inputs(153));
    layer0_outputs(3578) <= (inputs(137)) or (inputs(221));
    layer0_outputs(3579) <= inputs(70);
    layer0_outputs(3580) <= not(inputs(167)) or (inputs(32));
    layer0_outputs(3581) <= not((inputs(119)) xor (inputs(4)));
    layer0_outputs(3582) <= not(inputs(83)) or (inputs(18));
    layer0_outputs(3583) <= inputs(24);
    layer0_outputs(3584) <= inputs(41);
    layer0_outputs(3585) <= (inputs(104)) and not (inputs(35));
    layer0_outputs(3586) <= (inputs(253)) or (inputs(183));
    layer0_outputs(3587) <= not(inputs(82));
    layer0_outputs(3588) <= (inputs(50)) or (inputs(236));
    layer0_outputs(3589) <= not(inputs(155)) or (inputs(0));
    layer0_outputs(3590) <= (inputs(43)) and not (inputs(51));
    layer0_outputs(3591) <= (inputs(66)) or (inputs(212));
    layer0_outputs(3592) <= inputs(56);
    layer0_outputs(3593) <= (inputs(15)) or (inputs(9));
    layer0_outputs(3594) <= inputs(205);
    layer0_outputs(3595) <= not(inputs(46));
    layer0_outputs(3596) <= inputs(222);
    layer0_outputs(3597) <= inputs(234);
    layer0_outputs(3598) <= not((inputs(156)) xor (inputs(250)));
    layer0_outputs(3599) <= (inputs(165)) xor (inputs(163));
    layer0_outputs(3600) <= (inputs(197)) xor (inputs(222));
    layer0_outputs(3601) <= not(inputs(194));
    layer0_outputs(3602) <= not(inputs(52)) or (inputs(39));
    layer0_outputs(3603) <= (inputs(138)) and not (inputs(11));
    layer0_outputs(3604) <= not(inputs(230));
    layer0_outputs(3605) <= not((inputs(222)) xor (inputs(203)));
    layer0_outputs(3606) <= (inputs(161)) or (inputs(62));
    layer0_outputs(3607) <= inputs(184);
    layer0_outputs(3608) <= not((inputs(33)) or (inputs(67)));
    layer0_outputs(3609) <= (inputs(49)) and not (inputs(14));
    layer0_outputs(3610) <= (inputs(173)) and (inputs(88));
    layer0_outputs(3611) <= (inputs(199)) or (inputs(32));
    layer0_outputs(3612) <= not(inputs(186)) or (inputs(22));
    layer0_outputs(3613) <= not((inputs(95)) or (inputs(74)));
    layer0_outputs(3614) <= inputs(2);
    layer0_outputs(3615) <= not(inputs(193));
    layer0_outputs(3616) <= inputs(156);
    layer0_outputs(3617) <= not(inputs(114)) or (inputs(225));
    layer0_outputs(3618) <= not(inputs(56));
    layer0_outputs(3619) <= inputs(241);
    layer0_outputs(3620) <= '1';
    layer0_outputs(3621) <= not((inputs(162)) or (inputs(222)));
    layer0_outputs(3622) <= (inputs(97)) and (inputs(225));
    layer0_outputs(3623) <= not((inputs(179)) xor (inputs(138)));
    layer0_outputs(3624) <= not((inputs(165)) xor (inputs(236)));
    layer0_outputs(3625) <= inputs(46);
    layer0_outputs(3626) <= not((inputs(142)) xor (inputs(250)));
    layer0_outputs(3627) <= '0';
    layer0_outputs(3628) <= not((inputs(47)) xor (inputs(15)));
    layer0_outputs(3629) <= not((inputs(94)) xor (inputs(179)));
    layer0_outputs(3630) <= inputs(97);
    layer0_outputs(3631) <= not(inputs(63));
    layer0_outputs(3632) <= not((inputs(114)) and (inputs(243)));
    layer0_outputs(3633) <= not(inputs(246)) or (inputs(83));
    layer0_outputs(3634) <= inputs(82);
    layer0_outputs(3635) <= not((inputs(241)) or (inputs(248)));
    layer0_outputs(3636) <= (inputs(70)) and not (inputs(220));
    layer0_outputs(3637) <= (inputs(28)) and not (inputs(110));
    layer0_outputs(3638) <= (inputs(18)) xor (inputs(80));
    layer0_outputs(3639) <= not(inputs(78));
    layer0_outputs(3640) <= (inputs(120)) and not (inputs(158));
    layer0_outputs(3641) <= not((inputs(232)) or (inputs(186)));
    layer0_outputs(3642) <= (inputs(22)) and not (inputs(216));
    layer0_outputs(3643) <= not(inputs(0)) or (inputs(161));
    layer0_outputs(3644) <= not((inputs(254)) or (inputs(146)));
    layer0_outputs(3645) <= inputs(167);
    layer0_outputs(3646) <= inputs(195);
    layer0_outputs(3647) <= (inputs(116)) and not (inputs(209));
    layer0_outputs(3648) <= (inputs(43)) and not (inputs(207));
    layer0_outputs(3649) <= not((inputs(71)) xor (inputs(110)));
    layer0_outputs(3650) <= (inputs(20)) xor (inputs(53));
    layer0_outputs(3651) <= inputs(98);
    layer0_outputs(3652) <= not(inputs(200));
    layer0_outputs(3653) <= (inputs(164)) or (inputs(7));
    layer0_outputs(3654) <= not(inputs(118)) or (inputs(141));
    layer0_outputs(3655) <= (inputs(60)) or (inputs(239));
    layer0_outputs(3656) <= not(inputs(88));
    layer0_outputs(3657) <= not((inputs(218)) and (inputs(188)));
    layer0_outputs(3658) <= (inputs(182)) or (inputs(160));
    layer0_outputs(3659) <= (inputs(60)) and not (inputs(242));
    layer0_outputs(3660) <= not((inputs(253)) or (inputs(34)));
    layer0_outputs(3661) <= not(inputs(220)) or (inputs(127));
    layer0_outputs(3662) <= not(inputs(171));
    layer0_outputs(3663) <= not(inputs(119));
    layer0_outputs(3664) <= (inputs(134)) or (inputs(190));
    layer0_outputs(3665) <= not((inputs(111)) or (inputs(194)));
    layer0_outputs(3666) <= (inputs(16)) xor (inputs(238));
    layer0_outputs(3667) <= (inputs(155)) xor (inputs(37));
    layer0_outputs(3668) <= (inputs(40)) and not (inputs(228));
    layer0_outputs(3669) <= inputs(228);
    layer0_outputs(3670) <= not(inputs(183)) or (inputs(143));
    layer0_outputs(3671) <= (inputs(182)) and (inputs(25));
    layer0_outputs(3672) <= (inputs(164)) xor (inputs(203));
    layer0_outputs(3673) <= not(inputs(39)) or (inputs(176));
    layer0_outputs(3674) <= (inputs(88)) xor (inputs(108));
    layer0_outputs(3675) <= not((inputs(98)) or (inputs(119)));
    layer0_outputs(3676) <= inputs(167);
    layer0_outputs(3677) <= inputs(76);
    layer0_outputs(3678) <= (inputs(220)) and not (inputs(194));
    layer0_outputs(3679) <= (inputs(111)) xor (inputs(48));
    layer0_outputs(3680) <= not(inputs(164));
    layer0_outputs(3681) <= not((inputs(41)) xor (inputs(9)));
    layer0_outputs(3682) <= (inputs(140)) and not (inputs(152));
    layer0_outputs(3683) <= (inputs(252)) or (inputs(100));
    layer0_outputs(3684) <= inputs(121);
    layer0_outputs(3685) <= (inputs(6)) or (inputs(94));
    layer0_outputs(3686) <= (inputs(124)) xor (inputs(243));
    layer0_outputs(3687) <= not(inputs(194)) or (inputs(130));
    layer0_outputs(3688) <= inputs(20);
    layer0_outputs(3689) <= not(inputs(74));
    layer0_outputs(3690) <= (inputs(227)) or (inputs(132));
    layer0_outputs(3691) <= (inputs(145)) or (inputs(233));
    layer0_outputs(3692) <= (inputs(37)) and not (inputs(174));
    layer0_outputs(3693) <= (inputs(127)) or (inputs(20));
    layer0_outputs(3694) <= inputs(99);
    layer0_outputs(3695) <= inputs(51);
    layer0_outputs(3696) <= inputs(192);
    layer0_outputs(3697) <= not(inputs(84));
    layer0_outputs(3698) <= not(inputs(66));
    layer0_outputs(3699) <= not((inputs(153)) or (inputs(247)));
    layer0_outputs(3700) <= inputs(174);
    layer0_outputs(3701) <= (inputs(229)) xor (inputs(182));
    layer0_outputs(3702) <= inputs(3);
    layer0_outputs(3703) <= inputs(196);
    layer0_outputs(3704) <= (inputs(79)) xor (inputs(216));
    layer0_outputs(3705) <= not((inputs(33)) and (inputs(52)));
    layer0_outputs(3706) <= (inputs(33)) xor (inputs(94));
    layer0_outputs(3707) <= not((inputs(150)) xor (inputs(19)));
    layer0_outputs(3708) <= (inputs(248)) xor (inputs(177));
    layer0_outputs(3709) <= not(inputs(197));
    layer0_outputs(3710) <= not(inputs(34));
    layer0_outputs(3711) <= not(inputs(200));
    layer0_outputs(3712) <= inputs(211);
    layer0_outputs(3713) <= '1';
    layer0_outputs(3714) <= not(inputs(55));
    layer0_outputs(3715) <= not((inputs(156)) xor (inputs(207)));
    layer0_outputs(3716) <= not(inputs(114));
    layer0_outputs(3717) <= inputs(84);
    layer0_outputs(3718) <= (inputs(150)) xor (inputs(211));
    layer0_outputs(3719) <= not((inputs(244)) and (inputs(56)));
    layer0_outputs(3720) <= (inputs(71)) and not (inputs(176));
    layer0_outputs(3721) <= not(inputs(144)) or (inputs(95));
    layer0_outputs(3722) <= (inputs(33)) xor (inputs(100));
    layer0_outputs(3723) <= not(inputs(87));
    layer0_outputs(3724) <= not(inputs(249));
    layer0_outputs(3725) <= (inputs(208)) xor (inputs(170));
    layer0_outputs(3726) <= not((inputs(7)) or (inputs(67)));
    layer0_outputs(3727) <= inputs(218);
    layer0_outputs(3728) <= not((inputs(44)) xor (inputs(228)));
    layer0_outputs(3729) <= not(inputs(149)) or (inputs(77));
    layer0_outputs(3730) <= '1';
    layer0_outputs(3731) <= not((inputs(146)) or (inputs(117)));
    layer0_outputs(3732) <= '1';
    layer0_outputs(3733) <= (inputs(4)) or (inputs(245));
    layer0_outputs(3734) <= inputs(103);
    layer0_outputs(3735) <= not(inputs(99));
    layer0_outputs(3736) <= inputs(224);
    layer0_outputs(3737) <= (inputs(187)) or (inputs(33));
    layer0_outputs(3738) <= (inputs(92)) or (inputs(80));
    layer0_outputs(3739) <= not((inputs(171)) and (inputs(234)));
    layer0_outputs(3740) <= not(inputs(221)) or (inputs(114));
    layer0_outputs(3741) <= '0';
    layer0_outputs(3742) <= not(inputs(247)) or (inputs(111));
    layer0_outputs(3743) <= (inputs(51)) and not (inputs(171));
    layer0_outputs(3744) <= not(inputs(207));
    layer0_outputs(3745) <= not(inputs(133)) or (inputs(51));
    layer0_outputs(3746) <= not((inputs(240)) or (inputs(106)));
    layer0_outputs(3747) <= not(inputs(176));
    layer0_outputs(3748) <= inputs(162);
    layer0_outputs(3749) <= not(inputs(79));
    layer0_outputs(3750) <= (inputs(13)) or (inputs(129));
    layer0_outputs(3751) <= (inputs(174)) and not (inputs(255));
    layer0_outputs(3752) <= not(inputs(228)) or (inputs(3));
    layer0_outputs(3753) <= inputs(202);
    layer0_outputs(3754) <= not(inputs(136));
    layer0_outputs(3755) <= not((inputs(162)) or (inputs(42)));
    layer0_outputs(3756) <= not((inputs(66)) or (inputs(105)));
    layer0_outputs(3757) <= (inputs(143)) or (inputs(161));
    layer0_outputs(3758) <= inputs(188);
    layer0_outputs(3759) <= not(inputs(180));
    layer0_outputs(3760) <= not((inputs(78)) or (inputs(40)));
    layer0_outputs(3761) <= inputs(83);
    layer0_outputs(3762) <= not((inputs(162)) or (inputs(214)));
    layer0_outputs(3763) <= (inputs(171)) or (inputs(27));
    layer0_outputs(3764) <= not(inputs(168));
    layer0_outputs(3765) <= not(inputs(166));
    layer0_outputs(3766) <= not(inputs(68));
    layer0_outputs(3767) <= (inputs(39)) and not (inputs(46));
    layer0_outputs(3768) <= (inputs(115)) or (inputs(121));
    layer0_outputs(3769) <= inputs(126);
    layer0_outputs(3770) <= inputs(66);
    layer0_outputs(3771) <= (inputs(148)) and not (inputs(48));
    layer0_outputs(3772) <= (inputs(139)) or (inputs(159));
    layer0_outputs(3773) <= (inputs(19)) or (inputs(142));
    layer0_outputs(3774) <= not(inputs(99));
    layer0_outputs(3775) <= not(inputs(166));
    layer0_outputs(3776) <= not(inputs(51)) or (inputs(157));
    layer0_outputs(3777) <= (inputs(74)) xor (inputs(161));
    layer0_outputs(3778) <= (inputs(153)) or (inputs(252));
    layer0_outputs(3779) <= (inputs(170)) and not (inputs(79));
    layer0_outputs(3780) <= (inputs(42)) or (inputs(4));
    layer0_outputs(3781) <= not(inputs(162));
    layer0_outputs(3782) <= not((inputs(65)) xor (inputs(90)));
    layer0_outputs(3783) <= inputs(99);
    layer0_outputs(3784) <= not((inputs(90)) xor (inputs(129)));
    layer0_outputs(3785) <= (inputs(97)) or (inputs(121));
    layer0_outputs(3786) <= inputs(150);
    layer0_outputs(3787) <= inputs(128);
    layer0_outputs(3788) <= not(inputs(46));
    layer0_outputs(3789) <= inputs(117);
    layer0_outputs(3790) <= inputs(21);
    layer0_outputs(3791) <= not(inputs(37));
    layer0_outputs(3792) <= inputs(110);
    layer0_outputs(3793) <= (inputs(79)) or (inputs(46));
    layer0_outputs(3794) <= not(inputs(83)) or (inputs(159));
    layer0_outputs(3795) <= inputs(16);
    layer0_outputs(3796) <= (inputs(189)) or (inputs(99));
    layer0_outputs(3797) <= not(inputs(164));
    layer0_outputs(3798) <= inputs(226);
    layer0_outputs(3799) <= (inputs(135)) xor (inputs(157));
    layer0_outputs(3800) <= not(inputs(78)) or (inputs(213));
    layer0_outputs(3801) <= inputs(167);
    layer0_outputs(3802) <= (inputs(165)) and (inputs(138));
    layer0_outputs(3803) <= (inputs(230)) or (inputs(7));
    layer0_outputs(3804) <= (inputs(209)) or (inputs(95));
    layer0_outputs(3805) <= (inputs(180)) xor (inputs(208));
    layer0_outputs(3806) <= not(inputs(89));
    layer0_outputs(3807) <= inputs(209);
    layer0_outputs(3808) <= not((inputs(111)) or (inputs(218)));
    layer0_outputs(3809) <= inputs(41);
    layer0_outputs(3810) <= not((inputs(210)) or (inputs(177)));
    layer0_outputs(3811) <= inputs(9);
    layer0_outputs(3812) <= not(inputs(183)) or (inputs(189));
    layer0_outputs(3813) <= (inputs(55)) and (inputs(158));
    layer0_outputs(3814) <= not(inputs(54)) or (inputs(56));
    layer0_outputs(3815) <= not((inputs(132)) xor (inputs(242)));
    layer0_outputs(3816) <= (inputs(169)) and not (inputs(38));
    layer0_outputs(3817) <= inputs(6);
    layer0_outputs(3818) <= (inputs(203)) xor (inputs(201));
    layer0_outputs(3819) <= not((inputs(101)) xor (inputs(237)));
    layer0_outputs(3820) <= (inputs(25)) and not (inputs(152));
    layer0_outputs(3821) <= inputs(231);
    layer0_outputs(3822) <= inputs(181);
    layer0_outputs(3823) <= (inputs(200)) xor (inputs(28));
    layer0_outputs(3824) <= (inputs(68)) or (inputs(156));
    layer0_outputs(3825) <= (inputs(168)) and not (inputs(61));
    layer0_outputs(3826) <= '0';
    layer0_outputs(3827) <= not((inputs(177)) xor (inputs(133)));
    layer0_outputs(3828) <= inputs(15);
    layer0_outputs(3829) <= (inputs(179)) and not (inputs(16));
    layer0_outputs(3830) <= not(inputs(41));
    layer0_outputs(3831) <= (inputs(99)) xor (inputs(54));
    layer0_outputs(3832) <= not((inputs(89)) xor (inputs(59)));
    layer0_outputs(3833) <= not((inputs(51)) or (inputs(16)));
    layer0_outputs(3834) <= '0';
    layer0_outputs(3835) <= not((inputs(177)) or (inputs(165)));
    layer0_outputs(3836) <= not(inputs(106)) or (inputs(242));
    layer0_outputs(3837) <= '0';
    layer0_outputs(3838) <= not(inputs(64)) or (inputs(124));
    layer0_outputs(3839) <= inputs(228);
    layer0_outputs(3840) <= inputs(151);
    layer0_outputs(3841) <= (inputs(164)) or (inputs(194));
    layer0_outputs(3842) <= (inputs(68)) xor (inputs(81));
    layer0_outputs(3843) <= not(inputs(200)) or (inputs(106));
    layer0_outputs(3844) <= (inputs(5)) xor (inputs(159));
    layer0_outputs(3845) <= inputs(211);
    layer0_outputs(3846) <= not((inputs(34)) xor (inputs(199)));
    layer0_outputs(3847) <= not((inputs(185)) and (inputs(246)));
    layer0_outputs(3848) <= not(inputs(92));
    layer0_outputs(3849) <= not(inputs(227)) or (inputs(93));
    layer0_outputs(3850) <= (inputs(170)) and (inputs(183));
    layer0_outputs(3851) <= not((inputs(255)) or (inputs(118)));
    layer0_outputs(3852) <= inputs(130);
    layer0_outputs(3853) <= not((inputs(219)) xor (inputs(161)));
    layer0_outputs(3854) <= not(inputs(87)) or (inputs(207));
    layer0_outputs(3855) <= not((inputs(194)) xor (inputs(48)));
    layer0_outputs(3856) <= not((inputs(194)) or (inputs(15)));
    layer0_outputs(3857) <= not((inputs(250)) or (inputs(37)));
    layer0_outputs(3858) <= (inputs(18)) or (inputs(174));
    layer0_outputs(3859) <= not(inputs(234));
    layer0_outputs(3860) <= not((inputs(135)) or (inputs(82)));
    layer0_outputs(3861) <= not((inputs(84)) or (inputs(213)));
    layer0_outputs(3862) <= not(inputs(247));
    layer0_outputs(3863) <= (inputs(218)) or (inputs(250));
    layer0_outputs(3864) <= (inputs(42)) xor (inputs(8));
    layer0_outputs(3865) <= (inputs(42)) and not (inputs(82));
    layer0_outputs(3866) <= not(inputs(9));
    layer0_outputs(3867) <= (inputs(0)) xor (inputs(230));
    layer0_outputs(3868) <= not((inputs(226)) or (inputs(43)));
    layer0_outputs(3869) <= (inputs(74)) and not (inputs(160));
    layer0_outputs(3870) <= not(inputs(40));
    layer0_outputs(3871) <= not(inputs(203)) or (inputs(75));
    layer0_outputs(3872) <= not((inputs(149)) and (inputs(222)));
    layer0_outputs(3873) <= (inputs(216)) and not (inputs(103));
    layer0_outputs(3874) <= not((inputs(244)) or (inputs(72)));
    layer0_outputs(3875) <= (inputs(4)) and not (inputs(96));
    layer0_outputs(3876) <= (inputs(85)) xor (inputs(132));
    layer0_outputs(3877) <= inputs(93);
    layer0_outputs(3878) <= not((inputs(93)) xor (inputs(206)));
    layer0_outputs(3879) <= (inputs(207)) xor (inputs(194));
    layer0_outputs(3880) <= not((inputs(169)) or (inputs(164)));
    layer0_outputs(3881) <= (inputs(117)) and not (inputs(205));
    layer0_outputs(3882) <= (inputs(104)) or (inputs(253));
    layer0_outputs(3883) <= not(inputs(244));
    layer0_outputs(3884) <= not((inputs(155)) xor (inputs(73)));
    layer0_outputs(3885) <= (inputs(208)) or (inputs(211));
    layer0_outputs(3886) <= (inputs(242)) xor (inputs(181));
    layer0_outputs(3887) <= inputs(192);
    layer0_outputs(3888) <= not(inputs(62)) or (inputs(104));
    layer0_outputs(3889) <= (inputs(212)) xor (inputs(222));
    layer0_outputs(3890) <= not((inputs(251)) or (inputs(137)));
    layer0_outputs(3891) <= not(inputs(146));
    layer0_outputs(3892) <= not((inputs(191)) and (inputs(177)));
    layer0_outputs(3893) <= (inputs(200)) and not (inputs(89));
    layer0_outputs(3894) <= not(inputs(177));
    layer0_outputs(3895) <= not(inputs(212));
    layer0_outputs(3896) <= not((inputs(23)) and (inputs(10)));
    layer0_outputs(3897) <= not(inputs(99));
    layer0_outputs(3898) <= (inputs(137)) and not (inputs(44));
    layer0_outputs(3899) <= not(inputs(229));
    layer0_outputs(3900) <= inputs(217);
    layer0_outputs(3901) <= (inputs(59)) or (inputs(253));
    layer0_outputs(3902) <= not(inputs(101));
    layer0_outputs(3903) <= (inputs(25)) and not (inputs(177));
    layer0_outputs(3904) <= inputs(113);
    layer0_outputs(3905) <= inputs(94);
    layer0_outputs(3906) <= not(inputs(40)) or (inputs(254));
    layer0_outputs(3907) <= (inputs(151)) or (inputs(147));
    layer0_outputs(3908) <= (inputs(86)) or (inputs(166));
    layer0_outputs(3909) <= inputs(51);
    layer0_outputs(3910) <= not((inputs(193)) or (inputs(191)));
    layer0_outputs(3911) <= not(inputs(112));
    layer0_outputs(3912) <= inputs(219);
    layer0_outputs(3913) <= not(inputs(199));
    layer0_outputs(3914) <= not((inputs(153)) xor (inputs(58)));
    layer0_outputs(3915) <= not(inputs(48)) or (inputs(207));
    layer0_outputs(3916) <= not((inputs(20)) or (inputs(202)));
    layer0_outputs(3917) <= not((inputs(238)) or (inputs(73)));
    layer0_outputs(3918) <= not((inputs(138)) or (inputs(97)));
    layer0_outputs(3919) <= not((inputs(252)) or (inputs(34)));
    layer0_outputs(3920) <= (inputs(193)) xor (inputs(179));
    layer0_outputs(3921) <= inputs(184);
    layer0_outputs(3922) <= (inputs(36)) or (inputs(107));
    layer0_outputs(3923) <= inputs(85);
    layer0_outputs(3924) <= (inputs(121)) and not (inputs(161));
    layer0_outputs(3925) <= not((inputs(39)) xor (inputs(232)));
    layer0_outputs(3926) <= not((inputs(55)) or (inputs(158)));
    layer0_outputs(3927) <= inputs(155);
    layer0_outputs(3928) <= inputs(120);
    layer0_outputs(3929) <= (inputs(64)) or (inputs(142));
    layer0_outputs(3930) <= (inputs(153)) and not (inputs(36));
    layer0_outputs(3931) <= not(inputs(119)) or (inputs(37));
    layer0_outputs(3932) <= not(inputs(24)) or (inputs(173));
    layer0_outputs(3933) <= not((inputs(17)) or (inputs(40)));
    layer0_outputs(3934) <= (inputs(209)) and not (inputs(128));
    layer0_outputs(3935) <= (inputs(226)) or (inputs(48));
    layer0_outputs(3936) <= not(inputs(224)) or (inputs(83));
    layer0_outputs(3937) <= inputs(30);
    layer0_outputs(3938) <= not(inputs(165));
    layer0_outputs(3939) <= inputs(54);
    layer0_outputs(3940) <= inputs(28);
    layer0_outputs(3941) <= not(inputs(3));
    layer0_outputs(3942) <= (inputs(251)) or (inputs(241));
    layer0_outputs(3943) <= not((inputs(18)) xor (inputs(168)));
    layer0_outputs(3944) <= (inputs(167)) and not (inputs(43));
    layer0_outputs(3945) <= (inputs(27)) and not (inputs(25));
    layer0_outputs(3946) <= not((inputs(215)) or (inputs(95)));
    layer0_outputs(3947) <= (inputs(184)) and (inputs(220));
    layer0_outputs(3948) <= not(inputs(219));
    layer0_outputs(3949) <= not(inputs(168));
    layer0_outputs(3950) <= not(inputs(26)) or (inputs(165));
    layer0_outputs(3951) <= not((inputs(236)) xor (inputs(9)));
    layer0_outputs(3952) <= not(inputs(123));
    layer0_outputs(3953) <= not(inputs(45));
    layer0_outputs(3954) <= (inputs(178)) and not (inputs(48));
    layer0_outputs(3955) <= not(inputs(211)) or (inputs(122));
    layer0_outputs(3956) <= not((inputs(154)) or (inputs(198)));
    layer0_outputs(3957) <= not((inputs(205)) xor (inputs(109)));
    layer0_outputs(3958) <= not((inputs(118)) or (inputs(26)));
    layer0_outputs(3959) <= not((inputs(210)) and (inputs(154)));
    layer0_outputs(3960) <= (inputs(66)) and (inputs(35));
    layer0_outputs(3961) <= not(inputs(176));
    layer0_outputs(3962) <= inputs(152);
    layer0_outputs(3963) <= (inputs(206)) or (inputs(239));
    layer0_outputs(3964) <= not(inputs(12));
    layer0_outputs(3965) <= (inputs(48)) or (inputs(192));
    layer0_outputs(3966) <= inputs(3);
    layer0_outputs(3967) <= not((inputs(52)) or (inputs(84)));
    layer0_outputs(3968) <= not(inputs(100));
    layer0_outputs(3969) <= not((inputs(194)) or (inputs(65)));
    layer0_outputs(3970) <= (inputs(80)) xor (inputs(86));
    layer0_outputs(3971) <= inputs(52);
    layer0_outputs(3972) <= (inputs(22)) or (inputs(206));
    layer0_outputs(3973) <= not(inputs(137)) or (inputs(48));
    layer0_outputs(3974) <= not(inputs(111));
    layer0_outputs(3975) <= (inputs(147)) xor (inputs(182));
    layer0_outputs(3976) <= not((inputs(20)) or (inputs(171)));
    layer0_outputs(3977) <= not((inputs(17)) xor (inputs(243)));
    layer0_outputs(3978) <= (inputs(27)) or (inputs(52));
    layer0_outputs(3979) <= (inputs(121)) and not (inputs(21));
    layer0_outputs(3980) <= not(inputs(55));
    layer0_outputs(3981) <= not((inputs(48)) xor (inputs(9)));
    layer0_outputs(3982) <= not(inputs(230));
    layer0_outputs(3983) <= not((inputs(122)) and (inputs(187)));
    layer0_outputs(3984) <= (inputs(166)) and not (inputs(209));
    layer0_outputs(3985) <= not(inputs(151)) or (inputs(252));
    layer0_outputs(3986) <= not((inputs(131)) and (inputs(115)));
    layer0_outputs(3987) <= not((inputs(144)) or (inputs(235)));
    layer0_outputs(3988) <= not((inputs(7)) or (inputs(223)));
    layer0_outputs(3989) <= (inputs(178)) or (inputs(20));
    layer0_outputs(3990) <= not((inputs(249)) or (inputs(127)));
    layer0_outputs(3991) <= not(inputs(12)) or (inputs(108));
    layer0_outputs(3992) <= inputs(247);
    layer0_outputs(3993) <= (inputs(5)) and not (inputs(254));
    layer0_outputs(3994) <= (inputs(245)) or (inputs(158));
    layer0_outputs(3995) <= inputs(137);
    layer0_outputs(3996) <= (inputs(126)) and not (inputs(239));
    layer0_outputs(3997) <= (inputs(27)) and (inputs(169));
    layer0_outputs(3998) <= inputs(98);
    layer0_outputs(3999) <= not((inputs(237)) xor (inputs(101)));
    layer0_outputs(4000) <= '1';
    layer0_outputs(4001) <= inputs(238);
    layer0_outputs(4002) <= not((inputs(188)) xor (inputs(8)));
    layer0_outputs(4003) <= not(inputs(213)) or (inputs(6));
    layer0_outputs(4004) <= not(inputs(179));
    layer0_outputs(4005) <= (inputs(148)) xor (inputs(102));
    layer0_outputs(4006) <= (inputs(239)) or (inputs(66));
    layer0_outputs(4007) <= inputs(183);
    layer0_outputs(4008) <= not(inputs(197));
    layer0_outputs(4009) <= (inputs(126)) xor (inputs(190));
    layer0_outputs(4010) <= (inputs(101)) and not (inputs(238));
    layer0_outputs(4011) <= not(inputs(11)) or (inputs(43));
    layer0_outputs(4012) <= (inputs(147)) or (inputs(34));
    layer0_outputs(4013) <= '1';
    layer0_outputs(4014) <= not((inputs(10)) or (inputs(248)));
    layer0_outputs(4015) <= not((inputs(159)) or (inputs(216)));
    layer0_outputs(4016) <= (inputs(139)) and not (inputs(66));
    layer0_outputs(4017) <= not(inputs(150));
    layer0_outputs(4018) <= not(inputs(103));
    layer0_outputs(4019) <= not((inputs(5)) xor (inputs(93)));
    layer0_outputs(4020) <= not((inputs(129)) xor (inputs(40)));
    layer0_outputs(4021) <= not((inputs(126)) or (inputs(185)));
    layer0_outputs(4022) <= (inputs(245)) and not (inputs(38));
    layer0_outputs(4023) <= (inputs(205)) xor (inputs(10));
    layer0_outputs(4024) <= not(inputs(194));
    layer0_outputs(4025) <= (inputs(36)) and not (inputs(87));
    layer0_outputs(4026) <= not(inputs(145));
    layer0_outputs(4027) <= not(inputs(170)) or (inputs(17));
    layer0_outputs(4028) <= not((inputs(247)) and (inputs(188)));
    layer0_outputs(4029) <= not(inputs(74)) or (inputs(144));
    layer0_outputs(4030) <= not((inputs(45)) xor (inputs(27)));
    layer0_outputs(4031) <= (inputs(74)) and not (inputs(254));
    layer0_outputs(4032) <= not(inputs(116));
    layer0_outputs(4033) <= (inputs(128)) or (inputs(7));
    layer0_outputs(4034) <= not((inputs(31)) or (inputs(234)));
    layer0_outputs(4035) <= not(inputs(179));
    layer0_outputs(4036) <= (inputs(24)) xor (inputs(74));
    layer0_outputs(4037) <= not(inputs(74));
    layer0_outputs(4038) <= not((inputs(33)) or (inputs(201)));
    layer0_outputs(4039) <= not((inputs(251)) xor (inputs(208)));
    layer0_outputs(4040) <= not(inputs(196)) or (inputs(46));
    layer0_outputs(4041) <= (inputs(51)) and not (inputs(0));
    layer0_outputs(4042) <= not(inputs(169));
    layer0_outputs(4043) <= not(inputs(182)) or (inputs(75));
    layer0_outputs(4044) <= not((inputs(18)) or (inputs(79)));
    layer0_outputs(4045) <= not((inputs(27)) xor (inputs(135)));
    layer0_outputs(4046) <= not((inputs(195)) or (inputs(42)));
    layer0_outputs(4047) <= (inputs(86)) and (inputs(104));
    layer0_outputs(4048) <= (inputs(85)) xor (inputs(66));
    layer0_outputs(4049) <= (inputs(18)) and (inputs(163));
    layer0_outputs(4050) <= (inputs(121)) xor (inputs(103));
    layer0_outputs(4051) <= not((inputs(83)) xor (inputs(81)));
    layer0_outputs(4052) <= not(inputs(90)) or (inputs(238));
    layer0_outputs(4053) <= not((inputs(78)) xor (inputs(63)));
    layer0_outputs(4054) <= not((inputs(102)) xor (inputs(100)));
    layer0_outputs(4055) <= not(inputs(154));
    layer0_outputs(4056) <= not(inputs(2)) or (inputs(64));
    layer0_outputs(4057) <= (inputs(84)) or (inputs(12));
    layer0_outputs(4058) <= not(inputs(136));
    layer0_outputs(4059) <= not((inputs(158)) or (inputs(247)));
    layer0_outputs(4060) <= inputs(86);
    layer0_outputs(4061) <= (inputs(2)) xor (inputs(109));
    layer0_outputs(4062) <= (inputs(151)) or (inputs(146));
    layer0_outputs(4063) <= not(inputs(248));
    layer0_outputs(4064) <= not(inputs(194)) or (inputs(142));
    layer0_outputs(4065) <= not((inputs(102)) xor (inputs(175)));
    layer0_outputs(4066) <= not((inputs(85)) or (inputs(84)));
    layer0_outputs(4067) <= (inputs(182)) and not (inputs(67));
    layer0_outputs(4068) <= (inputs(173)) or (inputs(101));
    layer0_outputs(4069) <= not(inputs(90));
    layer0_outputs(4070) <= (inputs(87)) and not (inputs(188));
    layer0_outputs(4071) <= (inputs(174)) xor (inputs(68));
    layer0_outputs(4072) <= (inputs(235)) and not (inputs(123));
    layer0_outputs(4073) <= not((inputs(240)) xor (inputs(22)));
    layer0_outputs(4074) <= inputs(187);
    layer0_outputs(4075) <= not((inputs(208)) xor (inputs(248)));
    layer0_outputs(4076) <= (inputs(7)) or (inputs(66));
    layer0_outputs(4077) <= '1';
    layer0_outputs(4078) <= not(inputs(206)) or (inputs(214));
    layer0_outputs(4079) <= (inputs(127)) or (inputs(147));
    layer0_outputs(4080) <= not((inputs(73)) xor (inputs(22)));
    layer0_outputs(4081) <= inputs(12);
    layer0_outputs(4082) <= not((inputs(180)) or (inputs(184)));
    layer0_outputs(4083) <= not((inputs(19)) or (inputs(237)));
    layer0_outputs(4084) <= not((inputs(89)) xor (inputs(223)));
    layer0_outputs(4085) <= inputs(226);
    layer0_outputs(4086) <= not((inputs(154)) or (inputs(137)));
    layer0_outputs(4087) <= not(inputs(150));
    layer0_outputs(4088) <= (inputs(88)) xor (inputs(182));
    layer0_outputs(4089) <= (inputs(128)) or (inputs(146));
    layer0_outputs(4090) <= (inputs(191)) or (inputs(133));
    layer0_outputs(4091) <= (inputs(224)) xor (inputs(205));
    layer0_outputs(4092) <= (inputs(145)) xor (inputs(128));
    layer0_outputs(4093) <= not(inputs(244)) or (inputs(82));
    layer0_outputs(4094) <= not((inputs(247)) or (inputs(202)));
    layer0_outputs(4095) <= not((inputs(87)) or (inputs(246)));
    layer0_outputs(4096) <= not((inputs(153)) or (inputs(187)));
    layer0_outputs(4097) <= not((inputs(204)) xor (inputs(179)));
    layer0_outputs(4098) <= not((inputs(146)) xor (inputs(241)));
    layer0_outputs(4099) <= not((inputs(178)) or (inputs(70)));
    layer0_outputs(4100) <= (inputs(160)) xor (inputs(49));
    layer0_outputs(4101) <= not(inputs(71)) or (inputs(149));
    layer0_outputs(4102) <= not(inputs(201)) or (inputs(52));
    layer0_outputs(4103) <= inputs(255);
    layer0_outputs(4104) <= (inputs(219)) or (inputs(243));
    layer0_outputs(4105) <= not(inputs(129));
    layer0_outputs(4106) <= (inputs(77)) and not (inputs(136));
    layer0_outputs(4107) <= not((inputs(190)) or (inputs(118)));
    layer0_outputs(4108) <= not(inputs(40));
    layer0_outputs(4109) <= (inputs(157)) and not (inputs(55));
    layer0_outputs(4110) <= inputs(72);
    layer0_outputs(4111) <= not(inputs(222));
    layer0_outputs(4112) <= (inputs(100)) and not (inputs(201));
    layer0_outputs(4113) <= (inputs(26)) or (inputs(41));
    layer0_outputs(4114) <= (inputs(33)) or (inputs(197));
    layer0_outputs(4115) <= (inputs(138)) and not (inputs(245));
    layer0_outputs(4116) <= (inputs(230)) and not (inputs(49));
    layer0_outputs(4117) <= not(inputs(36));
    layer0_outputs(4118) <= (inputs(62)) xor (inputs(125));
    layer0_outputs(4119) <= (inputs(129)) xor (inputs(118));
    layer0_outputs(4120) <= (inputs(254)) or (inputs(7));
    layer0_outputs(4121) <= not(inputs(3)) or (inputs(96));
    layer0_outputs(4122) <= not(inputs(165));
    layer0_outputs(4123) <= (inputs(20)) and not (inputs(178));
    layer0_outputs(4124) <= (inputs(120)) xor (inputs(203));
    layer0_outputs(4125) <= (inputs(47)) xor (inputs(8));
    layer0_outputs(4126) <= not(inputs(194));
    layer0_outputs(4127) <= inputs(79);
    layer0_outputs(4128) <= (inputs(87)) or (inputs(73));
    layer0_outputs(4129) <= (inputs(95)) and not (inputs(237));
    layer0_outputs(4130) <= inputs(81);
    layer0_outputs(4131) <= (inputs(23)) xor (inputs(73));
    layer0_outputs(4132) <= not((inputs(48)) or (inputs(154)));
    layer0_outputs(4133) <= not(inputs(228)) or (inputs(211));
    layer0_outputs(4134) <= not(inputs(186));
    layer0_outputs(4135) <= inputs(192);
    layer0_outputs(4136) <= not(inputs(39)) or (inputs(144));
    layer0_outputs(4137) <= not(inputs(212)) or (inputs(87));
    layer0_outputs(4138) <= (inputs(181)) and not (inputs(98));
    layer0_outputs(4139) <= inputs(5);
    layer0_outputs(4140) <= (inputs(182)) and not (inputs(54));
    layer0_outputs(4141) <= inputs(94);
    layer0_outputs(4142) <= (inputs(76)) and not (inputs(127));
    layer0_outputs(4143) <= (inputs(11)) xor (inputs(16));
    layer0_outputs(4144) <= not(inputs(227));
    layer0_outputs(4145) <= (inputs(116)) or (inputs(146));
    layer0_outputs(4146) <= (inputs(91)) or (inputs(72));
    layer0_outputs(4147) <= not((inputs(3)) or (inputs(176)));
    layer0_outputs(4148) <= not((inputs(18)) or (inputs(119)));
    layer0_outputs(4149) <= (inputs(69)) and not (inputs(223));
    layer0_outputs(4150) <= '1';
    layer0_outputs(4151) <= (inputs(15)) or (inputs(194));
    layer0_outputs(4152) <= (inputs(35)) or (inputs(17));
    layer0_outputs(4153) <= inputs(38);
    layer0_outputs(4154) <= (inputs(151)) or (inputs(222));
    layer0_outputs(4155) <= (inputs(100)) or (inputs(156));
    layer0_outputs(4156) <= not((inputs(169)) xor (inputs(224)));
    layer0_outputs(4157) <= inputs(136);
    layer0_outputs(4158) <= inputs(10);
    layer0_outputs(4159) <= (inputs(4)) xor (inputs(77));
    layer0_outputs(4160) <= (inputs(220)) xor (inputs(71));
    layer0_outputs(4161) <= inputs(102);
    layer0_outputs(4162) <= not(inputs(30)) or (inputs(16));
    layer0_outputs(4163) <= (inputs(164)) and not (inputs(62));
    layer0_outputs(4164) <= (inputs(124)) and (inputs(83));
    layer0_outputs(4165) <= (inputs(97)) or (inputs(9));
    layer0_outputs(4166) <= (inputs(156)) or (inputs(102));
    layer0_outputs(4167) <= not(inputs(222));
    layer0_outputs(4168) <= (inputs(202)) or (inputs(174));
    layer0_outputs(4169) <= not(inputs(84)) or (inputs(47));
    layer0_outputs(4170) <= not(inputs(203));
    layer0_outputs(4171) <= (inputs(102)) or (inputs(146));
    layer0_outputs(4172) <= not(inputs(164));
    layer0_outputs(4173) <= (inputs(199)) and not (inputs(96));
    layer0_outputs(4174) <= inputs(80);
    layer0_outputs(4175) <= inputs(230);
    layer0_outputs(4176) <= not(inputs(69));
    layer0_outputs(4177) <= not(inputs(131));
    layer0_outputs(4178) <= (inputs(194)) xor (inputs(24));
    layer0_outputs(4179) <= (inputs(123)) and not (inputs(163));
    layer0_outputs(4180) <= not(inputs(71)) or (inputs(80));
    layer0_outputs(4181) <= (inputs(99)) xor (inputs(11));
    layer0_outputs(4182) <= not(inputs(104));
    layer0_outputs(4183) <= not(inputs(73));
    layer0_outputs(4184) <= not(inputs(213)) or (inputs(13));
    layer0_outputs(4185) <= (inputs(114)) and not (inputs(65));
    layer0_outputs(4186) <= (inputs(60)) or (inputs(155));
    layer0_outputs(4187) <= (inputs(169)) and not (inputs(187));
    layer0_outputs(4188) <= inputs(202);
    layer0_outputs(4189) <= (inputs(227)) or (inputs(253));
    layer0_outputs(4190) <= not(inputs(99)) or (inputs(31));
    layer0_outputs(4191) <= inputs(246);
    layer0_outputs(4192) <= (inputs(210)) and not (inputs(112));
    layer0_outputs(4193) <= (inputs(84)) and not (inputs(229));
    layer0_outputs(4194) <= (inputs(243)) xor (inputs(177));
    layer0_outputs(4195) <= inputs(136);
    layer0_outputs(4196) <= (inputs(149)) and not (inputs(123));
    layer0_outputs(4197) <= (inputs(227)) or (inputs(178));
    layer0_outputs(4198) <= (inputs(19)) and not (inputs(129));
    layer0_outputs(4199) <= not(inputs(1));
    layer0_outputs(4200) <= not(inputs(26));
    layer0_outputs(4201) <= not(inputs(101));
    layer0_outputs(4202) <= inputs(134);
    layer0_outputs(4203) <= (inputs(24)) and not (inputs(189));
    layer0_outputs(4204) <= '1';
    layer0_outputs(4205) <= (inputs(152)) or (inputs(56));
    layer0_outputs(4206) <= not(inputs(136));
    layer0_outputs(4207) <= not(inputs(100)) or (inputs(193));
    layer0_outputs(4208) <= (inputs(93)) xor (inputs(64));
    layer0_outputs(4209) <= (inputs(233)) and (inputs(3));
    layer0_outputs(4210) <= not((inputs(97)) or (inputs(125)));
    layer0_outputs(4211) <= not((inputs(50)) or (inputs(3)));
    layer0_outputs(4212) <= not(inputs(235)) or (inputs(139));
    layer0_outputs(4213) <= not(inputs(233)) or (inputs(15));
    layer0_outputs(4214) <= not((inputs(232)) or (inputs(79)));
    layer0_outputs(4215) <= inputs(23);
    layer0_outputs(4216) <= not(inputs(53));
    layer0_outputs(4217) <= not(inputs(24)) or (inputs(245));
    layer0_outputs(4218) <= inputs(109);
    layer0_outputs(4219) <= (inputs(156)) or (inputs(243));
    layer0_outputs(4220) <= (inputs(93)) or (inputs(242));
    layer0_outputs(4221) <= not(inputs(209));
    layer0_outputs(4222) <= not(inputs(213));
    layer0_outputs(4223) <= inputs(232);
    layer0_outputs(4224) <= (inputs(10)) and not (inputs(187));
    layer0_outputs(4225) <= inputs(212);
    layer0_outputs(4226) <= not(inputs(23));
    layer0_outputs(4227) <= not(inputs(74));
    layer0_outputs(4228) <= '0';
    layer0_outputs(4229) <= (inputs(196)) xor (inputs(238));
    layer0_outputs(4230) <= not(inputs(25));
    layer0_outputs(4231) <= not(inputs(101));
    layer0_outputs(4232) <= not(inputs(59)) or (inputs(127));
    layer0_outputs(4233) <= not(inputs(119)) or (inputs(155));
    layer0_outputs(4234) <= (inputs(225)) xor (inputs(78));
    layer0_outputs(4235) <= not((inputs(74)) xor (inputs(187)));
    layer0_outputs(4236) <= (inputs(24)) and not (inputs(244));
    layer0_outputs(4237) <= (inputs(210)) or (inputs(191));
    layer0_outputs(4238) <= inputs(166);
    layer0_outputs(4239) <= (inputs(228)) or (inputs(230));
    layer0_outputs(4240) <= (inputs(195)) xor (inputs(63));
    layer0_outputs(4241) <= inputs(185);
    layer0_outputs(4242) <= (inputs(255)) or (inputs(170));
    layer0_outputs(4243) <= not(inputs(42)) or (inputs(145));
    layer0_outputs(4244) <= not(inputs(98)) or (inputs(199));
    layer0_outputs(4245) <= inputs(11);
    layer0_outputs(4246) <= not((inputs(255)) or (inputs(50)));
    layer0_outputs(4247) <= (inputs(109)) or (inputs(63));
    layer0_outputs(4248) <= not((inputs(221)) xor (inputs(251)));
    layer0_outputs(4249) <= not(inputs(5)) or (inputs(52));
    layer0_outputs(4250) <= not(inputs(55));
    layer0_outputs(4251) <= (inputs(238)) and not (inputs(116));
    layer0_outputs(4252) <= not((inputs(233)) or (inputs(227)));
    layer0_outputs(4253) <= not((inputs(121)) xor (inputs(61)));
    layer0_outputs(4254) <= (inputs(125)) and not (inputs(37));
    layer0_outputs(4255) <= not((inputs(48)) and (inputs(17)));
    layer0_outputs(4256) <= '1';
    layer0_outputs(4257) <= (inputs(179)) or (inputs(105));
    layer0_outputs(4258) <= inputs(19);
    layer0_outputs(4259) <= inputs(70);
    layer0_outputs(4260) <= not((inputs(197)) or (inputs(157)));
    layer0_outputs(4261) <= not(inputs(136)) or (inputs(15));
    layer0_outputs(4262) <= not(inputs(74));
    layer0_outputs(4263) <= not((inputs(172)) or (inputs(143)));
    layer0_outputs(4264) <= not((inputs(111)) xor (inputs(140)));
    layer0_outputs(4265) <= (inputs(42)) xor (inputs(77));
    layer0_outputs(4266) <= (inputs(229)) xor (inputs(48));
    layer0_outputs(4267) <= (inputs(180)) xor (inputs(215));
    layer0_outputs(4268) <= not((inputs(147)) and (inputs(219)));
    layer0_outputs(4269) <= not(inputs(201));
    layer0_outputs(4270) <= inputs(1);
    layer0_outputs(4271) <= (inputs(163)) and not (inputs(172));
    layer0_outputs(4272) <= not(inputs(231)) or (inputs(84));
    layer0_outputs(4273) <= (inputs(180)) xor (inputs(217));
    layer0_outputs(4274) <= (inputs(68)) and not (inputs(254));
    layer0_outputs(4275) <= (inputs(49)) or (inputs(186));
    layer0_outputs(4276) <= inputs(246);
    layer0_outputs(4277) <= (inputs(228)) xor (inputs(172));
    layer0_outputs(4278) <= inputs(141);
    layer0_outputs(4279) <= inputs(117);
    layer0_outputs(4280) <= not(inputs(67)) or (inputs(216));
    layer0_outputs(4281) <= not(inputs(246)) or (inputs(223));
    layer0_outputs(4282) <= not((inputs(213)) and (inputs(163)));
    layer0_outputs(4283) <= (inputs(130)) or (inputs(182));
    layer0_outputs(4284) <= not((inputs(188)) or (inputs(157)));
    layer0_outputs(4285) <= inputs(96);
    layer0_outputs(4286) <= (inputs(213)) and not (inputs(30));
    layer0_outputs(4287) <= inputs(94);
    layer0_outputs(4288) <= inputs(178);
    layer0_outputs(4289) <= '1';
    layer0_outputs(4290) <= not(inputs(225)) or (inputs(48));
    layer0_outputs(4291) <= (inputs(243)) xor (inputs(175));
    layer0_outputs(4292) <= not(inputs(71));
    layer0_outputs(4293) <= not(inputs(148));
    layer0_outputs(4294) <= (inputs(21)) or (inputs(142));
    layer0_outputs(4295) <= not(inputs(145));
    layer0_outputs(4296) <= inputs(254);
    layer0_outputs(4297) <= inputs(135);
    layer0_outputs(4298) <= not(inputs(146));
    layer0_outputs(4299) <= (inputs(12)) and not (inputs(242));
    layer0_outputs(4300) <= not(inputs(142));
    layer0_outputs(4301) <= (inputs(232)) and (inputs(191));
    layer0_outputs(4302) <= inputs(230);
    layer0_outputs(4303) <= not(inputs(204)) or (inputs(65));
    layer0_outputs(4304) <= inputs(167);
    layer0_outputs(4305) <= (inputs(158)) and not (inputs(83));
    layer0_outputs(4306) <= (inputs(138)) or (inputs(19));
    layer0_outputs(4307) <= (inputs(241)) and (inputs(111));
    layer0_outputs(4308) <= (inputs(199)) or (inputs(1));
    layer0_outputs(4309) <= inputs(109);
    layer0_outputs(4310) <= (inputs(46)) and (inputs(28));
    layer0_outputs(4311) <= inputs(50);
    layer0_outputs(4312) <= (inputs(125)) xor (inputs(174));
    layer0_outputs(4313) <= not((inputs(34)) or (inputs(205)));
    layer0_outputs(4314) <= not((inputs(244)) or (inputs(242)));
    layer0_outputs(4315) <= not((inputs(50)) or (inputs(12)));
    layer0_outputs(4316) <= not(inputs(179)) or (inputs(35));
    layer0_outputs(4317) <= not((inputs(58)) xor (inputs(43)));
    layer0_outputs(4318) <= not((inputs(208)) or (inputs(214)));
    layer0_outputs(4319) <= not(inputs(127)) or (inputs(239));
    layer0_outputs(4320) <= not(inputs(121));
    layer0_outputs(4321) <= inputs(21);
    layer0_outputs(4322) <= not((inputs(24)) or (inputs(28)));
    layer0_outputs(4323) <= inputs(121);
    layer0_outputs(4324) <= not(inputs(27));
    layer0_outputs(4325) <= (inputs(20)) xor (inputs(53));
    layer0_outputs(4326) <= not(inputs(59)) or (inputs(121));
    layer0_outputs(4327) <= not(inputs(169)) or (inputs(133));
    layer0_outputs(4328) <= not((inputs(86)) xor (inputs(121)));
    layer0_outputs(4329) <= not(inputs(66));
    layer0_outputs(4330) <= (inputs(136)) xor (inputs(89));
    layer0_outputs(4331) <= not((inputs(5)) or (inputs(216)));
    layer0_outputs(4332) <= not(inputs(229)) or (inputs(170));
    layer0_outputs(4333) <= inputs(207);
    layer0_outputs(4334) <= not(inputs(178));
    layer0_outputs(4335) <= not(inputs(103));
    layer0_outputs(4336) <= not((inputs(110)) or (inputs(49)));
    layer0_outputs(4337) <= (inputs(177)) xor (inputs(26));
    layer0_outputs(4338) <= (inputs(120)) xor (inputs(98));
    layer0_outputs(4339) <= not((inputs(50)) or (inputs(217)));
    layer0_outputs(4340) <= inputs(165);
    layer0_outputs(4341) <= inputs(210);
    layer0_outputs(4342) <= (inputs(212)) or (inputs(159));
    layer0_outputs(4343) <= inputs(140);
    layer0_outputs(4344) <= not(inputs(90));
    layer0_outputs(4345) <= not(inputs(102));
    layer0_outputs(4346) <= (inputs(195)) and not (inputs(170));
    layer0_outputs(4347) <= not((inputs(227)) xor (inputs(130)));
    layer0_outputs(4348) <= not((inputs(134)) xor (inputs(152)));
    layer0_outputs(4349) <= (inputs(120)) and not (inputs(145));
    layer0_outputs(4350) <= not(inputs(67));
    layer0_outputs(4351) <= not((inputs(216)) or (inputs(106)));
    layer0_outputs(4352) <= (inputs(117)) and not (inputs(173));
    layer0_outputs(4353) <= not((inputs(178)) or (inputs(12)));
    layer0_outputs(4354) <= (inputs(42)) and not (inputs(145));
    layer0_outputs(4355) <= not(inputs(230));
    layer0_outputs(4356) <= not((inputs(156)) or (inputs(11)));
    layer0_outputs(4357) <= not(inputs(165));
    layer0_outputs(4358) <= not(inputs(211)) or (inputs(6));
    layer0_outputs(4359) <= not(inputs(181));
    layer0_outputs(4360) <= inputs(76);
    layer0_outputs(4361) <= not((inputs(223)) xor (inputs(87)));
    layer0_outputs(4362) <= (inputs(182)) or (inputs(196));
    layer0_outputs(4363) <= not((inputs(222)) or (inputs(205)));
    layer0_outputs(4364) <= not(inputs(136));
    layer0_outputs(4365) <= not(inputs(165));
    layer0_outputs(4366) <= not(inputs(91));
    layer0_outputs(4367) <= not((inputs(152)) or (inputs(73)));
    layer0_outputs(4368) <= not((inputs(92)) or (inputs(8)));
    layer0_outputs(4369) <= inputs(133);
    layer0_outputs(4370) <= not(inputs(196)) or (inputs(117));
    layer0_outputs(4371) <= (inputs(61)) xor (inputs(108));
    layer0_outputs(4372) <= (inputs(180)) and not (inputs(94));
    layer0_outputs(4373) <= not(inputs(33)) or (inputs(135));
    layer0_outputs(4374) <= not((inputs(167)) or (inputs(110)));
    layer0_outputs(4375) <= not(inputs(56));
    layer0_outputs(4376) <= not(inputs(148));
    layer0_outputs(4377) <= inputs(136);
    layer0_outputs(4378) <= not((inputs(156)) or (inputs(133)));
    layer0_outputs(4379) <= inputs(135);
    layer0_outputs(4380) <= (inputs(89)) or (inputs(21));
    layer0_outputs(4381) <= (inputs(168)) xor (inputs(130));
    layer0_outputs(4382) <= (inputs(52)) and not (inputs(113));
    layer0_outputs(4383) <= inputs(132);
    layer0_outputs(4384) <= inputs(193);
    layer0_outputs(4385) <= (inputs(96)) and (inputs(238));
    layer0_outputs(4386) <= not(inputs(126));
    layer0_outputs(4387) <= not(inputs(5));
    layer0_outputs(4388) <= (inputs(45)) or (inputs(13));
    layer0_outputs(4389) <= not(inputs(127));
    layer0_outputs(4390) <= not((inputs(73)) xor (inputs(123)));
    layer0_outputs(4391) <= not(inputs(46)) or (inputs(253));
    layer0_outputs(4392) <= not(inputs(235));
    layer0_outputs(4393) <= inputs(195);
    layer0_outputs(4394) <= not(inputs(145));
    layer0_outputs(4395) <= inputs(39);
    layer0_outputs(4396) <= not(inputs(212));
    layer0_outputs(4397) <= not((inputs(68)) xor (inputs(221)));
    layer0_outputs(4398) <= not((inputs(2)) xor (inputs(130)));
    layer0_outputs(4399) <= not(inputs(227));
    layer0_outputs(4400) <= not(inputs(155));
    layer0_outputs(4401) <= inputs(171);
    layer0_outputs(4402) <= (inputs(87)) xor (inputs(41));
    layer0_outputs(4403) <= not(inputs(166));
    layer0_outputs(4404) <= (inputs(76)) and not (inputs(204));
    layer0_outputs(4405) <= not((inputs(147)) xor (inputs(197)));
    layer0_outputs(4406) <= inputs(97);
    layer0_outputs(4407) <= (inputs(229)) and not (inputs(65));
    layer0_outputs(4408) <= not(inputs(253));
    layer0_outputs(4409) <= not((inputs(18)) or (inputs(224)));
    layer0_outputs(4410) <= (inputs(27)) and not (inputs(253));
    layer0_outputs(4411) <= not(inputs(30));
    layer0_outputs(4412) <= (inputs(35)) and not (inputs(143));
    layer0_outputs(4413) <= (inputs(252)) and not (inputs(249));
    layer0_outputs(4414) <= not(inputs(210));
    layer0_outputs(4415) <= (inputs(17)) xor (inputs(144));
    layer0_outputs(4416) <= inputs(85);
    layer0_outputs(4417) <= inputs(56);
    layer0_outputs(4418) <= not((inputs(3)) or (inputs(165)));
    layer0_outputs(4419) <= (inputs(225)) xor (inputs(168));
    layer0_outputs(4420) <= (inputs(149)) and not (inputs(81));
    layer0_outputs(4421) <= not(inputs(252)) or (inputs(219));
    layer0_outputs(4422) <= inputs(52);
    layer0_outputs(4423) <= not(inputs(244));
    layer0_outputs(4424) <= not((inputs(253)) xor (inputs(151)));
    layer0_outputs(4425) <= not(inputs(254));
    layer0_outputs(4426) <= inputs(78);
    layer0_outputs(4427) <= not((inputs(170)) or (inputs(60)));
    layer0_outputs(4428) <= not((inputs(78)) or (inputs(43)));
    layer0_outputs(4429) <= (inputs(62)) xor (inputs(59));
    layer0_outputs(4430) <= not(inputs(226)) or (inputs(132));
    layer0_outputs(4431) <= not(inputs(56));
    layer0_outputs(4432) <= (inputs(35)) and not (inputs(78));
    layer0_outputs(4433) <= inputs(116);
    layer0_outputs(4434) <= (inputs(3)) and not (inputs(254));
    layer0_outputs(4435) <= not((inputs(83)) or (inputs(11)));
    layer0_outputs(4436) <= not(inputs(188)) or (inputs(50));
    layer0_outputs(4437) <= not(inputs(101));
    layer0_outputs(4438) <= inputs(161);
    layer0_outputs(4439) <= (inputs(28)) or (inputs(5));
    layer0_outputs(4440) <= inputs(145);
    layer0_outputs(4441) <= not(inputs(57)) or (inputs(193));
    layer0_outputs(4442) <= not(inputs(7)) or (inputs(70));
    layer0_outputs(4443) <= not((inputs(162)) or (inputs(99)));
    layer0_outputs(4444) <= not((inputs(119)) or (inputs(244)));
    layer0_outputs(4445) <= (inputs(58)) xor (inputs(55));
    layer0_outputs(4446) <= inputs(161);
    layer0_outputs(4447) <= not((inputs(47)) or (inputs(18)));
    layer0_outputs(4448) <= inputs(233);
    layer0_outputs(4449) <= inputs(107);
    layer0_outputs(4450) <= (inputs(86)) or (inputs(1));
    layer0_outputs(4451) <= '1';
    layer0_outputs(4452) <= not((inputs(88)) or (inputs(66)));
    layer0_outputs(4453) <= not(inputs(132));
    layer0_outputs(4454) <= inputs(23);
    layer0_outputs(4455) <= (inputs(75)) and not (inputs(167));
    layer0_outputs(4456) <= (inputs(22)) or (inputs(79));
    layer0_outputs(4457) <= inputs(8);
    layer0_outputs(4458) <= not((inputs(231)) or (inputs(40)));
    layer0_outputs(4459) <= not((inputs(134)) xor (inputs(12)));
    layer0_outputs(4460) <= (inputs(209)) or (inputs(187));
    layer0_outputs(4461) <= (inputs(225)) or (inputs(220));
    layer0_outputs(4462) <= (inputs(113)) or (inputs(112));
    layer0_outputs(4463) <= inputs(14);
    layer0_outputs(4464) <= not(inputs(84)) or (inputs(228));
    layer0_outputs(4465) <= (inputs(51)) or (inputs(125));
    layer0_outputs(4466) <= inputs(71);
    layer0_outputs(4467) <= not((inputs(53)) or (inputs(98)));
    layer0_outputs(4468) <= not(inputs(58));
    layer0_outputs(4469) <= not((inputs(175)) xor (inputs(88)));
    layer0_outputs(4470) <= inputs(42);
    layer0_outputs(4471) <= not((inputs(81)) xor (inputs(219)));
    layer0_outputs(4472) <= (inputs(97)) and not (inputs(30));
    layer0_outputs(4473) <= (inputs(119)) and not (inputs(50));
    layer0_outputs(4474) <= '0';
    layer0_outputs(4475) <= not(inputs(93));
    layer0_outputs(4476) <= not(inputs(188));
    layer0_outputs(4477) <= (inputs(9)) xor (inputs(247));
    layer0_outputs(4478) <= not(inputs(155));
    layer0_outputs(4479) <= inputs(167);
    layer0_outputs(4480) <= not(inputs(152));
    layer0_outputs(4481) <= not(inputs(68)) or (inputs(2));
    layer0_outputs(4482) <= (inputs(106)) or (inputs(67));
    layer0_outputs(4483) <= not((inputs(153)) or (inputs(250)));
    layer0_outputs(4484) <= inputs(64);
    layer0_outputs(4485) <= (inputs(72)) and not (inputs(181));
    layer0_outputs(4486) <= (inputs(121)) or (inputs(102));
    layer0_outputs(4487) <= (inputs(158)) and not (inputs(189));
    layer0_outputs(4488) <= not((inputs(181)) xor (inputs(227)));
    layer0_outputs(4489) <= inputs(7);
    layer0_outputs(4490) <= not((inputs(119)) or (inputs(181)));
    layer0_outputs(4491) <= not(inputs(115));
    layer0_outputs(4492) <= (inputs(200)) or (inputs(128));
    layer0_outputs(4493) <= (inputs(24)) or (inputs(80));
    layer0_outputs(4494) <= not(inputs(40));
    layer0_outputs(4495) <= not(inputs(93)) or (inputs(33));
    layer0_outputs(4496) <= inputs(30);
    layer0_outputs(4497) <= inputs(198);
    layer0_outputs(4498) <= (inputs(98)) or (inputs(189));
    layer0_outputs(4499) <= (inputs(163)) or (inputs(141));
    layer0_outputs(4500) <= not(inputs(132)) or (inputs(64));
    layer0_outputs(4501) <= not(inputs(198)) or (inputs(39));
    layer0_outputs(4502) <= (inputs(79)) and not (inputs(118));
    layer0_outputs(4503) <= (inputs(120)) and not (inputs(196));
    layer0_outputs(4504) <= not((inputs(239)) xor (inputs(90)));
    layer0_outputs(4505) <= not((inputs(124)) xor (inputs(86)));
    layer0_outputs(4506) <= not((inputs(67)) xor (inputs(104)));
    layer0_outputs(4507) <= inputs(60);
    layer0_outputs(4508) <= not(inputs(185)) or (inputs(174));
    layer0_outputs(4509) <= not((inputs(25)) or (inputs(25)));
    layer0_outputs(4510) <= not((inputs(87)) xor (inputs(206)));
    layer0_outputs(4511) <= not((inputs(5)) or (inputs(31)));
    layer0_outputs(4512) <= not(inputs(113)) or (inputs(87));
    layer0_outputs(4513) <= not((inputs(224)) xor (inputs(33)));
    layer0_outputs(4514) <= not(inputs(73));
    layer0_outputs(4515) <= not(inputs(179));
    layer0_outputs(4516) <= inputs(193);
    layer0_outputs(4517) <= not((inputs(62)) xor (inputs(205)));
    layer0_outputs(4518) <= (inputs(73)) and not (inputs(185));
    layer0_outputs(4519) <= '0';
    layer0_outputs(4520) <= (inputs(36)) or (inputs(55));
    layer0_outputs(4521) <= (inputs(135)) and not (inputs(43));
    layer0_outputs(4522) <= not((inputs(125)) or (inputs(168)));
    layer0_outputs(4523) <= not(inputs(17));
    layer0_outputs(4524) <= (inputs(67)) and not (inputs(236));
    layer0_outputs(4525) <= (inputs(167)) xor (inputs(178));
    layer0_outputs(4526) <= inputs(110);
    layer0_outputs(4527) <= not(inputs(136));
    layer0_outputs(4528) <= (inputs(97)) and not (inputs(112));
    layer0_outputs(4529) <= not((inputs(114)) or (inputs(2)));
    layer0_outputs(4530) <= not(inputs(35));
    layer0_outputs(4531) <= inputs(141);
    layer0_outputs(4532) <= (inputs(199)) or (inputs(151));
    layer0_outputs(4533) <= '1';
    layer0_outputs(4534) <= (inputs(197)) xor (inputs(81));
    layer0_outputs(4535) <= not((inputs(95)) xor (inputs(242)));
    layer0_outputs(4536) <= not(inputs(82)) or (inputs(158));
    layer0_outputs(4537) <= (inputs(204)) xor (inputs(95));
    layer0_outputs(4538) <= not((inputs(168)) or (inputs(65)));
    layer0_outputs(4539) <= (inputs(197)) and not (inputs(111));
    layer0_outputs(4540) <= not((inputs(33)) or (inputs(209)));
    layer0_outputs(4541) <= '0';
    layer0_outputs(4542) <= (inputs(144)) and not (inputs(11));
    layer0_outputs(4543) <= not(inputs(108));
    layer0_outputs(4544) <= inputs(13);
    layer0_outputs(4545) <= (inputs(249)) and not (inputs(19));
    layer0_outputs(4546) <= (inputs(237)) or (inputs(248));
    layer0_outputs(4547) <= not((inputs(218)) xor (inputs(132)));
    layer0_outputs(4548) <= not(inputs(98)) or (inputs(134));
    layer0_outputs(4549) <= (inputs(215)) or (inputs(142));
    layer0_outputs(4550) <= not((inputs(13)) xor (inputs(192)));
    layer0_outputs(4551) <= (inputs(179)) and not (inputs(29));
    layer0_outputs(4552) <= (inputs(18)) or (inputs(187));
    layer0_outputs(4553) <= not(inputs(158));
    layer0_outputs(4554) <= (inputs(139)) or (inputs(44));
    layer0_outputs(4555) <= not(inputs(143)) or (inputs(205));
    layer0_outputs(4556) <= not(inputs(188));
    layer0_outputs(4557) <= (inputs(50)) or (inputs(51));
    layer0_outputs(4558) <= not(inputs(233));
    layer0_outputs(4559) <= (inputs(165)) and not (inputs(214));
    layer0_outputs(4560) <= (inputs(249)) and not (inputs(253));
    layer0_outputs(4561) <= not((inputs(232)) xor (inputs(95)));
    layer0_outputs(4562) <= (inputs(74)) and not (inputs(194));
    layer0_outputs(4563) <= not(inputs(119));
    layer0_outputs(4564) <= not(inputs(56));
    layer0_outputs(4565) <= (inputs(113)) xor (inputs(83));
    layer0_outputs(4566) <= '0';
    layer0_outputs(4567) <= inputs(101);
    layer0_outputs(4568) <= (inputs(235)) or (inputs(249));
    layer0_outputs(4569) <= (inputs(30)) or (inputs(17));
    layer0_outputs(4570) <= (inputs(118)) or (inputs(220));
    layer0_outputs(4571) <= inputs(146);
    layer0_outputs(4572) <= not((inputs(64)) or (inputs(194)));
    layer0_outputs(4573) <= (inputs(183)) or (inputs(118));
    layer0_outputs(4574) <= (inputs(25)) and not (inputs(198));
    layer0_outputs(4575) <= inputs(179);
    layer0_outputs(4576) <= '0';
    layer0_outputs(4577) <= not((inputs(6)) xor (inputs(221)));
    layer0_outputs(4578) <= not((inputs(241)) or (inputs(9)));
    layer0_outputs(4579) <= (inputs(149)) and not (inputs(141));
    layer0_outputs(4580) <= (inputs(227)) xor (inputs(153));
    layer0_outputs(4581) <= not((inputs(12)) xor (inputs(208)));
    layer0_outputs(4582) <= (inputs(159)) or (inputs(223));
    layer0_outputs(4583) <= (inputs(141)) or (inputs(132));
    layer0_outputs(4584) <= not((inputs(72)) or (inputs(32)));
    layer0_outputs(4585) <= (inputs(91)) and not (inputs(96));
    layer0_outputs(4586) <= (inputs(49)) or (inputs(32));
    layer0_outputs(4587) <= (inputs(224)) or (inputs(7));
    layer0_outputs(4588) <= '1';
    layer0_outputs(4589) <= not(inputs(177)) or (inputs(113));
    layer0_outputs(4590) <= not(inputs(242)) or (inputs(178));
    layer0_outputs(4591) <= inputs(113);
    layer0_outputs(4592) <= (inputs(208)) xor (inputs(96));
    layer0_outputs(4593) <= inputs(247);
    layer0_outputs(4594) <= inputs(215);
    layer0_outputs(4595) <= not(inputs(61));
    layer0_outputs(4596) <= (inputs(247)) and not (inputs(139));
    layer0_outputs(4597) <= not(inputs(243));
    layer0_outputs(4598) <= not((inputs(86)) xor (inputs(0)));
    layer0_outputs(4599) <= not(inputs(125));
    layer0_outputs(4600) <= '1';
    layer0_outputs(4601) <= (inputs(48)) xor (inputs(211));
    layer0_outputs(4602) <= not(inputs(70));
    layer0_outputs(4603) <= not((inputs(96)) xor (inputs(68)));
    layer0_outputs(4604) <= not(inputs(110));
    layer0_outputs(4605) <= not((inputs(132)) xor (inputs(161)));
    layer0_outputs(4606) <= not(inputs(120));
    layer0_outputs(4607) <= (inputs(131)) and not (inputs(205));
    layer0_outputs(4608) <= (inputs(176)) and not (inputs(78));
    layer0_outputs(4609) <= (inputs(203)) xor (inputs(96));
    layer0_outputs(4610) <= not(inputs(77));
    layer0_outputs(4611) <= inputs(76);
    layer0_outputs(4612) <= not(inputs(210)) or (inputs(203));
    layer0_outputs(4613) <= inputs(74);
    layer0_outputs(4614) <= not((inputs(108)) or (inputs(32)));
    layer0_outputs(4615) <= not((inputs(20)) xor (inputs(240)));
    layer0_outputs(4616) <= not(inputs(231));
    layer0_outputs(4617) <= inputs(67);
    layer0_outputs(4618) <= not((inputs(228)) xor (inputs(222)));
    layer0_outputs(4619) <= (inputs(154)) or (inputs(98));
    layer0_outputs(4620) <= not((inputs(68)) or (inputs(197)));
    layer0_outputs(4621) <= '0';
    layer0_outputs(4622) <= (inputs(254)) and not (inputs(46));
    layer0_outputs(4623) <= not(inputs(155)) or (inputs(63));
    layer0_outputs(4624) <= not(inputs(225)) or (inputs(14));
    layer0_outputs(4625) <= (inputs(236)) or (inputs(208));
    layer0_outputs(4626) <= not((inputs(144)) xor (inputs(152)));
    layer0_outputs(4627) <= (inputs(251)) and not (inputs(2));
    layer0_outputs(4628) <= not((inputs(91)) xor (inputs(115)));
    layer0_outputs(4629) <= (inputs(104)) and not (inputs(179));
    layer0_outputs(4630) <= (inputs(237)) or (inputs(243));
    layer0_outputs(4631) <= not((inputs(124)) xor (inputs(138)));
    layer0_outputs(4632) <= inputs(101);
    layer0_outputs(4633) <= not((inputs(86)) or (inputs(225)));
    layer0_outputs(4634) <= not(inputs(235)) or (inputs(53));
    layer0_outputs(4635) <= (inputs(118)) or (inputs(235));
    layer0_outputs(4636) <= not(inputs(40));
    layer0_outputs(4637) <= inputs(97);
    layer0_outputs(4638) <= inputs(229);
    layer0_outputs(4639) <= inputs(78);
    layer0_outputs(4640) <= not(inputs(131)) or (inputs(48));
    layer0_outputs(4641) <= not((inputs(103)) or (inputs(226)));
    layer0_outputs(4642) <= inputs(27);
    layer0_outputs(4643) <= inputs(215);
    layer0_outputs(4644) <= (inputs(224)) xor (inputs(216));
    layer0_outputs(4645) <= not(inputs(231));
    layer0_outputs(4646) <= not((inputs(207)) and (inputs(207)));
    layer0_outputs(4647) <= '1';
    layer0_outputs(4648) <= (inputs(224)) xor (inputs(247));
    layer0_outputs(4649) <= (inputs(220)) or (inputs(160));
    layer0_outputs(4650) <= inputs(219);
    layer0_outputs(4651) <= inputs(238);
    layer0_outputs(4652) <= (inputs(178)) and not (inputs(92));
    layer0_outputs(4653) <= (inputs(53)) and not (inputs(175));
    layer0_outputs(4654) <= '0';
    layer0_outputs(4655) <= inputs(163);
    layer0_outputs(4656) <= not(inputs(202));
    layer0_outputs(4657) <= not((inputs(96)) or (inputs(216)));
    layer0_outputs(4658) <= not((inputs(116)) or (inputs(20)));
    layer0_outputs(4659) <= not(inputs(99)) or (inputs(2));
    layer0_outputs(4660) <= (inputs(210)) xor (inputs(218));
    layer0_outputs(4661) <= not(inputs(107)) or (inputs(62));
    layer0_outputs(4662) <= '1';
    layer0_outputs(4663) <= (inputs(113)) or (inputs(196));
    layer0_outputs(4664) <= (inputs(168)) or (inputs(239));
    layer0_outputs(4665) <= not((inputs(141)) xor (inputs(235)));
    layer0_outputs(4666) <= not(inputs(29));
    layer0_outputs(4667) <= inputs(78);
    layer0_outputs(4668) <= (inputs(150)) xor (inputs(168));
    layer0_outputs(4669) <= not(inputs(22));
    layer0_outputs(4670) <= inputs(141);
    layer0_outputs(4671) <= inputs(232);
    layer0_outputs(4672) <= inputs(198);
    layer0_outputs(4673) <= not(inputs(172));
    layer0_outputs(4674) <= (inputs(105)) and not (inputs(196));
    layer0_outputs(4675) <= not(inputs(26));
    layer0_outputs(4676) <= not((inputs(24)) or (inputs(230)));
    layer0_outputs(4677) <= (inputs(156)) xor (inputs(136));
    layer0_outputs(4678) <= (inputs(54)) and (inputs(57));
    layer0_outputs(4679) <= not(inputs(92)) or (inputs(105));
    layer0_outputs(4680) <= not((inputs(75)) and (inputs(154)));
    layer0_outputs(4681) <= (inputs(194)) or (inputs(213));
    layer0_outputs(4682) <= not((inputs(96)) or (inputs(217)));
    layer0_outputs(4683) <= not(inputs(79));
    layer0_outputs(4684) <= not(inputs(231)) or (inputs(240));
    layer0_outputs(4685) <= (inputs(208)) and (inputs(169));
    layer0_outputs(4686) <= not((inputs(131)) or (inputs(9)));
    layer0_outputs(4687) <= (inputs(133)) and not (inputs(111));
    layer0_outputs(4688) <= (inputs(86)) xor (inputs(133));
    layer0_outputs(4689) <= not(inputs(146));
    layer0_outputs(4690) <= (inputs(198)) and not (inputs(206));
    layer0_outputs(4691) <= (inputs(221)) and not (inputs(249));
    layer0_outputs(4692) <= not((inputs(254)) or (inputs(103)));
    layer0_outputs(4693) <= not(inputs(111));
    layer0_outputs(4694) <= (inputs(217)) or (inputs(235));
    layer0_outputs(4695) <= not((inputs(253)) xor (inputs(43)));
    layer0_outputs(4696) <= (inputs(192)) xor (inputs(145));
    layer0_outputs(4697) <= (inputs(134)) or (inputs(97));
    layer0_outputs(4698) <= (inputs(153)) xor (inputs(139));
    layer0_outputs(4699) <= (inputs(225)) or (inputs(108));
    layer0_outputs(4700) <= inputs(76);
    layer0_outputs(4701) <= (inputs(255)) xor (inputs(137));
    layer0_outputs(4702) <= inputs(217);
    layer0_outputs(4703) <= not(inputs(48)) or (inputs(150));
    layer0_outputs(4704) <= not((inputs(141)) or (inputs(43)));
    layer0_outputs(4705) <= not(inputs(93));
    layer0_outputs(4706) <= '1';
    layer0_outputs(4707) <= inputs(164);
    layer0_outputs(4708) <= not((inputs(114)) xor (inputs(160)));
    layer0_outputs(4709) <= inputs(28);
    layer0_outputs(4710) <= inputs(24);
    layer0_outputs(4711) <= not(inputs(196)) or (inputs(16));
    layer0_outputs(4712) <= (inputs(26)) and not (inputs(129));
    layer0_outputs(4713) <= not((inputs(219)) or (inputs(92)));
    layer0_outputs(4714) <= not(inputs(60));
    layer0_outputs(4715) <= not((inputs(62)) or (inputs(168)));
    layer0_outputs(4716) <= not((inputs(195)) xor (inputs(37)));
    layer0_outputs(4717) <= (inputs(252)) and not (inputs(191));
    layer0_outputs(4718) <= not(inputs(248));
    layer0_outputs(4719) <= (inputs(20)) and not (inputs(157));
    layer0_outputs(4720) <= (inputs(39)) and not (inputs(10));
    layer0_outputs(4721) <= not(inputs(134)) or (inputs(107));
    layer0_outputs(4722) <= not(inputs(248)) or (inputs(3));
    layer0_outputs(4723) <= not((inputs(251)) or (inputs(199)));
    layer0_outputs(4724) <= not((inputs(35)) xor (inputs(95)));
    layer0_outputs(4725) <= not((inputs(226)) or (inputs(50)));
    layer0_outputs(4726) <= not(inputs(135));
    layer0_outputs(4727) <= not(inputs(107)) or (inputs(6));
    layer0_outputs(4728) <= not(inputs(231)) or (inputs(165));
    layer0_outputs(4729) <= inputs(113);
    layer0_outputs(4730) <= inputs(74);
    layer0_outputs(4731) <= (inputs(213)) and not (inputs(66));
    layer0_outputs(4732) <= not((inputs(255)) or (inputs(8)));
    layer0_outputs(4733) <= not(inputs(95));
    layer0_outputs(4734) <= inputs(135);
    layer0_outputs(4735) <= '1';
    layer0_outputs(4736) <= inputs(41);
    layer0_outputs(4737) <= not(inputs(10));
    layer0_outputs(4738) <= not(inputs(130));
    layer0_outputs(4739) <= not(inputs(205));
    layer0_outputs(4740) <= (inputs(246)) or (inputs(155));
    layer0_outputs(4741) <= not(inputs(39));
    layer0_outputs(4742) <= (inputs(8)) and not (inputs(233));
    layer0_outputs(4743) <= inputs(83);
    layer0_outputs(4744) <= not(inputs(254));
    layer0_outputs(4745) <= not((inputs(91)) or (inputs(207)));
    layer0_outputs(4746) <= not(inputs(117));
    layer0_outputs(4747) <= (inputs(145)) or (inputs(77));
    layer0_outputs(4748) <= not(inputs(2)) or (inputs(168));
    layer0_outputs(4749) <= not((inputs(226)) xor (inputs(166)));
    layer0_outputs(4750) <= (inputs(98)) or (inputs(69));
    layer0_outputs(4751) <= (inputs(37)) xor (inputs(200));
    layer0_outputs(4752) <= not(inputs(35));
    layer0_outputs(4753) <= '1';
    layer0_outputs(4754) <= (inputs(91)) and not (inputs(79));
    layer0_outputs(4755) <= not((inputs(14)) xor (inputs(143)));
    layer0_outputs(4756) <= inputs(228);
    layer0_outputs(4757) <= (inputs(141)) and not (inputs(152));
    layer0_outputs(4758) <= (inputs(203)) and not (inputs(46));
    layer0_outputs(4759) <= (inputs(84)) and not (inputs(4));
    layer0_outputs(4760) <= not(inputs(244));
    layer0_outputs(4761) <= (inputs(208)) and not (inputs(200));
    layer0_outputs(4762) <= not(inputs(249));
    layer0_outputs(4763) <= not(inputs(239));
    layer0_outputs(4764) <= inputs(118);
    layer0_outputs(4765) <= (inputs(183)) and not (inputs(128));
    layer0_outputs(4766) <= not((inputs(180)) xor (inputs(128)));
    layer0_outputs(4767) <= (inputs(100)) xor (inputs(73));
    layer0_outputs(4768) <= not(inputs(135));
    layer0_outputs(4769) <= not(inputs(200));
    layer0_outputs(4770) <= (inputs(237)) and (inputs(17));
    layer0_outputs(4771) <= not(inputs(92));
    layer0_outputs(4772) <= (inputs(185)) and not (inputs(16));
    layer0_outputs(4773) <= not((inputs(69)) xor (inputs(5)));
    layer0_outputs(4774) <= not((inputs(178)) and (inputs(205)));
    layer0_outputs(4775) <= (inputs(38)) and not (inputs(213));
    layer0_outputs(4776) <= (inputs(64)) or (inputs(146));
    layer0_outputs(4777) <= inputs(252);
    layer0_outputs(4778) <= (inputs(126)) or (inputs(35));
    layer0_outputs(4779) <= not(inputs(243));
    layer0_outputs(4780) <= not(inputs(84)) or (inputs(9));
    layer0_outputs(4781) <= not(inputs(181)) or (inputs(78));
    layer0_outputs(4782) <= (inputs(19)) and not (inputs(100));
    layer0_outputs(4783) <= not(inputs(69)) or (inputs(253));
    layer0_outputs(4784) <= not(inputs(210)) or (inputs(212));
    layer0_outputs(4785) <= inputs(59);
    layer0_outputs(4786) <= (inputs(82)) or (inputs(50));
    layer0_outputs(4787) <= inputs(113);
    layer0_outputs(4788) <= inputs(98);
    layer0_outputs(4789) <= not(inputs(139));
    layer0_outputs(4790) <= (inputs(99)) and (inputs(3));
    layer0_outputs(4791) <= inputs(122);
    layer0_outputs(4792) <= not((inputs(23)) xor (inputs(60)));
    layer0_outputs(4793) <= (inputs(9)) or (inputs(206));
    layer0_outputs(4794) <= inputs(22);
    layer0_outputs(4795) <= (inputs(244)) and not (inputs(67));
    layer0_outputs(4796) <= not((inputs(233)) xor (inputs(17)));
    layer0_outputs(4797) <= not(inputs(53));
    layer0_outputs(4798) <= not((inputs(7)) or (inputs(100)));
    layer0_outputs(4799) <= not((inputs(10)) and (inputs(108)));
    layer0_outputs(4800) <= inputs(164);
    layer0_outputs(4801) <= (inputs(216)) and not (inputs(49));
    layer0_outputs(4802) <= not(inputs(92));
    layer0_outputs(4803) <= inputs(111);
    layer0_outputs(4804) <= inputs(52);
    layer0_outputs(4805) <= not((inputs(147)) xor (inputs(169)));
    layer0_outputs(4806) <= (inputs(174)) or (inputs(154));
    layer0_outputs(4807) <= (inputs(101)) or (inputs(146));
    layer0_outputs(4808) <= inputs(154);
    layer0_outputs(4809) <= not((inputs(127)) or (inputs(127)));
    layer0_outputs(4810) <= not(inputs(43)) or (inputs(160));
    layer0_outputs(4811) <= not((inputs(146)) or (inputs(66)));
    layer0_outputs(4812) <= not((inputs(219)) xor (inputs(107)));
    layer0_outputs(4813) <= (inputs(7)) and not (inputs(112));
    layer0_outputs(4814) <= not(inputs(177));
    layer0_outputs(4815) <= not(inputs(26));
    layer0_outputs(4816) <= not(inputs(19)) or (inputs(220));
    layer0_outputs(4817) <= inputs(148);
    layer0_outputs(4818) <= not((inputs(162)) or (inputs(234)));
    layer0_outputs(4819) <= (inputs(36)) and not (inputs(140));
    layer0_outputs(4820) <= not(inputs(9)) or (inputs(15));
    layer0_outputs(4821) <= inputs(82);
    layer0_outputs(4822) <= not((inputs(110)) or (inputs(41)));
    layer0_outputs(4823) <= (inputs(85)) xor (inputs(56));
    layer0_outputs(4824) <= not((inputs(27)) xor (inputs(37)));
    layer0_outputs(4825) <= not((inputs(213)) or (inputs(44)));
    layer0_outputs(4826) <= inputs(85);
    layer0_outputs(4827) <= not(inputs(189));
    layer0_outputs(4828) <= (inputs(143)) or (inputs(52));
    layer0_outputs(4829) <= not(inputs(114));
    layer0_outputs(4830) <= (inputs(128)) xor (inputs(76));
    layer0_outputs(4831) <= not(inputs(238)) or (inputs(251));
    layer0_outputs(4832) <= inputs(166);
    layer0_outputs(4833) <= not((inputs(94)) or (inputs(255)));
    layer0_outputs(4834) <= (inputs(204)) and not (inputs(139));
    layer0_outputs(4835) <= not((inputs(212)) or (inputs(41)));
    layer0_outputs(4836) <= (inputs(231)) and not (inputs(46));
    layer0_outputs(4837) <= (inputs(178)) and not (inputs(122));
    layer0_outputs(4838) <= (inputs(160)) and (inputs(135));
    layer0_outputs(4839) <= (inputs(102)) and not (inputs(79));
    layer0_outputs(4840) <= (inputs(201)) or (inputs(157));
    layer0_outputs(4841) <= not((inputs(216)) or (inputs(211)));
    layer0_outputs(4842) <= not((inputs(200)) xor (inputs(31)));
    layer0_outputs(4843) <= (inputs(41)) and (inputs(159));
    layer0_outputs(4844) <= (inputs(88)) xor (inputs(171));
    layer0_outputs(4845) <= (inputs(254)) or (inputs(86));
    layer0_outputs(4846) <= not((inputs(75)) or (inputs(224)));
    layer0_outputs(4847) <= not(inputs(193));
    layer0_outputs(4848) <= (inputs(141)) or (inputs(85));
    layer0_outputs(4849) <= not(inputs(141));
    layer0_outputs(4850) <= not(inputs(246)) or (inputs(131));
    layer0_outputs(4851) <= (inputs(130)) or (inputs(75));
    layer0_outputs(4852) <= not((inputs(189)) xor (inputs(229)));
    layer0_outputs(4853) <= (inputs(201)) or (inputs(132));
    layer0_outputs(4854) <= not((inputs(88)) or (inputs(186)));
    layer0_outputs(4855) <= (inputs(93)) xor (inputs(159));
    layer0_outputs(4856) <= not((inputs(205)) or (inputs(128)));
    layer0_outputs(4857) <= not(inputs(222)) or (inputs(195));
    layer0_outputs(4858) <= (inputs(56)) and (inputs(201));
    layer0_outputs(4859) <= (inputs(179)) and (inputs(170));
    layer0_outputs(4860) <= (inputs(188)) or (inputs(173));
    layer0_outputs(4861) <= inputs(97);
    layer0_outputs(4862) <= not(inputs(170));
    layer0_outputs(4863) <= not(inputs(109));
    layer0_outputs(4864) <= inputs(74);
    layer0_outputs(4865) <= not(inputs(11)) or (inputs(224));
    layer0_outputs(4866) <= not((inputs(161)) or (inputs(40)));
    layer0_outputs(4867) <= not((inputs(20)) xor (inputs(26)));
    layer0_outputs(4868) <= not(inputs(190)) or (inputs(184));
    layer0_outputs(4869) <= (inputs(79)) or (inputs(156));
    layer0_outputs(4870) <= (inputs(219)) and not (inputs(86));
    layer0_outputs(4871) <= not(inputs(135)) or (inputs(138));
    layer0_outputs(4872) <= (inputs(139)) xor (inputs(91));
    layer0_outputs(4873) <= (inputs(160)) or (inputs(175));
    layer0_outputs(4874) <= not((inputs(105)) and (inputs(168)));
    layer0_outputs(4875) <= '1';
    layer0_outputs(4876) <= (inputs(21)) or (inputs(150));
    layer0_outputs(4877) <= (inputs(67)) or (inputs(94));
    layer0_outputs(4878) <= not((inputs(117)) or (inputs(116)));
    layer0_outputs(4879) <= not(inputs(110)) or (inputs(33));
    layer0_outputs(4880) <= '1';
    layer0_outputs(4881) <= (inputs(203)) and not (inputs(47));
    layer0_outputs(4882) <= inputs(135);
    layer0_outputs(4883) <= (inputs(10)) or (inputs(168));
    layer0_outputs(4884) <= not((inputs(252)) or (inputs(96)));
    layer0_outputs(4885) <= (inputs(11)) xor (inputs(45));
    layer0_outputs(4886) <= not((inputs(68)) xor (inputs(173)));
    layer0_outputs(4887) <= (inputs(57)) and not (inputs(232));
    layer0_outputs(4888) <= (inputs(119)) or (inputs(122));
    layer0_outputs(4889) <= not(inputs(126));
    layer0_outputs(4890) <= inputs(221);
    layer0_outputs(4891) <= not(inputs(68));
    layer0_outputs(4892) <= (inputs(50)) or (inputs(180));
    layer0_outputs(4893) <= not((inputs(65)) xor (inputs(22)));
    layer0_outputs(4894) <= not(inputs(10));
    layer0_outputs(4895) <= (inputs(1)) or (inputs(109));
    layer0_outputs(4896) <= (inputs(54)) and not (inputs(16));
    layer0_outputs(4897) <= (inputs(71)) and not (inputs(0));
    layer0_outputs(4898) <= not(inputs(135));
    layer0_outputs(4899) <= not(inputs(120));
    layer0_outputs(4900) <= inputs(212);
    layer0_outputs(4901) <= not(inputs(84)) or (inputs(162));
    layer0_outputs(4902) <= (inputs(164)) xor (inputs(240));
    layer0_outputs(4903) <= not((inputs(147)) or (inputs(175)));
    layer0_outputs(4904) <= (inputs(1)) or (inputs(13));
    layer0_outputs(4905) <= inputs(56);
    layer0_outputs(4906) <= not(inputs(69)) or (inputs(128));
    layer0_outputs(4907) <= not((inputs(149)) xor (inputs(117)));
    layer0_outputs(4908) <= not((inputs(249)) or (inputs(245)));
    layer0_outputs(4909) <= not(inputs(195)) or (inputs(254));
    layer0_outputs(4910) <= not(inputs(191)) or (inputs(145));
    layer0_outputs(4911) <= not((inputs(213)) and (inputs(226)));
    layer0_outputs(4912) <= not(inputs(76));
    layer0_outputs(4913) <= not(inputs(132)) or (inputs(4));
    layer0_outputs(4914) <= (inputs(174)) or (inputs(24));
    layer0_outputs(4915) <= not(inputs(134)) or (inputs(96));
    layer0_outputs(4916) <= (inputs(1)) xor (inputs(25));
    layer0_outputs(4917) <= inputs(9);
    layer0_outputs(4918) <= '0';
    layer0_outputs(4919) <= inputs(230);
    layer0_outputs(4920) <= (inputs(28)) and not (inputs(174));
    layer0_outputs(4921) <= (inputs(103)) or (inputs(132));
    layer0_outputs(4922) <= (inputs(226)) and not (inputs(252));
    layer0_outputs(4923) <= (inputs(27)) xor (inputs(44));
    layer0_outputs(4924) <= (inputs(151)) and not (inputs(223));
    layer0_outputs(4925) <= not((inputs(56)) and (inputs(43)));
    layer0_outputs(4926) <= not((inputs(11)) and (inputs(19)));
    layer0_outputs(4927) <= not(inputs(191)) or (inputs(69));
    layer0_outputs(4928) <= inputs(34);
    layer0_outputs(4929) <= (inputs(76)) and not (inputs(0));
    layer0_outputs(4930) <= '0';
    layer0_outputs(4931) <= (inputs(100)) and not (inputs(235));
    layer0_outputs(4932) <= not(inputs(151));
    layer0_outputs(4933) <= not((inputs(59)) xor (inputs(58)));
    layer0_outputs(4934) <= not((inputs(45)) or (inputs(4)));
    layer0_outputs(4935) <= not((inputs(60)) and (inputs(1)));
    layer0_outputs(4936) <= not(inputs(120)) or (inputs(1));
    layer0_outputs(4937) <= (inputs(139)) or (inputs(85));
    layer0_outputs(4938) <= (inputs(90)) and not (inputs(194));
    layer0_outputs(4939) <= (inputs(16)) or (inputs(26));
    layer0_outputs(4940) <= not(inputs(55)) or (inputs(101));
    layer0_outputs(4941) <= not((inputs(79)) or (inputs(225)));
    layer0_outputs(4942) <= (inputs(247)) and not (inputs(44));
    layer0_outputs(4943) <= (inputs(128)) or (inputs(84));
    layer0_outputs(4944) <= not(inputs(2)) or (inputs(175));
    layer0_outputs(4945) <= inputs(10);
    layer0_outputs(4946) <= (inputs(230)) or (inputs(15));
    layer0_outputs(4947) <= inputs(80);
    layer0_outputs(4948) <= (inputs(114)) or (inputs(145));
    layer0_outputs(4949) <= inputs(169);
    layer0_outputs(4950) <= (inputs(0)) xor (inputs(84));
    layer0_outputs(4951) <= (inputs(119)) or (inputs(173));
    layer0_outputs(4952) <= (inputs(226)) xor (inputs(176));
    layer0_outputs(4953) <= not((inputs(197)) xor (inputs(139)));
    layer0_outputs(4954) <= not(inputs(100));
    layer0_outputs(4955) <= not((inputs(180)) or (inputs(227)));
    layer0_outputs(4956) <= inputs(82);
    layer0_outputs(4957) <= inputs(21);
    layer0_outputs(4958) <= not((inputs(21)) or (inputs(32)));
    layer0_outputs(4959) <= not(inputs(243)) or (inputs(245));
    layer0_outputs(4960) <= (inputs(7)) or (inputs(49));
    layer0_outputs(4961) <= (inputs(172)) and not (inputs(168));
    layer0_outputs(4962) <= not((inputs(1)) or (inputs(153)));
    layer0_outputs(4963) <= not(inputs(147)) or (inputs(21));
    layer0_outputs(4964) <= not((inputs(177)) or (inputs(17)));
    layer0_outputs(4965) <= inputs(96);
    layer0_outputs(4966) <= not((inputs(32)) or (inputs(19)));
    layer0_outputs(4967) <= inputs(129);
    layer0_outputs(4968) <= not((inputs(186)) xor (inputs(218)));
    layer0_outputs(4969) <= (inputs(245)) xor (inputs(227));
    layer0_outputs(4970) <= not((inputs(32)) xor (inputs(33)));
    layer0_outputs(4971) <= not(inputs(248));
    layer0_outputs(4972) <= (inputs(180)) or (inputs(130));
    layer0_outputs(4973) <= (inputs(121)) and not (inputs(166));
    layer0_outputs(4974) <= (inputs(85)) xor (inputs(112));
    layer0_outputs(4975) <= (inputs(43)) and not (inputs(238));
    layer0_outputs(4976) <= inputs(183);
    layer0_outputs(4977) <= not(inputs(21));
    layer0_outputs(4978) <= (inputs(84)) and not (inputs(25));
    layer0_outputs(4979) <= (inputs(149)) or (inputs(231));
    layer0_outputs(4980) <= (inputs(104)) or (inputs(206));
    layer0_outputs(4981) <= inputs(90);
    layer0_outputs(4982) <= (inputs(49)) xor (inputs(162));
    layer0_outputs(4983) <= not((inputs(119)) and (inputs(164)));
    layer0_outputs(4984) <= not(inputs(83));
    layer0_outputs(4985) <= not(inputs(175));
    layer0_outputs(4986) <= '1';
    layer0_outputs(4987) <= not(inputs(146));
    layer0_outputs(4988) <= not(inputs(201)) or (inputs(168));
    layer0_outputs(4989) <= not(inputs(67));
    layer0_outputs(4990) <= (inputs(98)) or (inputs(226));
    layer0_outputs(4991) <= not(inputs(152));
    layer0_outputs(4992) <= not(inputs(248));
    layer0_outputs(4993) <= inputs(4);
    layer0_outputs(4994) <= not((inputs(243)) or (inputs(233)));
    layer0_outputs(4995) <= inputs(13);
    layer0_outputs(4996) <= inputs(125);
    layer0_outputs(4997) <= not(inputs(231));
    layer0_outputs(4998) <= not(inputs(73)) or (inputs(17));
    layer0_outputs(4999) <= (inputs(50)) xor (inputs(6));
    layer0_outputs(5000) <= (inputs(164)) or (inputs(255));
    layer0_outputs(5001) <= inputs(172);
    layer0_outputs(5002) <= not(inputs(116)) or (inputs(254));
    layer0_outputs(5003) <= not((inputs(136)) xor (inputs(151)));
    layer0_outputs(5004) <= (inputs(191)) xor (inputs(147));
    layer0_outputs(5005) <= not(inputs(231)) or (inputs(45));
    layer0_outputs(5006) <= inputs(198);
    layer0_outputs(5007) <= not(inputs(6)) or (inputs(131));
    layer0_outputs(5008) <= not(inputs(34)) or (inputs(167));
    layer0_outputs(5009) <= (inputs(21)) or (inputs(10));
    layer0_outputs(5010) <= not(inputs(202)) or (inputs(69));
    layer0_outputs(5011) <= (inputs(133)) and (inputs(134));
    layer0_outputs(5012) <= not(inputs(250));
    layer0_outputs(5013) <= not(inputs(236)) or (inputs(144));
    layer0_outputs(5014) <= not((inputs(17)) or (inputs(52)));
    layer0_outputs(5015) <= not((inputs(233)) xor (inputs(199)));
    layer0_outputs(5016) <= inputs(23);
    layer0_outputs(5017) <= inputs(180);
    layer0_outputs(5018) <= inputs(249);
    layer0_outputs(5019) <= (inputs(140)) and not (inputs(84));
    layer0_outputs(5020) <= (inputs(166)) and not (inputs(17));
    layer0_outputs(5021) <= not((inputs(47)) or (inputs(195)));
    layer0_outputs(5022) <= (inputs(170)) xor (inputs(123));
    layer0_outputs(5023) <= (inputs(96)) xor (inputs(104));
    layer0_outputs(5024) <= not((inputs(40)) xor (inputs(46)));
    layer0_outputs(5025) <= (inputs(136)) and not (inputs(114));
    layer0_outputs(5026) <= (inputs(83)) xor (inputs(93));
    layer0_outputs(5027) <= not(inputs(178)) or (inputs(103));
    layer0_outputs(5028) <= inputs(153);
    layer0_outputs(5029) <= (inputs(214)) or (inputs(24));
    layer0_outputs(5030) <= (inputs(199)) xor (inputs(6));
    layer0_outputs(5031) <= not(inputs(183)) or (inputs(11));
    layer0_outputs(5032) <= (inputs(71)) or (inputs(6));
    layer0_outputs(5033) <= inputs(1);
    layer0_outputs(5034) <= not((inputs(110)) or (inputs(79)));
    layer0_outputs(5035) <= not(inputs(201)) or (inputs(30));
    layer0_outputs(5036) <= (inputs(70)) xor (inputs(129));
    layer0_outputs(5037) <= (inputs(77)) and (inputs(149));
    layer0_outputs(5038) <= (inputs(129)) xor (inputs(89));
    layer0_outputs(5039) <= not((inputs(3)) or (inputs(75)));
    layer0_outputs(5040) <= not(inputs(145)) or (inputs(28));
    layer0_outputs(5041) <= not((inputs(132)) xor (inputs(204)));
    layer0_outputs(5042) <= inputs(188);
    layer0_outputs(5043) <= not(inputs(60));
    layer0_outputs(5044) <= not((inputs(55)) xor (inputs(116)));
    layer0_outputs(5045) <= '0';
    layer0_outputs(5046) <= inputs(36);
    layer0_outputs(5047) <= not(inputs(145));
    layer0_outputs(5048) <= not((inputs(120)) xor (inputs(91)));
    layer0_outputs(5049) <= inputs(140);
    layer0_outputs(5050) <= (inputs(34)) or (inputs(247));
    layer0_outputs(5051) <= not((inputs(9)) and (inputs(243)));
    layer0_outputs(5052) <= (inputs(192)) and not (inputs(128));
    layer0_outputs(5053) <= (inputs(6)) and not (inputs(6));
    layer0_outputs(5054) <= (inputs(91)) xor (inputs(179));
    layer0_outputs(5055) <= inputs(40);
    layer0_outputs(5056) <= (inputs(140)) or (inputs(164));
    layer0_outputs(5057) <= (inputs(111)) or (inputs(186));
    layer0_outputs(5058) <= (inputs(135)) xor (inputs(196));
    layer0_outputs(5059) <= inputs(151);
    layer0_outputs(5060) <= not(inputs(60)) or (inputs(14));
    layer0_outputs(5061) <= not((inputs(128)) xor (inputs(100)));
    layer0_outputs(5062) <= not(inputs(209));
    layer0_outputs(5063) <= inputs(14);
    layer0_outputs(5064) <= not(inputs(163));
    layer0_outputs(5065) <= not((inputs(113)) or (inputs(121)));
    layer0_outputs(5066) <= inputs(45);
    layer0_outputs(5067) <= not(inputs(83)) or (inputs(164));
    layer0_outputs(5068) <= not(inputs(12)) or (inputs(253));
    layer0_outputs(5069) <= (inputs(205)) xor (inputs(225));
    layer0_outputs(5070) <= (inputs(214)) xor (inputs(191));
    layer0_outputs(5071) <= not((inputs(211)) or (inputs(76)));
    layer0_outputs(5072) <= inputs(136);
    layer0_outputs(5073) <= (inputs(58)) xor (inputs(55));
    layer0_outputs(5074) <= not((inputs(113)) or (inputs(104)));
    layer0_outputs(5075) <= not((inputs(94)) or (inputs(138)));
    layer0_outputs(5076) <= not((inputs(211)) or (inputs(224)));
    layer0_outputs(5077) <= (inputs(45)) xor (inputs(157));
    layer0_outputs(5078) <= (inputs(101)) xor (inputs(136));
    layer0_outputs(5079) <= inputs(103);
    layer0_outputs(5080) <= inputs(134);
    layer0_outputs(5081) <= not(inputs(116));
    layer0_outputs(5082) <= (inputs(233)) and (inputs(81));
    layer0_outputs(5083) <= not((inputs(94)) or (inputs(80)));
    layer0_outputs(5084) <= not(inputs(27));
    layer0_outputs(5085) <= not((inputs(199)) xor (inputs(230)));
    layer0_outputs(5086) <= not((inputs(134)) or (inputs(196)));
    layer0_outputs(5087) <= (inputs(102)) or (inputs(173));
    layer0_outputs(5088) <= not(inputs(166));
    layer0_outputs(5089) <= not((inputs(218)) xor (inputs(22)));
    layer0_outputs(5090) <= '1';
    layer0_outputs(5091) <= (inputs(86)) and not (inputs(223));
    layer0_outputs(5092) <= not(inputs(25));
    layer0_outputs(5093) <= (inputs(74)) and not (inputs(204));
    layer0_outputs(5094) <= inputs(101);
    layer0_outputs(5095) <= not(inputs(219)) or (inputs(34));
    layer0_outputs(5096) <= (inputs(209)) xor (inputs(11));
    layer0_outputs(5097) <= not((inputs(249)) or (inputs(159)));
    layer0_outputs(5098) <= not((inputs(33)) xor (inputs(206)));
    layer0_outputs(5099) <= (inputs(218)) and not (inputs(48));
    layer0_outputs(5100) <= not((inputs(171)) or (inputs(208)));
    layer0_outputs(5101) <= not(inputs(199));
    layer0_outputs(5102) <= not(inputs(183));
    layer0_outputs(5103) <= (inputs(124)) and not (inputs(206));
    layer0_outputs(5104) <= (inputs(218)) and not (inputs(87));
    layer0_outputs(5105) <= (inputs(90)) and not (inputs(16));
    layer0_outputs(5106) <= not(inputs(202));
    layer0_outputs(5107) <= (inputs(138)) and not (inputs(70));
    layer0_outputs(5108) <= not((inputs(140)) or (inputs(156)));
    layer0_outputs(5109) <= not(inputs(87));
    layer0_outputs(5110) <= (inputs(198)) xor (inputs(238));
    layer0_outputs(5111) <= not(inputs(184)) or (inputs(85));
    layer0_outputs(5112) <= not(inputs(233)) or (inputs(239));
    layer0_outputs(5113) <= inputs(114);
    layer0_outputs(5114) <= not((inputs(33)) or (inputs(67)));
    layer0_outputs(5115) <= (inputs(172)) and (inputs(42));
    layer0_outputs(5116) <= not((inputs(82)) xor (inputs(96)));
    layer0_outputs(5117) <= not(inputs(147));
    layer0_outputs(5118) <= (inputs(211)) xor (inputs(243));
    layer0_outputs(5119) <= not((inputs(31)) or (inputs(255)));
    layer0_outputs(5120) <= not(inputs(80)) or (inputs(112));
    layer0_outputs(5121) <= not(inputs(186));
    layer0_outputs(5122) <= not((inputs(33)) or (inputs(220)));
    layer0_outputs(5123) <= (inputs(89)) or (inputs(161));
    layer0_outputs(5124) <= inputs(231);
    layer0_outputs(5125) <= inputs(182);
    layer0_outputs(5126) <= not(inputs(231));
    layer0_outputs(5127) <= not((inputs(168)) xor (inputs(162)));
    layer0_outputs(5128) <= not(inputs(56));
    layer0_outputs(5129) <= (inputs(220)) xor (inputs(174));
    layer0_outputs(5130) <= inputs(246);
    layer0_outputs(5131) <= inputs(244);
    layer0_outputs(5132) <= (inputs(21)) xor (inputs(66));
    layer0_outputs(5133) <= not((inputs(197)) xor (inputs(145)));
    layer0_outputs(5134) <= not(inputs(179));
    layer0_outputs(5135) <= not(inputs(250));
    layer0_outputs(5136) <= not(inputs(218));
    layer0_outputs(5137) <= not(inputs(41));
    layer0_outputs(5138) <= not((inputs(243)) or (inputs(218)));
    layer0_outputs(5139) <= not(inputs(120));
    layer0_outputs(5140) <= (inputs(110)) or (inputs(30));
    layer0_outputs(5141) <= not(inputs(74));
    layer0_outputs(5142) <= not(inputs(207)) or (inputs(198));
    layer0_outputs(5143) <= (inputs(110)) and (inputs(57));
    layer0_outputs(5144) <= (inputs(44)) or (inputs(77));
    layer0_outputs(5145) <= not((inputs(165)) or (inputs(251)));
    layer0_outputs(5146) <= not((inputs(44)) xor (inputs(195)));
    layer0_outputs(5147) <= (inputs(235)) or (inputs(192));
    layer0_outputs(5148) <= not(inputs(209));
    layer0_outputs(5149) <= (inputs(76)) or (inputs(0));
    layer0_outputs(5150) <= not((inputs(85)) and (inputs(151)));
    layer0_outputs(5151) <= (inputs(0)) xor (inputs(235));
    layer0_outputs(5152) <= inputs(214);
    layer0_outputs(5153) <= '1';
    layer0_outputs(5154) <= (inputs(91)) and not (inputs(177));
    layer0_outputs(5155) <= (inputs(191)) or (inputs(194));
    layer0_outputs(5156) <= not((inputs(254)) or (inputs(37)));
    layer0_outputs(5157) <= not((inputs(147)) xor (inputs(81)));
    layer0_outputs(5158) <= inputs(250);
    layer0_outputs(5159) <= not(inputs(114));
    layer0_outputs(5160) <= not(inputs(150));
    layer0_outputs(5161) <= not((inputs(48)) or (inputs(140)));
    layer0_outputs(5162) <= not((inputs(252)) xor (inputs(164)));
    layer0_outputs(5163) <= (inputs(202)) and (inputs(228));
    layer0_outputs(5164) <= not((inputs(155)) xor (inputs(134)));
    layer0_outputs(5165) <= inputs(227);
    layer0_outputs(5166) <= (inputs(243)) xor (inputs(67));
    layer0_outputs(5167) <= not(inputs(58)) or (inputs(50));
    layer0_outputs(5168) <= '0';
    layer0_outputs(5169) <= not(inputs(251)) or (inputs(191));
    layer0_outputs(5170) <= not(inputs(157)) or (inputs(68));
    layer0_outputs(5171) <= not((inputs(79)) xor (inputs(42)));
    layer0_outputs(5172) <= not(inputs(226));
    layer0_outputs(5173) <= not((inputs(167)) or (inputs(44)));
    layer0_outputs(5174) <= not((inputs(227)) xor (inputs(20)));
    layer0_outputs(5175) <= inputs(158);
    layer0_outputs(5176) <= inputs(144);
    layer0_outputs(5177) <= (inputs(31)) xor (inputs(191));
    layer0_outputs(5178) <= not(inputs(245));
    layer0_outputs(5179) <= (inputs(74)) and (inputs(23));
    layer0_outputs(5180) <= not((inputs(234)) xor (inputs(59)));
    layer0_outputs(5181) <= not((inputs(123)) or (inputs(81)));
    layer0_outputs(5182) <= not((inputs(199)) xor (inputs(195)));
    layer0_outputs(5183) <= not((inputs(44)) xor (inputs(91)));
    layer0_outputs(5184) <= (inputs(235)) and not (inputs(47));
    layer0_outputs(5185) <= not((inputs(234)) and (inputs(131)));
    layer0_outputs(5186) <= (inputs(134)) xor (inputs(241));
    layer0_outputs(5187) <= not((inputs(216)) and (inputs(70)));
    layer0_outputs(5188) <= not((inputs(221)) xor (inputs(229)));
    layer0_outputs(5189) <= not(inputs(30));
    layer0_outputs(5190) <= inputs(131);
    layer0_outputs(5191) <= not(inputs(237)) or (inputs(129));
    layer0_outputs(5192) <= inputs(136);
    layer0_outputs(5193) <= (inputs(203)) xor (inputs(170));
    layer0_outputs(5194) <= not(inputs(252)) or (inputs(34));
    layer0_outputs(5195) <= '1';
    layer0_outputs(5196) <= (inputs(244)) and not (inputs(96));
    layer0_outputs(5197) <= not(inputs(76));
    layer0_outputs(5198) <= (inputs(85)) and not (inputs(71));
    layer0_outputs(5199) <= (inputs(237)) or (inputs(239));
    layer0_outputs(5200) <= (inputs(249)) and not (inputs(79));
    layer0_outputs(5201) <= not((inputs(30)) xor (inputs(157)));
    layer0_outputs(5202) <= not(inputs(228));
    layer0_outputs(5203) <= (inputs(84)) xor (inputs(86));
    layer0_outputs(5204) <= (inputs(86)) and (inputs(10));
    layer0_outputs(5205) <= not(inputs(82)) or (inputs(252));
    layer0_outputs(5206) <= (inputs(7)) xor (inputs(89));
    layer0_outputs(5207) <= (inputs(203)) or (inputs(108));
    layer0_outputs(5208) <= not((inputs(114)) xor (inputs(246)));
    layer0_outputs(5209) <= not(inputs(211)) or (inputs(80));
    layer0_outputs(5210) <= not(inputs(177));
    layer0_outputs(5211) <= (inputs(57)) or (inputs(205));
    layer0_outputs(5212) <= not(inputs(202)) or (inputs(191));
    layer0_outputs(5213) <= (inputs(47)) and not (inputs(220));
    layer0_outputs(5214) <= not((inputs(32)) or (inputs(219)));
    layer0_outputs(5215) <= not((inputs(98)) or (inputs(101)));
    layer0_outputs(5216) <= (inputs(134)) xor (inputs(88));
    layer0_outputs(5217) <= (inputs(189)) xor (inputs(193));
    layer0_outputs(5218) <= (inputs(214)) or (inputs(243));
    layer0_outputs(5219) <= not(inputs(164));
    layer0_outputs(5220) <= not(inputs(217)) or (inputs(112));
    layer0_outputs(5221) <= (inputs(68)) or (inputs(197));
    layer0_outputs(5222) <= not(inputs(81)) or (inputs(181));
    layer0_outputs(5223) <= inputs(109);
    layer0_outputs(5224) <= not(inputs(166)) or (inputs(38));
    layer0_outputs(5225) <= not((inputs(242)) and (inputs(175)));
    layer0_outputs(5226) <= (inputs(49)) or (inputs(164));
    layer0_outputs(5227) <= not(inputs(226));
    layer0_outputs(5228) <= not((inputs(40)) xor (inputs(220)));
    layer0_outputs(5229) <= not((inputs(176)) or (inputs(22)));
    layer0_outputs(5230) <= inputs(120);
    layer0_outputs(5231) <= (inputs(89)) and (inputs(7));
    layer0_outputs(5232) <= not((inputs(44)) xor (inputs(101)));
    layer0_outputs(5233) <= inputs(219);
    layer0_outputs(5234) <= not((inputs(229)) and (inputs(179)));
    layer0_outputs(5235) <= inputs(224);
    layer0_outputs(5236) <= not(inputs(139)) or (inputs(33));
    layer0_outputs(5237) <= not(inputs(184)) or (inputs(125));
    layer0_outputs(5238) <= (inputs(124)) or (inputs(43));
    layer0_outputs(5239) <= inputs(195);
    layer0_outputs(5240) <= inputs(136);
    layer0_outputs(5241) <= not(inputs(249));
    layer0_outputs(5242) <= not(inputs(186));
    layer0_outputs(5243) <= not(inputs(46)) or (inputs(141));
    layer0_outputs(5244) <= inputs(178);
    layer0_outputs(5245) <= not(inputs(183)) or (inputs(129));
    layer0_outputs(5246) <= not(inputs(2)) or (inputs(127));
    layer0_outputs(5247) <= (inputs(32)) or (inputs(24));
    layer0_outputs(5248) <= not(inputs(249)) or (inputs(139));
    layer0_outputs(5249) <= inputs(162);
    layer0_outputs(5250) <= not((inputs(6)) and (inputs(24)));
    layer0_outputs(5251) <= (inputs(130)) xor (inputs(20));
    layer0_outputs(5252) <= not(inputs(166)) or (inputs(143));
    layer0_outputs(5253) <= inputs(228);
    layer0_outputs(5254) <= not((inputs(179)) xor (inputs(11)));
    layer0_outputs(5255) <= (inputs(22)) and not (inputs(113));
    layer0_outputs(5256) <= not((inputs(82)) or (inputs(95)));
    layer0_outputs(5257) <= (inputs(72)) xor (inputs(208));
    layer0_outputs(5258) <= (inputs(45)) and not (inputs(166));
    layer0_outputs(5259) <= not((inputs(240)) xor (inputs(8)));
    layer0_outputs(5260) <= (inputs(160)) or (inputs(6));
    layer0_outputs(5261) <= not((inputs(108)) and (inputs(63)));
    layer0_outputs(5262) <= not(inputs(183)) or (inputs(121));
    layer0_outputs(5263) <= inputs(98);
    layer0_outputs(5264) <= not(inputs(205));
    layer0_outputs(5265) <= not((inputs(178)) xor (inputs(198)));
    layer0_outputs(5266) <= (inputs(155)) xor (inputs(3));
    layer0_outputs(5267) <= inputs(61);
    layer0_outputs(5268) <= not(inputs(104)) or (inputs(147));
    layer0_outputs(5269) <= not((inputs(26)) or (inputs(36)));
    layer0_outputs(5270) <= (inputs(162)) or (inputs(70));
    layer0_outputs(5271) <= not(inputs(141));
    layer0_outputs(5272) <= inputs(126);
    layer0_outputs(5273) <= (inputs(11)) xor (inputs(74));
    layer0_outputs(5274) <= not(inputs(61));
    layer0_outputs(5275) <= inputs(8);
    layer0_outputs(5276) <= not(inputs(140));
    layer0_outputs(5277) <= not((inputs(77)) xor (inputs(67)));
    layer0_outputs(5278) <= inputs(122);
    layer0_outputs(5279) <= (inputs(18)) xor (inputs(176));
    layer0_outputs(5280) <= not(inputs(141));
    layer0_outputs(5281) <= (inputs(139)) or (inputs(32));
    layer0_outputs(5282) <= (inputs(140)) xor (inputs(232));
    layer0_outputs(5283) <= not(inputs(19));
    layer0_outputs(5284) <= not(inputs(216)) or (inputs(77));
    layer0_outputs(5285) <= not(inputs(53));
    layer0_outputs(5286) <= not(inputs(137));
    layer0_outputs(5287) <= not((inputs(95)) xor (inputs(30)));
    layer0_outputs(5288) <= not((inputs(207)) or (inputs(247)));
    layer0_outputs(5289) <= not((inputs(185)) xor (inputs(198)));
    layer0_outputs(5290) <= inputs(148);
    layer0_outputs(5291) <= (inputs(211)) or (inputs(232));
    layer0_outputs(5292) <= (inputs(86)) xor (inputs(9));
    layer0_outputs(5293) <= not((inputs(67)) xor (inputs(161)));
    layer0_outputs(5294) <= (inputs(192)) xor (inputs(180));
    layer0_outputs(5295) <= not(inputs(231));
    layer0_outputs(5296) <= '0';
    layer0_outputs(5297) <= (inputs(186)) or (inputs(161));
    layer0_outputs(5298) <= not((inputs(71)) xor (inputs(117)));
    layer0_outputs(5299) <= not(inputs(170));
    layer0_outputs(5300) <= (inputs(95)) or (inputs(69));
    layer0_outputs(5301) <= (inputs(44)) or (inputs(169));
    layer0_outputs(5302) <= not(inputs(180)) or (inputs(34));
    layer0_outputs(5303) <= '0';
    layer0_outputs(5304) <= not((inputs(138)) xor (inputs(96)));
    layer0_outputs(5305) <= (inputs(148)) or (inputs(117));
    layer0_outputs(5306) <= not(inputs(121)) or (inputs(232));
    layer0_outputs(5307) <= not(inputs(29)) or (inputs(157));
    layer0_outputs(5308) <= not(inputs(186)) or (inputs(1));
    layer0_outputs(5309) <= not(inputs(99));
    layer0_outputs(5310) <= not((inputs(31)) or (inputs(44)));
    layer0_outputs(5311) <= not((inputs(33)) or (inputs(40)));
    layer0_outputs(5312) <= (inputs(175)) xor (inputs(222));
    layer0_outputs(5313) <= (inputs(216)) or (inputs(222));
    layer0_outputs(5314) <= (inputs(249)) or (inputs(46));
    layer0_outputs(5315) <= not((inputs(255)) or (inputs(48)));
    layer0_outputs(5316) <= not(inputs(33)) or (inputs(144));
    layer0_outputs(5317) <= not((inputs(16)) xor (inputs(210)));
    layer0_outputs(5318) <= inputs(115);
    layer0_outputs(5319) <= (inputs(235)) or (inputs(166));
    layer0_outputs(5320) <= not(inputs(21)) or (inputs(112));
    layer0_outputs(5321) <= not(inputs(161)) or (inputs(7));
    layer0_outputs(5322) <= not((inputs(74)) or (inputs(239)));
    layer0_outputs(5323) <= not(inputs(103)) or (inputs(19));
    layer0_outputs(5324) <= not(inputs(75)) or (inputs(96));
    layer0_outputs(5325) <= (inputs(41)) xor (inputs(10));
    layer0_outputs(5326) <= inputs(91);
    layer0_outputs(5327) <= not((inputs(138)) or (inputs(175)));
    layer0_outputs(5328) <= (inputs(24)) or (inputs(78));
    layer0_outputs(5329) <= (inputs(106)) or (inputs(35));
    layer0_outputs(5330) <= (inputs(22)) xor (inputs(77));
    layer0_outputs(5331) <= not(inputs(200));
    layer0_outputs(5332) <= (inputs(212)) and not (inputs(110));
    layer0_outputs(5333) <= inputs(62);
    layer0_outputs(5334) <= inputs(140);
    layer0_outputs(5335) <= not(inputs(244));
    layer0_outputs(5336) <= not(inputs(6));
    layer0_outputs(5337) <= (inputs(219)) or (inputs(111));
    layer0_outputs(5338) <= (inputs(90)) and not (inputs(201));
    layer0_outputs(5339) <= not(inputs(65));
    layer0_outputs(5340) <= '1';
    layer0_outputs(5341) <= not((inputs(239)) or (inputs(40)));
    layer0_outputs(5342) <= inputs(110);
    layer0_outputs(5343) <= (inputs(233)) xor (inputs(205));
    layer0_outputs(5344) <= not(inputs(10));
    layer0_outputs(5345) <= not((inputs(14)) xor (inputs(61)));
    layer0_outputs(5346) <= not(inputs(103));
    layer0_outputs(5347) <= (inputs(185)) xor (inputs(149));
    layer0_outputs(5348) <= (inputs(184)) or (inputs(145));
    layer0_outputs(5349) <= (inputs(53)) or (inputs(27));
    layer0_outputs(5350) <= '0';
    layer0_outputs(5351) <= not(inputs(58));
    layer0_outputs(5352) <= not(inputs(65));
    layer0_outputs(5353) <= inputs(6);
    layer0_outputs(5354) <= inputs(149);
    layer0_outputs(5355) <= not(inputs(12)) or (inputs(96));
    layer0_outputs(5356) <= (inputs(36)) and (inputs(42));
    layer0_outputs(5357) <= inputs(149);
    layer0_outputs(5358) <= (inputs(63)) and not (inputs(73));
    layer0_outputs(5359) <= inputs(224);
    layer0_outputs(5360) <= not((inputs(32)) xor (inputs(202)));
    layer0_outputs(5361) <= (inputs(112)) or (inputs(247));
    layer0_outputs(5362) <= not(inputs(215));
    layer0_outputs(5363) <= not((inputs(39)) xor (inputs(67)));
    layer0_outputs(5364) <= inputs(160);
    layer0_outputs(5365) <= not(inputs(25));
    layer0_outputs(5366) <= not(inputs(219)) or (inputs(113));
    layer0_outputs(5367) <= (inputs(197)) and (inputs(209));
    layer0_outputs(5368) <= not(inputs(215));
    layer0_outputs(5369) <= inputs(214);
    layer0_outputs(5370) <= (inputs(245)) or (inputs(238));
    layer0_outputs(5371) <= (inputs(135)) and not (inputs(101));
    layer0_outputs(5372) <= (inputs(39)) or (inputs(60));
    layer0_outputs(5373) <= not(inputs(233));
    layer0_outputs(5374) <= inputs(225);
    layer0_outputs(5375) <= not((inputs(68)) and (inputs(110)));
    layer0_outputs(5376) <= not((inputs(108)) and (inputs(158)));
    layer0_outputs(5377) <= not(inputs(148));
    layer0_outputs(5378) <= not((inputs(23)) xor (inputs(62)));
    layer0_outputs(5379) <= not(inputs(66));
    layer0_outputs(5380) <= (inputs(155)) or (inputs(209));
    layer0_outputs(5381) <= not(inputs(81)) or (inputs(87));
    layer0_outputs(5382) <= not((inputs(153)) and (inputs(197)));
    layer0_outputs(5383) <= not((inputs(35)) xor (inputs(229)));
    layer0_outputs(5384) <= not((inputs(110)) xor (inputs(17)));
    layer0_outputs(5385) <= not(inputs(41)) or (inputs(119));
    layer0_outputs(5386) <= not(inputs(131));
    layer0_outputs(5387) <= not((inputs(157)) or (inputs(227)));
    layer0_outputs(5388) <= inputs(166);
    layer0_outputs(5389) <= (inputs(140)) and not (inputs(6));
    layer0_outputs(5390) <= not(inputs(195));
    layer0_outputs(5391) <= not(inputs(231)) or (inputs(35));
    layer0_outputs(5392) <= (inputs(74)) and (inputs(204));
    layer0_outputs(5393) <= not(inputs(74));
    layer0_outputs(5394) <= (inputs(141)) xor (inputs(249));
    layer0_outputs(5395) <= not((inputs(206)) xor (inputs(237)));
    layer0_outputs(5396) <= inputs(231);
    layer0_outputs(5397) <= not(inputs(232)) or (inputs(46));
    layer0_outputs(5398) <= (inputs(31)) xor (inputs(47));
    layer0_outputs(5399) <= not(inputs(137)) or (inputs(158));
    layer0_outputs(5400) <= inputs(165);
    layer0_outputs(5401) <= inputs(41);
    layer0_outputs(5402) <= inputs(114);
    layer0_outputs(5403) <= not(inputs(195));
    layer0_outputs(5404) <= (inputs(5)) and not (inputs(160));
    layer0_outputs(5405) <= not((inputs(69)) or (inputs(206)));
    layer0_outputs(5406) <= (inputs(5)) xor (inputs(249));
    layer0_outputs(5407) <= not(inputs(61)) or (inputs(206));
    layer0_outputs(5408) <= not(inputs(110)) or (inputs(179));
    layer0_outputs(5409) <= not(inputs(213)) or (inputs(19));
    layer0_outputs(5410) <= not(inputs(58)) or (inputs(100));
    layer0_outputs(5411) <= inputs(251);
    layer0_outputs(5412) <= not(inputs(101));
    layer0_outputs(5413) <= not((inputs(67)) or (inputs(140)));
    layer0_outputs(5414) <= (inputs(90)) xor (inputs(231));
    layer0_outputs(5415) <= (inputs(150)) xor (inputs(144));
    layer0_outputs(5416) <= '1';
    layer0_outputs(5417) <= not(inputs(8)) or (inputs(97));
    layer0_outputs(5418) <= (inputs(91)) and not (inputs(247));
    layer0_outputs(5419) <= inputs(218);
    layer0_outputs(5420) <= not(inputs(59));
    layer0_outputs(5421) <= inputs(195);
    layer0_outputs(5422) <= inputs(128);
    layer0_outputs(5423) <= not(inputs(114));
    layer0_outputs(5424) <= inputs(74);
    layer0_outputs(5425) <= not(inputs(152)) or (inputs(193));
    layer0_outputs(5426) <= (inputs(43)) and (inputs(139));
    layer0_outputs(5427) <= not(inputs(69));
    layer0_outputs(5428) <= (inputs(198)) and not (inputs(50));
    layer0_outputs(5429) <= (inputs(111)) or (inputs(168));
    layer0_outputs(5430) <= not((inputs(3)) xor (inputs(31)));
    layer0_outputs(5431) <= not(inputs(59));
    layer0_outputs(5432) <= not(inputs(183)) or (inputs(207));
    layer0_outputs(5433) <= (inputs(89)) and not (inputs(67));
    layer0_outputs(5434) <= inputs(102);
    layer0_outputs(5435) <= (inputs(191)) and not (inputs(254));
    layer0_outputs(5436) <= (inputs(90)) xor (inputs(188));
    layer0_outputs(5437) <= inputs(154);
    layer0_outputs(5438) <= inputs(157);
    layer0_outputs(5439) <= inputs(166);
    layer0_outputs(5440) <= not((inputs(247)) or (inputs(160)));
    layer0_outputs(5441) <= (inputs(72)) xor (inputs(220));
    layer0_outputs(5442) <= (inputs(93)) or (inputs(105));
    layer0_outputs(5443) <= '1';
    layer0_outputs(5444) <= not((inputs(188)) xor (inputs(157)));
    layer0_outputs(5445) <= not((inputs(187)) or (inputs(19)));
    layer0_outputs(5446) <= (inputs(86)) or (inputs(187));
    layer0_outputs(5447) <= not((inputs(89)) or (inputs(133)));
    layer0_outputs(5448) <= not((inputs(189)) xor (inputs(53)));
    layer0_outputs(5449) <= not(inputs(118));
    layer0_outputs(5450) <= (inputs(53)) xor (inputs(187));
    layer0_outputs(5451) <= (inputs(211)) or (inputs(51));
    layer0_outputs(5452) <= (inputs(154)) or (inputs(237));
    layer0_outputs(5453) <= not(inputs(68)) or (inputs(234));
    layer0_outputs(5454) <= not(inputs(132)) or (inputs(194));
    layer0_outputs(5455) <= not(inputs(77));
    layer0_outputs(5456) <= not((inputs(196)) xor (inputs(202)));
    layer0_outputs(5457) <= not((inputs(152)) xor (inputs(207)));
    layer0_outputs(5458) <= (inputs(105)) and not (inputs(38));
    layer0_outputs(5459) <= not((inputs(221)) or (inputs(190)));
    layer0_outputs(5460) <= not((inputs(208)) and (inputs(108)));
    layer0_outputs(5461) <= not(inputs(77));
    layer0_outputs(5462) <= not(inputs(189));
    layer0_outputs(5463) <= not((inputs(7)) and (inputs(248)));
    layer0_outputs(5464) <= not(inputs(206));
    layer0_outputs(5465) <= (inputs(174)) xor (inputs(196));
    layer0_outputs(5466) <= not(inputs(120));
    layer0_outputs(5467) <= not(inputs(252));
    layer0_outputs(5468) <= not(inputs(250)) or (inputs(172));
    layer0_outputs(5469) <= not(inputs(194));
    layer0_outputs(5470) <= not(inputs(47));
    layer0_outputs(5471) <= inputs(221);
    layer0_outputs(5472) <= (inputs(42)) and not (inputs(251));
    layer0_outputs(5473) <= not(inputs(119)) or (inputs(26));
    layer0_outputs(5474) <= (inputs(149)) or (inputs(106));
    layer0_outputs(5475) <= (inputs(80)) or (inputs(83));
    layer0_outputs(5476) <= (inputs(181)) and not (inputs(123));
    layer0_outputs(5477) <= not((inputs(118)) or (inputs(141)));
    layer0_outputs(5478) <= inputs(83);
    layer0_outputs(5479) <= not(inputs(109));
    layer0_outputs(5480) <= not((inputs(89)) or (inputs(240)));
    layer0_outputs(5481) <= not((inputs(173)) or (inputs(208)));
    layer0_outputs(5482) <= (inputs(41)) or (inputs(178));
    layer0_outputs(5483) <= not((inputs(211)) or (inputs(120)));
    layer0_outputs(5484) <= inputs(164);
    layer0_outputs(5485) <= not((inputs(55)) or (inputs(42)));
    layer0_outputs(5486) <= (inputs(215)) xor (inputs(133));
    layer0_outputs(5487) <= '0';
    layer0_outputs(5488) <= (inputs(121)) xor (inputs(204));
    layer0_outputs(5489) <= not(inputs(86));
    layer0_outputs(5490) <= not(inputs(196));
    layer0_outputs(5491) <= (inputs(183)) and not (inputs(111));
    layer0_outputs(5492) <= not((inputs(82)) xor (inputs(84)));
    layer0_outputs(5493) <= not((inputs(249)) or (inputs(212)));
    layer0_outputs(5494) <= inputs(171);
    layer0_outputs(5495) <= not((inputs(11)) or (inputs(47)));
    layer0_outputs(5496) <= (inputs(114)) and not (inputs(188));
    layer0_outputs(5497) <= (inputs(149)) and not (inputs(247));
    layer0_outputs(5498) <= not((inputs(159)) xor (inputs(22)));
    layer0_outputs(5499) <= not(inputs(211)) or (inputs(13));
    layer0_outputs(5500) <= (inputs(9)) and not (inputs(204));
    layer0_outputs(5501) <= not(inputs(118)) or (inputs(225));
    layer0_outputs(5502) <= inputs(179);
    layer0_outputs(5503) <= (inputs(85)) xor (inputs(23));
    layer0_outputs(5504) <= (inputs(95)) or (inputs(25));
    layer0_outputs(5505) <= inputs(6);
    layer0_outputs(5506) <= not(inputs(26));
    layer0_outputs(5507) <= inputs(43);
    layer0_outputs(5508) <= not(inputs(57)) or (inputs(15));
    layer0_outputs(5509) <= inputs(24);
    layer0_outputs(5510) <= inputs(151);
    layer0_outputs(5511) <= not((inputs(126)) or (inputs(208)));
    layer0_outputs(5512) <= not(inputs(113)) or (inputs(139));
    layer0_outputs(5513) <= not((inputs(176)) or (inputs(42)));
    layer0_outputs(5514) <= (inputs(18)) xor (inputs(26));
    layer0_outputs(5515) <= (inputs(99)) or (inputs(234));
    layer0_outputs(5516) <= inputs(38);
    layer0_outputs(5517) <= (inputs(224)) or (inputs(29));
    layer0_outputs(5518) <= (inputs(23)) xor (inputs(194));
    layer0_outputs(5519) <= not((inputs(149)) or (inputs(227)));
    layer0_outputs(5520) <= not(inputs(187));
    layer0_outputs(5521) <= (inputs(237)) and not (inputs(84));
    layer0_outputs(5522) <= (inputs(47)) or (inputs(219));
    layer0_outputs(5523) <= not(inputs(194));
    layer0_outputs(5524) <= inputs(244);
    layer0_outputs(5525) <= (inputs(46)) xor (inputs(22));
    layer0_outputs(5526) <= inputs(20);
    layer0_outputs(5527) <= not((inputs(10)) or (inputs(110)));
    layer0_outputs(5528) <= (inputs(139)) or (inputs(188));
    layer0_outputs(5529) <= '0';
    layer0_outputs(5530) <= (inputs(152)) and not (inputs(111));
    layer0_outputs(5531) <= (inputs(223)) xor (inputs(75));
    layer0_outputs(5532) <= inputs(150);
    layer0_outputs(5533) <= not(inputs(163));
    layer0_outputs(5534) <= inputs(4);
    layer0_outputs(5535) <= inputs(97);
    layer0_outputs(5536) <= (inputs(20)) and (inputs(117));
    layer0_outputs(5537) <= not(inputs(153));
    layer0_outputs(5538) <= not(inputs(180)) or (inputs(66));
    layer0_outputs(5539) <= not((inputs(147)) and (inputs(178)));
    layer0_outputs(5540) <= not((inputs(173)) or (inputs(54)));
    layer0_outputs(5541) <= (inputs(19)) xor (inputs(144));
    layer0_outputs(5542) <= not(inputs(0)) or (inputs(177));
    layer0_outputs(5543) <= inputs(248);
    layer0_outputs(5544) <= not((inputs(5)) and (inputs(150)));
    layer0_outputs(5545) <= (inputs(67)) xor (inputs(37));
    layer0_outputs(5546) <= (inputs(25)) xor (inputs(169));
    layer0_outputs(5547) <= (inputs(177)) xor (inputs(181));
    layer0_outputs(5548) <= inputs(93);
    layer0_outputs(5549) <= (inputs(47)) or (inputs(99));
    layer0_outputs(5550) <= not(inputs(45));
    layer0_outputs(5551) <= not((inputs(65)) xor (inputs(219)));
    layer0_outputs(5552) <= (inputs(247)) and not (inputs(48));
    layer0_outputs(5553) <= inputs(98);
    layer0_outputs(5554) <= inputs(103);
    layer0_outputs(5555) <= (inputs(137)) and not (inputs(166));
    layer0_outputs(5556) <= not(inputs(163)) or (inputs(82));
    layer0_outputs(5557) <= not(inputs(247));
    layer0_outputs(5558) <= inputs(115);
    layer0_outputs(5559) <= (inputs(229)) and not (inputs(121));
    layer0_outputs(5560) <= (inputs(29)) and (inputs(220));
    layer0_outputs(5561) <= not(inputs(178));
    layer0_outputs(5562) <= inputs(10);
    layer0_outputs(5563) <= inputs(151);
    layer0_outputs(5564) <= (inputs(75)) and not (inputs(15));
    layer0_outputs(5565) <= (inputs(15)) or (inputs(180));
    layer0_outputs(5566) <= not((inputs(57)) or (inputs(167)));
    layer0_outputs(5567) <= not((inputs(57)) or (inputs(218)));
    layer0_outputs(5568) <= not((inputs(207)) or (inputs(152)));
    layer0_outputs(5569) <= (inputs(236)) or (inputs(125));
    layer0_outputs(5570) <= not(inputs(59));
    layer0_outputs(5571) <= inputs(58);
    layer0_outputs(5572) <= not((inputs(64)) xor (inputs(18)));
    layer0_outputs(5573) <= not((inputs(56)) or (inputs(245)));
    layer0_outputs(5574) <= inputs(119);
    layer0_outputs(5575) <= (inputs(169)) and not (inputs(105));
    layer0_outputs(5576) <= (inputs(23)) and not (inputs(177));
    layer0_outputs(5577) <= not(inputs(109));
    layer0_outputs(5578) <= (inputs(50)) or (inputs(139));
    layer0_outputs(5579) <= inputs(232);
    layer0_outputs(5580) <= (inputs(92)) xor (inputs(78));
    layer0_outputs(5581) <= not((inputs(78)) or (inputs(28)));
    layer0_outputs(5582) <= not((inputs(171)) and (inputs(186)));
    layer0_outputs(5583) <= not((inputs(63)) or (inputs(32)));
    layer0_outputs(5584) <= (inputs(192)) and not (inputs(234));
    layer0_outputs(5585) <= (inputs(175)) or (inputs(117));
    layer0_outputs(5586) <= inputs(185);
    layer0_outputs(5587) <= not(inputs(75));
    layer0_outputs(5588) <= (inputs(213)) and (inputs(172));
    layer0_outputs(5589) <= not(inputs(229));
    layer0_outputs(5590) <= (inputs(179)) and not (inputs(93));
    layer0_outputs(5591) <= inputs(161);
    layer0_outputs(5592) <= (inputs(191)) and (inputs(114));
    layer0_outputs(5593) <= not(inputs(105));
    layer0_outputs(5594) <= not(inputs(103));
    layer0_outputs(5595) <= not(inputs(135));
    layer0_outputs(5596) <= not((inputs(37)) and (inputs(19)));
    layer0_outputs(5597) <= not((inputs(51)) or (inputs(88)));
    layer0_outputs(5598) <= (inputs(190)) or (inputs(115));
    layer0_outputs(5599) <= inputs(161);
    layer0_outputs(5600) <= not((inputs(18)) xor (inputs(71)));
    layer0_outputs(5601) <= inputs(198);
    layer0_outputs(5602) <= not(inputs(31)) or (inputs(127));
    layer0_outputs(5603) <= (inputs(107)) and not (inputs(167));
    layer0_outputs(5604) <= inputs(110);
    layer0_outputs(5605) <= not(inputs(165));
    layer0_outputs(5606) <= '1';
    layer0_outputs(5607) <= not((inputs(207)) xor (inputs(32)));
    layer0_outputs(5608) <= not((inputs(19)) xor (inputs(51)));
    layer0_outputs(5609) <= (inputs(227)) and not (inputs(93));
    layer0_outputs(5610) <= (inputs(239)) or (inputs(28));
    layer0_outputs(5611) <= (inputs(159)) and (inputs(102));
    layer0_outputs(5612) <= not((inputs(64)) or (inputs(90)));
    layer0_outputs(5613) <= not(inputs(103));
    layer0_outputs(5614) <= not(inputs(164)) or (inputs(107));
    layer0_outputs(5615) <= (inputs(148)) or (inputs(169));
    layer0_outputs(5616) <= (inputs(88)) xor (inputs(93));
    layer0_outputs(5617) <= inputs(143);
    layer0_outputs(5618) <= not(inputs(244)) or (inputs(245));
    layer0_outputs(5619) <= (inputs(197)) or (inputs(176));
    layer0_outputs(5620) <= (inputs(155)) xor (inputs(173));
    layer0_outputs(5621) <= inputs(213);
    layer0_outputs(5622) <= (inputs(39)) and not (inputs(200));
    layer0_outputs(5623) <= not(inputs(18));
    layer0_outputs(5624) <= inputs(71);
    layer0_outputs(5625) <= inputs(176);
    layer0_outputs(5626) <= (inputs(63)) and (inputs(206));
    layer0_outputs(5627) <= (inputs(115)) or (inputs(111));
    layer0_outputs(5628) <= (inputs(214)) or (inputs(200));
    layer0_outputs(5629) <= inputs(229);
    layer0_outputs(5630) <= inputs(42);
    layer0_outputs(5631) <= (inputs(170)) or (inputs(19));
    layer0_outputs(5632) <= not(inputs(12)) or (inputs(223));
    layer0_outputs(5633) <= not(inputs(233));
    layer0_outputs(5634) <= not(inputs(175));
    layer0_outputs(5635) <= (inputs(93)) xor (inputs(28));
    layer0_outputs(5636) <= (inputs(87)) xor (inputs(139));
    layer0_outputs(5637) <= not((inputs(65)) or (inputs(120)));
    layer0_outputs(5638) <= not(inputs(19)) or (inputs(252));
    layer0_outputs(5639) <= (inputs(4)) xor (inputs(26));
    layer0_outputs(5640) <= (inputs(64)) and not (inputs(145));
    layer0_outputs(5641) <= (inputs(162)) or (inputs(235));
    layer0_outputs(5642) <= (inputs(68)) and (inputs(85));
    layer0_outputs(5643) <= (inputs(213)) and not (inputs(156));
    layer0_outputs(5644) <= not((inputs(13)) or (inputs(182)));
    layer0_outputs(5645) <= (inputs(238)) xor (inputs(191));
    layer0_outputs(5646) <= inputs(39);
    layer0_outputs(5647) <= (inputs(10)) xor (inputs(6));
    layer0_outputs(5648) <= inputs(167);
    layer0_outputs(5649) <= inputs(120);
    layer0_outputs(5650) <= not(inputs(40)) or (inputs(85));
    layer0_outputs(5651) <= not(inputs(244)) or (inputs(255));
    layer0_outputs(5652) <= inputs(83);
    layer0_outputs(5653) <= not((inputs(207)) or (inputs(186)));
    layer0_outputs(5654) <= (inputs(179)) or (inputs(158));
    layer0_outputs(5655) <= not(inputs(232)) or (inputs(1));
    layer0_outputs(5656) <= not(inputs(114)) or (inputs(138));
    layer0_outputs(5657) <= not((inputs(42)) or (inputs(162)));
    layer0_outputs(5658) <= (inputs(243)) or (inputs(148));
    layer0_outputs(5659) <= (inputs(77)) and not (inputs(222));
    layer0_outputs(5660) <= not((inputs(76)) or (inputs(51)));
    layer0_outputs(5661) <= (inputs(15)) or (inputs(123));
    layer0_outputs(5662) <= inputs(183);
    layer0_outputs(5663) <= (inputs(23)) xor (inputs(232));
    layer0_outputs(5664) <= not(inputs(230));
    layer0_outputs(5665) <= not((inputs(134)) or (inputs(58)));
    layer0_outputs(5666) <= (inputs(138)) and not (inputs(227));
    layer0_outputs(5667) <= inputs(6);
    layer0_outputs(5668) <= not(inputs(188));
    layer0_outputs(5669) <= inputs(143);
    layer0_outputs(5670) <= not(inputs(20));
    layer0_outputs(5671) <= not((inputs(59)) xor (inputs(16)));
    layer0_outputs(5672) <= inputs(211);
    layer0_outputs(5673) <= not(inputs(234));
    layer0_outputs(5674) <= not((inputs(143)) or (inputs(235)));
    layer0_outputs(5675) <= (inputs(197)) xor (inputs(32));
    layer0_outputs(5676) <= not((inputs(206)) or (inputs(57)));
    layer0_outputs(5677) <= (inputs(246)) and not (inputs(132));
    layer0_outputs(5678) <= not((inputs(50)) xor (inputs(3)));
    layer0_outputs(5679) <= inputs(98);
    layer0_outputs(5680) <= not(inputs(8)) or (inputs(239));
    layer0_outputs(5681) <= inputs(252);
    layer0_outputs(5682) <= not((inputs(151)) and (inputs(57)));
    layer0_outputs(5683) <= not(inputs(226)) or (inputs(47));
    layer0_outputs(5684) <= (inputs(174)) and not (inputs(29));
    layer0_outputs(5685) <= (inputs(144)) xor (inputs(16));
    layer0_outputs(5686) <= not(inputs(83));
    layer0_outputs(5687) <= not((inputs(106)) xor (inputs(167)));
    layer0_outputs(5688) <= (inputs(197)) and not (inputs(89));
    layer0_outputs(5689) <= not((inputs(244)) or (inputs(207)));
    layer0_outputs(5690) <= not(inputs(75));
    layer0_outputs(5691) <= not((inputs(61)) or (inputs(150)));
    layer0_outputs(5692) <= not(inputs(17)) or (inputs(82));
    layer0_outputs(5693) <= not(inputs(119));
    layer0_outputs(5694) <= not(inputs(93));
    layer0_outputs(5695) <= inputs(6);
    layer0_outputs(5696) <= (inputs(77)) or (inputs(121));
    layer0_outputs(5697) <= (inputs(90)) xor (inputs(253));
    layer0_outputs(5698) <= inputs(73);
    layer0_outputs(5699) <= '1';
    layer0_outputs(5700) <= (inputs(250)) and (inputs(152));
    layer0_outputs(5701) <= not((inputs(208)) or (inputs(114)));
    layer0_outputs(5702) <= not(inputs(40));
    layer0_outputs(5703) <= inputs(252);
    layer0_outputs(5704) <= not(inputs(149));
    layer0_outputs(5705) <= not(inputs(63)) or (inputs(129));
    layer0_outputs(5706) <= not(inputs(180));
    layer0_outputs(5707) <= not(inputs(221)) or (inputs(206));
    layer0_outputs(5708) <= not(inputs(4)) or (inputs(53));
    layer0_outputs(5709) <= not(inputs(74));
    layer0_outputs(5710) <= (inputs(178)) and not (inputs(119));
    layer0_outputs(5711) <= inputs(43);
    layer0_outputs(5712) <= (inputs(250)) and not (inputs(49));
    layer0_outputs(5713) <= (inputs(35)) or (inputs(53));
    layer0_outputs(5714) <= not(inputs(88)) or (inputs(49));
    layer0_outputs(5715) <= inputs(155);
    layer0_outputs(5716) <= not(inputs(130));
    layer0_outputs(5717) <= (inputs(43)) xor (inputs(93));
    layer0_outputs(5718) <= not(inputs(211)) or (inputs(125));
    layer0_outputs(5719) <= not((inputs(255)) or (inputs(47)));
    layer0_outputs(5720) <= not((inputs(201)) or (inputs(124)));
    layer0_outputs(5721) <= not((inputs(119)) or (inputs(158)));
    layer0_outputs(5722) <= inputs(122);
    layer0_outputs(5723) <= not((inputs(82)) xor (inputs(170)));
    layer0_outputs(5724) <= not(inputs(234)) or (inputs(123));
    layer0_outputs(5725) <= inputs(155);
    layer0_outputs(5726) <= not(inputs(213)) or (inputs(93));
    layer0_outputs(5727) <= not((inputs(142)) or (inputs(222)));
    layer0_outputs(5728) <= not(inputs(99)) or (inputs(251));
    layer0_outputs(5729) <= not(inputs(254));
    layer0_outputs(5730) <= not((inputs(56)) or (inputs(104)));
    layer0_outputs(5731) <= inputs(212);
    layer0_outputs(5732) <= inputs(180);
    layer0_outputs(5733) <= (inputs(249)) xor (inputs(236));
    layer0_outputs(5734) <= not(inputs(215));
    layer0_outputs(5735) <= not(inputs(112));
    layer0_outputs(5736) <= not((inputs(8)) or (inputs(54)));
    layer0_outputs(5737) <= (inputs(155)) or (inputs(41));
    layer0_outputs(5738) <= not(inputs(214)) or (inputs(67));
    layer0_outputs(5739) <= inputs(186);
    layer0_outputs(5740) <= (inputs(224)) or (inputs(149));
    layer0_outputs(5741) <= (inputs(247)) xor (inputs(243));
    layer0_outputs(5742) <= not((inputs(34)) xor (inputs(244)));
    layer0_outputs(5743) <= inputs(94);
    layer0_outputs(5744) <= not((inputs(41)) xor (inputs(175)));
    layer0_outputs(5745) <= (inputs(203)) and not (inputs(5));
    layer0_outputs(5746) <= not((inputs(212)) and (inputs(132)));
    layer0_outputs(5747) <= inputs(69);
    layer0_outputs(5748) <= not(inputs(36));
    layer0_outputs(5749) <= not((inputs(253)) and (inputs(173)));
    layer0_outputs(5750) <= inputs(198);
    layer0_outputs(5751) <= inputs(85);
    layer0_outputs(5752) <= (inputs(68)) or (inputs(165));
    layer0_outputs(5753) <= (inputs(205)) xor (inputs(64));
    layer0_outputs(5754) <= not((inputs(252)) xor (inputs(175)));
    layer0_outputs(5755) <= (inputs(69)) xor (inputs(52));
    layer0_outputs(5756) <= not(inputs(130)) or (inputs(152));
    layer0_outputs(5757) <= (inputs(146)) or (inputs(182));
    layer0_outputs(5758) <= (inputs(96)) xor (inputs(185));
    layer0_outputs(5759) <= not(inputs(189)) or (inputs(93));
    layer0_outputs(5760) <= (inputs(204)) and not (inputs(29));
    layer0_outputs(5761) <= inputs(59);
    layer0_outputs(5762) <= not(inputs(218));
    layer0_outputs(5763) <= inputs(206);
    layer0_outputs(5764) <= not((inputs(97)) or (inputs(149)));
    layer0_outputs(5765) <= not(inputs(124));
    layer0_outputs(5766) <= (inputs(206)) or (inputs(162));
    layer0_outputs(5767) <= not((inputs(154)) and (inputs(83)));
    layer0_outputs(5768) <= inputs(10);
    layer0_outputs(5769) <= (inputs(122)) xor (inputs(204));
    layer0_outputs(5770) <= not(inputs(24));
    layer0_outputs(5771) <= not((inputs(31)) xor (inputs(109)));
    layer0_outputs(5772) <= '1';
    layer0_outputs(5773) <= not(inputs(79)) or (inputs(208));
    layer0_outputs(5774) <= inputs(122);
    layer0_outputs(5775) <= (inputs(89)) and not (inputs(35));
    layer0_outputs(5776) <= (inputs(125)) or (inputs(130));
    layer0_outputs(5777) <= not(inputs(7));
    layer0_outputs(5778) <= (inputs(201)) or (inputs(61));
    layer0_outputs(5779) <= not(inputs(115));
    layer0_outputs(5780) <= (inputs(11)) and not (inputs(237));
    layer0_outputs(5781) <= inputs(81);
    layer0_outputs(5782) <= not((inputs(76)) or (inputs(77)));
    layer0_outputs(5783) <= not((inputs(211)) or (inputs(187)));
    layer0_outputs(5784) <= not((inputs(97)) or (inputs(8)));
    layer0_outputs(5785) <= inputs(46);
    layer0_outputs(5786) <= '1';
    layer0_outputs(5787) <= not((inputs(223)) xor (inputs(53)));
    layer0_outputs(5788) <= (inputs(197)) xor (inputs(217));
    layer0_outputs(5789) <= not((inputs(196)) xor (inputs(42)));
    layer0_outputs(5790) <= not(inputs(204)) or (inputs(126));
    layer0_outputs(5791) <= not(inputs(179)) or (inputs(15));
    layer0_outputs(5792) <= '1';
    layer0_outputs(5793) <= not((inputs(82)) or (inputs(78)));
    layer0_outputs(5794) <= inputs(23);
    layer0_outputs(5795) <= (inputs(217)) and not (inputs(33));
    layer0_outputs(5796) <= (inputs(249)) or (inputs(27));
    layer0_outputs(5797) <= (inputs(83)) and not (inputs(254));
    layer0_outputs(5798) <= not(inputs(246));
    layer0_outputs(5799) <= not(inputs(122));
    layer0_outputs(5800) <= (inputs(173)) or (inputs(229));
    layer0_outputs(5801) <= (inputs(142)) and not (inputs(197));
    layer0_outputs(5802) <= inputs(22);
    layer0_outputs(5803) <= (inputs(123)) or (inputs(245));
    layer0_outputs(5804) <= (inputs(132)) or (inputs(65));
    layer0_outputs(5805) <= not((inputs(243)) or (inputs(17)));
    layer0_outputs(5806) <= not(inputs(13));
    layer0_outputs(5807) <= (inputs(100)) or (inputs(118));
    layer0_outputs(5808) <= (inputs(176)) and not (inputs(45));
    layer0_outputs(5809) <= inputs(216);
    layer0_outputs(5810) <= not((inputs(115)) xor (inputs(248)));
    layer0_outputs(5811) <= (inputs(75)) and (inputs(122));
    layer0_outputs(5812) <= inputs(206);
    layer0_outputs(5813) <= not(inputs(68));
    layer0_outputs(5814) <= inputs(113);
    layer0_outputs(5815) <= (inputs(38)) and not (inputs(102));
    layer0_outputs(5816) <= not((inputs(16)) or (inputs(249)));
    layer0_outputs(5817) <= not(inputs(216)) or (inputs(17));
    layer0_outputs(5818) <= (inputs(225)) and not (inputs(253));
    layer0_outputs(5819) <= not(inputs(150));
    layer0_outputs(5820) <= not((inputs(42)) xor (inputs(90)));
    layer0_outputs(5821) <= inputs(14);
    layer0_outputs(5822) <= (inputs(223)) and not (inputs(111));
    layer0_outputs(5823) <= (inputs(127)) and not (inputs(89));
    layer0_outputs(5824) <= not(inputs(44));
    layer0_outputs(5825) <= (inputs(120)) xor (inputs(130));
    layer0_outputs(5826) <= not(inputs(186)) or (inputs(3));
    layer0_outputs(5827) <= not((inputs(106)) and (inputs(95)));
    layer0_outputs(5828) <= not(inputs(43));
    layer0_outputs(5829) <= not((inputs(49)) or (inputs(234)));
    layer0_outputs(5830) <= (inputs(53)) and not (inputs(225));
    layer0_outputs(5831) <= (inputs(48)) xor (inputs(247));
    layer0_outputs(5832) <= not(inputs(120)) or (inputs(235));
    layer0_outputs(5833) <= (inputs(238)) or (inputs(35));
    layer0_outputs(5834) <= not(inputs(199));
    layer0_outputs(5835) <= (inputs(235)) and not (inputs(7));
    layer0_outputs(5836) <= inputs(179);
    layer0_outputs(5837) <= (inputs(214)) and not (inputs(113));
    layer0_outputs(5838) <= inputs(120);
    layer0_outputs(5839) <= '1';
    layer0_outputs(5840) <= (inputs(138)) or (inputs(252));
    layer0_outputs(5841) <= (inputs(67)) xor (inputs(163));
    layer0_outputs(5842) <= not(inputs(120)) or (inputs(80));
    layer0_outputs(5843) <= (inputs(31)) or (inputs(4));
    layer0_outputs(5844) <= not(inputs(59));
    layer0_outputs(5845) <= not((inputs(26)) and (inputs(89)));
    layer0_outputs(5846) <= not((inputs(128)) or (inputs(246)));
    layer0_outputs(5847) <= (inputs(230)) and not (inputs(64));
    layer0_outputs(5848) <= not(inputs(226));
    layer0_outputs(5849) <= not(inputs(66));
    layer0_outputs(5850) <= not(inputs(91));
    layer0_outputs(5851) <= (inputs(126)) and not (inputs(218));
    layer0_outputs(5852) <= not(inputs(230));
    layer0_outputs(5853) <= not(inputs(124)) or (inputs(224));
    layer0_outputs(5854) <= not(inputs(44));
    layer0_outputs(5855) <= not((inputs(219)) xor (inputs(60)));
    layer0_outputs(5856) <= not((inputs(125)) xor (inputs(17)));
    layer0_outputs(5857) <= not((inputs(225)) xor (inputs(80)));
    layer0_outputs(5858) <= not((inputs(47)) or (inputs(214)));
    layer0_outputs(5859) <= inputs(99);
    layer0_outputs(5860) <= (inputs(32)) or (inputs(36));
    layer0_outputs(5861) <= (inputs(113)) or (inputs(72));
    layer0_outputs(5862) <= (inputs(134)) or (inputs(101));
    layer0_outputs(5863) <= not(inputs(184)) or (inputs(106));
    layer0_outputs(5864) <= not((inputs(7)) or (inputs(31)));
    layer0_outputs(5865) <= (inputs(3)) and (inputs(239));
    layer0_outputs(5866) <= not(inputs(9));
    layer0_outputs(5867) <= not(inputs(178)) or (inputs(169));
    layer0_outputs(5868) <= not((inputs(147)) xor (inputs(86)));
    layer0_outputs(5869) <= not(inputs(171));
    layer0_outputs(5870) <= not((inputs(118)) or (inputs(224)));
    layer0_outputs(5871) <= not(inputs(243));
    layer0_outputs(5872) <= not(inputs(138)) or (inputs(72));
    layer0_outputs(5873) <= inputs(152);
    layer0_outputs(5874) <= (inputs(142)) or (inputs(111));
    layer0_outputs(5875) <= (inputs(84)) or (inputs(19));
    layer0_outputs(5876) <= not((inputs(75)) xor (inputs(79)));
    layer0_outputs(5877) <= not(inputs(189)) or (inputs(68));
    layer0_outputs(5878) <= '0';
    layer0_outputs(5879) <= inputs(194);
    layer0_outputs(5880) <= not(inputs(55));
    layer0_outputs(5881) <= not(inputs(78));
    layer0_outputs(5882) <= (inputs(129)) and not (inputs(174));
    layer0_outputs(5883) <= not((inputs(45)) or (inputs(200)));
    layer0_outputs(5884) <= not((inputs(57)) xor (inputs(72)));
    layer0_outputs(5885) <= not(inputs(87));
    layer0_outputs(5886) <= (inputs(35)) xor (inputs(172));
    layer0_outputs(5887) <= not((inputs(8)) or (inputs(21)));
    layer0_outputs(5888) <= not((inputs(220)) and (inputs(106)));
    layer0_outputs(5889) <= not((inputs(37)) xor (inputs(61)));
    layer0_outputs(5890) <= (inputs(242)) or (inputs(82));
    layer0_outputs(5891) <= (inputs(159)) or (inputs(241));
    layer0_outputs(5892) <= not(inputs(18));
    layer0_outputs(5893) <= inputs(122);
    layer0_outputs(5894) <= not(inputs(56)) or (inputs(18));
    layer0_outputs(5895) <= not(inputs(221));
    layer0_outputs(5896) <= inputs(85);
    layer0_outputs(5897) <= not(inputs(61));
    layer0_outputs(5898) <= not(inputs(21)) or (inputs(188));
    layer0_outputs(5899) <= (inputs(178)) and not (inputs(77));
    layer0_outputs(5900) <= inputs(99);
    layer0_outputs(5901) <= not(inputs(50)) or (inputs(208));
    layer0_outputs(5902) <= (inputs(123)) xor (inputs(232));
    layer0_outputs(5903) <= (inputs(53)) xor (inputs(46));
    layer0_outputs(5904) <= not((inputs(184)) xor (inputs(142)));
    layer0_outputs(5905) <= (inputs(203)) and not (inputs(17));
    layer0_outputs(5906) <= not((inputs(94)) xor (inputs(6)));
    layer0_outputs(5907) <= not((inputs(237)) or (inputs(195)));
    layer0_outputs(5908) <= (inputs(229)) and not (inputs(47));
    layer0_outputs(5909) <= inputs(30);
    layer0_outputs(5910) <= (inputs(230)) or (inputs(78));
    layer0_outputs(5911) <= not(inputs(122));
    layer0_outputs(5912) <= (inputs(181)) and not (inputs(59));
    layer0_outputs(5913) <= not(inputs(195)) or (inputs(137));
    layer0_outputs(5914) <= (inputs(147)) xor (inputs(234));
    layer0_outputs(5915) <= (inputs(180)) or (inputs(229));
    layer0_outputs(5916) <= not(inputs(57));
    layer0_outputs(5917) <= (inputs(98)) xor (inputs(209));
    layer0_outputs(5918) <= not(inputs(82));
    layer0_outputs(5919) <= not(inputs(25));
    layer0_outputs(5920) <= not((inputs(63)) xor (inputs(243)));
    layer0_outputs(5921) <= not(inputs(140));
    layer0_outputs(5922) <= (inputs(166)) xor (inputs(94));
    layer0_outputs(5923) <= not((inputs(44)) or (inputs(141)));
    layer0_outputs(5924) <= inputs(174);
    layer0_outputs(5925) <= not((inputs(147)) or (inputs(164)));
    layer0_outputs(5926) <= not((inputs(72)) or (inputs(91)));
    layer0_outputs(5927) <= (inputs(5)) or (inputs(22));
    layer0_outputs(5928) <= not(inputs(188));
    layer0_outputs(5929) <= inputs(25);
    layer0_outputs(5930) <= inputs(2);
    layer0_outputs(5931) <= not(inputs(114));
    layer0_outputs(5932) <= not((inputs(177)) or (inputs(89)));
    layer0_outputs(5933) <= '0';
    layer0_outputs(5934) <= inputs(177);
    layer0_outputs(5935) <= not(inputs(139));
    layer0_outputs(5936) <= not(inputs(7)) or (inputs(227));
    layer0_outputs(5937) <= not((inputs(155)) and (inputs(135)));
    layer0_outputs(5938) <= not((inputs(40)) xor (inputs(23)));
    layer0_outputs(5939) <= not((inputs(78)) or (inputs(145)));
    layer0_outputs(5940) <= (inputs(65)) and not (inputs(38));
    layer0_outputs(5941) <= not(inputs(182));
    layer0_outputs(5942) <= (inputs(65)) or (inputs(255));
    layer0_outputs(5943) <= not(inputs(49)) or (inputs(158));
    layer0_outputs(5944) <= inputs(246);
    layer0_outputs(5945) <= not((inputs(148)) or (inputs(183)));
    layer0_outputs(5946) <= (inputs(189)) or (inputs(31));
    layer0_outputs(5947) <= not((inputs(170)) or (inputs(205)));
    layer0_outputs(5948) <= not((inputs(12)) xor (inputs(111)));
    layer0_outputs(5949) <= not(inputs(64));
    layer0_outputs(5950) <= inputs(111);
    layer0_outputs(5951) <= not(inputs(3)) or (inputs(14));
    layer0_outputs(5952) <= (inputs(130)) and not (inputs(28));
    layer0_outputs(5953) <= not(inputs(87));
    layer0_outputs(5954) <= not(inputs(204)) or (inputs(127));
    layer0_outputs(5955) <= (inputs(57)) xor (inputs(27));
    layer0_outputs(5956) <= (inputs(67)) and not (inputs(206));
    layer0_outputs(5957) <= (inputs(240)) or (inputs(219));
    layer0_outputs(5958) <= (inputs(92)) and (inputs(81));
    layer0_outputs(5959) <= (inputs(150)) xor (inputs(129));
    layer0_outputs(5960) <= not((inputs(181)) xor (inputs(77)));
    layer0_outputs(5961) <= not((inputs(226)) or (inputs(32)));
    layer0_outputs(5962) <= (inputs(3)) or (inputs(38));
    layer0_outputs(5963) <= inputs(57);
    layer0_outputs(5964) <= inputs(13);
    layer0_outputs(5965) <= (inputs(218)) xor (inputs(254));
    layer0_outputs(5966) <= not(inputs(207));
    layer0_outputs(5967) <= inputs(178);
    layer0_outputs(5968) <= not((inputs(20)) xor (inputs(209)));
    layer0_outputs(5969) <= not((inputs(3)) xor (inputs(130)));
    layer0_outputs(5970) <= (inputs(40)) and (inputs(41));
    layer0_outputs(5971) <= not(inputs(99));
    layer0_outputs(5972) <= (inputs(46)) or (inputs(184));
    layer0_outputs(5973) <= not(inputs(241)) or (inputs(179));
    layer0_outputs(5974) <= (inputs(138)) and (inputs(125));
    layer0_outputs(5975) <= not(inputs(222)) or (inputs(95));
    layer0_outputs(5976) <= (inputs(195)) or (inputs(232));
    layer0_outputs(5977) <= (inputs(19)) xor (inputs(222));
    layer0_outputs(5978) <= (inputs(21)) xor (inputs(46));
    layer0_outputs(5979) <= (inputs(63)) and not (inputs(18));
    layer0_outputs(5980) <= inputs(91);
    layer0_outputs(5981) <= not((inputs(119)) xor (inputs(54)));
    layer0_outputs(5982) <= (inputs(163)) or (inputs(110));
    layer0_outputs(5983) <= not(inputs(226)) or (inputs(129));
    layer0_outputs(5984) <= not(inputs(152));
    layer0_outputs(5985) <= not(inputs(249)) or (inputs(13));
    layer0_outputs(5986) <= not(inputs(178));
    layer0_outputs(5987) <= inputs(105);
    layer0_outputs(5988) <= not((inputs(36)) xor (inputs(156)));
    layer0_outputs(5989) <= inputs(248);
    layer0_outputs(5990) <= (inputs(92)) and not (inputs(105));
    layer0_outputs(5991) <= inputs(119);
    layer0_outputs(5992) <= (inputs(60)) and not (inputs(131));
    layer0_outputs(5993) <= (inputs(178)) or (inputs(194));
    layer0_outputs(5994) <= inputs(107);
    layer0_outputs(5995) <= (inputs(162)) xor (inputs(58));
    layer0_outputs(5996) <= not(inputs(147));
    layer0_outputs(5997) <= not((inputs(63)) or (inputs(246)));
    layer0_outputs(5998) <= '1';
    layer0_outputs(5999) <= not((inputs(181)) xor (inputs(89)));
    layer0_outputs(6000) <= (inputs(60)) xor (inputs(245));
    layer0_outputs(6001) <= not(inputs(1));
    layer0_outputs(6002) <= (inputs(157)) and not (inputs(80));
    layer0_outputs(6003) <= not(inputs(140));
    layer0_outputs(6004) <= (inputs(86)) xor (inputs(94));
    layer0_outputs(6005) <= not((inputs(241)) xor (inputs(147)));
    layer0_outputs(6006) <= not(inputs(131));
    layer0_outputs(6007) <= not((inputs(187)) xor (inputs(136)));
    layer0_outputs(6008) <= not((inputs(38)) xor (inputs(74)));
    layer0_outputs(6009) <= (inputs(15)) or (inputs(196));
    layer0_outputs(6010) <= not((inputs(63)) or (inputs(39)));
    layer0_outputs(6011) <= not((inputs(206)) or (inputs(92)));
    layer0_outputs(6012) <= not((inputs(228)) and (inputs(228)));
    layer0_outputs(6013) <= not(inputs(8));
    layer0_outputs(6014) <= not(inputs(29));
    layer0_outputs(6015) <= not(inputs(232));
    layer0_outputs(6016) <= not((inputs(113)) xor (inputs(100)));
    layer0_outputs(6017) <= inputs(153);
    layer0_outputs(6018) <= not((inputs(107)) xor (inputs(65)));
    layer0_outputs(6019) <= not(inputs(117)) or (inputs(55));
    layer0_outputs(6020) <= not((inputs(145)) and (inputs(210)));
    layer0_outputs(6021) <= (inputs(184)) xor (inputs(248));
    layer0_outputs(6022) <= inputs(7);
    layer0_outputs(6023) <= not((inputs(86)) xor (inputs(18)));
    layer0_outputs(6024) <= not(inputs(132));
    layer0_outputs(6025) <= (inputs(66)) or (inputs(249));
    layer0_outputs(6026) <= inputs(49);
    layer0_outputs(6027) <= not(inputs(218)) or (inputs(49));
    layer0_outputs(6028) <= '1';
    layer0_outputs(6029) <= inputs(163);
    layer0_outputs(6030) <= not((inputs(44)) xor (inputs(63)));
    layer0_outputs(6031) <= not((inputs(255)) or (inputs(88)));
    layer0_outputs(6032) <= inputs(211);
    layer0_outputs(6033) <= inputs(124);
    layer0_outputs(6034) <= not((inputs(24)) xor (inputs(175)));
    layer0_outputs(6035) <= not(inputs(93));
    layer0_outputs(6036) <= (inputs(22)) and not (inputs(29));
    layer0_outputs(6037) <= not(inputs(220)) or (inputs(48));
    layer0_outputs(6038) <= inputs(153);
    layer0_outputs(6039) <= not(inputs(136));
    layer0_outputs(6040) <= not(inputs(234)) or (inputs(66));
    layer0_outputs(6041) <= (inputs(30)) and (inputs(240));
    layer0_outputs(6042) <= not((inputs(150)) xor (inputs(64)));
    layer0_outputs(6043) <= inputs(105);
    layer0_outputs(6044) <= not(inputs(244)) or (inputs(7));
    layer0_outputs(6045) <= not((inputs(203)) or (inputs(170)));
    layer0_outputs(6046) <= (inputs(108)) xor (inputs(143));
    layer0_outputs(6047) <= (inputs(61)) and not (inputs(223));
    layer0_outputs(6048) <= inputs(7);
    layer0_outputs(6049) <= inputs(170);
    layer0_outputs(6050) <= inputs(179);
    layer0_outputs(6051) <= not(inputs(72));
    layer0_outputs(6052) <= not((inputs(179)) or (inputs(142)));
    layer0_outputs(6053) <= inputs(196);
    layer0_outputs(6054) <= (inputs(178)) xor (inputs(173));
    layer0_outputs(6055) <= not(inputs(91));
    layer0_outputs(6056) <= (inputs(94)) or (inputs(25));
    layer0_outputs(6057) <= not(inputs(47));
    layer0_outputs(6058) <= '0';
    layer0_outputs(6059) <= '1';
    layer0_outputs(6060) <= (inputs(230)) and not (inputs(91));
    layer0_outputs(6061) <= not((inputs(236)) xor (inputs(203)));
    layer0_outputs(6062) <= '0';
    layer0_outputs(6063) <= inputs(213);
    layer0_outputs(6064) <= not((inputs(100)) or (inputs(113)));
    layer0_outputs(6065) <= not(inputs(162)) or (inputs(253));
    layer0_outputs(6066) <= not((inputs(53)) or (inputs(254)));
    layer0_outputs(6067) <= inputs(83);
    layer0_outputs(6068) <= not(inputs(244));
    layer0_outputs(6069) <= inputs(197);
    layer0_outputs(6070) <= not((inputs(117)) xor (inputs(208)));
    layer0_outputs(6071) <= not(inputs(70)) or (inputs(109));
    layer0_outputs(6072) <= inputs(99);
    layer0_outputs(6073) <= not(inputs(190));
    layer0_outputs(6074) <= not(inputs(123)) or (inputs(251));
    layer0_outputs(6075) <= not(inputs(71)) or (inputs(143));
    layer0_outputs(6076) <= (inputs(118)) xor (inputs(210));
    layer0_outputs(6077) <= (inputs(93)) or (inputs(233));
    layer0_outputs(6078) <= not((inputs(11)) or (inputs(248)));
    layer0_outputs(6079) <= not((inputs(71)) or (inputs(239)));
    layer0_outputs(6080) <= not(inputs(31));
    layer0_outputs(6081) <= (inputs(145)) and (inputs(211));
    layer0_outputs(6082) <= not(inputs(232));
    layer0_outputs(6083) <= not((inputs(9)) and (inputs(26)));
    layer0_outputs(6084) <= not(inputs(197));
    layer0_outputs(6085) <= (inputs(188)) or (inputs(26));
    layer0_outputs(6086) <= not(inputs(120)) or (inputs(2));
    layer0_outputs(6087) <= not((inputs(211)) or (inputs(134)));
    layer0_outputs(6088) <= inputs(14);
    layer0_outputs(6089) <= (inputs(205)) or (inputs(75));
    layer0_outputs(6090) <= not(inputs(240)) or (inputs(184));
    layer0_outputs(6091) <= not(inputs(133));
    layer0_outputs(6092) <= (inputs(73)) and not (inputs(237));
    layer0_outputs(6093) <= inputs(103);
    layer0_outputs(6094) <= (inputs(217)) and not (inputs(123));
    layer0_outputs(6095) <= not((inputs(175)) or (inputs(143)));
    layer0_outputs(6096) <= not((inputs(31)) or (inputs(102)));
    layer0_outputs(6097) <= not(inputs(135));
    layer0_outputs(6098) <= not((inputs(150)) or (inputs(50)));
    layer0_outputs(6099) <= (inputs(87)) xor (inputs(244));
    layer0_outputs(6100) <= inputs(94);
    layer0_outputs(6101) <= (inputs(100)) and not (inputs(48));
    layer0_outputs(6102) <= not(inputs(230)) or (inputs(14));
    layer0_outputs(6103) <= not((inputs(103)) or (inputs(70)));
    layer0_outputs(6104) <= not((inputs(80)) and (inputs(238)));
    layer0_outputs(6105) <= not((inputs(61)) and (inputs(57)));
    layer0_outputs(6106) <= not(inputs(183)) or (inputs(20));
    layer0_outputs(6107) <= not((inputs(204)) or (inputs(194)));
    layer0_outputs(6108) <= not(inputs(142)) or (inputs(142));
    layer0_outputs(6109) <= not((inputs(221)) and (inputs(85)));
    layer0_outputs(6110) <= not((inputs(201)) xor (inputs(226)));
    layer0_outputs(6111) <= not(inputs(57)) or (inputs(49));
    layer0_outputs(6112) <= (inputs(51)) xor (inputs(176));
    layer0_outputs(6113) <= not((inputs(43)) or (inputs(253)));
    layer0_outputs(6114) <= not((inputs(253)) or (inputs(26)));
    layer0_outputs(6115) <= '0';
    layer0_outputs(6116) <= not(inputs(41));
    layer0_outputs(6117) <= not(inputs(62)) or (inputs(206));
    layer0_outputs(6118) <= not(inputs(118)) or (inputs(13));
    layer0_outputs(6119) <= not((inputs(66)) xor (inputs(133)));
    layer0_outputs(6120) <= (inputs(188)) xor (inputs(142));
    layer0_outputs(6121) <= (inputs(102)) and not (inputs(191));
    layer0_outputs(6122) <= not(inputs(164));
    layer0_outputs(6123) <= not((inputs(167)) xor (inputs(54)));
    layer0_outputs(6124) <= (inputs(26)) and not (inputs(87));
    layer0_outputs(6125) <= (inputs(142)) and not (inputs(78));
    layer0_outputs(6126) <= not(inputs(220));
    layer0_outputs(6127) <= (inputs(249)) xor (inputs(44));
    layer0_outputs(6128) <= not((inputs(209)) or (inputs(20)));
    layer0_outputs(6129) <= not(inputs(176));
    layer0_outputs(6130) <= not((inputs(90)) xor (inputs(79)));
    layer0_outputs(6131) <= not(inputs(233)) or (inputs(16));
    layer0_outputs(6132) <= not((inputs(225)) and (inputs(24)));
    layer0_outputs(6133) <= (inputs(153)) and not (inputs(78));
    layer0_outputs(6134) <= (inputs(216)) and not (inputs(87));
    layer0_outputs(6135) <= (inputs(7)) or (inputs(160));
    layer0_outputs(6136) <= not((inputs(184)) xor (inputs(166)));
    layer0_outputs(6137) <= (inputs(46)) and not (inputs(152));
    layer0_outputs(6138) <= (inputs(168)) and not (inputs(107));
    layer0_outputs(6139) <= (inputs(215)) or (inputs(178));
    layer0_outputs(6140) <= (inputs(76)) or (inputs(47));
    layer0_outputs(6141) <= not((inputs(126)) xor (inputs(121)));
    layer0_outputs(6142) <= not(inputs(211)) or (inputs(109));
    layer0_outputs(6143) <= not(inputs(106));
    layer0_outputs(6144) <= not(inputs(44)) or (inputs(243));
    layer0_outputs(6145) <= not(inputs(118)) or (inputs(238));
    layer0_outputs(6146) <= inputs(124);
    layer0_outputs(6147) <= (inputs(19)) or (inputs(241));
    layer0_outputs(6148) <= not((inputs(194)) or (inputs(144)));
    layer0_outputs(6149) <= (inputs(228)) and not (inputs(150));
    layer0_outputs(6150) <= inputs(140);
    layer0_outputs(6151) <= (inputs(131)) and not (inputs(174));
    layer0_outputs(6152) <= not((inputs(189)) or (inputs(108)));
    layer0_outputs(6153) <= not((inputs(8)) or (inputs(201)));
    layer0_outputs(6154) <= not(inputs(181));
    layer0_outputs(6155) <= not(inputs(201));
    layer0_outputs(6156) <= (inputs(252)) or (inputs(19));
    layer0_outputs(6157) <= (inputs(109)) xor (inputs(107));
    layer0_outputs(6158) <= not((inputs(96)) or (inputs(231)));
    layer0_outputs(6159) <= not(inputs(24));
    layer0_outputs(6160) <= (inputs(67)) xor (inputs(21));
    layer0_outputs(6161) <= not(inputs(214));
    layer0_outputs(6162) <= (inputs(121)) and (inputs(108));
    layer0_outputs(6163) <= (inputs(148)) or (inputs(163));
    layer0_outputs(6164) <= (inputs(134)) xor (inputs(118));
    layer0_outputs(6165) <= not((inputs(78)) or (inputs(222)));
    layer0_outputs(6166) <= not((inputs(194)) xor (inputs(39)));
    layer0_outputs(6167) <= (inputs(117)) or (inputs(255));
    layer0_outputs(6168) <= (inputs(141)) and not (inputs(49));
    layer0_outputs(6169) <= (inputs(180)) xor (inputs(236));
    layer0_outputs(6170) <= inputs(162);
    layer0_outputs(6171) <= (inputs(203)) xor (inputs(233));
    layer0_outputs(6172) <= not(inputs(159));
    layer0_outputs(6173) <= not((inputs(84)) or (inputs(128)));
    layer0_outputs(6174) <= not((inputs(74)) or (inputs(176)));
    layer0_outputs(6175) <= not(inputs(75));
    layer0_outputs(6176) <= inputs(146);
    layer0_outputs(6177) <= inputs(149);
    layer0_outputs(6178) <= (inputs(126)) and not (inputs(223));
    layer0_outputs(6179) <= (inputs(239)) xor (inputs(103));
    layer0_outputs(6180) <= not((inputs(128)) or (inputs(207)));
    layer0_outputs(6181) <= (inputs(145)) or (inputs(169));
    layer0_outputs(6182) <= inputs(70);
    layer0_outputs(6183) <= not((inputs(141)) or (inputs(2)));
    layer0_outputs(6184) <= not((inputs(210)) and (inputs(64)));
    layer0_outputs(6185) <= (inputs(212)) and not (inputs(72));
    layer0_outputs(6186) <= '0';
    layer0_outputs(6187) <= not(inputs(231));
    layer0_outputs(6188) <= not(inputs(193));
    layer0_outputs(6189) <= (inputs(170)) and not (inputs(228));
    layer0_outputs(6190) <= not(inputs(163)) or (inputs(113));
    layer0_outputs(6191) <= inputs(179);
    layer0_outputs(6192) <= '0';
    layer0_outputs(6193) <= inputs(112);
    layer0_outputs(6194) <= (inputs(220)) xor (inputs(220));
    layer0_outputs(6195) <= (inputs(165)) xor (inputs(211));
    layer0_outputs(6196) <= (inputs(245)) or (inputs(40));
    layer0_outputs(6197) <= not(inputs(118)) or (inputs(237));
    layer0_outputs(6198) <= not(inputs(146));
    layer0_outputs(6199) <= inputs(157);
    layer0_outputs(6200) <= not((inputs(175)) xor (inputs(26)));
    layer0_outputs(6201) <= not(inputs(103));
    layer0_outputs(6202) <= (inputs(113)) or (inputs(233));
    layer0_outputs(6203) <= inputs(247);
    layer0_outputs(6204) <= not((inputs(46)) xor (inputs(68)));
    layer0_outputs(6205) <= not(inputs(229));
    layer0_outputs(6206) <= (inputs(32)) or (inputs(94));
    layer0_outputs(6207) <= not(inputs(104)) or (inputs(19));
    layer0_outputs(6208) <= not(inputs(212));
    layer0_outputs(6209) <= not(inputs(213));
    layer0_outputs(6210) <= '1';
    layer0_outputs(6211) <= inputs(109);
    layer0_outputs(6212) <= not((inputs(114)) or (inputs(138)));
    layer0_outputs(6213) <= not(inputs(12)) or (inputs(206));
    layer0_outputs(6214) <= not(inputs(226)) or (inputs(64));
    layer0_outputs(6215) <= inputs(58);
    layer0_outputs(6216) <= not((inputs(61)) or (inputs(36)));
    layer0_outputs(6217) <= (inputs(174)) or (inputs(206));
    layer0_outputs(6218) <= (inputs(155)) xor (inputs(144));
    layer0_outputs(6219) <= (inputs(8)) or (inputs(1));
    layer0_outputs(6220) <= not(inputs(194));
    layer0_outputs(6221) <= (inputs(165)) or (inputs(237));
    layer0_outputs(6222) <= not(inputs(140)) or (inputs(247));
    layer0_outputs(6223) <= not((inputs(81)) xor (inputs(20)));
    layer0_outputs(6224) <= inputs(214);
    layer0_outputs(6225) <= not(inputs(202));
    layer0_outputs(6226) <= (inputs(32)) xor (inputs(58));
    layer0_outputs(6227) <= inputs(74);
    layer0_outputs(6228) <= not(inputs(201)) or (inputs(109));
    layer0_outputs(6229) <= not((inputs(234)) or (inputs(208)));
    layer0_outputs(6230) <= not(inputs(48));
    layer0_outputs(6231) <= (inputs(185)) xor (inputs(161));
    layer0_outputs(6232) <= (inputs(124)) xor (inputs(132));
    layer0_outputs(6233) <= inputs(5);
    layer0_outputs(6234) <= not((inputs(187)) xor (inputs(36)));
    layer0_outputs(6235) <= (inputs(45)) or (inputs(63));
    layer0_outputs(6236) <= not((inputs(154)) and (inputs(140)));
    layer0_outputs(6237) <= (inputs(243)) and not (inputs(255));
    layer0_outputs(6238) <= (inputs(154)) and not (inputs(81));
    layer0_outputs(6239) <= not(inputs(187));
    layer0_outputs(6240) <= not(inputs(197));
    layer0_outputs(6241) <= not(inputs(128));
    layer0_outputs(6242) <= not(inputs(41));
    layer0_outputs(6243) <= (inputs(45)) or (inputs(44));
    layer0_outputs(6244) <= not(inputs(250));
    layer0_outputs(6245) <= (inputs(57)) and not (inputs(16));
    layer0_outputs(6246) <= (inputs(243)) xor (inputs(235));
    layer0_outputs(6247) <= '1';
    layer0_outputs(6248) <= inputs(197);
    layer0_outputs(6249) <= (inputs(166)) or (inputs(236));
    layer0_outputs(6250) <= (inputs(32)) or (inputs(240));
    layer0_outputs(6251) <= (inputs(210)) and (inputs(146));
    layer0_outputs(6252) <= (inputs(127)) or (inputs(60));
    layer0_outputs(6253) <= not((inputs(228)) or (inputs(146)));
    layer0_outputs(6254) <= (inputs(194)) or (inputs(116));
    layer0_outputs(6255) <= (inputs(53)) and not (inputs(189));
    layer0_outputs(6256) <= not((inputs(248)) xor (inputs(114)));
    layer0_outputs(6257) <= not((inputs(96)) or (inputs(230)));
    layer0_outputs(6258) <= (inputs(72)) and not (inputs(46));
    layer0_outputs(6259) <= (inputs(198)) xor (inputs(249));
    layer0_outputs(6260) <= not(inputs(149));
    layer0_outputs(6261) <= inputs(137);
    layer0_outputs(6262) <= (inputs(104)) or (inputs(1));
    layer0_outputs(6263) <= not(inputs(245));
    layer0_outputs(6264) <= not((inputs(130)) xor (inputs(150)));
    layer0_outputs(6265) <= inputs(164);
    layer0_outputs(6266) <= (inputs(135)) and not (inputs(56));
    layer0_outputs(6267) <= (inputs(151)) or (inputs(250));
    layer0_outputs(6268) <= not(inputs(119));
    layer0_outputs(6269) <= not(inputs(83)) or (inputs(142));
    layer0_outputs(6270) <= (inputs(200)) or (inputs(145));
    layer0_outputs(6271) <= (inputs(167)) and (inputs(181));
    layer0_outputs(6272) <= (inputs(212)) or (inputs(234));
    layer0_outputs(6273) <= not(inputs(164));
    layer0_outputs(6274) <= not((inputs(108)) or (inputs(132)));
    layer0_outputs(6275) <= not(inputs(148)) or (inputs(2));
    layer0_outputs(6276) <= not(inputs(184));
    layer0_outputs(6277) <= (inputs(58)) xor (inputs(140));
    layer0_outputs(6278) <= (inputs(76)) xor (inputs(17));
    layer0_outputs(6279) <= inputs(247);
    layer0_outputs(6280) <= not(inputs(204));
    layer0_outputs(6281) <= inputs(150);
    layer0_outputs(6282) <= (inputs(39)) and not (inputs(188));
    layer0_outputs(6283) <= not((inputs(131)) or (inputs(9)));
    layer0_outputs(6284) <= (inputs(171)) or (inputs(159));
    layer0_outputs(6285) <= not(inputs(130));
    layer0_outputs(6286) <= not(inputs(152));
    layer0_outputs(6287) <= inputs(180);
    layer0_outputs(6288) <= not(inputs(75)) or (inputs(197));
    layer0_outputs(6289) <= not((inputs(27)) xor (inputs(232)));
    layer0_outputs(6290) <= (inputs(84)) and not (inputs(94));
    layer0_outputs(6291) <= not((inputs(183)) or (inputs(177)));
    layer0_outputs(6292) <= inputs(211);
    layer0_outputs(6293) <= (inputs(214)) or (inputs(51));
    layer0_outputs(6294) <= not((inputs(119)) xor (inputs(252)));
    layer0_outputs(6295) <= not(inputs(169));
    layer0_outputs(6296) <= not((inputs(193)) xor (inputs(221)));
    layer0_outputs(6297) <= (inputs(174)) and not (inputs(111));
    layer0_outputs(6298) <= not(inputs(157));
    layer0_outputs(6299) <= (inputs(191)) xor (inputs(123));
    layer0_outputs(6300) <= not(inputs(75));
    layer0_outputs(6301) <= not((inputs(205)) xor (inputs(145)));
    layer0_outputs(6302) <= (inputs(34)) or (inputs(25));
    layer0_outputs(6303) <= not(inputs(112));
    layer0_outputs(6304) <= (inputs(189)) and not (inputs(18));
    layer0_outputs(6305) <= (inputs(153)) xor (inputs(192));
    layer0_outputs(6306) <= (inputs(134)) xor (inputs(168));
    layer0_outputs(6307) <= inputs(214);
    layer0_outputs(6308) <= (inputs(151)) or (inputs(90));
    layer0_outputs(6309) <= (inputs(253)) or (inputs(136));
    layer0_outputs(6310) <= not((inputs(18)) or (inputs(230)));
    layer0_outputs(6311) <= not((inputs(150)) xor (inputs(163)));
    layer0_outputs(6312) <= not(inputs(41)) or (inputs(252));
    layer0_outputs(6313) <= inputs(67);
    layer0_outputs(6314) <= not((inputs(177)) or (inputs(197)));
    layer0_outputs(6315) <= inputs(152);
    layer0_outputs(6316) <= (inputs(48)) xor (inputs(52));
    layer0_outputs(6317) <= inputs(167);
    layer0_outputs(6318) <= (inputs(166)) and (inputs(231));
    layer0_outputs(6319) <= (inputs(212)) and not (inputs(58));
    layer0_outputs(6320) <= inputs(105);
    layer0_outputs(6321) <= not((inputs(65)) or (inputs(50)));
    layer0_outputs(6322) <= (inputs(74)) and not (inputs(127));
    layer0_outputs(6323) <= not(inputs(183));
    layer0_outputs(6324) <= not((inputs(114)) and (inputs(137)));
    layer0_outputs(6325) <= inputs(226);
    layer0_outputs(6326) <= inputs(169);
    layer0_outputs(6327) <= not(inputs(245)) or (inputs(90));
    layer0_outputs(6328) <= not(inputs(214)) or (inputs(167));
    layer0_outputs(6329) <= inputs(69);
    layer0_outputs(6330) <= inputs(66);
    layer0_outputs(6331) <= (inputs(98)) or (inputs(144));
    layer0_outputs(6332) <= (inputs(95)) and (inputs(254));
    layer0_outputs(6333) <= (inputs(179)) and not (inputs(29));
    layer0_outputs(6334) <= not(inputs(212));
    layer0_outputs(6335) <= not((inputs(205)) xor (inputs(155)));
    layer0_outputs(6336) <= (inputs(29)) xor (inputs(45));
    layer0_outputs(6337) <= not(inputs(221));
    layer0_outputs(6338) <= not((inputs(37)) or (inputs(141)));
    layer0_outputs(6339) <= not((inputs(145)) or (inputs(144)));
    layer0_outputs(6340) <= not((inputs(100)) xor (inputs(192)));
    layer0_outputs(6341) <= not((inputs(31)) or (inputs(85)));
    layer0_outputs(6342) <= not((inputs(201)) or (inputs(2)));
    layer0_outputs(6343) <= not((inputs(246)) or (inputs(233)));
    layer0_outputs(6344) <= not(inputs(80)) or (inputs(238));
    layer0_outputs(6345) <= inputs(56);
    layer0_outputs(6346) <= not(inputs(193)) or (inputs(31));
    layer0_outputs(6347) <= not((inputs(208)) xor (inputs(174)));
    layer0_outputs(6348) <= (inputs(21)) and not (inputs(187));
    layer0_outputs(6349) <= not(inputs(29));
    layer0_outputs(6350) <= not(inputs(0)) or (inputs(195));
    layer0_outputs(6351) <= not((inputs(52)) xor (inputs(38)));
    layer0_outputs(6352) <= (inputs(73)) xor (inputs(55));
    layer0_outputs(6353) <= not((inputs(161)) or (inputs(167)));
    layer0_outputs(6354) <= inputs(69);
    layer0_outputs(6355) <= inputs(15);
    layer0_outputs(6356) <= not(inputs(40)) or (inputs(127));
    layer0_outputs(6357) <= not(inputs(67));
    layer0_outputs(6358) <= not(inputs(62));
    layer0_outputs(6359) <= inputs(63);
    layer0_outputs(6360) <= not(inputs(93));
    layer0_outputs(6361) <= (inputs(140)) or (inputs(248));
    layer0_outputs(6362) <= not(inputs(1)) or (inputs(1));
    layer0_outputs(6363) <= inputs(135);
    layer0_outputs(6364) <= (inputs(148)) and not (inputs(92));
    layer0_outputs(6365) <= not(inputs(133));
    layer0_outputs(6366) <= not(inputs(228));
    layer0_outputs(6367) <= not((inputs(159)) or (inputs(188)));
    layer0_outputs(6368) <= inputs(165);
    layer0_outputs(6369) <= inputs(246);
    layer0_outputs(6370) <= not(inputs(22)) or (inputs(95));
    layer0_outputs(6371) <= (inputs(241)) xor (inputs(232));
    layer0_outputs(6372) <= not((inputs(232)) xor (inputs(75)));
    layer0_outputs(6373) <= not(inputs(32));
    layer0_outputs(6374) <= '1';
    layer0_outputs(6375) <= not(inputs(101));
    layer0_outputs(6376) <= inputs(56);
    layer0_outputs(6377) <= not(inputs(56)) or (inputs(14));
    layer0_outputs(6378) <= not((inputs(39)) or (inputs(251)));
    layer0_outputs(6379) <= (inputs(232)) or (inputs(107));
    layer0_outputs(6380) <= not((inputs(94)) or (inputs(78)));
    layer0_outputs(6381) <= (inputs(104)) xor (inputs(159));
    layer0_outputs(6382) <= (inputs(106)) xor (inputs(7));
    layer0_outputs(6383) <= inputs(141);
    layer0_outputs(6384) <= (inputs(228)) and not (inputs(28));
    layer0_outputs(6385) <= (inputs(66)) and not (inputs(244));
    layer0_outputs(6386) <= not((inputs(188)) and (inputs(54)));
    layer0_outputs(6387) <= inputs(82);
    layer0_outputs(6388) <= (inputs(134)) and not (inputs(176));
    layer0_outputs(6389) <= not((inputs(115)) xor (inputs(86)));
    layer0_outputs(6390) <= (inputs(113)) or (inputs(115));
    layer0_outputs(6391) <= (inputs(168)) or (inputs(142));
    layer0_outputs(6392) <= (inputs(95)) and not (inputs(127));
    layer0_outputs(6393) <= not((inputs(66)) or (inputs(174)));
    layer0_outputs(6394) <= not((inputs(27)) xor (inputs(6)));
    layer0_outputs(6395) <= not(inputs(213));
    layer0_outputs(6396) <= not((inputs(12)) or (inputs(142)));
    layer0_outputs(6397) <= inputs(109);
    layer0_outputs(6398) <= not(inputs(235)) or (inputs(151));
    layer0_outputs(6399) <= inputs(183);
    layer0_outputs(6400) <= not(inputs(202));
    layer0_outputs(6401) <= not(inputs(200)) or (inputs(140));
    layer0_outputs(6402) <= (inputs(22)) or (inputs(24));
    layer0_outputs(6403) <= inputs(246);
    layer0_outputs(6404) <= (inputs(239)) and not (inputs(46));
    layer0_outputs(6405) <= (inputs(131)) or (inputs(39));
    layer0_outputs(6406) <= not(inputs(26)) or (inputs(35));
    layer0_outputs(6407) <= not((inputs(91)) xor (inputs(189)));
    layer0_outputs(6408) <= (inputs(177)) or (inputs(181));
    layer0_outputs(6409) <= not(inputs(83));
    layer0_outputs(6410) <= (inputs(54)) and not (inputs(248));
    layer0_outputs(6411) <= not((inputs(76)) xor (inputs(47)));
    layer0_outputs(6412) <= not((inputs(185)) xor (inputs(83)));
    layer0_outputs(6413) <= (inputs(113)) and not (inputs(254));
    layer0_outputs(6414) <= inputs(195);
    layer0_outputs(6415) <= (inputs(239)) or (inputs(240));
    layer0_outputs(6416) <= (inputs(239)) and not (inputs(160));
    layer0_outputs(6417) <= not(inputs(210)) or (inputs(201));
    layer0_outputs(6418) <= (inputs(185)) xor (inputs(224));
    layer0_outputs(6419) <= not((inputs(95)) xor (inputs(255)));
    layer0_outputs(6420) <= inputs(132);
    layer0_outputs(6421) <= not(inputs(220));
    layer0_outputs(6422) <= not(inputs(25));
    layer0_outputs(6423) <= not((inputs(180)) or (inputs(59)));
    layer0_outputs(6424) <= not(inputs(155));
    layer0_outputs(6425) <= not(inputs(100));
    layer0_outputs(6426) <= (inputs(147)) or (inputs(8));
    layer0_outputs(6427) <= (inputs(254)) and (inputs(233));
    layer0_outputs(6428) <= inputs(197);
    layer0_outputs(6429) <= inputs(193);
    layer0_outputs(6430) <= not((inputs(210)) xor (inputs(61)));
    layer0_outputs(6431) <= inputs(158);
    layer0_outputs(6432) <= not((inputs(67)) xor (inputs(39)));
    layer0_outputs(6433) <= not(inputs(146));
    layer0_outputs(6434) <= (inputs(245)) and not (inputs(152));
    layer0_outputs(6435) <= not(inputs(12)) or (inputs(252));
    layer0_outputs(6436) <= '0';
    layer0_outputs(6437) <= inputs(115);
    layer0_outputs(6438) <= not((inputs(245)) or (inputs(41)));
    layer0_outputs(6439) <= (inputs(184)) or (inputs(248));
    layer0_outputs(6440) <= (inputs(52)) or (inputs(21));
    layer0_outputs(6441) <= not(inputs(178));
    layer0_outputs(6442) <= inputs(89);
    layer0_outputs(6443) <= inputs(177);
    layer0_outputs(6444) <= not(inputs(114));
    layer0_outputs(6445) <= (inputs(171)) or (inputs(51));
    layer0_outputs(6446) <= (inputs(54)) and not (inputs(0));
    layer0_outputs(6447) <= (inputs(214)) and not (inputs(119));
    layer0_outputs(6448) <= (inputs(13)) and (inputs(101));
    layer0_outputs(6449) <= (inputs(160)) and (inputs(81));
    layer0_outputs(6450) <= inputs(141);
    layer0_outputs(6451) <= not((inputs(187)) or (inputs(35)));
    layer0_outputs(6452) <= (inputs(73)) xor (inputs(201));
    layer0_outputs(6453) <= not((inputs(224)) or (inputs(75)));
    layer0_outputs(6454) <= inputs(167);
    layer0_outputs(6455) <= (inputs(220)) or (inputs(176));
    layer0_outputs(6456) <= (inputs(215)) or (inputs(207));
    layer0_outputs(6457) <= inputs(238);
    layer0_outputs(6458) <= inputs(123);
    layer0_outputs(6459) <= not(inputs(99));
    layer0_outputs(6460) <= not(inputs(136));
    layer0_outputs(6461) <= inputs(97);
    layer0_outputs(6462) <= not(inputs(12)) or (inputs(240));
    layer0_outputs(6463) <= inputs(104);
    layer0_outputs(6464) <= not(inputs(139)) or (inputs(22));
    layer0_outputs(6465) <= (inputs(103)) or (inputs(246));
    layer0_outputs(6466) <= not(inputs(137)) or (inputs(49));
    layer0_outputs(6467) <= not(inputs(164));
    layer0_outputs(6468) <= (inputs(29)) and not (inputs(166));
    layer0_outputs(6469) <= inputs(102);
    layer0_outputs(6470) <= (inputs(246)) and not (inputs(1));
    layer0_outputs(6471) <= not(inputs(27)) or (inputs(134));
    layer0_outputs(6472) <= inputs(45);
    layer0_outputs(6473) <= not(inputs(117));
    layer0_outputs(6474) <= (inputs(151)) and not (inputs(40));
    layer0_outputs(6475) <= not((inputs(105)) and (inputs(36)));
    layer0_outputs(6476) <= inputs(59);
    layer0_outputs(6477) <= (inputs(139)) xor (inputs(133));
    layer0_outputs(6478) <= not(inputs(137));
    layer0_outputs(6479) <= not(inputs(210)) or (inputs(28));
    layer0_outputs(6480) <= (inputs(57)) and not (inputs(120));
    layer0_outputs(6481) <= '1';
    layer0_outputs(6482) <= (inputs(11)) xor (inputs(108));
    layer0_outputs(6483) <= inputs(84);
    layer0_outputs(6484) <= (inputs(239)) xor (inputs(207));
    layer0_outputs(6485) <= (inputs(22)) and not (inputs(114));
    layer0_outputs(6486) <= (inputs(22)) xor (inputs(119));
    layer0_outputs(6487) <= (inputs(97)) or (inputs(108));
    layer0_outputs(6488) <= (inputs(190)) or (inputs(13));
    layer0_outputs(6489) <= inputs(214);
    layer0_outputs(6490) <= (inputs(102)) or (inputs(203));
    layer0_outputs(6491) <= not((inputs(159)) or (inputs(92)));
    layer0_outputs(6492) <= not(inputs(242));
    layer0_outputs(6493) <= inputs(150);
    layer0_outputs(6494) <= (inputs(76)) xor (inputs(78));
    layer0_outputs(6495) <= (inputs(126)) and not (inputs(56));
    layer0_outputs(6496) <= not((inputs(234)) or (inputs(9)));
    layer0_outputs(6497) <= inputs(65);
    layer0_outputs(6498) <= (inputs(84)) and not (inputs(93));
    layer0_outputs(6499) <= (inputs(244)) and not (inputs(112));
    layer0_outputs(6500) <= not((inputs(174)) or (inputs(250)));
    layer0_outputs(6501) <= (inputs(99)) xor (inputs(118));
    layer0_outputs(6502) <= not((inputs(205)) or (inputs(91)));
    layer0_outputs(6503) <= not(inputs(185));
    layer0_outputs(6504) <= not(inputs(59)) or (inputs(236));
    layer0_outputs(6505) <= (inputs(172)) xor (inputs(79));
    layer0_outputs(6506) <= not(inputs(233)) or (inputs(2));
    layer0_outputs(6507) <= not(inputs(231)) or (inputs(41));
    layer0_outputs(6508) <= inputs(101);
    layer0_outputs(6509) <= not(inputs(157)) or (inputs(80));
    layer0_outputs(6510) <= inputs(135);
    layer0_outputs(6511) <= not((inputs(216)) or (inputs(200)));
    layer0_outputs(6512) <= (inputs(207)) xor (inputs(87));
    layer0_outputs(6513) <= (inputs(36)) and not (inputs(188));
    layer0_outputs(6514) <= not(inputs(163));
    layer0_outputs(6515) <= not(inputs(72));
    layer0_outputs(6516) <= inputs(162);
    layer0_outputs(6517) <= not(inputs(209)) or (inputs(159));
    layer0_outputs(6518) <= not((inputs(248)) or (inputs(211)));
    layer0_outputs(6519) <= not((inputs(56)) or (inputs(231)));
    layer0_outputs(6520) <= not(inputs(149));
    layer0_outputs(6521) <= not(inputs(99));
    layer0_outputs(6522) <= inputs(160);
    layer0_outputs(6523) <= not((inputs(92)) or (inputs(100)));
    layer0_outputs(6524) <= (inputs(63)) or (inputs(9));
    layer0_outputs(6525) <= (inputs(6)) xor (inputs(52));
    layer0_outputs(6526) <= inputs(21);
    layer0_outputs(6527) <= not((inputs(94)) xor (inputs(181)));
    layer0_outputs(6528) <= inputs(65);
    layer0_outputs(6529) <= not((inputs(244)) xor (inputs(150)));
    layer0_outputs(6530) <= not(inputs(97));
    layer0_outputs(6531) <= (inputs(80)) xor (inputs(43));
    layer0_outputs(6532) <= not(inputs(215)) or (inputs(253));
    layer0_outputs(6533) <= (inputs(57)) or (inputs(212));
    layer0_outputs(6534) <= inputs(57);
    layer0_outputs(6535) <= not(inputs(74));
    layer0_outputs(6536) <= not(inputs(220)) or (inputs(72));
    layer0_outputs(6537) <= inputs(236);
    layer0_outputs(6538) <= '1';
    layer0_outputs(6539) <= not(inputs(149));
    layer0_outputs(6540) <= not(inputs(199)) or (inputs(190));
    layer0_outputs(6541) <= not((inputs(80)) or (inputs(54)));
    layer0_outputs(6542) <= not(inputs(249));
    layer0_outputs(6543) <= (inputs(103)) xor (inputs(162));
    layer0_outputs(6544) <= not(inputs(204));
    layer0_outputs(6545) <= (inputs(121)) and not (inputs(196));
    layer0_outputs(6546) <= not(inputs(216)) or (inputs(64));
    layer0_outputs(6547) <= not(inputs(116));
    layer0_outputs(6548) <= (inputs(101)) xor (inputs(66));
    layer0_outputs(6549) <= not((inputs(25)) xor (inputs(76)));
    layer0_outputs(6550) <= (inputs(247)) xor (inputs(207));
    layer0_outputs(6551) <= inputs(195);
    layer0_outputs(6552) <= not((inputs(0)) xor (inputs(204)));
    layer0_outputs(6553) <= not(inputs(134));
    layer0_outputs(6554) <= not((inputs(189)) or (inputs(204)));
    layer0_outputs(6555) <= not(inputs(133)) or (inputs(36));
    layer0_outputs(6556) <= (inputs(176)) or (inputs(118));
    layer0_outputs(6557) <= inputs(251);
    layer0_outputs(6558) <= (inputs(45)) or (inputs(58));
    layer0_outputs(6559) <= (inputs(71)) or (inputs(108));
    layer0_outputs(6560) <= not((inputs(71)) xor (inputs(64)));
    layer0_outputs(6561) <= (inputs(4)) or (inputs(231));
    layer0_outputs(6562) <= not(inputs(231)) or (inputs(125));
    layer0_outputs(6563) <= (inputs(198)) xor (inputs(199));
    layer0_outputs(6564) <= (inputs(167)) and not (inputs(31));
    layer0_outputs(6565) <= (inputs(119)) or (inputs(243));
    layer0_outputs(6566) <= not(inputs(232)) or (inputs(15));
    layer0_outputs(6567) <= '1';
    layer0_outputs(6568) <= not((inputs(138)) xor (inputs(120)));
    layer0_outputs(6569) <= not((inputs(247)) xor (inputs(169)));
    layer0_outputs(6570) <= not(inputs(153));
    layer0_outputs(6571) <= (inputs(108)) and not (inputs(32));
    layer0_outputs(6572) <= not(inputs(86));
    layer0_outputs(6573) <= not((inputs(209)) xor (inputs(144)));
    layer0_outputs(6574) <= not((inputs(157)) or (inputs(250)));
    layer0_outputs(6575) <= (inputs(109)) and not (inputs(47));
    layer0_outputs(6576) <= not(inputs(63));
    layer0_outputs(6577) <= not(inputs(195)) or (inputs(122));
    layer0_outputs(6578) <= (inputs(22)) xor (inputs(64));
    layer0_outputs(6579) <= (inputs(244)) and not (inputs(66));
    layer0_outputs(6580) <= not((inputs(137)) xor (inputs(108)));
    layer0_outputs(6581) <= (inputs(162)) and not (inputs(151));
    layer0_outputs(6582) <= not((inputs(68)) or (inputs(229)));
    layer0_outputs(6583) <= (inputs(76)) xor (inputs(73));
    layer0_outputs(6584) <= not(inputs(39)) or (inputs(3));
    layer0_outputs(6585) <= inputs(151);
    layer0_outputs(6586) <= (inputs(122)) and not (inputs(240));
    layer0_outputs(6587) <= (inputs(238)) xor (inputs(36));
    layer0_outputs(6588) <= inputs(42);
    layer0_outputs(6589) <= not(inputs(20)) or (inputs(173));
    layer0_outputs(6590) <= (inputs(36)) or (inputs(253));
    layer0_outputs(6591) <= inputs(138);
    layer0_outputs(6592) <= not((inputs(129)) or (inputs(12)));
    layer0_outputs(6593) <= not((inputs(36)) xor (inputs(178)));
    layer0_outputs(6594) <= inputs(136);
    layer0_outputs(6595) <= not(inputs(107)) or (inputs(81));
    layer0_outputs(6596) <= '0';
    layer0_outputs(6597) <= '0';
    layer0_outputs(6598) <= not(inputs(247)) or (inputs(147));
    layer0_outputs(6599) <= not(inputs(41)) or (inputs(235));
    layer0_outputs(6600) <= not((inputs(168)) and (inputs(213)));
    layer0_outputs(6601) <= not((inputs(110)) or (inputs(110)));
    layer0_outputs(6602) <= (inputs(250)) xor (inputs(164));
    layer0_outputs(6603) <= not(inputs(147));
    layer0_outputs(6604) <= (inputs(253)) xor (inputs(143));
    layer0_outputs(6605) <= (inputs(188)) or (inputs(204));
    layer0_outputs(6606) <= not(inputs(237));
    layer0_outputs(6607) <= (inputs(122)) xor (inputs(237));
    layer0_outputs(6608) <= (inputs(123)) xor (inputs(12));
    layer0_outputs(6609) <= not((inputs(155)) xor (inputs(117)));
    layer0_outputs(6610) <= (inputs(72)) or (inputs(136));
    layer0_outputs(6611) <= inputs(255);
    layer0_outputs(6612) <= not(inputs(140));
    layer0_outputs(6613) <= (inputs(230)) xor (inputs(40));
    layer0_outputs(6614) <= inputs(163);
    layer0_outputs(6615) <= inputs(134);
    layer0_outputs(6616) <= not(inputs(253)) or (inputs(34));
    layer0_outputs(6617) <= (inputs(104)) xor (inputs(68));
    layer0_outputs(6618) <= not(inputs(140)) or (inputs(34));
    layer0_outputs(6619) <= (inputs(90)) xor (inputs(137));
    layer0_outputs(6620) <= not((inputs(35)) xor (inputs(154)));
    layer0_outputs(6621) <= inputs(179);
    layer0_outputs(6622) <= not(inputs(90));
    layer0_outputs(6623) <= not((inputs(7)) xor (inputs(76)));
    layer0_outputs(6624) <= (inputs(69)) or (inputs(155));
    layer0_outputs(6625) <= not(inputs(88));
    layer0_outputs(6626) <= not((inputs(189)) or (inputs(88)));
    layer0_outputs(6627) <= inputs(182);
    layer0_outputs(6628) <= inputs(228);
    layer0_outputs(6629) <= inputs(8);
    layer0_outputs(6630) <= not((inputs(116)) and (inputs(67)));
    layer0_outputs(6631) <= not(inputs(198));
    layer0_outputs(6632) <= not(inputs(196));
    layer0_outputs(6633) <= (inputs(86)) and not (inputs(144));
    layer0_outputs(6634) <= not(inputs(83));
    layer0_outputs(6635) <= not(inputs(212));
    layer0_outputs(6636) <= not(inputs(230)) or (inputs(254));
    layer0_outputs(6637) <= not(inputs(139)) or (inputs(49));
    layer0_outputs(6638) <= (inputs(140)) and not (inputs(185));
    layer0_outputs(6639) <= (inputs(14)) or (inputs(143));
    layer0_outputs(6640) <= not((inputs(234)) or (inputs(191)));
    layer0_outputs(6641) <= not(inputs(135)) or (inputs(144));
    layer0_outputs(6642) <= inputs(225);
    layer0_outputs(6643) <= (inputs(101)) xor (inputs(128));
    layer0_outputs(6644) <= inputs(131);
    layer0_outputs(6645) <= (inputs(6)) or (inputs(215));
    layer0_outputs(6646) <= not(inputs(133)) or (inputs(6));
    layer0_outputs(6647) <= (inputs(158)) or (inputs(67));
    layer0_outputs(6648) <= (inputs(202)) and (inputs(215));
    layer0_outputs(6649) <= not(inputs(83)) or (inputs(23));
    layer0_outputs(6650) <= not((inputs(246)) or (inputs(106)));
    layer0_outputs(6651) <= not(inputs(58));
    layer0_outputs(6652) <= (inputs(94)) and not (inputs(65));
    layer0_outputs(6653) <= (inputs(102)) xor (inputs(241));
    layer0_outputs(6654) <= (inputs(220)) or (inputs(32));
    layer0_outputs(6655) <= not(inputs(229));
    layer0_outputs(6656) <= (inputs(90)) and (inputs(88));
    layer0_outputs(6657) <= inputs(173);
    layer0_outputs(6658) <= not((inputs(164)) or (inputs(85)));
    layer0_outputs(6659) <= not(inputs(25)) or (inputs(222));
    layer0_outputs(6660) <= (inputs(7)) and not (inputs(126));
    layer0_outputs(6661) <= not(inputs(190));
    layer0_outputs(6662) <= (inputs(69)) or (inputs(100));
    layer0_outputs(6663) <= (inputs(108)) xor (inputs(178));
    layer0_outputs(6664) <= inputs(26);
    layer0_outputs(6665) <= not((inputs(136)) xor (inputs(147)));
    layer0_outputs(6666) <= (inputs(63)) or (inputs(93));
    layer0_outputs(6667) <= (inputs(13)) and not (inputs(226));
    layer0_outputs(6668) <= not((inputs(92)) xor (inputs(30)));
    layer0_outputs(6669) <= (inputs(152)) xor (inputs(186));
    layer0_outputs(6670) <= (inputs(168)) and (inputs(197));
    layer0_outputs(6671) <= not((inputs(29)) and (inputs(235)));
    layer0_outputs(6672) <= '0';
    layer0_outputs(6673) <= not((inputs(60)) or (inputs(95)));
    layer0_outputs(6674) <= not((inputs(123)) xor (inputs(173)));
    layer0_outputs(6675) <= inputs(212);
    layer0_outputs(6676) <= (inputs(58)) or (inputs(4));
    layer0_outputs(6677) <= not(inputs(165)) or (inputs(49));
    layer0_outputs(6678) <= not((inputs(52)) or (inputs(77)));
    layer0_outputs(6679) <= not((inputs(50)) xor (inputs(131)));
    layer0_outputs(6680) <= not((inputs(152)) xor (inputs(129)));
    layer0_outputs(6681) <= not(inputs(61));
    layer0_outputs(6682) <= (inputs(80)) or (inputs(118));
    layer0_outputs(6683) <= not((inputs(168)) or (inputs(125)));
    layer0_outputs(6684) <= not(inputs(59)) or (inputs(47));
    layer0_outputs(6685) <= (inputs(147)) xor (inputs(55));
    layer0_outputs(6686) <= (inputs(203)) xor (inputs(67));
    layer0_outputs(6687) <= (inputs(34)) xor (inputs(208));
    layer0_outputs(6688) <= not(inputs(219));
    layer0_outputs(6689) <= not(inputs(75));
    layer0_outputs(6690) <= (inputs(111)) xor (inputs(62));
    layer0_outputs(6691) <= inputs(56);
    layer0_outputs(6692) <= not((inputs(42)) xor (inputs(191)));
    layer0_outputs(6693) <= inputs(52);
    layer0_outputs(6694) <= not((inputs(223)) xor (inputs(172)));
    layer0_outputs(6695) <= not(inputs(23));
    layer0_outputs(6696) <= (inputs(58)) xor (inputs(212));
    layer0_outputs(6697) <= not(inputs(254));
    layer0_outputs(6698) <= (inputs(137)) and not (inputs(188));
    layer0_outputs(6699) <= not(inputs(228)) or (inputs(129));
    layer0_outputs(6700) <= not((inputs(116)) or (inputs(49)));
    layer0_outputs(6701) <= not((inputs(115)) or (inputs(50)));
    layer0_outputs(6702) <= (inputs(178)) and not (inputs(180));
    layer0_outputs(6703) <= (inputs(35)) xor (inputs(93));
    layer0_outputs(6704) <= not(inputs(227));
    layer0_outputs(6705) <= (inputs(223)) or (inputs(22));
    layer0_outputs(6706) <= (inputs(181)) and not (inputs(79));
    layer0_outputs(6707) <= (inputs(217)) or (inputs(216));
    layer0_outputs(6708) <= (inputs(101)) or (inputs(146));
    layer0_outputs(6709) <= (inputs(134)) or (inputs(98));
    layer0_outputs(6710) <= not((inputs(168)) xor (inputs(134)));
    layer0_outputs(6711) <= not((inputs(113)) and (inputs(144)));
    layer0_outputs(6712) <= not((inputs(156)) or (inputs(38)));
    layer0_outputs(6713) <= not((inputs(18)) xor (inputs(198)));
    layer0_outputs(6714) <= inputs(20);
    layer0_outputs(6715) <= (inputs(249)) or (inputs(209));
    layer0_outputs(6716) <= inputs(232);
    layer0_outputs(6717) <= not(inputs(55));
    layer0_outputs(6718) <= not((inputs(222)) or (inputs(121)));
    layer0_outputs(6719) <= (inputs(69)) or (inputs(50));
    layer0_outputs(6720) <= (inputs(182)) and not (inputs(218));
    layer0_outputs(6721) <= (inputs(42)) and not (inputs(102));
    layer0_outputs(6722) <= not((inputs(185)) xor (inputs(182)));
    layer0_outputs(6723) <= not((inputs(245)) or (inputs(196)));
    layer0_outputs(6724) <= inputs(228);
    layer0_outputs(6725) <= (inputs(127)) and not (inputs(190));
    layer0_outputs(6726) <= inputs(67);
    layer0_outputs(6727) <= inputs(233);
    layer0_outputs(6728) <= not(inputs(190)) or (inputs(223));
    layer0_outputs(6729) <= not(inputs(248));
    layer0_outputs(6730) <= (inputs(23)) and not (inputs(188));
    layer0_outputs(6731) <= inputs(142);
    layer0_outputs(6732) <= not(inputs(123));
    layer0_outputs(6733) <= not((inputs(212)) xor (inputs(178)));
    layer0_outputs(6734) <= not(inputs(180));
    layer0_outputs(6735) <= not(inputs(120)) or (inputs(179));
    layer0_outputs(6736) <= (inputs(137)) or (inputs(143));
    layer0_outputs(6737) <= not((inputs(107)) xor (inputs(114)));
    layer0_outputs(6738) <= not((inputs(34)) or (inputs(151)));
    layer0_outputs(6739) <= (inputs(24)) xor (inputs(69));
    layer0_outputs(6740) <= not((inputs(231)) xor (inputs(146)));
    layer0_outputs(6741) <= inputs(95);
    layer0_outputs(6742) <= (inputs(138)) xor (inputs(190));
    layer0_outputs(6743) <= inputs(227);
    layer0_outputs(6744) <= inputs(37);
    layer0_outputs(6745) <= (inputs(210)) and not (inputs(144));
    layer0_outputs(6746) <= not(inputs(68)) or (inputs(161));
    layer0_outputs(6747) <= (inputs(124)) or (inputs(53));
    layer0_outputs(6748) <= not(inputs(22));
    layer0_outputs(6749) <= not((inputs(32)) or (inputs(27)));
    layer0_outputs(6750) <= inputs(90);
    layer0_outputs(6751) <= (inputs(232)) and not (inputs(16));
    layer0_outputs(6752) <= (inputs(43)) and (inputs(92));
    layer0_outputs(6753) <= (inputs(4)) or (inputs(154));
    layer0_outputs(6754) <= (inputs(11)) and not (inputs(155));
    layer0_outputs(6755) <= not(inputs(99));
    layer0_outputs(6756) <= inputs(108);
    layer0_outputs(6757) <= not(inputs(55)) or (inputs(92));
    layer0_outputs(6758) <= not((inputs(137)) or (inputs(31)));
    layer0_outputs(6759) <= (inputs(52)) and not (inputs(234));
    layer0_outputs(6760) <= (inputs(7)) and not (inputs(196));
    layer0_outputs(6761) <= not(inputs(233)) or (inputs(238));
    layer0_outputs(6762) <= not(inputs(70)) or (inputs(188));
    layer0_outputs(6763) <= inputs(145);
    layer0_outputs(6764) <= (inputs(68)) or (inputs(169));
    layer0_outputs(6765) <= (inputs(5)) or (inputs(30));
    layer0_outputs(6766) <= (inputs(89)) and not (inputs(83));
    layer0_outputs(6767) <= not((inputs(174)) xor (inputs(57)));
    layer0_outputs(6768) <= (inputs(121)) xor (inputs(52));
    layer0_outputs(6769) <= (inputs(96)) xor (inputs(172));
    layer0_outputs(6770) <= (inputs(67)) or (inputs(86));
    layer0_outputs(6771) <= (inputs(246)) and not (inputs(30));
    layer0_outputs(6772) <= (inputs(26)) or (inputs(10));
    layer0_outputs(6773) <= (inputs(164)) or (inputs(82));
    layer0_outputs(6774) <= not(inputs(177));
    layer0_outputs(6775) <= not((inputs(20)) or (inputs(125)));
    layer0_outputs(6776) <= not((inputs(219)) xor (inputs(38)));
    layer0_outputs(6777) <= not(inputs(108)) or (inputs(14));
    layer0_outputs(6778) <= not((inputs(232)) or (inputs(75)));
    layer0_outputs(6779) <= not((inputs(157)) or (inputs(175)));
    layer0_outputs(6780) <= (inputs(182)) xor (inputs(33));
    layer0_outputs(6781) <= inputs(47);
    layer0_outputs(6782) <= inputs(165);
    layer0_outputs(6783) <= (inputs(61)) and not (inputs(255));
    layer0_outputs(6784) <= (inputs(137)) xor (inputs(170));
    layer0_outputs(6785) <= not((inputs(253)) xor (inputs(246)));
    layer0_outputs(6786) <= not(inputs(169)) or (inputs(78));
    layer0_outputs(6787) <= not((inputs(195)) or (inputs(178)));
    layer0_outputs(6788) <= (inputs(37)) xor (inputs(13));
    layer0_outputs(6789) <= inputs(119);
    layer0_outputs(6790) <= not(inputs(218));
    layer0_outputs(6791) <= '0';
    layer0_outputs(6792) <= inputs(146);
    layer0_outputs(6793) <= not(inputs(13));
    layer0_outputs(6794) <= (inputs(18)) xor (inputs(251));
    layer0_outputs(6795) <= not(inputs(89)) or (inputs(150));
    layer0_outputs(6796) <= inputs(219);
    layer0_outputs(6797) <= (inputs(133)) and not (inputs(242));
    layer0_outputs(6798) <= inputs(198);
    layer0_outputs(6799) <= not(inputs(254));
    layer0_outputs(6800) <= not((inputs(148)) xor (inputs(209)));
    layer0_outputs(6801) <= inputs(217);
    layer0_outputs(6802) <= (inputs(219)) xor (inputs(187));
    layer0_outputs(6803) <= not((inputs(140)) or (inputs(100)));
    layer0_outputs(6804) <= (inputs(162)) xor (inputs(116));
    layer0_outputs(6805) <= '0';
    layer0_outputs(6806) <= not(inputs(177));
    layer0_outputs(6807) <= not((inputs(1)) or (inputs(62)));
    layer0_outputs(6808) <= (inputs(218)) xor (inputs(78));
    layer0_outputs(6809) <= inputs(210);
    layer0_outputs(6810) <= (inputs(245)) or (inputs(35));
    layer0_outputs(6811) <= inputs(163);
    layer0_outputs(6812) <= inputs(165);
    layer0_outputs(6813) <= (inputs(29)) and not (inputs(210));
    layer0_outputs(6814) <= not(inputs(125)) or (inputs(34));
    layer0_outputs(6815) <= not(inputs(85)) or (inputs(127));
    layer0_outputs(6816) <= '0';
    layer0_outputs(6817) <= not(inputs(217)) or (inputs(43));
    layer0_outputs(6818) <= inputs(75);
    layer0_outputs(6819) <= (inputs(223)) or (inputs(173));
    layer0_outputs(6820) <= not((inputs(236)) or (inputs(6)));
    layer0_outputs(6821) <= (inputs(184)) or (inputs(45));
    layer0_outputs(6822) <= (inputs(168)) xor (inputs(246));
    layer0_outputs(6823) <= (inputs(36)) and not (inputs(9));
    layer0_outputs(6824) <= (inputs(91)) and not (inputs(64));
    layer0_outputs(6825) <= not((inputs(82)) or (inputs(53)));
    layer0_outputs(6826) <= (inputs(77)) and not (inputs(240));
    layer0_outputs(6827) <= not((inputs(101)) xor (inputs(49)));
    layer0_outputs(6828) <= not((inputs(48)) or (inputs(176)));
    layer0_outputs(6829) <= not((inputs(204)) xor (inputs(170)));
    layer0_outputs(6830) <= not(inputs(117));
    layer0_outputs(6831) <= (inputs(178)) or (inputs(56));
    layer0_outputs(6832) <= not(inputs(246)) or (inputs(225));
    layer0_outputs(6833) <= '1';
    layer0_outputs(6834) <= not((inputs(38)) or (inputs(155)));
    layer0_outputs(6835) <= not(inputs(118));
    layer0_outputs(6836) <= (inputs(72)) and not (inputs(8));
    layer0_outputs(6837) <= not(inputs(148)) or (inputs(240));
    layer0_outputs(6838) <= inputs(148);
    layer0_outputs(6839) <= (inputs(65)) or (inputs(213));
    layer0_outputs(6840) <= inputs(233);
    layer0_outputs(6841) <= not(inputs(2));
    layer0_outputs(6842) <= (inputs(149)) and (inputs(31));
    layer0_outputs(6843) <= inputs(213);
    layer0_outputs(6844) <= not((inputs(63)) and (inputs(65)));
    layer0_outputs(6845) <= not(inputs(29)) or (inputs(10));
    layer0_outputs(6846) <= not((inputs(197)) xor (inputs(244)));
    layer0_outputs(6847) <= (inputs(120)) and not (inputs(191));
    layer0_outputs(6848) <= (inputs(132)) and not (inputs(80));
    layer0_outputs(6849) <= '0';
    layer0_outputs(6850) <= not(inputs(102));
    layer0_outputs(6851) <= not((inputs(4)) xor (inputs(142)));
    layer0_outputs(6852) <= not(inputs(197));
    layer0_outputs(6853) <= not(inputs(144)) or (inputs(171));
    layer0_outputs(6854) <= not(inputs(199));
    layer0_outputs(6855) <= (inputs(79)) and not (inputs(50));
    layer0_outputs(6856) <= not(inputs(133)) or (inputs(17));
    layer0_outputs(6857) <= (inputs(174)) or (inputs(199));
    layer0_outputs(6858) <= (inputs(56)) and not (inputs(27));
    layer0_outputs(6859) <= not((inputs(60)) xor (inputs(155)));
    layer0_outputs(6860) <= inputs(157);
    layer0_outputs(6861) <= (inputs(17)) xor (inputs(36));
    layer0_outputs(6862) <= (inputs(31)) or (inputs(159));
    layer0_outputs(6863) <= (inputs(218)) and not (inputs(3));
    layer0_outputs(6864) <= (inputs(127)) and not (inputs(207));
    layer0_outputs(6865) <= not(inputs(112));
    layer0_outputs(6866) <= not((inputs(22)) xor (inputs(217)));
    layer0_outputs(6867) <= not((inputs(47)) or (inputs(196)));
    layer0_outputs(6868) <= '0';
    layer0_outputs(6869) <= inputs(72);
    layer0_outputs(6870) <= (inputs(92)) and (inputs(212));
    layer0_outputs(6871) <= not((inputs(228)) or (inputs(52)));
    layer0_outputs(6872) <= inputs(72);
    layer0_outputs(6873) <= (inputs(29)) or (inputs(184));
    layer0_outputs(6874) <= not(inputs(222));
    layer0_outputs(6875) <= not(inputs(11));
    layer0_outputs(6876) <= (inputs(79)) and not (inputs(251));
    layer0_outputs(6877) <= (inputs(182)) and not (inputs(53));
    layer0_outputs(6878) <= (inputs(250)) or (inputs(186));
    layer0_outputs(6879) <= not((inputs(42)) or (inputs(15)));
    layer0_outputs(6880) <= (inputs(250)) or (inputs(244));
    layer0_outputs(6881) <= inputs(183);
    layer0_outputs(6882) <= (inputs(200)) and (inputs(195));
    layer0_outputs(6883) <= not(inputs(26)) or (inputs(255));
    layer0_outputs(6884) <= not((inputs(9)) xor (inputs(207)));
    layer0_outputs(6885) <= not(inputs(69)) or (inputs(168));
    layer0_outputs(6886) <= not(inputs(189)) or (inputs(1));
    layer0_outputs(6887) <= not(inputs(43)) or (inputs(35));
    layer0_outputs(6888) <= not(inputs(255));
    layer0_outputs(6889) <= not(inputs(158));
    layer0_outputs(6890) <= not((inputs(208)) xor (inputs(124)));
    layer0_outputs(6891) <= not((inputs(144)) or (inputs(239)));
    layer0_outputs(6892) <= (inputs(246)) and not (inputs(59));
    layer0_outputs(6893) <= not((inputs(248)) or (inputs(94)));
    layer0_outputs(6894) <= inputs(90);
    layer0_outputs(6895) <= not(inputs(22));
    layer0_outputs(6896) <= not(inputs(91));
    layer0_outputs(6897) <= not((inputs(195)) xor (inputs(77)));
    layer0_outputs(6898) <= not((inputs(194)) xor (inputs(28)));
    layer0_outputs(6899) <= (inputs(30)) and (inputs(14));
    layer0_outputs(6900) <= not(inputs(117)) or (inputs(225));
    layer0_outputs(6901) <= inputs(63);
    layer0_outputs(6902) <= not(inputs(210));
    layer0_outputs(6903) <= not((inputs(228)) and (inputs(92)));
    layer0_outputs(6904) <= (inputs(15)) or (inputs(99));
    layer0_outputs(6905) <= inputs(126);
    layer0_outputs(6906) <= not(inputs(165)) or (inputs(224));
    layer0_outputs(6907) <= not((inputs(102)) xor (inputs(8)));
    layer0_outputs(6908) <= (inputs(86)) and not (inputs(97));
    layer0_outputs(6909) <= (inputs(189)) xor (inputs(88));
    layer0_outputs(6910) <= (inputs(230)) and not (inputs(107));
    layer0_outputs(6911) <= (inputs(116)) and not (inputs(197));
    layer0_outputs(6912) <= not((inputs(76)) or (inputs(20)));
    layer0_outputs(6913) <= not((inputs(29)) or (inputs(87)));
    layer0_outputs(6914) <= not(inputs(123)) or (inputs(218));
    layer0_outputs(6915) <= inputs(150);
    layer0_outputs(6916) <= not(inputs(71)) or (inputs(177));
    layer0_outputs(6917) <= inputs(198);
    layer0_outputs(6918) <= not((inputs(225)) or (inputs(237)));
    layer0_outputs(6919) <= (inputs(33)) or (inputs(167));
    layer0_outputs(6920) <= not(inputs(132));
    layer0_outputs(6921) <= (inputs(151)) and not (inputs(144));
    layer0_outputs(6922) <= (inputs(34)) xor (inputs(45));
    layer0_outputs(6923) <= inputs(68);
    layer0_outputs(6924) <= not((inputs(207)) xor (inputs(188)));
    layer0_outputs(6925) <= (inputs(84)) and not (inputs(31));
    layer0_outputs(6926) <= inputs(37);
    layer0_outputs(6927) <= inputs(137);
    layer0_outputs(6928) <= not(inputs(60));
    layer0_outputs(6929) <= (inputs(85)) or (inputs(29));
    layer0_outputs(6930) <= inputs(110);
    layer0_outputs(6931) <= (inputs(184)) or (inputs(110));
    layer0_outputs(6932) <= inputs(102);
    layer0_outputs(6933) <= inputs(233);
    layer0_outputs(6934) <= not(inputs(181));
    layer0_outputs(6935) <= (inputs(194)) or (inputs(242));
    layer0_outputs(6936) <= not((inputs(5)) or (inputs(175)));
    layer0_outputs(6937) <= not(inputs(26)) or (inputs(199));
    layer0_outputs(6938) <= (inputs(177)) or (inputs(225));
    layer0_outputs(6939) <= (inputs(221)) or (inputs(245));
    layer0_outputs(6940) <= not((inputs(139)) xor (inputs(219)));
    layer0_outputs(6941) <= (inputs(126)) or (inputs(83));
    layer0_outputs(6942) <= inputs(102);
    layer0_outputs(6943) <= (inputs(22)) xor (inputs(94));
    layer0_outputs(6944) <= inputs(165);
    layer0_outputs(6945) <= inputs(18);
    layer0_outputs(6946) <= (inputs(245)) xor (inputs(94));
    layer0_outputs(6947) <= not((inputs(20)) or (inputs(140)));
    layer0_outputs(6948) <= (inputs(219)) xor (inputs(45));
    layer0_outputs(6949) <= not(inputs(176));
    layer0_outputs(6950) <= not(inputs(63));
    layer0_outputs(6951) <= '0';
    layer0_outputs(6952) <= (inputs(228)) xor (inputs(177));
    layer0_outputs(6953) <= (inputs(176)) or (inputs(28));
    layer0_outputs(6954) <= not((inputs(113)) or (inputs(246)));
    layer0_outputs(6955) <= not(inputs(233));
    layer0_outputs(6956) <= not(inputs(181)) or (inputs(33));
    layer0_outputs(6957) <= (inputs(111)) or (inputs(26));
    layer0_outputs(6958) <= not(inputs(35));
    layer0_outputs(6959) <= inputs(114);
    layer0_outputs(6960) <= '0';
    layer0_outputs(6961) <= not(inputs(29));
    layer0_outputs(6962) <= not(inputs(37));
    layer0_outputs(6963) <= inputs(40);
    layer0_outputs(6964) <= not((inputs(35)) or (inputs(176)));
    layer0_outputs(6965) <= not(inputs(18));
    layer0_outputs(6966) <= (inputs(34)) and not (inputs(193));
    layer0_outputs(6967) <= (inputs(5)) and not (inputs(171));
    layer0_outputs(6968) <= not(inputs(49)) or (inputs(81));
    layer0_outputs(6969) <= (inputs(80)) or (inputs(212));
    layer0_outputs(6970) <= not(inputs(106));
    layer0_outputs(6971) <= not(inputs(169));
    layer0_outputs(6972) <= (inputs(131)) and (inputs(233));
    layer0_outputs(6973) <= not((inputs(33)) or (inputs(57)));
    layer0_outputs(6974) <= (inputs(149)) xor (inputs(200));
    layer0_outputs(6975) <= not((inputs(51)) or (inputs(90)));
    layer0_outputs(6976) <= (inputs(224)) and not (inputs(187));
    layer0_outputs(6977) <= inputs(146);
    layer0_outputs(6978) <= (inputs(189)) xor (inputs(191));
    layer0_outputs(6979) <= not(inputs(153)) or (inputs(9));
    layer0_outputs(6980) <= not(inputs(47));
    layer0_outputs(6981) <= (inputs(77)) or (inputs(170));
    layer0_outputs(6982) <= not((inputs(186)) xor (inputs(153)));
    layer0_outputs(6983) <= not(inputs(89)) or (inputs(185));
    layer0_outputs(6984) <= (inputs(64)) and (inputs(27));
    layer0_outputs(6985) <= not((inputs(40)) and (inputs(42)));
    layer0_outputs(6986) <= (inputs(92)) and (inputs(122));
    layer0_outputs(6987) <= (inputs(5)) or (inputs(253));
    layer0_outputs(6988) <= not(inputs(199)) or (inputs(108));
    layer0_outputs(6989) <= inputs(183);
    layer0_outputs(6990) <= inputs(97);
    layer0_outputs(6991) <= (inputs(58)) xor (inputs(106));
    layer0_outputs(6992) <= inputs(145);
    layer0_outputs(6993) <= not(inputs(140)) or (inputs(22));
    layer0_outputs(6994) <= not((inputs(161)) xor (inputs(181)));
    layer0_outputs(6995) <= not((inputs(180)) or (inputs(197)));
    layer0_outputs(6996) <= inputs(62);
    layer0_outputs(6997) <= not(inputs(248));
    layer0_outputs(6998) <= (inputs(108)) and not (inputs(190));
    layer0_outputs(6999) <= not((inputs(46)) or (inputs(126)));
    layer0_outputs(7000) <= (inputs(150)) or (inputs(153));
    layer0_outputs(7001) <= (inputs(31)) or (inputs(212));
    layer0_outputs(7002) <= not(inputs(197));
    layer0_outputs(7003) <= (inputs(5)) and not (inputs(21));
    layer0_outputs(7004) <= not(inputs(120));
    layer0_outputs(7005) <= not(inputs(30));
    layer0_outputs(7006) <= (inputs(121)) or (inputs(86));
    layer0_outputs(7007) <= not(inputs(116));
    layer0_outputs(7008) <= not((inputs(118)) or (inputs(18)));
    layer0_outputs(7009) <= not(inputs(21));
    layer0_outputs(7010) <= inputs(107);
    layer0_outputs(7011) <= (inputs(229)) or (inputs(159));
    layer0_outputs(7012) <= not(inputs(154)) or (inputs(174));
    layer0_outputs(7013) <= not((inputs(12)) xor (inputs(39)));
    layer0_outputs(7014) <= not((inputs(144)) xor (inputs(163)));
    layer0_outputs(7015) <= (inputs(103)) and (inputs(87));
    layer0_outputs(7016) <= not(inputs(213));
    layer0_outputs(7017) <= inputs(91);
    layer0_outputs(7018) <= inputs(230);
    layer0_outputs(7019) <= not(inputs(25));
    layer0_outputs(7020) <= inputs(105);
    layer0_outputs(7021) <= not((inputs(118)) xor (inputs(97)));
    layer0_outputs(7022) <= (inputs(62)) and not (inputs(128));
    layer0_outputs(7023) <= (inputs(213)) xor (inputs(211));
    layer0_outputs(7024) <= not(inputs(71)) or (inputs(11));
    layer0_outputs(7025) <= not(inputs(136)) or (inputs(128));
    layer0_outputs(7026) <= not((inputs(185)) xor (inputs(51)));
    layer0_outputs(7027) <= not(inputs(9));
    layer0_outputs(7028) <= not(inputs(42));
    layer0_outputs(7029) <= (inputs(90)) and (inputs(122));
    layer0_outputs(7030) <= not((inputs(184)) xor (inputs(120)));
    layer0_outputs(7031) <= not((inputs(94)) or (inputs(184)));
    layer0_outputs(7032) <= inputs(148);
    layer0_outputs(7033) <= not(inputs(197)) or (inputs(34));
    layer0_outputs(7034) <= '0';
    layer0_outputs(7035) <= (inputs(25)) xor (inputs(71));
    layer0_outputs(7036) <= '1';
    layer0_outputs(7037) <= inputs(230);
    layer0_outputs(7038) <= not((inputs(189)) or (inputs(180)));
    layer0_outputs(7039) <= (inputs(250)) or (inputs(232));
    layer0_outputs(7040) <= not(inputs(105)) or (inputs(81));
    layer0_outputs(7041) <= not(inputs(42));
    layer0_outputs(7042) <= inputs(105);
    layer0_outputs(7043) <= not(inputs(35));
    layer0_outputs(7044) <= inputs(211);
    layer0_outputs(7045) <= not(inputs(55)) or (inputs(64));
    layer0_outputs(7046) <= (inputs(166)) or (inputs(110));
    layer0_outputs(7047) <= not(inputs(52));
    layer0_outputs(7048) <= not((inputs(238)) or (inputs(255)));
    layer0_outputs(7049) <= (inputs(119)) and not (inputs(58));
    layer0_outputs(7050) <= (inputs(197)) xor (inputs(107));
    layer0_outputs(7051) <= not((inputs(251)) or (inputs(184)));
    layer0_outputs(7052) <= not((inputs(5)) xor (inputs(36)));
    layer0_outputs(7053) <= (inputs(59)) and not (inputs(15));
    layer0_outputs(7054) <= not(inputs(231));
    layer0_outputs(7055) <= (inputs(233)) and (inputs(247));
    layer0_outputs(7056) <= '1';
    layer0_outputs(7057) <= not(inputs(125)) or (inputs(113));
    layer0_outputs(7058) <= not(inputs(181));
    layer0_outputs(7059) <= (inputs(184)) and not (inputs(225));
    layer0_outputs(7060) <= not(inputs(213));
    layer0_outputs(7061) <= '1';
    layer0_outputs(7062) <= inputs(66);
    layer0_outputs(7063) <= (inputs(108)) and (inputs(76));
    layer0_outputs(7064) <= (inputs(132)) and not (inputs(6));
    layer0_outputs(7065) <= (inputs(151)) and not (inputs(255));
    layer0_outputs(7066) <= (inputs(140)) and not (inputs(227));
    layer0_outputs(7067) <= not(inputs(26)) or (inputs(93));
    layer0_outputs(7068) <= not(inputs(188));
    layer0_outputs(7069) <= not(inputs(206));
    layer0_outputs(7070) <= not(inputs(13));
    layer0_outputs(7071) <= (inputs(176)) and (inputs(97));
    layer0_outputs(7072) <= not((inputs(160)) or (inputs(204)));
    layer0_outputs(7073) <= (inputs(58)) and not (inputs(203));
    layer0_outputs(7074) <= (inputs(20)) and not (inputs(254));
    layer0_outputs(7075) <= inputs(176);
    layer0_outputs(7076) <= (inputs(164)) xor (inputs(167));
    layer0_outputs(7077) <= (inputs(45)) xor (inputs(225));
    layer0_outputs(7078) <= not(inputs(112));
    layer0_outputs(7079) <= (inputs(134)) or (inputs(3));
    layer0_outputs(7080) <= not((inputs(78)) xor (inputs(175)));
    layer0_outputs(7081) <= not(inputs(107));
    layer0_outputs(7082) <= not(inputs(215));
    layer0_outputs(7083) <= (inputs(134)) and not (inputs(187));
    layer0_outputs(7084) <= inputs(9);
    layer0_outputs(7085) <= not(inputs(42));
    layer0_outputs(7086) <= not((inputs(28)) and (inputs(229)));
    layer0_outputs(7087) <= not((inputs(117)) xor (inputs(148)));
    layer0_outputs(7088) <= (inputs(125)) or (inputs(30));
    layer0_outputs(7089) <= not(inputs(10));
    layer0_outputs(7090) <= (inputs(73)) xor (inputs(36));
    layer0_outputs(7091) <= (inputs(99)) or (inputs(98));
    layer0_outputs(7092) <= not(inputs(200)) or (inputs(53));
    layer0_outputs(7093) <= not((inputs(151)) xor (inputs(75)));
    layer0_outputs(7094) <= not((inputs(174)) xor (inputs(148)));
    layer0_outputs(7095) <= (inputs(6)) and not (inputs(242));
    layer0_outputs(7096) <= not((inputs(229)) or (inputs(95)));
    layer0_outputs(7097) <= not((inputs(220)) or (inputs(118)));
    layer0_outputs(7098) <= '1';
    layer0_outputs(7099) <= not(inputs(188)) or (inputs(141));
    layer0_outputs(7100) <= not((inputs(105)) xor (inputs(23)));
    layer0_outputs(7101) <= not(inputs(76));
    layer0_outputs(7102) <= inputs(52);
    layer0_outputs(7103) <= (inputs(213)) xor (inputs(110));
    layer0_outputs(7104) <= not(inputs(23)) or (inputs(183));
    layer0_outputs(7105) <= inputs(115);
    layer0_outputs(7106) <= (inputs(18)) or (inputs(112));
    layer0_outputs(7107) <= (inputs(29)) or (inputs(115));
    layer0_outputs(7108) <= inputs(53);
    layer0_outputs(7109) <= (inputs(247)) and not (inputs(121));
    layer0_outputs(7110) <= not(inputs(51));
    layer0_outputs(7111) <= not((inputs(229)) xor (inputs(60)));
    layer0_outputs(7112) <= not((inputs(191)) xor (inputs(41)));
    layer0_outputs(7113) <= (inputs(137)) xor (inputs(200));
    layer0_outputs(7114) <= not((inputs(159)) or (inputs(210)));
    layer0_outputs(7115) <= inputs(8);
    layer0_outputs(7116) <= '1';
    layer0_outputs(7117) <= not(inputs(161)) or (inputs(245));
    layer0_outputs(7118) <= not((inputs(224)) xor (inputs(174)));
    layer0_outputs(7119) <= '0';
    layer0_outputs(7120) <= (inputs(78)) or (inputs(103));
    layer0_outputs(7121) <= not(inputs(100));
    layer0_outputs(7122) <= not((inputs(61)) xor (inputs(51)));
    layer0_outputs(7123) <= inputs(233);
    layer0_outputs(7124) <= not((inputs(204)) xor (inputs(197)));
    layer0_outputs(7125) <= not((inputs(90)) or (inputs(167)));
    layer0_outputs(7126) <= not((inputs(88)) xor (inputs(190)));
    layer0_outputs(7127) <= inputs(44);
    layer0_outputs(7128) <= (inputs(6)) xor (inputs(50));
    layer0_outputs(7129) <= (inputs(19)) xor (inputs(101));
    layer0_outputs(7130) <= (inputs(59)) and not (inputs(253));
    layer0_outputs(7131) <= inputs(160);
    layer0_outputs(7132) <= not((inputs(72)) xor (inputs(24)));
    layer0_outputs(7133) <= not((inputs(195)) xor (inputs(128)));
    layer0_outputs(7134) <= (inputs(124)) xor (inputs(21));
    layer0_outputs(7135) <= (inputs(38)) or (inputs(23));
    layer0_outputs(7136) <= not((inputs(153)) xor (inputs(181)));
    layer0_outputs(7137) <= (inputs(66)) and not (inputs(32));
    layer0_outputs(7138) <= (inputs(112)) xor (inputs(104));
    layer0_outputs(7139) <= not((inputs(50)) xor (inputs(242)));
    layer0_outputs(7140) <= inputs(138);
    layer0_outputs(7141) <= inputs(114);
    layer0_outputs(7142) <= (inputs(78)) or (inputs(140));
    layer0_outputs(7143) <= (inputs(134)) and not (inputs(217));
    layer0_outputs(7144) <= (inputs(186)) or (inputs(172));
    layer0_outputs(7145) <= inputs(135);
    layer0_outputs(7146) <= (inputs(208)) or (inputs(61));
    layer0_outputs(7147) <= inputs(97);
    layer0_outputs(7148) <= inputs(113);
    layer0_outputs(7149) <= (inputs(181)) xor (inputs(196));
    layer0_outputs(7150) <= (inputs(127)) or (inputs(125));
    layer0_outputs(7151) <= not((inputs(104)) xor (inputs(238)));
    layer0_outputs(7152) <= not(inputs(25));
    layer0_outputs(7153) <= (inputs(200)) and (inputs(237));
    layer0_outputs(7154) <= not(inputs(182));
    layer0_outputs(7155) <= not((inputs(224)) xor (inputs(133)));
    layer0_outputs(7156) <= inputs(144);
    layer0_outputs(7157) <= inputs(85);
    layer0_outputs(7158) <= not((inputs(247)) or (inputs(223)));
    layer0_outputs(7159) <= not((inputs(133)) xor (inputs(141)));
    layer0_outputs(7160) <= (inputs(59)) and not (inputs(30));
    layer0_outputs(7161) <= not(inputs(166)) or (inputs(173));
    layer0_outputs(7162) <= (inputs(151)) xor (inputs(184));
    layer0_outputs(7163) <= (inputs(242)) xor (inputs(88));
    layer0_outputs(7164) <= inputs(79);
    layer0_outputs(7165) <= not(inputs(193));
    layer0_outputs(7166) <= (inputs(164)) or (inputs(80));
    layer0_outputs(7167) <= inputs(100);
    layer0_outputs(7168) <= not(inputs(53));
    layer0_outputs(7169) <= not((inputs(71)) xor (inputs(128)));
    layer0_outputs(7170) <= (inputs(138)) and not (inputs(213));
    layer0_outputs(7171) <= (inputs(182)) and not (inputs(82));
    layer0_outputs(7172) <= not(inputs(171)) or (inputs(22));
    layer0_outputs(7173) <= not(inputs(89)) or (inputs(112));
    layer0_outputs(7174) <= not((inputs(15)) or (inputs(241)));
    layer0_outputs(7175) <= not((inputs(221)) xor (inputs(7)));
    layer0_outputs(7176) <= not(inputs(119)) or (inputs(19));
    layer0_outputs(7177) <= (inputs(196)) and not (inputs(91));
    layer0_outputs(7178) <= not((inputs(224)) xor (inputs(222)));
    layer0_outputs(7179) <= not(inputs(20));
    layer0_outputs(7180) <= (inputs(74)) and not (inputs(188));
    layer0_outputs(7181) <= inputs(248);
    layer0_outputs(7182) <= inputs(241);
    layer0_outputs(7183) <= not((inputs(213)) and (inputs(64)));
    layer0_outputs(7184) <= not((inputs(232)) or (inputs(17)));
    layer0_outputs(7185) <= not(inputs(232));
    layer0_outputs(7186) <= not((inputs(124)) and (inputs(166)));
    layer0_outputs(7187) <= (inputs(213)) and (inputs(158));
    layer0_outputs(7188) <= not(inputs(104)) or (inputs(226));
    layer0_outputs(7189) <= not((inputs(141)) xor (inputs(236)));
    layer0_outputs(7190) <= (inputs(165)) or (inputs(50));
    layer0_outputs(7191) <= not((inputs(228)) and (inputs(175)));
    layer0_outputs(7192) <= (inputs(106)) and not (inputs(221));
    layer0_outputs(7193) <= not((inputs(11)) xor (inputs(61)));
    layer0_outputs(7194) <= not(inputs(229)) or (inputs(15));
    layer0_outputs(7195) <= '0';
    layer0_outputs(7196) <= not((inputs(37)) xor (inputs(197)));
    layer0_outputs(7197) <= not((inputs(204)) and (inputs(101)));
    layer0_outputs(7198) <= (inputs(193)) xor (inputs(39));
    layer0_outputs(7199) <= (inputs(230)) xor (inputs(36));
    layer0_outputs(7200) <= inputs(14);
    layer0_outputs(7201) <= inputs(85);
    layer0_outputs(7202) <= not((inputs(125)) xor (inputs(44)));
    layer0_outputs(7203) <= not((inputs(135)) xor (inputs(148)));
    layer0_outputs(7204) <= (inputs(166)) xor (inputs(131));
    layer0_outputs(7205) <= not((inputs(85)) xor (inputs(25)));
    layer0_outputs(7206) <= (inputs(196)) and not (inputs(86));
    layer0_outputs(7207) <= not(inputs(102));
    layer0_outputs(7208) <= inputs(191);
    layer0_outputs(7209) <= not((inputs(137)) or (inputs(123)));
    layer0_outputs(7210) <= inputs(177);
    layer0_outputs(7211) <= inputs(46);
    layer0_outputs(7212) <= not(inputs(181));
    layer0_outputs(7213) <= not((inputs(206)) xor (inputs(64)));
    layer0_outputs(7214) <= not((inputs(218)) or (inputs(178)));
    layer0_outputs(7215) <= (inputs(77)) xor (inputs(159));
    layer0_outputs(7216) <= not(inputs(185));
    layer0_outputs(7217) <= '0';
    layer0_outputs(7218) <= (inputs(104)) xor (inputs(190));
    layer0_outputs(7219) <= not((inputs(99)) or (inputs(233)));
    layer0_outputs(7220) <= not((inputs(133)) or (inputs(72)));
    layer0_outputs(7221) <= inputs(133);
    layer0_outputs(7222) <= inputs(217);
    layer0_outputs(7223) <= not(inputs(87)) or (inputs(111));
    layer0_outputs(7224) <= (inputs(3)) and (inputs(21));
    layer0_outputs(7225) <= not(inputs(2)) or (inputs(220));
    layer0_outputs(7226) <= (inputs(119)) and not (inputs(57));
    layer0_outputs(7227) <= inputs(105);
    layer0_outputs(7228) <= (inputs(79)) or (inputs(193));
    layer0_outputs(7229) <= '1';
    layer0_outputs(7230) <= (inputs(53)) xor (inputs(174));
    layer0_outputs(7231) <= not((inputs(201)) or (inputs(225)));
    layer0_outputs(7232) <= inputs(82);
    layer0_outputs(7233) <= (inputs(163)) or (inputs(51));
    layer0_outputs(7234) <= (inputs(113)) or (inputs(140));
    layer0_outputs(7235) <= not(inputs(217));
    layer0_outputs(7236) <= not((inputs(242)) xor (inputs(197)));
    layer0_outputs(7237) <= '0';
    layer0_outputs(7238) <= not((inputs(63)) or (inputs(218)));
    layer0_outputs(7239) <= not(inputs(106)) or (inputs(225));
    layer0_outputs(7240) <= (inputs(72)) or (inputs(110));
    layer0_outputs(7241) <= (inputs(221)) or (inputs(63));
    layer0_outputs(7242) <= (inputs(244)) or (inputs(4));
    layer0_outputs(7243) <= not(inputs(248));
    layer0_outputs(7244) <= not((inputs(127)) and (inputs(105)));
    layer0_outputs(7245) <= not((inputs(114)) or (inputs(83)));
    layer0_outputs(7246) <= not((inputs(148)) or (inputs(112)));
    layer0_outputs(7247) <= inputs(60);
    layer0_outputs(7248) <= not(inputs(243)) or (inputs(62));
    layer0_outputs(7249) <= '0';
    layer0_outputs(7250) <= not(inputs(25));
    layer0_outputs(7251) <= '1';
    layer0_outputs(7252) <= (inputs(200)) and not (inputs(143));
    layer0_outputs(7253) <= (inputs(221)) or (inputs(194));
    layer0_outputs(7254) <= not((inputs(204)) xor (inputs(70)));
    layer0_outputs(7255) <= (inputs(134)) and not (inputs(142));
    layer0_outputs(7256) <= inputs(84);
    layer0_outputs(7257) <= not(inputs(147));
    layer0_outputs(7258) <= '0';
    layer0_outputs(7259) <= not(inputs(221)) or (inputs(30));
    layer0_outputs(7260) <= not(inputs(116));
    layer0_outputs(7261) <= not((inputs(250)) or (inputs(165)));
    layer0_outputs(7262) <= (inputs(219)) or (inputs(184));
    layer0_outputs(7263) <= not(inputs(152)) or (inputs(227));
    layer0_outputs(7264) <= not(inputs(143));
    layer0_outputs(7265) <= inputs(155);
    layer0_outputs(7266) <= not((inputs(238)) or (inputs(80)));
    layer0_outputs(7267) <= (inputs(217)) or (inputs(130));
    layer0_outputs(7268) <= not((inputs(227)) or (inputs(10)));
    layer0_outputs(7269) <= not(inputs(100));
    layer0_outputs(7270) <= (inputs(52)) or (inputs(211));
    layer0_outputs(7271) <= not(inputs(69)) or (inputs(157));
    layer0_outputs(7272) <= (inputs(135)) and not (inputs(69));
    layer0_outputs(7273) <= (inputs(67)) and not (inputs(38));
    layer0_outputs(7274) <= inputs(104);
    layer0_outputs(7275) <= (inputs(92)) and not (inputs(221));
    layer0_outputs(7276) <= (inputs(107)) xor (inputs(26));
    layer0_outputs(7277) <= not((inputs(166)) xor (inputs(204)));
    layer0_outputs(7278) <= inputs(7);
    layer0_outputs(7279) <= inputs(154);
    layer0_outputs(7280) <= (inputs(52)) and not (inputs(158));
    layer0_outputs(7281) <= not(inputs(43));
    layer0_outputs(7282) <= not(inputs(227));
    layer0_outputs(7283) <= '1';
    layer0_outputs(7284) <= inputs(167);
    layer0_outputs(7285) <= not(inputs(11)) or (inputs(240));
    layer0_outputs(7286) <= inputs(153);
    layer0_outputs(7287) <= not((inputs(154)) xor (inputs(172)));
    layer0_outputs(7288) <= inputs(196);
    layer0_outputs(7289) <= not((inputs(228)) xor (inputs(203)));
    layer0_outputs(7290) <= (inputs(24)) and not (inputs(82));
    layer0_outputs(7291) <= inputs(223);
    layer0_outputs(7292) <= inputs(137);
    layer0_outputs(7293) <= (inputs(23)) and not (inputs(227));
    layer0_outputs(7294) <= (inputs(24)) and not (inputs(112));
    layer0_outputs(7295) <= not(inputs(111));
    layer0_outputs(7296) <= not((inputs(34)) or (inputs(151)));
    layer0_outputs(7297) <= not(inputs(142));
    layer0_outputs(7298) <= not(inputs(13));
    layer0_outputs(7299) <= not(inputs(212));
    layer0_outputs(7300) <= (inputs(152)) and not (inputs(61));
    layer0_outputs(7301) <= inputs(115);
    layer0_outputs(7302) <= (inputs(147)) xor (inputs(113));
    layer0_outputs(7303) <= not(inputs(28));
    layer0_outputs(7304) <= not(inputs(57)) or (inputs(171));
    layer0_outputs(7305) <= inputs(144);
    layer0_outputs(7306) <= not((inputs(50)) xor (inputs(7)));
    layer0_outputs(7307) <= not((inputs(189)) xor (inputs(69)));
    layer0_outputs(7308) <= not((inputs(158)) or (inputs(2)));
    layer0_outputs(7309) <= not((inputs(81)) or (inputs(77)));
    layer0_outputs(7310) <= (inputs(37)) and not (inputs(99));
    layer0_outputs(7311) <= (inputs(218)) and not (inputs(167));
    layer0_outputs(7312) <= inputs(146);
    layer0_outputs(7313) <= not((inputs(220)) or (inputs(238)));
    layer0_outputs(7314) <= not((inputs(77)) or (inputs(53)));
    layer0_outputs(7315) <= not(inputs(121));
    layer0_outputs(7316) <= not((inputs(20)) xor (inputs(109)));
    layer0_outputs(7317) <= not(inputs(163));
    layer0_outputs(7318) <= (inputs(212)) and not (inputs(15));
    layer0_outputs(7319) <= inputs(110);
    layer0_outputs(7320) <= not((inputs(138)) or (inputs(191)));
    layer0_outputs(7321) <= not((inputs(129)) xor (inputs(106)));
    layer0_outputs(7322) <= (inputs(157)) xor (inputs(159));
    layer0_outputs(7323) <= (inputs(226)) or (inputs(241));
    layer0_outputs(7324) <= '1';
    layer0_outputs(7325) <= inputs(165);
    layer0_outputs(7326) <= '0';
    layer0_outputs(7327) <= inputs(228);
    layer0_outputs(7328) <= (inputs(40)) xor (inputs(208));
    layer0_outputs(7329) <= not(inputs(18));
    layer0_outputs(7330) <= not((inputs(143)) or (inputs(13)));
    layer0_outputs(7331) <= inputs(25);
    layer0_outputs(7332) <= not(inputs(100));
    layer0_outputs(7333) <= not(inputs(139)) or (inputs(74));
    layer0_outputs(7334) <= not(inputs(151)) or (inputs(237));
    layer0_outputs(7335) <= (inputs(93)) and not (inputs(97));
    layer0_outputs(7336) <= inputs(74);
    layer0_outputs(7337) <= not((inputs(29)) and (inputs(207)));
    layer0_outputs(7338) <= (inputs(56)) and not (inputs(194));
    layer0_outputs(7339) <= not((inputs(211)) or (inputs(166)));
    layer0_outputs(7340) <= inputs(121);
    layer0_outputs(7341) <= not((inputs(94)) or (inputs(140)));
    layer0_outputs(7342) <= inputs(20);
    layer0_outputs(7343) <= not((inputs(40)) xor (inputs(13)));
    layer0_outputs(7344) <= not(inputs(229)) or (inputs(24));
    layer0_outputs(7345) <= not((inputs(207)) or (inputs(191)));
    layer0_outputs(7346) <= (inputs(229)) and not (inputs(107));
    layer0_outputs(7347) <= not(inputs(218)) or (inputs(81));
    layer0_outputs(7348) <= (inputs(140)) xor (inputs(138));
    layer0_outputs(7349) <= inputs(240);
    layer0_outputs(7350) <= not(inputs(52)) or (inputs(113));
    layer0_outputs(7351) <= inputs(78);
    layer0_outputs(7352) <= not(inputs(120));
    layer0_outputs(7353) <= not((inputs(167)) and (inputs(198)));
    layer0_outputs(7354) <= (inputs(75)) or (inputs(81));
    layer0_outputs(7355) <= inputs(37);
    layer0_outputs(7356) <= not(inputs(161));
    layer0_outputs(7357) <= not((inputs(16)) and (inputs(65)));
    layer0_outputs(7358) <= not((inputs(182)) xor (inputs(161)));
    layer0_outputs(7359) <= not(inputs(97));
    layer0_outputs(7360) <= not(inputs(156)) or (inputs(96));
    layer0_outputs(7361) <= (inputs(212)) and not (inputs(77));
    layer0_outputs(7362) <= not((inputs(78)) xor (inputs(110)));
    layer0_outputs(7363) <= (inputs(74)) and not (inputs(185));
    layer0_outputs(7364) <= (inputs(254)) or (inputs(138));
    layer0_outputs(7365) <= inputs(201);
    layer0_outputs(7366) <= (inputs(217)) or (inputs(39));
    layer0_outputs(7367) <= (inputs(223)) and not (inputs(15));
    layer0_outputs(7368) <= (inputs(161)) or (inputs(44));
    layer0_outputs(7369) <= (inputs(158)) and not (inputs(172));
    layer0_outputs(7370) <= (inputs(28)) or (inputs(201));
    layer0_outputs(7371) <= not((inputs(191)) or (inputs(248)));
    layer0_outputs(7372) <= (inputs(146)) and not (inputs(73));
    layer0_outputs(7373) <= not((inputs(33)) xor (inputs(172)));
    layer0_outputs(7374) <= (inputs(6)) xor (inputs(214));
    layer0_outputs(7375) <= '1';
    layer0_outputs(7376) <= (inputs(70)) xor (inputs(96));
    layer0_outputs(7377) <= (inputs(53)) xor (inputs(71));
    layer0_outputs(7378) <= inputs(238);
    layer0_outputs(7379) <= not(inputs(62));
    layer0_outputs(7380) <= inputs(181);
    layer0_outputs(7381) <= '1';
    layer0_outputs(7382) <= not(inputs(85));
    layer0_outputs(7383) <= not(inputs(79));
    layer0_outputs(7384) <= not((inputs(177)) xor (inputs(242)));
    layer0_outputs(7385) <= inputs(14);
    layer0_outputs(7386) <= not(inputs(76));
    layer0_outputs(7387) <= (inputs(36)) and not (inputs(189));
    layer0_outputs(7388) <= (inputs(252)) or (inputs(145));
    layer0_outputs(7389) <= not((inputs(83)) xor (inputs(132)));
    layer0_outputs(7390) <= not(inputs(142));
    layer0_outputs(7391) <= (inputs(185)) and (inputs(163));
    layer0_outputs(7392) <= not((inputs(189)) or (inputs(15)));
    layer0_outputs(7393) <= inputs(35);
    layer0_outputs(7394) <= not((inputs(242)) xor (inputs(227)));
    layer0_outputs(7395) <= (inputs(87)) and not (inputs(46));
    layer0_outputs(7396) <= not(inputs(21)) or (inputs(241));
    layer0_outputs(7397) <= (inputs(108)) and not (inputs(79));
    layer0_outputs(7398) <= not(inputs(91));
    layer0_outputs(7399) <= not((inputs(63)) xor (inputs(24)));
    layer0_outputs(7400) <= (inputs(122)) xor (inputs(48));
    layer0_outputs(7401) <= not((inputs(127)) or (inputs(163)));
    layer0_outputs(7402) <= (inputs(64)) and not (inputs(79));
    layer0_outputs(7403) <= (inputs(43)) or (inputs(41));
    layer0_outputs(7404) <= not(inputs(226)) or (inputs(81));
    layer0_outputs(7405) <= (inputs(192)) xor (inputs(29));
    layer0_outputs(7406) <= not(inputs(92));
    layer0_outputs(7407) <= not(inputs(235));
    layer0_outputs(7408) <= inputs(148);
    layer0_outputs(7409) <= (inputs(99)) and not (inputs(190));
    layer0_outputs(7410) <= not(inputs(35));
    layer0_outputs(7411) <= not(inputs(215)) or (inputs(93));
    layer0_outputs(7412) <= not(inputs(193));
    layer0_outputs(7413) <= not(inputs(22));
    layer0_outputs(7414) <= (inputs(132)) xor (inputs(175));
    layer0_outputs(7415) <= (inputs(99)) and not (inputs(60));
    layer0_outputs(7416) <= (inputs(79)) and not (inputs(238));
    layer0_outputs(7417) <= not(inputs(76)) or (inputs(253));
    layer0_outputs(7418) <= inputs(170);
    layer0_outputs(7419) <= (inputs(99)) and not (inputs(243));
    layer0_outputs(7420) <= not((inputs(249)) or (inputs(218)));
    layer0_outputs(7421) <= inputs(91);
    layer0_outputs(7422) <= not(inputs(151)) or (inputs(54));
    layer0_outputs(7423) <= inputs(176);
    layer0_outputs(7424) <= not(inputs(181));
    layer0_outputs(7425) <= inputs(109);
    layer0_outputs(7426) <= not(inputs(131)) or (inputs(193));
    layer0_outputs(7427) <= (inputs(74)) and not (inputs(65));
    layer0_outputs(7428) <= not((inputs(201)) xor (inputs(143)));
    layer0_outputs(7429) <= inputs(8);
    layer0_outputs(7430) <= not(inputs(151));
    layer0_outputs(7431) <= not((inputs(37)) or (inputs(253)));
    layer0_outputs(7432) <= (inputs(24)) and not (inputs(251));
    layer0_outputs(7433) <= not((inputs(103)) or (inputs(89)));
    layer0_outputs(7434) <= (inputs(153)) and not (inputs(7));
    layer0_outputs(7435) <= (inputs(187)) xor (inputs(10));
    layer0_outputs(7436) <= (inputs(199)) xor (inputs(185));
    layer0_outputs(7437) <= (inputs(132)) or (inputs(46));
    layer0_outputs(7438) <= (inputs(205)) or (inputs(183));
    layer0_outputs(7439) <= '0';
    layer0_outputs(7440) <= inputs(226);
    layer0_outputs(7441) <= (inputs(45)) and (inputs(163));
    layer0_outputs(7442) <= not(inputs(57));
    layer0_outputs(7443) <= inputs(141);
    layer0_outputs(7444) <= (inputs(234)) and not (inputs(130));
    layer0_outputs(7445) <= (inputs(20)) xor (inputs(123));
    layer0_outputs(7446) <= not((inputs(160)) xor (inputs(170)));
    layer0_outputs(7447) <= inputs(73);
    layer0_outputs(7448) <= inputs(99);
    layer0_outputs(7449) <= (inputs(45)) and not (inputs(94));
    layer0_outputs(7450) <= (inputs(2)) or (inputs(24));
    layer0_outputs(7451) <= (inputs(165)) xor (inputs(62));
    layer0_outputs(7452) <= not(inputs(250)) or (inputs(76));
    layer0_outputs(7453) <= not(inputs(28));
    layer0_outputs(7454) <= (inputs(59)) xor (inputs(34));
    layer0_outputs(7455) <= inputs(208);
    layer0_outputs(7456) <= inputs(69);
    layer0_outputs(7457) <= (inputs(128)) or (inputs(199));
    layer0_outputs(7458) <= not((inputs(109)) or (inputs(38)));
    layer0_outputs(7459) <= not((inputs(115)) or (inputs(155)));
    layer0_outputs(7460) <= (inputs(198)) and (inputs(197));
    layer0_outputs(7461) <= not(inputs(181)) or (inputs(63));
    layer0_outputs(7462) <= not(inputs(5));
    layer0_outputs(7463) <= not(inputs(57));
    layer0_outputs(7464) <= not((inputs(119)) or (inputs(104)));
    layer0_outputs(7465) <= (inputs(187)) xor (inputs(185));
    layer0_outputs(7466) <= (inputs(218)) and not (inputs(86));
    layer0_outputs(7467) <= not((inputs(117)) xor (inputs(66)));
    layer0_outputs(7468) <= not(inputs(171));
    layer0_outputs(7469) <= not(inputs(57));
    layer0_outputs(7470) <= not(inputs(33));
    layer0_outputs(7471) <= not((inputs(245)) xor (inputs(212)));
    layer0_outputs(7472) <= (inputs(133)) xor (inputs(26));
    layer0_outputs(7473) <= not((inputs(164)) or (inputs(209)));
    layer0_outputs(7474) <= not((inputs(202)) or (inputs(12)));
    layer0_outputs(7475) <= (inputs(242)) and not (inputs(78));
    layer0_outputs(7476) <= (inputs(96)) or (inputs(37));
    layer0_outputs(7477) <= not(inputs(195)) or (inputs(32));
    layer0_outputs(7478) <= not((inputs(74)) xor (inputs(87)));
    layer0_outputs(7479) <= not((inputs(53)) or (inputs(177)));
    layer0_outputs(7480) <= not(inputs(27)) or (inputs(234));
    layer0_outputs(7481) <= (inputs(182)) and not (inputs(209));
    layer0_outputs(7482) <= inputs(27);
    layer0_outputs(7483) <= not((inputs(72)) and (inputs(160)));
    layer0_outputs(7484) <= inputs(178);
    layer0_outputs(7485) <= (inputs(252)) xor (inputs(246));
    layer0_outputs(7486) <= not(inputs(169));
    layer0_outputs(7487) <= not((inputs(67)) xor (inputs(153)));
    layer0_outputs(7488) <= not(inputs(218));
    layer0_outputs(7489) <= (inputs(173)) xor (inputs(168));
    layer0_outputs(7490) <= not(inputs(225));
    layer0_outputs(7491) <= (inputs(77)) xor (inputs(154));
    layer0_outputs(7492) <= (inputs(37)) xor (inputs(126));
    layer0_outputs(7493) <= not((inputs(32)) or (inputs(1)));
    layer0_outputs(7494) <= (inputs(92)) and (inputs(119));
    layer0_outputs(7495) <= inputs(161);
    layer0_outputs(7496) <= (inputs(23)) and not (inputs(234));
    layer0_outputs(7497) <= (inputs(39)) xor (inputs(165));
    layer0_outputs(7498) <= not(inputs(70));
    layer0_outputs(7499) <= not((inputs(32)) xor (inputs(149)));
    layer0_outputs(7500) <= (inputs(215)) and not (inputs(112));
    layer0_outputs(7501) <= (inputs(244)) and not (inputs(5));
    layer0_outputs(7502) <= (inputs(201)) and not (inputs(92));
    layer0_outputs(7503) <= not((inputs(85)) xor (inputs(5)));
    layer0_outputs(7504) <= not(inputs(65));
    layer0_outputs(7505) <= inputs(59);
    layer0_outputs(7506) <= (inputs(24)) and not (inputs(170));
    layer0_outputs(7507) <= not((inputs(137)) xor (inputs(125)));
    layer0_outputs(7508) <= not(inputs(244)) or (inputs(103));
    layer0_outputs(7509) <= not((inputs(174)) or (inputs(166)));
    layer0_outputs(7510) <= not((inputs(53)) xor (inputs(67)));
    layer0_outputs(7511) <= (inputs(159)) xor (inputs(187));
    layer0_outputs(7512) <= not((inputs(248)) or (inputs(45)));
    layer0_outputs(7513) <= not(inputs(120));
    layer0_outputs(7514) <= not((inputs(186)) xor (inputs(236)));
    layer0_outputs(7515) <= not((inputs(182)) xor (inputs(178)));
    layer0_outputs(7516) <= (inputs(34)) or (inputs(126));
    layer0_outputs(7517) <= (inputs(102)) xor (inputs(162));
    layer0_outputs(7518) <= (inputs(19)) or (inputs(163));
    layer0_outputs(7519) <= (inputs(188)) xor (inputs(191));
    layer0_outputs(7520) <= (inputs(73)) or (inputs(47));
    layer0_outputs(7521) <= not((inputs(32)) xor (inputs(109)));
    layer0_outputs(7522) <= not((inputs(168)) xor (inputs(135)));
    layer0_outputs(7523) <= not(inputs(199));
    layer0_outputs(7524) <= not(inputs(117)) or (inputs(2));
    layer0_outputs(7525) <= not(inputs(18));
    layer0_outputs(7526) <= (inputs(38)) or (inputs(188));
    layer0_outputs(7527) <= (inputs(120)) and (inputs(39));
    layer0_outputs(7528) <= not((inputs(228)) or (inputs(152)));
    layer0_outputs(7529) <= '1';
    layer0_outputs(7530) <= (inputs(90)) xor (inputs(140));
    layer0_outputs(7531) <= not(inputs(236));
    layer0_outputs(7532) <= not(inputs(196)) or (inputs(28));
    layer0_outputs(7533) <= not((inputs(5)) xor (inputs(186)));
    layer0_outputs(7534) <= not(inputs(177));
    layer0_outputs(7535) <= not(inputs(25));
    layer0_outputs(7536) <= (inputs(147)) and not (inputs(34));
    layer0_outputs(7537) <= not((inputs(200)) xor (inputs(11)));
    layer0_outputs(7538) <= (inputs(165)) and not (inputs(239));
    layer0_outputs(7539) <= (inputs(113)) and not (inputs(13));
    layer0_outputs(7540) <= not(inputs(82));
    layer0_outputs(7541) <= inputs(165);
    layer0_outputs(7542) <= inputs(110);
    layer0_outputs(7543) <= (inputs(27)) xor (inputs(247));
    layer0_outputs(7544) <= inputs(212);
    layer0_outputs(7545) <= not((inputs(201)) and (inputs(132)));
    layer0_outputs(7546) <= not((inputs(150)) xor (inputs(241)));
    layer0_outputs(7547) <= (inputs(190)) xor (inputs(19));
    layer0_outputs(7548) <= (inputs(203)) or (inputs(171));
    layer0_outputs(7549) <= not(inputs(36)) or (inputs(111));
    layer0_outputs(7550) <= (inputs(159)) or (inputs(5));
    layer0_outputs(7551) <= not((inputs(18)) or (inputs(211)));
    layer0_outputs(7552) <= not(inputs(163));
    layer0_outputs(7553) <= not((inputs(37)) or (inputs(19)));
    layer0_outputs(7554) <= not(inputs(69)) or (inputs(179));
    layer0_outputs(7555) <= not(inputs(67)) or (inputs(221));
    layer0_outputs(7556) <= not(inputs(77));
    layer0_outputs(7557) <= not(inputs(153)) or (inputs(110));
    layer0_outputs(7558) <= (inputs(195)) xor (inputs(226));
    layer0_outputs(7559) <= inputs(90);
    layer0_outputs(7560) <= (inputs(73)) xor (inputs(20));
    layer0_outputs(7561) <= (inputs(233)) and (inputs(172));
    layer0_outputs(7562) <= (inputs(130)) or (inputs(220));
    layer0_outputs(7563) <= (inputs(147)) or (inputs(239));
    layer0_outputs(7564) <= inputs(152);
    layer0_outputs(7565) <= not(inputs(153)) or (inputs(225));
    layer0_outputs(7566) <= not(inputs(135));
    layer0_outputs(7567) <= (inputs(78)) or (inputs(189));
    layer0_outputs(7568) <= (inputs(108)) and not (inputs(192));
    layer0_outputs(7569) <= (inputs(189)) or (inputs(140));
    layer0_outputs(7570) <= inputs(6);
    layer0_outputs(7571) <= not(inputs(88));
    layer0_outputs(7572) <= not((inputs(102)) xor (inputs(42)));
    layer0_outputs(7573) <= inputs(85);
    layer0_outputs(7574) <= not(inputs(203));
    layer0_outputs(7575) <= not((inputs(148)) xor (inputs(170)));
    layer0_outputs(7576) <= (inputs(147)) or (inputs(101));
    layer0_outputs(7577) <= (inputs(188)) and not (inputs(62));
    layer0_outputs(7578) <= not(inputs(242)) or (inputs(74));
    layer0_outputs(7579) <= not(inputs(193));
    layer0_outputs(7580) <= not(inputs(235)) or (inputs(130));
    layer0_outputs(7581) <= not((inputs(103)) xor (inputs(44)));
    layer0_outputs(7582) <= (inputs(73)) xor (inputs(23));
    layer0_outputs(7583) <= not(inputs(216));
    layer0_outputs(7584) <= not(inputs(155));
    layer0_outputs(7585) <= not((inputs(240)) or (inputs(48)));
    layer0_outputs(7586) <= (inputs(213)) or (inputs(232));
    layer0_outputs(7587) <= (inputs(231)) and (inputs(92));
    layer0_outputs(7588) <= not(inputs(34));
    layer0_outputs(7589) <= not((inputs(76)) or (inputs(192)));
    layer0_outputs(7590) <= (inputs(149)) and not (inputs(251));
    layer0_outputs(7591) <= not(inputs(22));
    layer0_outputs(7592) <= not((inputs(29)) xor (inputs(76)));
    layer0_outputs(7593) <= (inputs(245)) and not (inputs(108));
    layer0_outputs(7594) <= not((inputs(139)) xor (inputs(121)));
    layer0_outputs(7595) <= not(inputs(231));
    layer0_outputs(7596) <= not(inputs(185));
    layer0_outputs(7597) <= (inputs(130)) and not (inputs(165));
    layer0_outputs(7598) <= inputs(29);
    layer0_outputs(7599) <= not(inputs(99));
    layer0_outputs(7600) <= (inputs(92)) xor (inputs(21));
    layer0_outputs(7601) <= not(inputs(67)) or (inputs(129));
    layer0_outputs(7602) <= not((inputs(241)) xor (inputs(190)));
    layer0_outputs(7603) <= not(inputs(124)) or (inputs(64));
    layer0_outputs(7604) <= not((inputs(254)) or (inputs(102)));
    layer0_outputs(7605) <= inputs(131);
    layer0_outputs(7606) <= (inputs(102)) or (inputs(229));
    layer0_outputs(7607) <= not(inputs(149)) or (inputs(78));
    layer0_outputs(7608) <= not((inputs(195)) xor (inputs(119)));
    layer0_outputs(7609) <= (inputs(79)) or (inputs(205));
    layer0_outputs(7610) <= (inputs(200)) or (inputs(182));
    layer0_outputs(7611) <= (inputs(209)) xor (inputs(232));
    layer0_outputs(7612) <= inputs(165);
    layer0_outputs(7613) <= (inputs(46)) or (inputs(49));
    layer0_outputs(7614) <= (inputs(90)) and not (inputs(180));
    layer0_outputs(7615) <= (inputs(82)) xor (inputs(210));
    layer0_outputs(7616) <= inputs(59);
    layer0_outputs(7617) <= not(inputs(114));
    layer0_outputs(7618) <= (inputs(27)) xor (inputs(195));
    layer0_outputs(7619) <= (inputs(32)) xor (inputs(49));
    layer0_outputs(7620) <= (inputs(118)) or (inputs(115));
    layer0_outputs(7621) <= (inputs(126)) xor (inputs(228));
    layer0_outputs(7622) <= not((inputs(238)) and (inputs(87)));
    layer0_outputs(7623) <= (inputs(210)) and (inputs(98));
    layer0_outputs(7624) <= not((inputs(71)) or (inputs(33)));
    layer0_outputs(7625) <= not(inputs(223)) or (inputs(102));
    layer0_outputs(7626) <= not((inputs(156)) xor (inputs(31)));
    layer0_outputs(7627) <= inputs(192);
    layer0_outputs(7628) <= not(inputs(143));
    layer0_outputs(7629) <= '1';
    layer0_outputs(7630) <= (inputs(113)) xor (inputs(217));
    layer0_outputs(7631) <= not(inputs(67)) or (inputs(38));
    layer0_outputs(7632) <= (inputs(19)) xor (inputs(94));
    layer0_outputs(7633) <= (inputs(234)) or (inputs(157));
    layer0_outputs(7634) <= not((inputs(151)) or (inputs(4)));
    layer0_outputs(7635) <= (inputs(157)) xor (inputs(93));
    layer0_outputs(7636) <= not((inputs(200)) and (inputs(198)));
    layer0_outputs(7637) <= not(inputs(21));
    layer0_outputs(7638) <= (inputs(53)) xor (inputs(131));
    layer0_outputs(7639) <= not(inputs(254)) or (inputs(208));
    layer0_outputs(7640) <= (inputs(56)) or (inputs(159));
    layer0_outputs(7641) <= not((inputs(122)) xor (inputs(12)));
    layer0_outputs(7642) <= inputs(23);
    layer0_outputs(7643) <= (inputs(40)) xor (inputs(232));
    layer0_outputs(7644) <= (inputs(111)) or (inputs(1));
    layer0_outputs(7645) <= not(inputs(111)) or (inputs(150));
    layer0_outputs(7646) <= (inputs(122)) and not (inputs(203));
    layer0_outputs(7647) <= (inputs(188)) and not (inputs(40));
    layer0_outputs(7648) <= not(inputs(132)) or (inputs(192));
    layer0_outputs(7649) <= (inputs(141)) and (inputs(249));
    layer0_outputs(7650) <= not((inputs(20)) xor (inputs(181)));
    layer0_outputs(7651) <= not(inputs(227)) or (inputs(125));
    layer0_outputs(7652) <= not((inputs(28)) xor (inputs(150)));
    layer0_outputs(7653) <= not((inputs(38)) xor (inputs(8)));
    layer0_outputs(7654) <= not(inputs(205));
    layer0_outputs(7655) <= not(inputs(52)) or (inputs(33));
    layer0_outputs(7656) <= inputs(165);
    layer0_outputs(7657) <= not((inputs(193)) or (inputs(79)));
    layer0_outputs(7658) <= inputs(233);
    layer0_outputs(7659) <= not(inputs(78));
    layer0_outputs(7660) <= inputs(112);
    layer0_outputs(7661) <= inputs(159);
    layer0_outputs(7662) <= (inputs(168)) and not (inputs(175));
    layer0_outputs(7663) <= not((inputs(198)) or (inputs(27)));
    layer0_outputs(7664) <= (inputs(124)) and not (inputs(151));
    layer0_outputs(7665) <= (inputs(182)) or (inputs(135));
    layer0_outputs(7666) <= not(inputs(246)) or (inputs(24));
    layer0_outputs(7667) <= not(inputs(158));
    layer0_outputs(7668) <= (inputs(181)) or (inputs(145));
    layer0_outputs(7669) <= (inputs(40)) and not (inputs(100));
    layer0_outputs(7670) <= (inputs(196)) or (inputs(126));
    layer0_outputs(7671) <= (inputs(208)) and not (inputs(155));
    layer0_outputs(7672) <= (inputs(156)) xor (inputs(158));
    layer0_outputs(7673) <= not((inputs(203)) or (inputs(89)));
    layer0_outputs(7674) <= not(inputs(201));
    layer0_outputs(7675) <= (inputs(136)) or (inputs(1));
    layer0_outputs(7676) <= not(inputs(42));
    layer0_outputs(7677) <= (inputs(201)) and not (inputs(33));
    layer0_outputs(7678) <= not((inputs(105)) xor (inputs(125)));
    layer0_outputs(7679) <= inputs(229);
    layer0_outputs(7680) <= (inputs(190)) xor (inputs(27));
    layer0_outputs(7681) <= not(inputs(24));
    layer0_outputs(7682) <= not((inputs(198)) xor (inputs(52)));
    layer0_outputs(7683) <= (inputs(16)) xor (inputs(136));
    layer0_outputs(7684) <= (inputs(52)) and not (inputs(92));
    layer0_outputs(7685) <= not(inputs(152)) or (inputs(208));
    layer0_outputs(7686) <= not((inputs(22)) or (inputs(149)));
    layer0_outputs(7687) <= inputs(114);
    layer0_outputs(7688) <= not((inputs(177)) or (inputs(202)));
    layer0_outputs(7689) <= not(inputs(249));
    layer0_outputs(7690) <= not(inputs(149));
    layer0_outputs(7691) <= not((inputs(171)) or (inputs(58)));
    layer0_outputs(7692) <= (inputs(128)) and (inputs(110));
    layer0_outputs(7693) <= not(inputs(23));
    layer0_outputs(7694) <= not((inputs(89)) xor (inputs(106)));
    layer0_outputs(7695) <= not(inputs(197));
    layer0_outputs(7696) <= (inputs(50)) and not (inputs(126));
    layer0_outputs(7697) <= (inputs(74)) or (inputs(123));
    layer0_outputs(7698) <= inputs(168);
    layer0_outputs(7699) <= not((inputs(163)) or (inputs(121)));
    layer0_outputs(7700) <= not(inputs(165)) or (inputs(94));
    layer0_outputs(7701) <= (inputs(239)) or (inputs(152));
    layer0_outputs(7702) <= (inputs(110)) xor (inputs(38));
    layer0_outputs(7703) <= not(inputs(213)) or (inputs(31));
    layer0_outputs(7704) <= (inputs(234)) and not (inputs(162));
    layer0_outputs(7705) <= not(inputs(62));
    layer0_outputs(7706) <= not(inputs(7));
    layer0_outputs(7707) <= not(inputs(213)) or (inputs(133));
    layer0_outputs(7708) <= not((inputs(231)) or (inputs(211)));
    layer0_outputs(7709) <= inputs(226);
    layer0_outputs(7710) <= not(inputs(186));
    layer0_outputs(7711) <= (inputs(63)) and (inputs(126));
    layer0_outputs(7712) <= not(inputs(250)) or (inputs(240));
    layer0_outputs(7713) <= not(inputs(64));
    layer0_outputs(7714) <= (inputs(194)) or (inputs(109));
    layer0_outputs(7715) <= not(inputs(187));
    layer0_outputs(7716) <= not((inputs(83)) or (inputs(132)));
    layer0_outputs(7717) <= (inputs(185)) xor (inputs(103));
    layer0_outputs(7718) <= not(inputs(75));
    layer0_outputs(7719) <= not(inputs(100));
    layer0_outputs(7720) <= inputs(236);
    layer0_outputs(7721) <= inputs(138);
    layer0_outputs(7722) <= inputs(153);
    layer0_outputs(7723) <= not(inputs(184));
    layer0_outputs(7724) <= (inputs(241)) and (inputs(117));
    layer0_outputs(7725) <= (inputs(141)) and not (inputs(81));
    layer0_outputs(7726) <= (inputs(109)) and not (inputs(10));
    layer0_outputs(7727) <= not(inputs(211)) or (inputs(114));
    layer0_outputs(7728) <= (inputs(88)) or (inputs(110));
    layer0_outputs(7729) <= not(inputs(178));
    layer0_outputs(7730) <= not((inputs(17)) or (inputs(39)));
    layer0_outputs(7731) <= '0';
    layer0_outputs(7732) <= not((inputs(114)) or (inputs(30)));
    layer0_outputs(7733) <= not(inputs(15));
    layer0_outputs(7734) <= not((inputs(233)) xor (inputs(185)));
    layer0_outputs(7735) <= not(inputs(82));
    layer0_outputs(7736) <= not(inputs(215));
    layer0_outputs(7737) <= not((inputs(2)) xor (inputs(231)));
    layer0_outputs(7738) <= not((inputs(199)) or (inputs(164)));
    layer0_outputs(7739) <= not((inputs(29)) or (inputs(131)));
    layer0_outputs(7740) <= not(inputs(109));
    layer0_outputs(7741) <= (inputs(20)) and not (inputs(226));
    layer0_outputs(7742) <= not(inputs(163));
    layer0_outputs(7743) <= not((inputs(133)) xor (inputs(117)));
    layer0_outputs(7744) <= (inputs(145)) and not (inputs(30));
    layer0_outputs(7745) <= not((inputs(42)) or (inputs(245)));
    layer0_outputs(7746) <= (inputs(224)) and (inputs(75));
    layer0_outputs(7747) <= (inputs(65)) and not (inputs(31));
    layer0_outputs(7748) <= not((inputs(89)) xor (inputs(75)));
    layer0_outputs(7749) <= not((inputs(57)) xor (inputs(30)));
    layer0_outputs(7750) <= (inputs(112)) or (inputs(172));
    layer0_outputs(7751) <= not(inputs(94)) or (inputs(201));
    layer0_outputs(7752) <= '1';
    layer0_outputs(7753) <= (inputs(233)) or (inputs(220));
    layer0_outputs(7754) <= (inputs(26)) or (inputs(62));
    layer0_outputs(7755) <= (inputs(166)) or (inputs(74));
    layer0_outputs(7756) <= not(inputs(103));
    layer0_outputs(7757) <= not((inputs(56)) xor (inputs(25)));
    layer0_outputs(7758) <= (inputs(199)) and (inputs(109));
    layer0_outputs(7759) <= (inputs(24)) or (inputs(68));
    layer0_outputs(7760) <= (inputs(20)) and not (inputs(110));
    layer0_outputs(7761) <= (inputs(155)) or (inputs(206));
    layer0_outputs(7762) <= (inputs(46)) and not (inputs(166));
    layer0_outputs(7763) <= (inputs(142)) or (inputs(149));
    layer0_outputs(7764) <= (inputs(61)) or (inputs(104));
    layer0_outputs(7765) <= not(inputs(185));
    layer0_outputs(7766) <= not((inputs(231)) xor (inputs(209)));
    layer0_outputs(7767) <= not(inputs(76));
    layer0_outputs(7768) <= not(inputs(178));
    layer0_outputs(7769) <= not(inputs(234));
    layer0_outputs(7770) <= not(inputs(118));
    layer0_outputs(7771) <= (inputs(192)) or (inputs(146));
    layer0_outputs(7772) <= not((inputs(110)) or (inputs(34)));
    layer0_outputs(7773) <= (inputs(115)) or (inputs(153));
    layer0_outputs(7774) <= not(inputs(2)) or (inputs(252));
    layer0_outputs(7775) <= (inputs(106)) or (inputs(220));
    layer0_outputs(7776) <= (inputs(11)) and (inputs(36));
    layer0_outputs(7777) <= (inputs(175)) and not (inputs(174));
    layer0_outputs(7778) <= not(inputs(77));
    layer0_outputs(7779) <= not(inputs(209));
    layer0_outputs(7780) <= not(inputs(227));
    layer0_outputs(7781) <= not((inputs(205)) or (inputs(101)));
    layer0_outputs(7782) <= not((inputs(135)) or (inputs(14)));
    layer0_outputs(7783) <= not((inputs(24)) xor (inputs(176)));
    layer0_outputs(7784) <= (inputs(58)) xor (inputs(134));
    layer0_outputs(7785) <= not((inputs(131)) or (inputs(193)));
    layer0_outputs(7786) <= not(inputs(126));
    layer0_outputs(7787) <= (inputs(217)) xor (inputs(161));
    layer0_outputs(7788) <= not(inputs(68));
    layer0_outputs(7789) <= (inputs(92)) and not (inputs(15));
    layer0_outputs(7790) <= not((inputs(102)) xor (inputs(85)));
    layer0_outputs(7791) <= not((inputs(141)) or (inputs(110)));
    layer0_outputs(7792) <= inputs(56);
    layer0_outputs(7793) <= not((inputs(196)) and (inputs(163)));
    layer0_outputs(7794) <= (inputs(118)) xor (inputs(134));
    layer0_outputs(7795) <= (inputs(219)) xor (inputs(232));
    layer0_outputs(7796) <= not(inputs(8)) or (inputs(232));
    layer0_outputs(7797) <= (inputs(171)) xor (inputs(112));
    layer0_outputs(7798) <= not((inputs(237)) or (inputs(255)));
    layer0_outputs(7799) <= (inputs(81)) xor (inputs(6));
    layer0_outputs(7800) <= (inputs(165)) xor (inputs(76));
    layer0_outputs(7801) <= inputs(101);
    layer0_outputs(7802) <= (inputs(34)) or (inputs(235));
    layer0_outputs(7803) <= not((inputs(72)) xor (inputs(201)));
    layer0_outputs(7804) <= not(inputs(237)) or (inputs(109));
    layer0_outputs(7805) <= (inputs(181)) xor (inputs(216));
    layer0_outputs(7806) <= inputs(240);
    layer0_outputs(7807) <= not((inputs(170)) or (inputs(59)));
    layer0_outputs(7808) <= (inputs(252)) or (inputs(154));
    layer0_outputs(7809) <= not(inputs(211)) or (inputs(70));
    layer0_outputs(7810) <= not((inputs(208)) or (inputs(49)));
    layer0_outputs(7811) <= not((inputs(203)) xor (inputs(49)));
    layer0_outputs(7812) <= not((inputs(14)) or (inputs(250)));
    layer0_outputs(7813) <= inputs(181);
    layer0_outputs(7814) <= '0';
    layer0_outputs(7815) <= not((inputs(152)) or (inputs(200)));
    layer0_outputs(7816) <= not((inputs(199)) xor (inputs(148)));
    layer0_outputs(7817) <= not(inputs(233)) or (inputs(31));
    layer0_outputs(7818) <= (inputs(192)) or (inputs(188));
    layer0_outputs(7819) <= not(inputs(37));
    layer0_outputs(7820) <= (inputs(112)) or (inputs(163));
    layer0_outputs(7821) <= (inputs(121)) or (inputs(122));
    layer0_outputs(7822) <= not(inputs(165));
    layer0_outputs(7823) <= not((inputs(26)) and (inputs(200)));
    layer0_outputs(7824) <= not((inputs(227)) or (inputs(20)));
    layer0_outputs(7825) <= (inputs(121)) or (inputs(20));
    layer0_outputs(7826) <= not((inputs(172)) or (inputs(237)));
    layer0_outputs(7827) <= not(inputs(213)) or (inputs(240));
    layer0_outputs(7828) <= (inputs(94)) or (inputs(41));
    layer0_outputs(7829) <= not(inputs(91));
    layer0_outputs(7830) <= inputs(116);
    layer0_outputs(7831) <= inputs(187);
    layer0_outputs(7832) <= inputs(163);
    layer0_outputs(7833) <= not(inputs(12));
    layer0_outputs(7834) <= not(inputs(66)) or (inputs(255));
    layer0_outputs(7835) <= not((inputs(7)) xor (inputs(70)));
    layer0_outputs(7836) <= not(inputs(184)) or (inputs(94));
    layer0_outputs(7837) <= not(inputs(7)) or (inputs(16));
    layer0_outputs(7838) <= not(inputs(174));
    layer0_outputs(7839) <= inputs(233);
    layer0_outputs(7840) <= (inputs(24)) and not (inputs(141));
    layer0_outputs(7841) <= inputs(97);
    layer0_outputs(7842) <= (inputs(217)) and not (inputs(76));
    layer0_outputs(7843) <= inputs(10);
    layer0_outputs(7844) <= (inputs(204)) or (inputs(145));
    layer0_outputs(7845) <= (inputs(200)) and (inputs(181));
    layer0_outputs(7846) <= not((inputs(154)) xor (inputs(184)));
    layer0_outputs(7847) <= not((inputs(64)) xor (inputs(122)));
    layer0_outputs(7848) <= (inputs(136)) and not (inputs(196));
    layer0_outputs(7849) <= (inputs(100)) and not (inputs(55));
    layer0_outputs(7850) <= (inputs(83)) or (inputs(65));
    layer0_outputs(7851) <= '1';
    layer0_outputs(7852) <= not((inputs(89)) and (inputs(90)));
    layer0_outputs(7853) <= not(inputs(178));
    layer0_outputs(7854) <= not((inputs(16)) and (inputs(75)));
    layer0_outputs(7855) <= not(inputs(119));
    layer0_outputs(7856) <= (inputs(88)) or (inputs(207));
    layer0_outputs(7857) <= (inputs(53)) and not (inputs(17));
    layer0_outputs(7858) <= not(inputs(81)) or (inputs(126));
    layer0_outputs(7859) <= inputs(124);
    layer0_outputs(7860) <= not(inputs(37)) or (inputs(200));
    layer0_outputs(7861) <= not((inputs(183)) xor (inputs(190)));
    layer0_outputs(7862) <= inputs(209);
    layer0_outputs(7863) <= not((inputs(129)) or (inputs(125)));
    layer0_outputs(7864) <= '0';
    layer0_outputs(7865) <= (inputs(188)) xor (inputs(154));
    layer0_outputs(7866) <= (inputs(65)) or (inputs(145));
    layer0_outputs(7867) <= (inputs(139)) and not (inputs(205));
    layer0_outputs(7868) <= (inputs(8)) xor (inputs(122));
    layer0_outputs(7869) <= not(inputs(89));
    layer0_outputs(7870) <= (inputs(42)) and not (inputs(95));
    layer0_outputs(7871) <= not(inputs(163));
    layer0_outputs(7872) <= not(inputs(181)) or (inputs(46));
    layer0_outputs(7873) <= inputs(168);
    layer0_outputs(7874) <= not(inputs(194)) or (inputs(2));
    layer0_outputs(7875) <= not(inputs(210));
    layer0_outputs(7876) <= inputs(236);
    layer0_outputs(7877) <= (inputs(74)) and not (inputs(176));
    layer0_outputs(7878) <= not((inputs(79)) xor (inputs(88)));
    layer0_outputs(7879) <= not(inputs(91));
    layer0_outputs(7880) <= not((inputs(70)) xor (inputs(18)));
    layer0_outputs(7881) <= not(inputs(88));
    layer0_outputs(7882) <= not((inputs(206)) or (inputs(181)));
    layer0_outputs(7883) <= inputs(113);
    layer0_outputs(7884) <= not((inputs(57)) or (inputs(96)));
    layer0_outputs(7885) <= (inputs(49)) or (inputs(144));
    layer0_outputs(7886) <= inputs(136);
    layer0_outputs(7887) <= not((inputs(73)) xor (inputs(209)));
    layer0_outputs(7888) <= not(inputs(98));
    layer0_outputs(7889) <= not((inputs(151)) or (inputs(115)));
    layer0_outputs(7890) <= inputs(132);
    layer0_outputs(7891) <= not(inputs(59));
    layer0_outputs(7892) <= not((inputs(68)) and (inputs(30)));
    layer0_outputs(7893) <= (inputs(122)) or (inputs(181));
    layer0_outputs(7894) <= (inputs(31)) or (inputs(213));
    layer0_outputs(7895) <= not((inputs(195)) or (inputs(111)));
    layer0_outputs(7896) <= inputs(188);
    layer0_outputs(7897) <= (inputs(129)) or (inputs(203));
    layer0_outputs(7898) <= (inputs(125)) or (inputs(4));
    layer0_outputs(7899) <= inputs(13);
    layer0_outputs(7900) <= not(inputs(236)) or (inputs(129));
    layer0_outputs(7901) <= not((inputs(204)) or (inputs(238)));
    layer0_outputs(7902) <= (inputs(94)) xor (inputs(90));
    layer0_outputs(7903) <= (inputs(131)) and not (inputs(98));
    layer0_outputs(7904) <= (inputs(119)) and not (inputs(122));
    layer0_outputs(7905) <= not(inputs(23));
    layer0_outputs(7906) <= inputs(188);
    layer0_outputs(7907) <= inputs(195);
    layer0_outputs(7908) <= inputs(65);
    layer0_outputs(7909) <= (inputs(62)) xor (inputs(125));
    layer0_outputs(7910) <= (inputs(23)) and not (inputs(32));
    layer0_outputs(7911) <= inputs(77);
    layer0_outputs(7912) <= (inputs(237)) or (inputs(202));
    layer0_outputs(7913) <= not((inputs(45)) xor (inputs(116)));
    layer0_outputs(7914) <= (inputs(41)) or (inputs(242));
    layer0_outputs(7915) <= not(inputs(229)) or (inputs(6));
    layer0_outputs(7916) <= not((inputs(86)) xor (inputs(117)));
    layer0_outputs(7917) <= inputs(76);
    layer0_outputs(7918) <= not(inputs(123));
    layer0_outputs(7919) <= not(inputs(89)) or (inputs(51));
    layer0_outputs(7920) <= inputs(161);
    layer0_outputs(7921) <= (inputs(119)) xor (inputs(103));
    layer0_outputs(7922) <= inputs(20);
    layer0_outputs(7923) <= (inputs(160)) xor (inputs(162));
    layer0_outputs(7924) <= inputs(17);
    layer0_outputs(7925) <= not((inputs(90)) or (inputs(64)));
    layer0_outputs(7926) <= not((inputs(31)) or (inputs(39)));
    layer0_outputs(7927) <= not((inputs(248)) or (inputs(228)));
    layer0_outputs(7928) <= not(inputs(167)) or (inputs(30));
    layer0_outputs(7929) <= not((inputs(97)) or (inputs(156)));
    layer0_outputs(7930) <= not(inputs(236));
    layer0_outputs(7931) <= (inputs(171)) or (inputs(219));
    layer0_outputs(7932) <= (inputs(221)) xor (inputs(115));
    layer0_outputs(7933) <= not((inputs(64)) xor (inputs(37)));
    layer0_outputs(7934) <= (inputs(184)) xor (inputs(147));
    layer0_outputs(7935) <= not(inputs(218));
    layer0_outputs(7936) <= not(inputs(157));
    layer0_outputs(7937) <= not((inputs(191)) or (inputs(73)));
    layer0_outputs(7938) <= not((inputs(203)) xor (inputs(253)));
    layer0_outputs(7939) <= not((inputs(174)) or (inputs(6)));
    layer0_outputs(7940) <= (inputs(51)) and not (inputs(96));
    layer0_outputs(7941) <= inputs(89);
    layer0_outputs(7942) <= inputs(164);
    layer0_outputs(7943) <= not(inputs(7));
    layer0_outputs(7944) <= not(inputs(28));
    layer0_outputs(7945) <= (inputs(41)) and not (inputs(194));
    layer0_outputs(7946) <= inputs(253);
    layer0_outputs(7947) <= not((inputs(223)) or (inputs(100)));
    layer0_outputs(7948) <= (inputs(205)) and not (inputs(186));
    layer0_outputs(7949) <= (inputs(218)) xor (inputs(163));
    layer0_outputs(7950) <= not((inputs(203)) xor (inputs(190)));
    layer0_outputs(7951) <= (inputs(229)) and not (inputs(104));
    layer0_outputs(7952) <= not(inputs(165)) or (inputs(15));
    layer0_outputs(7953) <= not((inputs(71)) and (inputs(67)));
    layer0_outputs(7954) <= (inputs(204)) and not (inputs(125));
    layer0_outputs(7955) <= (inputs(73)) and not (inputs(126));
    layer0_outputs(7956) <= (inputs(95)) xor (inputs(175));
    layer0_outputs(7957) <= not(inputs(105)) or (inputs(234));
    layer0_outputs(7958) <= not((inputs(202)) and (inputs(0)));
    layer0_outputs(7959) <= (inputs(216)) or (inputs(231));
    layer0_outputs(7960) <= (inputs(193)) or (inputs(107));
    layer0_outputs(7961) <= not(inputs(63));
    layer0_outputs(7962) <= (inputs(204)) or (inputs(140));
    layer0_outputs(7963) <= (inputs(34)) xor (inputs(188));
    layer0_outputs(7964) <= not((inputs(16)) xor (inputs(247)));
    layer0_outputs(7965) <= (inputs(134)) and not (inputs(95));
    layer0_outputs(7966) <= not(inputs(102));
    layer0_outputs(7967) <= (inputs(248)) xor (inputs(204));
    layer0_outputs(7968) <= not(inputs(43));
    layer0_outputs(7969) <= inputs(205);
    layer0_outputs(7970) <= not((inputs(244)) xor (inputs(247)));
    layer0_outputs(7971) <= not(inputs(62)) or (inputs(42));
    layer0_outputs(7972) <= inputs(241);
    layer0_outputs(7973) <= (inputs(170)) or (inputs(223));
    layer0_outputs(7974) <= not(inputs(222));
    layer0_outputs(7975) <= inputs(38);
    layer0_outputs(7976) <= not((inputs(223)) and (inputs(9)));
    layer0_outputs(7977) <= inputs(40);
    layer0_outputs(7978) <= (inputs(237)) and not (inputs(188));
    layer0_outputs(7979) <= (inputs(132)) and not (inputs(225));
    layer0_outputs(7980) <= inputs(178);
    layer0_outputs(7981) <= (inputs(193)) xor (inputs(133));
    layer0_outputs(7982) <= (inputs(50)) or (inputs(32));
    layer0_outputs(7983) <= inputs(196);
    layer0_outputs(7984) <= not(inputs(71));
    layer0_outputs(7985) <= (inputs(102)) or (inputs(81));
    layer0_outputs(7986) <= (inputs(25)) and not (inputs(251));
    layer0_outputs(7987) <= (inputs(154)) or (inputs(63));
    layer0_outputs(7988) <= (inputs(35)) and not (inputs(73));
    layer0_outputs(7989) <= (inputs(69)) and not (inputs(166));
    layer0_outputs(7990) <= not((inputs(173)) or (inputs(217)));
    layer0_outputs(7991) <= not(inputs(157));
    layer0_outputs(7992) <= (inputs(161)) and not (inputs(77));
    layer0_outputs(7993) <= not(inputs(122));
    layer0_outputs(7994) <= (inputs(17)) or (inputs(200));
    layer0_outputs(7995) <= not(inputs(243));
    layer0_outputs(7996) <= not((inputs(33)) xor (inputs(189)));
    layer0_outputs(7997) <= (inputs(59)) or (inputs(62));
    layer0_outputs(7998) <= not(inputs(130));
    layer0_outputs(7999) <= not((inputs(242)) or (inputs(142)));
    layer0_outputs(8000) <= not(inputs(149));
    layer0_outputs(8001) <= not(inputs(117)) or (inputs(29));
    layer0_outputs(8002) <= (inputs(94)) or (inputs(53));
    layer0_outputs(8003) <= (inputs(16)) and not (inputs(253));
    layer0_outputs(8004) <= inputs(186);
    layer0_outputs(8005) <= not(inputs(216));
    layer0_outputs(8006) <= inputs(23);
    layer0_outputs(8007) <= (inputs(138)) and (inputs(173));
    layer0_outputs(8008) <= inputs(166);
    layer0_outputs(8009) <= not((inputs(65)) or (inputs(114)));
    layer0_outputs(8010) <= (inputs(143)) or (inputs(225));
    layer0_outputs(8011) <= '1';
    layer0_outputs(8012) <= not(inputs(41));
    layer0_outputs(8013) <= inputs(9);
    layer0_outputs(8014) <= not(inputs(167)) or (inputs(223));
    layer0_outputs(8015) <= (inputs(151)) or (inputs(67));
    layer0_outputs(8016) <= not(inputs(157)) or (inputs(118));
    layer0_outputs(8017) <= not(inputs(156));
    layer0_outputs(8018) <= inputs(219);
    layer0_outputs(8019) <= not((inputs(123)) or (inputs(42)));
    layer0_outputs(8020) <= not(inputs(27)) or (inputs(143));
    layer0_outputs(8021) <= '1';
    layer0_outputs(8022) <= (inputs(220)) or (inputs(64));
    layer0_outputs(8023) <= (inputs(198)) and not (inputs(147));
    layer0_outputs(8024) <= (inputs(68)) and not (inputs(192));
    layer0_outputs(8025) <= (inputs(114)) and (inputs(227));
    layer0_outputs(8026) <= not(inputs(129));
    layer0_outputs(8027) <= not(inputs(137)) or (inputs(249));
    layer0_outputs(8028) <= (inputs(73)) and not (inputs(224));
    layer0_outputs(8029) <= not(inputs(243)) or (inputs(78));
    layer0_outputs(8030) <= not(inputs(204));
    layer0_outputs(8031) <= not(inputs(214)) or (inputs(4));
    layer0_outputs(8032) <= (inputs(218)) or (inputs(251));
    layer0_outputs(8033) <= (inputs(2)) or (inputs(200));
    layer0_outputs(8034) <= not(inputs(34)) or (inputs(144));
    layer0_outputs(8035) <= not(inputs(171)) or (inputs(77));
    layer0_outputs(8036) <= (inputs(183)) and not (inputs(172));
    layer0_outputs(8037) <= (inputs(149)) and not (inputs(138));
    layer0_outputs(8038) <= inputs(100);
    layer0_outputs(8039) <= (inputs(226)) xor (inputs(236));
    layer0_outputs(8040) <= (inputs(122)) and not (inputs(250));
    layer0_outputs(8041) <= inputs(5);
    layer0_outputs(8042) <= (inputs(162)) and not (inputs(18));
    layer0_outputs(8043) <= inputs(155);
    layer0_outputs(8044) <= not((inputs(211)) or (inputs(100)));
    layer0_outputs(8045) <= not(inputs(10));
    layer0_outputs(8046) <= (inputs(204)) or (inputs(229));
    layer0_outputs(8047) <= inputs(62);
    layer0_outputs(8048) <= not(inputs(20)) or (inputs(241));
    layer0_outputs(8049) <= not((inputs(163)) or (inputs(180)));
    layer0_outputs(8050) <= (inputs(206)) xor (inputs(219));
    layer0_outputs(8051) <= not(inputs(184)) or (inputs(107));
    layer0_outputs(8052) <= not((inputs(66)) or (inputs(47)));
    layer0_outputs(8053) <= (inputs(63)) and not (inputs(68));
    layer0_outputs(8054) <= inputs(142);
    layer0_outputs(8055) <= not((inputs(249)) or (inputs(142)));
    layer0_outputs(8056) <= not(inputs(181)) or (inputs(139));
    layer0_outputs(8057) <= (inputs(26)) xor (inputs(81));
    layer0_outputs(8058) <= not(inputs(116));
    layer0_outputs(8059) <= not(inputs(238));
    layer0_outputs(8060) <= inputs(218);
    layer0_outputs(8061) <= (inputs(197)) xor (inputs(23));
    layer0_outputs(8062) <= not(inputs(66));
    layer0_outputs(8063) <= inputs(171);
    layer0_outputs(8064) <= not(inputs(184)) or (inputs(123));
    layer0_outputs(8065) <= not((inputs(60)) xor (inputs(124)));
    layer0_outputs(8066) <= not((inputs(44)) or (inputs(81)));
    layer0_outputs(8067) <= (inputs(179)) or (inputs(203));
    layer0_outputs(8068) <= (inputs(101)) or (inputs(180));
    layer0_outputs(8069) <= (inputs(147)) or (inputs(84));
    layer0_outputs(8070) <= (inputs(227)) xor (inputs(205));
    layer0_outputs(8071) <= not((inputs(45)) or (inputs(248)));
    layer0_outputs(8072) <= inputs(208);
    layer0_outputs(8073) <= (inputs(208)) xor (inputs(175));
    layer0_outputs(8074) <= not(inputs(90));
    layer0_outputs(8075) <= not((inputs(207)) or (inputs(3)));
    layer0_outputs(8076) <= (inputs(133)) and not (inputs(126));
    layer0_outputs(8077) <= not(inputs(122));
    layer0_outputs(8078) <= (inputs(28)) and not (inputs(185));
    layer0_outputs(8079) <= not((inputs(128)) xor (inputs(11)));
    layer0_outputs(8080) <= inputs(109);
    layer0_outputs(8081) <= inputs(50);
    layer0_outputs(8082) <= not((inputs(175)) and (inputs(169)));
    layer0_outputs(8083) <= not((inputs(132)) xor (inputs(179)));
    layer0_outputs(8084) <= (inputs(57)) and not (inputs(225));
    layer0_outputs(8085) <= inputs(125);
    layer0_outputs(8086) <= '1';
    layer0_outputs(8087) <= not(inputs(162));
    layer0_outputs(8088) <= not(inputs(213));
    layer0_outputs(8089) <= (inputs(66)) or (inputs(50));
    layer0_outputs(8090) <= not(inputs(36));
    layer0_outputs(8091) <= (inputs(53)) and not (inputs(250));
    layer0_outputs(8092) <= not(inputs(75));
    layer0_outputs(8093) <= not((inputs(157)) or (inputs(247)));
    layer0_outputs(8094) <= (inputs(60)) xor (inputs(148));
    layer0_outputs(8095) <= not((inputs(72)) xor (inputs(115)));
    layer0_outputs(8096) <= not((inputs(216)) or (inputs(4)));
    layer0_outputs(8097) <= not((inputs(76)) or (inputs(36)));
    layer0_outputs(8098) <= not(inputs(186));
    layer0_outputs(8099) <= inputs(201);
    layer0_outputs(8100) <= inputs(54);
    layer0_outputs(8101) <= not((inputs(250)) or (inputs(234)));
    layer0_outputs(8102) <= not(inputs(148));
    layer0_outputs(8103) <= not((inputs(118)) xor (inputs(135)));
    layer0_outputs(8104) <= not(inputs(4)) or (inputs(112));
    layer0_outputs(8105) <= (inputs(48)) xor (inputs(150));
    layer0_outputs(8106) <= (inputs(37)) and not (inputs(235));
    layer0_outputs(8107) <= not((inputs(244)) or (inputs(9)));
    layer0_outputs(8108) <= inputs(134);
    layer0_outputs(8109) <= not(inputs(122));
    layer0_outputs(8110) <= not(inputs(171)) or (inputs(254));
    layer0_outputs(8111) <= (inputs(22)) and not (inputs(195));
    layer0_outputs(8112) <= inputs(92);
    layer0_outputs(8113) <= (inputs(218)) and not (inputs(3));
    layer0_outputs(8114) <= (inputs(183)) or (inputs(197));
    layer0_outputs(8115) <= not(inputs(231));
    layer0_outputs(8116) <= not((inputs(85)) xor (inputs(207)));
    layer0_outputs(8117) <= inputs(188);
    layer0_outputs(8118) <= (inputs(44)) or (inputs(210));
    layer0_outputs(8119) <= inputs(102);
    layer0_outputs(8120) <= (inputs(143)) and (inputs(77));
    layer0_outputs(8121) <= not(inputs(55));
    layer0_outputs(8122) <= inputs(200);
    layer0_outputs(8123) <= not((inputs(27)) xor (inputs(138)));
    layer0_outputs(8124) <= not((inputs(143)) or (inputs(132)));
    layer0_outputs(8125) <= not((inputs(147)) or (inputs(75)));
    layer0_outputs(8126) <= not(inputs(43)) or (inputs(239));
    layer0_outputs(8127) <= not((inputs(40)) or (inputs(194)));
    layer0_outputs(8128) <= not((inputs(222)) xor (inputs(99)));
    layer0_outputs(8129) <= (inputs(88)) xor (inputs(225));
    layer0_outputs(8130) <= (inputs(193)) xor (inputs(123));
    layer0_outputs(8131) <= not((inputs(123)) or (inputs(97)));
    layer0_outputs(8132) <= not(inputs(23)) or (inputs(95));
    layer0_outputs(8133) <= (inputs(218)) or (inputs(205));
    layer0_outputs(8134) <= (inputs(139)) xor (inputs(73));
    layer0_outputs(8135) <= (inputs(255)) xor (inputs(43));
    layer0_outputs(8136) <= not((inputs(183)) or (inputs(206)));
    layer0_outputs(8137) <= (inputs(143)) and not (inputs(240));
    layer0_outputs(8138) <= not(inputs(246)) or (inputs(16));
    layer0_outputs(8139) <= not((inputs(128)) and (inputs(145)));
    layer0_outputs(8140) <= inputs(230);
    layer0_outputs(8141) <= not((inputs(105)) xor (inputs(174)));
    layer0_outputs(8142) <= (inputs(246)) or (inputs(245));
    layer0_outputs(8143) <= (inputs(149)) or (inputs(175));
    layer0_outputs(8144) <= (inputs(108)) and (inputs(139));
    layer0_outputs(8145) <= not(inputs(220));
    layer0_outputs(8146) <= not((inputs(68)) or (inputs(120)));
    layer0_outputs(8147) <= not(inputs(179));
    layer0_outputs(8148) <= not((inputs(27)) xor (inputs(176)));
    layer0_outputs(8149) <= (inputs(82)) and not (inputs(240));
    layer0_outputs(8150) <= not((inputs(0)) xor (inputs(64)));
    layer0_outputs(8151) <= not(inputs(23)) or (inputs(162));
    layer0_outputs(8152) <= inputs(129);
    layer0_outputs(8153) <= not(inputs(231));
    layer0_outputs(8154) <= inputs(82);
    layer0_outputs(8155) <= (inputs(91)) and (inputs(217));
    layer0_outputs(8156) <= not((inputs(6)) or (inputs(0)));
    layer0_outputs(8157) <= not(inputs(192));
    layer0_outputs(8158) <= not(inputs(116)) or (inputs(216));
    layer0_outputs(8159) <= (inputs(178)) or (inputs(160));
    layer0_outputs(8160) <= (inputs(69)) xor (inputs(140));
    layer0_outputs(8161) <= (inputs(242)) xor (inputs(133));
    layer0_outputs(8162) <= not(inputs(215));
    layer0_outputs(8163) <= not(inputs(28));
    layer0_outputs(8164) <= (inputs(154)) or (inputs(75));
    layer0_outputs(8165) <= not(inputs(83)) or (inputs(207));
    layer0_outputs(8166) <= (inputs(55)) xor (inputs(252));
    layer0_outputs(8167) <= not(inputs(58)) or (inputs(225));
    layer0_outputs(8168) <= not(inputs(101)) or (inputs(235));
    layer0_outputs(8169) <= not(inputs(52));
    layer0_outputs(8170) <= not((inputs(3)) xor (inputs(116)));
    layer0_outputs(8171) <= inputs(180);
    layer0_outputs(8172) <= (inputs(233)) and (inputs(59));
    layer0_outputs(8173) <= not(inputs(10));
    layer0_outputs(8174) <= not(inputs(52));
    layer0_outputs(8175) <= (inputs(139)) and (inputs(228));
    layer0_outputs(8176) <= (inputs(23)) and (inputs(121));
    layer0_outputs(8177) <= (inputs(77)) xor (inputs(124));
    layer0_outputs(8178) <= not(inputs(107)) or (inputs(150));
    layer0_outputs(8179) <= not((inputs(152)) xor (inputs(56)));
    layer0_outputs(8180) <= (inputs(63)) or (inputs(221));
    layer0_outputs(8181) <= not((inputs(227)) or (inputs(86)));
    layer0_outputs(8182) <= not(inputs(112));
    layer0_outputs(8183) <= inputs(202);
    layer0_outputs(8184) <= not((inputs(79)) or (inputs(34)));
    layer0_outputs(8185) <= inputs(137);
    layer0_outputs(8186) <= inputs(215);
    layer0_outputs(8187) <= not(inputs(76));
    layer0_outputs(8188) <= (inputs(215)) and not (inputs(84));
    layer0_outputs(8189) <= inputs(179);
    layer0_outputs(8190) <= inputs(11);
    layer0_outputs(8191) <= not((inputs(220)) xor (inputs(210)));
    layer0_outputs(8192) <= not(inputs(69));
    layer0_outputs(8193) <= not(inputs(218)) or (inputs(61));
    layer0_outputs(8194) <= not(inputs(89));
    layer0_outputs(8195) <= (inputs(80)) or (inputs(179));
    layer0_outputs(8196) <= not((inputs(172)) xor (inputs(158)));
    layer0_outputs(8197) <= inputs(183);
    layer0_outputs(8198) <= not(inputs(145)) or (inputs(207));
    layer0_outputs(8199) <= not(inputs(55)) or (inputs(121));
    layer0_outputs(8200) <= (inputs(148)) and not (inputs(52));
    layer0_outputs(8201) <= (inputs(95)) xor (inputs(229));
    layer0_outputs(8202) <= (inputs(70)) and not (inputs(156));
    layer0_outputs(8203) <= (inputs(7)) or (inputs(166));
    layer0_outputs(8204) <= inputs(113);
    layer0_outputs(8205) <= not((inputs(195)) or (inputs(187)));
    layer0_outputs(8206) <= not(inputs(186)) or (inputs(159));
    layer0_outputs(8207) <= (inputs(62)) xor (inputs(46));
    layer0_outputs(8208) <= (inputs(85)) and not (inputs(33));
    layer0_outputs(8209) <= not(inputs(81));
    layer0_outputs(8210) <= not((inputs(58)) xor (inputs(221)));
    layer0_outputs(8211) <= not(inputs(181));
    layer0_outputs(8212) <= not(inputs(192));
    layer0_outputs(8213) <= not((inputs(252)) or (inputs(130)));
    layer0_outputs(8214) <= (inputs(121)) xor (inputs(119));
    layer0_outputs(8215) <= not(inputs(90));
    layer0_outputs(8216) <= (inputs(23)) or (inputs(252));
    layer0_outputs(8217) <= not((inputs(13)) or (inputs(148)));
    layer0_outputs(8218) <= '1';
    layer0_outputs(8219) <= (inputs(81)) or (inputs(111));
    layer0_outputs(8220) <= not(inputs(59));
    layer0_outputs(8221) <= (inputs(147)) and not (inputs(182));
    layer0_outputs(8222) <= inputs(205);
    layer0_outputs(8223) <= not(inputs(217)) or (inputs(49));
    layer0_outputs(8224) <= not((inputs(193)) or (inputs(99)));
    layer0_outputs(8225) <= inputs(211);
    layer0_outputs(8226) <= not(inputs(162));
    layer0_outputs(8227) <= not((inputs(47)) xor (inputs(222)));
    layer0_outputs(8228) <= inputs(22);
    layer0_outputs(8229) <= (inputs(75)) and (inputs(9));
    layer0_outputs(8230) <= inputs(126);
    layer0_outputs(8231) <= '0';
    layer0_outputs(8232) <= not(inputs(66));
    layer0_outputs(8233) <= not((inputs(145)) or (inputs(176)));
    layer0_outputs(8234) <= not((inputs(220)) or (inputs(68)));
    layer0_outputs(8235) <= (inputs(228)) and not (inputs(143));
    layer0_outputs(8236) <= not(inputs(212));
    layer0_outputs(8237) <= (inputs(97)) or (inputs(250));
    layer0_outputs(8238) <= (inputs(188)) and not (inputs(86));
    layer0_outputs(8239) <= not((inputs(9)) or (inputs(195)));
    layer0_outputs(8240) <= (inputs(137)) xor (inputs(80));
    layer0_outputs(8241) <= inputs(96);
    layer0_outputs(8242) <= not(inputs(91));
    layer0_outputs(8243) <= not((inputs(189)) xor (inputs(135)));
    layer0_outputs(8244) <= not((inputs(147)) or (inputs(109)));
    layer0_outputs(8245) <= (inputs(177)) xor (inputs(88));
    layer0_outputs(8246) <= (inputs(33)) xor (inputs(12));
    layer0_outputs(8247) <= not(inputs(162));
    layer0_outputs(8248) <= not(inputs(54));
    layer0_outputs(8249) <= inputs(91);
    layer0_outputs(8250) <= inputs(105);
    layer0_outputs(8251) <= not((inputs(206)) xor (inputs(199)));
    layer0_outputs(8252) <= (inputs(105)) or (inputs(30));
    layer0_outputs(8253) <= inputs(27);
    layer0_outputs(8254) <= not((inputs(2)) or (inputs(131)));
    layer0_outputs(8255) <= not(inputs(200));
    layer0_outputs(8256) <= not((inputs(69)) xor (inputs(81)));
    layer0_outputs(8257) <= not(inputs(30));
    layer0_outputs(8258) <= (inputs(21)) xor (inputs(162));
    layer0_outputs(8259) <= inputs(247);
    layer0_outputs(8260) <= not(inputs(247));
    layer0_outputs(8261) <= not(inputs(115));
    layer0_outputs(8262) <= (inputs(73)) or (inputs(60));
    layer0_outputs(8263) <= inputs(75);
    layer0_outputs(8264) <= not(inputs(12));
    layer0_outputs(8265) <= inputs(98);
    layer0_outputs(8266) <= not(inputs(89));
    layer0_outputs(8267) <= inputs(239);
    layer0_outputs(8268) <= not(inputs(38)) or (inputs(237));
    layer0_outputs(8269) <= (inputs(92)) and not (inputs(34));
    layer0_outputs(8270) <= inputs(154);
    layer0_outputs(8271) <= not((inputs(194)) or (inputs(49)));
    layer0_outputs(8272) <= '0';
    layer0_outputs(8273) <= not((inputs(5)) and (inputs(58)));
    layer0_outputs(8274) <= (inputs(213)) and not (inputs(13));
    layer0_outputs(8275) <= (inputs(217)) and not (inputs(97));
    layer0_outputs(8276) <= not((inputs(58)) xor (inputs(40)));
    layer0_outputs(8277) <= inputs(167);
    layer0_outputs(8278) <= not(inputs(183));
    layer0_outputs(8279) <= not((inputs(150)) or (inputs(190)));
    layer0_outputs(8280) <= (inputs(229)) and not (inputs(223));
    layer0_outputs(8281) <= (inputs(111)) xor (inputs(79));
    layer0_outputs(8282) <= inputs(167);
    layer0_outputs(8283) <= not(inputs(199));
    layer0_outputs(8284) <= not((inputs(245)) or (inputs(207)));
    layer0_outputs(8285) <= not(inputs(193)) or (inputs(123));
    layer0_outputs(8286) <= not(inputs(155));
    layer0_outputs(8287) <= (inputs(71)) and not (inputs(63));
    layer0_outputs(8288) <= inputs(123);
    layer0_outputs(8289) <= (inputs(72)) and not (inputs(143));
    layer0_outputs(8290) <= (inputs(255)) xor (inputs(133));
    layer0_outputs(8291) <= not((inputs(5)) or (inputs(113)));
    layer0_outputs(8292) <= not((inputs(23)) xor (inputs(237)));
    layer0_outputs(8293) <= not(inputs(38));
    layer0_outputs(8294) <= (inputs(244)) and not (inputs(63));
    layer0_outputs(8295) <= not(inputs(117)) or (inputs(240));
    layer0_outputs(8296) <= not(inputs(234));
    layer0_outputs(8297) <= not(inputs(203)) or (inputs(28));
    layer0_outputs(8298) <= (inputs(72)) xor (inputs(211));
    layer0_outputs(8299) <= '1';
    layer0_outputs(8300) <= not(inputs(106)) or (inputs(155));
    layer0_outputs(8301) <= not((inputs(112)) xor (inputs(124)));
    layer0_outputs(8302) <= not(inputs(10));
    layer0_outputs(8303) <= inputs(1);
    layer0_outputs(8304) <= not((inputs(128)) and (inputs(207)));
    layer0_outputs(8305) <= inputs(85);
    layer0_outputs(8306) <= (inputs(72)) and (inputs(119));
    layer0_outputs(8307) <= (inputs(170)) and (inputs(78));
    layer0_outputs(8308) <= not((inputs(40)) and (inputs(55)));
    layer0_outputs(8309) <= (inputs(3)) xor (inputs(103));
    layer0_outputs(8310) <= not((inputs(6)) or (inputs(209)));
    layer0_outputs(8311) <= not(inputs(214)) or (inputs(7));
    layer0_outputs(8312) <= (inputs(40)) and not (inputs(242));
    layer0_outputs(8313) <= (inputs(147)) and not (inputs(225));
    layer0_outputs(8314) <= inputs(151);
    layer0_outputs(8315) <= not(inputs(252)) or (inputs(48));
    layer0_outputs(8316) <= (inputs(183)) and not (inputs(150));
    layer0_outputs(8317) <= (inputs(142)) and not (inputs(113));
    layer0_outputs(8318) <= (inputs(247)) and not (inputs(239));
    layer0_outputs(8319) <= (inputs(183)) xor (inputs(76));
    layer0_outputs(8320) <= not((inputs(110)) xor (inputs(107)));
    layer0_outputs(8321) <= (inputs(41)) and (inputs(43));
    layer0_outputs(8322) <= (inputs(152)) and not (inputs(141));
    layer0_outputs(8323) <= not(inputs(135)) or (inputs(23));
    layer0_outputs(8324) <= not(inputs(193)) or (inputs(32));
    layer0_outputs(8325) <= (inputs(5)) xor (inputs(240));
    layer0_outputs(8326) <= (inputs(135)) or (inputs(254));
    layer0_outputs(8327) <= not(inputs(151)) or (inputs(75));
    layer0_outputs(8328) <= (inputs(30)) or (inputs(105));
    layer0_outputs(8329) <= not(inputs(164));
    layer0_outputs(8330) <= (inputs(184)) and not (inputs(76));
    layer0_outputs(8331) <= not((inputs(2)) or (inputs(127)));
    layer0_outputs(8332) <= (inputs(143)) or (inputs(189));
    layer0_outputs(8333) <= (inputs(188)) xor (inputs(190));
    layer0_outputs(8334) <= not(inputs(210));
    layer0_outputs(8335) <= inputs(72);
    layer0_outputs(8336) <= (inputs(178)) xor (inputs(202));
    layer0_outputs(8337) <= not(inputs(120)) or (inputs(202));
    layer0_outputs(8338) <= not(inputs(77)) or (inputs(15));
    layer0_outputs(8339) <= not((inputs(215)) or (inputs(131)));
    layer0_outputs(8340) <= not(inputs(114));
    layer0_outputs(8341) <= not(inputs(156));
    layer0_outputs(8342) <= inputs(165);
    layer0_outputs(8343) <= not((inputs(116)) or (inputs(50)));
    layer0_outputs(8344) <= (inputs(108)) xor (inputs(192));
    layer0_outputs(8345) <= (inputs(90)) and not (inputs(67));
    layer0_outputs(8346) <= not((inputs(123)) xor (inputs(130)));
    layer0_outputs(8347) <= not(inputs(141)) or (inputs(162));
    layer0_outputs(8348) <= not(inputs(177));
    layer0_outputs(8349) <= (inputs(73)) and (inputs(240));
    layer0_outputs(8350) <= not((inputs(180)) xor (inputs(192)));
    layer0_outputs(8351) <= (inputs(110)) and not (inputs(251));
    layer0_outputs(8352) <= not((inputs(137)) or (inputs(64)));
    layer0_outputs(8353) <= not(inputs(176));
    layer0_outputs(8354) <= not((inputs(2)) xor (inputs(168)));
    layer0_outputs(8355) <= (inputs(16)) or (inputs(21));
    layer0_outputs(8356) <= not(inputs(25));
    layer0_outputs(8357) <= (inputs(245)) or (inputs(74));
    layer0_outputs(8358) <= '1';
    layer0_outputs(8359) <= not(inputs(101));
    layer0_outputs(8360) <= not(inputs(218));
    layer0_outputs(8361) <= (inputs(119)) or (inputs(173));
    layer0_outputs(8362) <= not((inputs(203)) xor (inputs(162)));
    layer0_outputs(8363) <= inputs(94);
    layer0_outputs(8364) <= not((inputs(173)) or (inputs(234)));
    layer0_outputs(8365) <= not(inputs(19));
    layer0_outputs(8366) <= (inputs(164)) or (inputs(77));
    layer0_outputs(8367) <= inputs(106);
    layer0_outputs(8368) <= (inputs(52)) and (inputs(73));
    layer0_outputs(8369) <= (inputs(167)) or (inputs(11));
    layer0_outputs(8370) <= not((inputs(19)) xor (inputs(70)));
    layer0_outputs(8371) <= inputs(101);
    layer0_outputs(8372) <= not(inputs(216)) or (inputs(243));
    layer0_outputs(8373) <= inputs(218);
    layer0_outputs(8374) <= not(inputs(169)) or (inputs(123));
    layer0_outputs(8375) <= (inputs(18)) xor (inputs(78));
    layer0_outputs(8376) <= (inputs(148)) or (inputs(143));
    layer0_outputs(8377) <= not((inputs(154)) xor (inputs(186)));
    layer0_outputs(8378) <= not(inputs(90));
    layer0_outputs(8379) <= not((inputs(139)) xor (inputs(189)));
    layer0_outputs(8380) <= inputs(81);
    layer0_outputs(8381) <= '0';
    layer0_outputs(8382) <= not((inputs(82)) or (inputs(91)));
    layer0_outputs(8383) <= inputs(12);
    layer0_outputs(8384) <= not(inputs(114));
    layer0_outputs(8385) <= inputs(153);
    layer0_outputs(8386) <= not((inputs(165)) or (inputs(51)));
    layer0_outputs(8387) <= not((inputs(135)) xor (inputs(44)));
    layer0_outputs(8388) <= not(inputs(107)) or (inputs(88));
    layer0_outputs(8389) <= (inputs(249)) and not (inputs(81));
    layer0_outputs(8390) <= (inputs(164)) and not (inputs(46));
    layer0_outputs(8391) <= (inputs(115)) and not (inputs(47));
    layer0_outputs(8392) <= (inputs(128)) xor (inputs(193));
    layer0_outputs(8393) <= inputs(36);
    layer0_outputs(8394) <= (inputs(21)) and (inputs(23));
    layer0_outputs(8395) <= (inputs(213)) and not (inputs(254));
    layer0_outputs(8396) <= not(inputs(213));
    layer0_outputs(8397) <= '1';
    layer0_outputs(8398) <= not(inputs(9));
    layer0_outputs(8399) <= not((inputs(209)) xor (inputs(191)));
    layer0_outputs(8400) <= inputs(88);
    layer0_outputs(8401) <= inputs(151);
    layer0_outputs(8402) <= not((inputs(139)) or (inputs(206)));
    layer0_outputs(8403) <= (inputs(133)) xor (inputs(130));
    layer0_outputs(8404) <= (inputs(132)) and not (inputs(127));
    layer0_outputs(8405) <= not(inputs(21));
    layer0_outputs(8406) <= not((inputs(186)) xor (inputs(249)));
    layer0_outputs(8407) <= not((inputs(244)) or (inputs(58)));
    layer0_outputs(8408) <= (inputs(54)) or (inputs(172));
    layer0_outputs(8409) <= (inputs(22)) and not (inputs(84));
    layer0_outputs(8410) <= not(inputs(94));
    layer0_outputs(8411) <= inputs(44);
    layer0_outputs(8412) <= inputs(92);
    layer0_outputs(8413) <= (inputs(93)) and not (inputs(15));
    layer0_outputs(8414) <= inputs(90);
    layer0_outputs(8415) <= (inputs(59)) and not (inputs(215));
    layer0_outputs(8416) <= not((inputs(61)) xor (inputs(233)));
    layer0_outputs(8417) <= (inputs(114)) or (inputs(239));
    layer0_outputs(8418) <= inputs(36);
    layer0_outputs(8419) <= inputs(158);
    layer0_outputs(8420) <= '1';
    layer0_outputs(8421) <= not((inputs(160)) or (inputs(102)));
    layer0_outputs(8422) <= (inputs(227)) and not (inputs(181));
    layer0_outputs(8423) <= inputs(104);
    layer0_outputs(8424) <= (inputs(203)) or (inputs(16));
    layer0_outputs(8425) <= not(inputs(59));
    layer0_outputs(8426) <= not(inputs(222));
    layer0_outputs(8427) <= (inputs(60)) and (inputs(99));
    layer0_outputs(8428) <= not(inputs(27));
    layer0_outputs(8429) <= (inputs(122)) and not (inputs(18));
    layer0_outputs(8430) <= inputs(82);
    layer0_outputs(8431) <= (inputs(173)) or (inputs(48));
    layer0_outputs(8432) <= (inputs(190)) or (inputs(154));
    layer0_outputs(8433) <= (inputs(0)) xor (inputs(252));
    layer0_outputs(8434) <= not(inputs(36)) or (inputs(246));
    layer0_outputs(8435) <= (inputs(96)) and not (inputs(142));
    layer0_outputs(8436) <= (inputs(246)) and not (inputs(81));
    layer0_outputs(8437) <= (inputs(66)) or (inputs(100));
    layer0_outputs(8438) <= not(inputs(113)) or (inputs(240));
    layer0_outputs(8439) <= inputs(112);
    layer0_outputs(8440) <= inputs(54);
    layer0_outputs(8441) <= not(inputs(25));
    layer0_outputs(8442) <= not(inputs(154)) or (inputs(122));
    layer0_outputs(8443) <= not(inputs(180));
    layer0_outputs(8444) <= not((inputs(129)) xor (inputs(44)));
    layer0_outputs(8445) <= (inputs(186)) xor (inputs(201));
    layer0_outputs(8446) <= (inputs(54)) and not (inputs(139));
    layer0_outputs(8447) <= not((inputs(11)) xor (inputs(139)));
    layer0_outputs(8448) <= not(inputs(30)) or (inputs(245));
    layer0_outputs(8449) <= (inputs(205)) and (inputs(105));
    layer0_outputs(8450) <= inputs(212);
    layer0_outputs(8451) <= inputs(41);
    layer0_outputs(8452) <= inputs(118);
    layer0_outputs(8453) <= not((inputs(161)) or (inputs(47)));
    layer0_outputs(8454) <= not(inputs(117));
    layer0_outputs(8455) <= inputs(246);
    layer0_outputs(8456) <= not(inputs(249)) or (inputs(63));
    layer0_outputs(8457) <= not((inputs(86)) or (inputs(46)));
    layer0_outputs(8458) <= (inputs(82)) and (inputs(56));
    layer0_outputs(8459) <= (inputs(186)) and not (inputs(143));
    layer0_outputs(8460) <= not(inputs(126));
    layer0_outputs(8461) <= not(inputs(211)) or (inputs(112));
    layer0_outputs(8462) <= (inputs(90)) and not (inputs(101));
    layer0_outputs(8463) <= not(inputs(56));
    layer0_outputs(8464) <= not((inputs(17)) xor (inputs(144)));
    layer0_outputs(8465) <= (inputs(106)) and not (inputs(176));
    layer0_outputs(8466) <= not(inputs(76));
    layer0_outputs(8467) <= inputs(168);
    layer0_outputs(8468) <= (inputs(97)) and not (inputs(242));
    layer0_outputs(8469) <= not(inputs(43));
    layer0_outputs(8470) <= not((inputs(147)) or (inputs(126)));
    layer0_outputs(8471) <= (inputs(193)) or (inputs(202));
    layer0_outputs(8472) <= not((inputs(10)) xor (inputs(17)));
    layer0_outputs(8473) <= not(inputs(163));
    layer0_outputs(8474) <= not((inputs(125)) xor (inputs(3)));
    layer0_outputs(8475) <= not(inputs(98));
    layer0_outputs(8476) <= not(inputs(26)) or (inputs(231));
    layer0_outputs(8477) <= not((inputs(109)) xor (inputs(119)));
    layer0_outputs(8478) <= not(inputs(133)) or (inputs(193));
    layer0_outputs(8479) <= (inputs(184)) or (inputs(165));
    layer0_outputs(8480) <= inputs(39);
    layer0_outputs(8481) <= not(inputs(44));
    layer0_outputs(8482) <= (inputs(153)) and not (inputs(72));
    layer0_outputs(8483) <= (inputs(25)) and not (inputs(207));
    layer0_outputs(8484) <= not(inputs(166));
    layer0_outputs(8485) <= not(inputs(202));
    layer0_outputs(8486) <= not(inputs(210)) or (inputs(48));
    layer0_outputs(8487) <= not(inputs(148)) or (inputs(49));
    layer0_outputs(8488) <= not((inputs(94)) or (inputs(18)));
    layer0_outputs(8489) <= not(inputs(230));
    layer0_outputs(8490) <= (inputs(120)) and not (inputs(194));
    layer0_outputs(8491) <= inputs(104);
    layer0_outputs(8492) <= (inputs(209)) xor (inputs(164));
    layer0_outputs(8493) <= inputs(83);
    layer0_outputs(8494) <= (inputs(186)) and not (inputs(98));
    layer0_outputs(8495) <= not((inputs(218)) xor (inputs(64)));
    layer0_outputs(8496) <= (inputs(238)) or (inputs(142));
    layer0_outputs(8497) <= not(inputs(194));
    layer0_outputs(8498) <= inputs(145);
    layer0_outputs(8499) <= (inputs(174)) xor (inputs(90));
    layer0_outputs(8500) <= not(inputs(245));
    layer0_outputs(8501) <= not(inputs(85)) or (inputs(111));
    layer0_outputs(8502) <= (inputs(169)) or (inputs(126));
    layer0_outputs(8503) <= inputs(129);
    layer0_outputs(8504) <= not((inputs(153)) or (inputs(142)));
    layer0_outputs(8505) <= not(inputs(137)) or (inputs(192));
    layer0_outputs(8506) <= inputs(130);
    layer0_outputs(8507) <= inputs(121);
    layer0_outputs(8508) <= '1';
    layer0_outputs(8509) <= (inputs(175)) xor (inputs(21));
    layer0_outputs(8510) <= inputs(176);
    layer0_outputs(8511) <= (inputs(220)) or (inputs(75));
    layer0_outputs(8512) <= inputs(92);
    layer0_outputs(8513) <= not(inputs(43)) or (inputs(245));
    layer0_outputs(8514) <= not(inputs(91)) or (inputs(179));
    layer0_outputs(8515) <= (inputs(211)) and not (inputs(234));
    layer0_outputs(8516) <= not((inputs(19)) or (inputs(11)));
    layer0_outputs(8517) <= not((inputs(88)) xor (inputs(20)));
    layer0_outputs(8518) <= not(inputs(159)) or (inputs(239));
    layer0_outputs(8519) <= inputs(142);
    layer0_outputs(8520) <= (inputs(157)) or (inputs(145));
    layer0_outputs(8521) <= inputs(119);
    layer0_outputs(8522) <= (inputs(156)) or (inputs(155));
    layer0_outputs(8523) <= (inputs(109)) xor (inputs(33));
    layer0_outputs(8524) <= not(inputs(247)) or (inputs(1));
    layer0_outputs(8525) <= (inputs(105)) xor (inputs(158));
    layer0_outputs(8526) <= (inputs(251)) xor (inputs(151));
    layer0_outputs(8527) <= (inputs(116)) or (inputs(13));
    layer0_outputs(8528) <= not(inputs(30));
    layer0_outputs(8529) <= not((inputs(154)) xor (inputs(118)));
    layer0_outputs(8530) <= '1';
    layer0_outputs(8531) <= not(inputs(89)) or (inputs(163));
    layer0_outputs(8532) <= (inputs(107)) xor (inputs(136));
    layer0_outputs(8533) <= (inputs(17)) or (inputs(113));
    layer0_outputs(8534) <= (inputs(252)) xor (inputs(85));
    layer0_outputs(8535) <= not(inputs(9)) or (inputs(226));
    layer0_outputs(8536) <= (inputs(253)) or (inputs(184));
    layer0_outputs(8537) <= not(inputs(242)) or (inputs(155));
    layer0_outputs(8538) <= (inputs(108)) and not (inputs(59));
    layer0_outputs(8539) <= not((inputs(60)) or (inputs(78)));
    layer0_outputs(8540) <= (inputs(85)) and not (inputs(158));
    layer0_outputs(8541) <= not((inputs(32)) or (inputs(213)));
    layer0_outputs(8542) <= not(inputs(74)) or (inputs(3));
    layer0_outputs(8543) <= not((inputs(223)) xor (inputs(194)));
    layer0_outputs(8544) <= (inputs(84)) xor (inputs(7));
    layer0_outputs(8545) <= not(inputs(40));
    layer0_outputs(8546) <= not(inputs(86));
    layer0_outputs(8547) <= inputs(62);
    layer0_outputs(8548) <= not((inputs(216)) xor (inputs(119)));
    layer0_outputs(8549) <= (inputs(74)) or (inputs(211));
    layer0_outputs(8550) <= not((inputs(177)) or (inputs(162)));
    layer0_outputs(8551) <= (inputs(61)) and not (inputs(126));
    layer0_outputs(8552) <= not((inputs(24)) or (inputs(223)));
    layer0_outputs(8553) <= not(inputs(233));
    layer0_outputs(8554) <= not((inputs(99)) xor (inputs(186)));
    layer0_outputs(8555) <= inputs(236);
    layer0_outputs(8556) <= (inputs(205)) or (inputs(70));
    layer0_outputs(8557) <= (inputs(112)) xor (inputs(147));
    layer0_outputs(8558) <= inputs(69);
    layer0_outputs(8559) <= not((inputs(244)) xor (inputs(213)));
    layer0_outputs(8560) <= not(inputs(79)) or (inputs(254));
    layer0_outputs(8561) <= not((inputs(83)) or (inputs(243)));
    layer0_outputs(8562) <= (inputs(134)) and not (inputs(40));
    layer0_outputs(8563) <= (inputs(100)) and (inputs(117));
    layer0_outputs(8564) <= not((inputs(207)) or (inputs(193)));
    layer0_outputs(8565) <= not((inputs(180)) xor (inputs(73)));
    layer0_outputs(8566) <= not((inputs(212)) and (inputs(230)));
    layer0_outputs(8567) <= not((inputs(253)) or (inputs(70)));
    layer0_outputs(8568) <= not((inputs(163)) or (inputs(160)));
    layer0_outputs(8569) <= not(inputs(118));
    layer0_outputs(8570) <= (inputs(144)) and not (inputs(64));
    layer0_outputs(8571) <= inputs(78);
    layer0_outputs(8572) <= not(inputs(237)) or (inputs(254));
    layer0_outputs(8573) <= (inputs(181)) and not (inputs(114));
    layer0_outputs(8574) <= not((inputs(106)) xor (inputs(126)));
    layer0_outputs(8575) <= not((inputs(232)) or (inputs(28)));
    layer0_outputs(8576) <= inputs(74);
    layer0_outputs(8577) <= not(inputs(69));
    layer0_outputs(8578) <= inputs(221);
    layer0_outputs(8579) <= inputs(217);
    layer0_outputs(8580) <= inputs(85);
    layer0_outputs(8581) <= not(inputs(201)) or (inputs(45));
    layer0_outputs(8582) <= (inputs(32)) or (inputs(211));
    layer0_outputs(8583) <= not(inputs(4)) or (inputs(38));
    layer0_outputs(8584) <= (inputs(196)) xor (inputs(160));
    layer0_outputs(8585) <= inputs(144);
    layer0_outputs(8586) <= not((inputs(67)) or (inputs(160)));
    layer0_outputs(8587) <= inputs(48);
    layer0_outputs(8588) <= not((inputs(174)) xor (inputs(102)));
    layer0_outputs(8589) <= not(inputs(103));
    layer0_outputs(8590) <= (inputs(78)) or (inputs(86));
    layer0_outputs(8591) <= not(inputs(96));
    layer0_outputs(8592) <= not((inputs(52)) xor (inputs(164)));
    layer0_outputs(8593) <= not(inputs(27));
    layer0_outputs(8594) <= not((inputs(206)) or (inputs(15)));
    layer0_outputs(8595) <= not(inputs(138));
    layer0_outputs(8596) <= not(inputs(246)) or (inputs(47));
    layer0_outputs(8597) <= (inputs(110)) or (inputs(143));
    layer0_outputs(8598) <= (inputs(168)) and not (inputs(81));
    layer0_outputs(8599) <= (inputs(192)) and not (inputs(109));
    layer0_outputs(8600) <= inputs(27);
    layer0_outputs(8601) <= (inputs(76)) or (inputs(88));
    layer0_outputs(8602) <= inputs(109);
    layer0_outputs(8603) <= not((inputs(17)) xor (inputs(48)));
    layer0_outputs(8604) <= not(inputs(143)) or (inputs(18));
    layer0_outputs(8605) <= not(inputs(120)) or (inputs(158));
    layer0_outputs(8606) <= (inputs(89)) and not (inputs(11));
    layer0_outputs(8607) <= not((inputs(174)) xor (inputs(214)));
    layer0_outputs(8608) <= inputs(82);
    layer0_outputs(8609) <= not(inputs(118)) or (inputs(239));
    layer0_outputs(8610) <= (inputs(186)) xor (inputs(219));
    layer0_outputs(8611) <= (inputs(144)) xor (inputs(5));
    layer0_outputs(8612) <= not(inputs(153));
    layer0_outputs(8613) <= inputs(210);
    layer0_outputs(8614) <= not(inputs(91));
    layer0_outputs(8615) <= inputs(52);
    layer0_outputs(8616) <= inputs(167);
    layer0_outputs(8617) <= not((inputs(44)) or (inputs(176)));
    layer0_outputs(8618) <= not(inputs(125));
    layer0_outputs(8619) <= (inputs(0)) or (inputs(197));
    layer0_outputs(8620) <= (inputs(162)) xor (inputs(69));
    layer0_outputs(8621) <= (inputs(204)) xor (inputs(174));
    layer0_outputs(8622) <= not((inputs(51)) xor (inputs(103)));
    layer0_outputs(8623) <= (inputs(204)) and not (inputs(36));
    layer0_outputs(8624) <= not((inputs(93)) xor (inputs(105)));
    layer0_outputs(8625) <= inputs(119);
    layer0_outputs(8626) <= (inputs(159)) or (inputs(46));
    layer0_outputs(8627) <= not(inputs(167)) or (inputs(58));
    layer0_outputs(8628) <= inputs(251);
    layer0_outputs(8629) <= inputs(182);
    layer0_outputs(8630) <= not((inputs(158)) xor (inputs(106)));
    layer0_outputs(8631) <= not(inputs(246)) or (inputs(11));
    layer0_outputs(8632) <= (inputs(61)) or (inputs(175));
    layer0_outputs(8633) <= not(inputs(76));
    layer0_outputs(8634) <= (inputs(223)) or (inputs(69));
    layer0_outputs(8635) <= not((inputs(91)) or (inputs(78)));
    layer0_outputs(8636) <= inputs(182);
    layer0_outputs(8637) <= inputs(196);
    layer0_outputs(8638) <= (inputs(127)) and not (inputs(238));
    layer0_outputs(8639) <= inputs(146);
    layer0_outputs(8640) <= not(inputs(95));
    layer0_outputs(8641) <= (inputs(128)) xor (inputs(187));
    layer0_outputs(8642) <= (inputs(158)) and not (inputs(80));
    layer0_outputs(8643) <= inputs(114);
    layer0_outputs(8644) <= '1';
    layer0_outputs(8645) <= '1';
    layer0_outputs(8646) <= inputs(45);
    layer0_outputs(8647) <= (inputs(89)) and not (inputs(230));
    layer0_outputs(8648) <= not(inputs(3));
    layer0_outputs(8649) <= inputs(61);
    layer0_outputs(8650) <= not((inputs(96)) or (inputs(30)));
    layer0_outputs(8651) <= inputs(234);
    layer0_outputs(8652) <= not((inputs(66)) or (inputs(45)));
    layer0_outputs(8653) <= (inputs(227)) and not (inputs(86));
    layer0_outputs(8654) <= not(inputs(179));
    layer0_outputs(8655) <= (inputs(62)) xor (inputs(1));
    layer0_outputs(8656) <= not(inputs(232));
    layer0_outputs(8657) <= not(inputs(85));
    layer0_outputs(8658) <= inputs(0);
    layer0_outputs(8659) <= (inputs(23)) and not (inputs(181));
    layer0_outputs(8660) <= not((inputs(143)) or (inputs(40)));
    layer0_outputs(8661) <= not(inputs(181));
    layer0_outputs(8662) <= not((inputs(68)) and (inputs(90)));
    layer0_outputs(8663) <= inputs(182);
    layer0_outputs(8664) <= not(inputs(28)) or (inputs(193));
    layer0_outputs(8665) <= not(inputs(62));
    layer0_outputs(8666) <= (inputs(198)) and not (inputs(172));
    layer0_outputs(8667) <= (inputs(123)) and (inputs(124));
    layer0_outputs(8668) <= not((inputs(195)) or (inputs(65)));
    layer0_outputs(8669) <= (inputs(116)) or (inputs(140));
    layer0_outputs(8670) <= (inputs(71)) xor (inputs(22));
    layer0_outputs(8671) <= inputs(182);
    layer0_outputs(8672) <= not(inputs(7));
    layer0_outputs(8673) <= (inputs(226)) or (inputs(19));
    layer0_outputs(8674) <= not(inputs(83));
    layer0_outputs(8675) <= not(inputs(103));
    layer0_outputs(8676) <= (inputs(21)) or (inputs(143));
    layer0_outputs(8677) <= (inputs(141)) or (inputs(221));
    layer0_outputs(8678) <= inputs(220);
    layer0_outputs(8679) <= (inputs(134)) and (inputs(237));
    layer0_outputs(8680) <= (inputs(214)) xor (inputs(216));
    layer0_outputs(8681) <= not(inputs(108)) or (inputs(81));
    layer0_outputs(8682) <= not(inputs(44));
    layer0_outputs(8683) <= inputs(39);
    layer0_outputs(8684) <= (inputs(158)) xor (inputs(88));
    layer0_outputs(8685) <= (inputs(3)) xor (inputs(181));
    layer0_outputs(8686) <= (inputs(170)) or (inputs(159));
    layer0_outputs(8687) <= (inputs(231)) and not (inputs(64));
    layer0_outputs(8688) <= inputs(106);
    layer0_outputs(8689) <= (inputs(192)) or (inputs(116));
    layer0_outputs(8690) <= (inputs(178)) or (inputs(255));
    layer0_outputs(8691) <= (inputs(81)) or (inputs(136));
    layer0_outputs(8692) <= not(inputs(78)) or (inputs(255));
    layer0_outputs(8693) <= '1';
    layer0_outputs(8694) <= inputs(184);
    layer0_outputs(8695) <= not((inputs(132)) or (inputs(145)));
    layer0_outputs(8696) <= inputs(121);
    layer0_outputs(8697) <= not(inputs(23)) or (inputs(224));
    layer0_outputs(8698) <= inputs(127);
    layer0_outputs(8699) <= (inputs(68)) and not (inputs(49));
    layer0_outputs(8700) <= not(inputs(29)) or (inputs(115));
    layer0_outputs(8701) <= (inputs(190)) and not (inputs(12));
    layer0_outputs(8702) <= not((inputs(238)) xor (inputs(19)));
    layer0_outputs(8703) <= not((inputs(55)) xor (inputs(17)));
    layer0_outputs(8704) <= (inputs(68)) xor (inputs(133));
    layer0_outputs(8705) <= not((inputs(66)) or (inputs(63)));
    layer0_outputs(8706) <= not(inputs(69)) or (inputs(206));
    layer0_outputs(8707) <= not(inputs(198)) or (inputs(122));
    layer0_outputs(8708) <= (inputs(223)) xor (inputs(190));
    layer0_outputs(8709) <= (inputs(66)) xor (inputs(6));
    layer0_outputs(8710) <= (inputs(21)) xor (inputs(69));
    layer0_outputs(8711) <= inputs(102);
    layer0_outputs(8712) <= not((inputs(50)) or (inputs(167)));
    layer0_outputs(8713) <= not(inputs(172)) or (inputs(142));
    layer0_outputs(8714) <= not(inputs(99)) or (inputs(175));
    layer0_outputs(8715) <= inputs(182);
    layer0_outputs(8716) <= (inputs(55)) and not (inputs(255));
    layer0_outputs(8717) <= not((inputs(114)) or (inputs(171)));
    layer0_outputs(8718) <= inputs(150);
    layer0_outputs(8719) <= inputs(221);
    layer0_outputs(8720) <= (inputs(2)) or (inputs(10));
    layer0_outputs(8721) <= not(inputs(62));
    layer0_outputs(8722) <= inputs(78);
    layer0_outputs(8723) <= inputs(39);
    layer0_outputs(8724) <= (inputs(228)) and not (inputs(138));
    layer0_outputs(8725) <= (inputs(205)) or (inputs(144));
    layer0_outputs(8726) <= inputs(129);
    layer0_outputs(8727) <= not((inputs(38)) xor (inputs(109)));
    layer0_outputs(8728) <= not(inputs(130)) or (inputs(208));
    layer0_outputs(8729) <= not((inputs(32)) or (inputs(184)));
    layer0_outputs(8730) <= (inputs(228)) or (inputs(254));
    layer0_outputs(8731) <= not((inputs(192)) or (inputs(215)));
    layer0_outputs(8732) <= (inputs(195)) and not (inputs(153));
    layer0_outputs(8733) <= inputs(152);
    layer0_outputs(8734) <= inputs(182);
    layer0_outputs(8735) <= not(inputs(31));
    layer0_outputs(8736) <= not(inputs(61));
    layer0_outputs(8737) <= inputs(63);
    layer0_outputs(8738) <= not(inputs(40));
    layer0_outputs(8739) <= (inputs(186)) and not (inputs(59));
    layer0_outputs(8740) <= (inputs(229)) xor (inputs(198));
    layer0_outputs(8741) <= (inputs(12)) xor (inputs(71));
    layer0_outputs(8742) <= not((inputs(173)) or (inputs(149)));
    layer0_outputs(8743) <= inputs(229);
    layer0_outputs(8744) <= (inputs(61)) or (inputs(10));
    layer0_outputs(8745) <= (inputs(225)) or (inputs(15));
    layer0_outputs(8746) <= not(inputs(115));
    layer0_outputs(8747) <= not(inputs(182)) or (inputs(171));
    layer0_outputs(8748) <= not(inputs(228));
    layer0_outputs(8749) <= not(inputs(109));
    layer0_outputs(8750) <= not((inputs(3)) or (inputs(220)));
    layer0_outputs(8751) <= not((inputs(176)) or (inputs(67)));
    layer0_outputs(8752) <= not(inputs(105));
    layer0_outputs(8753) <= not((inputs(129)) xor (inputs(182)));
    layer0_outputs(8754) <= inputs(63);
    layer0_outputs(8755) <= (inputs(128)) or (inputs(30));
    layer0_outputs(8756) <= not((inputs(32)) or (inputs(48)));
    layer0_outputs(8757) <= inputs(140);
    layer0_outputs(8758) <= (inputs(101)) or (inputs(97));
    layer0_outputs(8759) <= not((inputs(38)) or (inputs(30)));
    layer0_outputs(8760) <= not((inputs(230)) or (inputs(225)));
    layer0_outputs(8761) <= not((inputs(87)) and (inputs(110)));
    layer0_outputs(8762) <= not((inputs(191)) xor (inputs(5)));
    layer0_outputs(8763) <= not(inputs(199));
    layer0_outputs(8764) <= inputs(104);
    layer0_outputs(8765) <= (inputs(190)) xor (inputs(223));
    layer0_outputs(8766) <= inputs(136);
    layer0_outputs(8767) <= (inputs(77)) and not (inputs(3));
    layer0_outputs(8768) <= not(inputs(212));
    layer0_outputs(8769) <= not((inputs(97)) or (inputs(255)));
    layer0_outputs(8770) <= inputs(228);
    layer0_outputs(8771) <= not((inputs(195)) or (inputs(248)));
    layer0_outputs(8772) <= inputs(3);
    layer0_outputs(8773) <= inputs(150);
    layer0_outputs(8774) <= not(inputs(164)) or (inputs(79));
    layer0_outputs(8775) <= not((inputs(112)) xor (inputs(133)));
    layer0_outputs(8776) <= not((inputs(123)) and (inputs(167)));
    layer0_outputs(8777) <= (inputs(113)) and (inputs(248));
    layer0_outputs(8778) <= not((inputs(168)) xor (inputs(196)));
    layer0_outputs(8779) <= inputs(18);
    layer0_outputs(8780) <= not((inputs(166)) xor (inputs(153)));
    layer0_outputs(8781) <= (inputs(143)) or (inputs(40));
    layer0_outputs(8782) <= not((inputs(130)) or (inputs(174)));
    layer0_outputs(8783) <= (inputs(196)) and not (inputs(78));
    layer0_outputs(8784) <= not((inputs(174)) or (inputs(163)));
    layer0_outputs(8785) <= not((inputs(145)) xor (inputs(115)));
    layer0_outputs(8786) <= (inputs(151)) and not (inputs(1));
    layer0_outputs(8787) <= inputs(43);
    layer0_outputs(8788) <= (inputs(10)) and not (inputs(207));
    layer0_outputs(8789) <= not((inputs(38)) xor (inputs(149)));
    layer0_outputs(8790) <= not((inputs(86)) or (inputs(134)));
    layer0_outputs(8791) <= inputs(230);
    layer0_outputs(8792) <= not((inputs(226)) and (inputs(72)));
    layer0_outputs(8793) <= inputs(101);
    layer0_outputs(8794) <= not((inputs(40)) or (inputs(243)));
    layer0_outputs(8795) <= not(inputs(103));
    layer0_outputs(8796) <= inputs(201);
    layer0_outputs(8797) <= not(inputs(216)) or (inputs(190));
    layer0_outputs(8798) <= (inputs(188)) or (inputs(2));
    layer0_outputs(8799) <= (inputs(35)) or (inputs(135));
    layer0_outputs(8800) <= (inputs(189)) and not (inputs(13));
    layer0_outputs(8801) <= not((inputs(15)) or (inputs(101)));
    layer0_outputs(8802) <= (inputs(242)) or (inputs(24));
    layer0_outputs(8803) <= not(inputs(119)) or (inputs(4));
    layer0_outputs(8804) <= (inputs(186)) or (inputs(224));
    layer0_outputs(8805) <= not(inputs(231));
    layer0_outputs(8806) <= (inputs(27)) or (inputs(111));
    layer0_outputs(8807) <= (inputs(67)) and not (inputs(178));
    layer0_outputs(8808) <= not((inputs(254)) xor (inputs(28)));
    layer0_outputs(8809) <= not((inputs(134)) xor (inputs(87)));
    layer0_outputs(8810) <= inputs(149);
    layer0_outputs(8811) <= (inputs(11)) xor (inputs(74));
    layer0_outputs(8812) <= not(inputs(87)) or (inputs(30));
    layer0_outputs(8813) <= not((inputs(36)) or (inputs(190)));
    layer0_outputs(8814) <= not((inputs(155)) or (inputs(95)));
    layer0_outputs(8815) <= inputs(87);
    layer0_outputs(8816) <= not((inputs(234)) or (inputs(217)));
    layer0_outputs(8817) <= not(inputs(62));
    layer0_outputs(8818) <= not((inputs(171)) xor (inputs(58)));
    layer0_outputs(8819) <= inputs(121);
    layer0_outputs(8820) <= not((inputs(151)) or (inputs(216)));
    layer0_outputs(8821) <= inputs(99);
    layer0_outputs(8822) <= not((inputs(26)) xor (inputs(28)));
    layer0_outputs(8823) <= not(inputs(89)) or (inputs(206));
    layer0_outputs(8824) <= not(inputs(243)) or (inputs(99));
    layer0_outputs(8825) <= not((inputs(146)) or (inputs(69)));
    layer0_outputs(8826) <= (inputs(122)) xor (inputs(14));
    layer0_outputs(8827) <= inputs(131);
    layer0_outputs(8828) <= '0';
    layer0_outputs(8829) <= not(inputs(27));
    layer0_outputs(8830) <= not((inputs(84)) xor (inputs(133)));
    layer0_outputs(8831) <= not(inputs(236));
    layer0_outputs(8832) <= not((inputs(122)) or (inputs(215)));
    layer0_outputs(8833) <= not(inputs(94)) or (inputs(12));
    layer0_outputs(8834) <= (inputs(68)) xor (inputs(20));
    layer0_outputs(8835) <= not(inputs(76));
    layer0_outputs(8836) <= (inputs(224)) or (inputs(117));
    layer0_outputs(8837) <= not(inputs(23));
    layer0_outputs(8838) <= (inputs(48)) or (inputs(79));
    layer0_outputs(8839) <= not((inputs(49)) xor (inputs(24)));
    layer0_outputs(8840) <= not((inputs(119)) or (inputs(62)));
    layer0_outputs(8841) <= (inputs(201)) and not (inputs(247));
    layer0_outputs(8842) <= not((inputs(134)) xor (inputs(183)));
    layer0_outputs(8843) <= inputs(227);
    layer0_outputs(8844) <= not((inputs(163)) or (inputs(17)));
    layer0_outputs(8845) <= inputs(154);
    layer0_outputs(8846) <= not((inputs(77)) xor (inputs(237)));
    layer0_outputs(8847) <= not((inputs(193)) or (inputs(226)));
    layer0_outputs(8848) <= (inputs(216)) and not (inputs(238));
    layer0_outputs(8849) <= (inputs(82)) or (inputs(98));
    layer0_outputs(8850) <= (inputs(94)) or (inputs(61));
    layer0_outputs(8851) <= not((inputs(246)) xor (inputs(74)));
    layer0_outputs(8852) <= not(inputs(24));
    layer0_outputs(8853) <= (inputs(219)) or (inputs(175));
    layer0_outputs(8854) <= inputs(33);
    layer0_outputs(8855) <= inputs(182);
    layer0_outputs(8856) <= not((inputs(36)) or (inputs(190)));
    layer0_outputs(8857) <= inputs(89);
    layer0_outputs(8858) <= not(inputs(230));
    layer0_outputs(8859) <= not((inputs(255)) or (inputs(182)));
    layer0_outputs(8860) <= not((inputs(43)) or (inputs(170)));
    layer0_outputs(8861) <= (inputs(125)) and not (inputs(16));
    layer0_outputs(8862) <= not(inputs(122)) or (inputs(76));
    layer0_outputs(8863) <= not(inputs(70));
    layer0_outputs(8864) <= not(inputs(60)) or (inputs(0));
    layer0_outputs(8865) <= inputs(34);
    layer0_outputs(8866) <= not((inputs(73)) xor (inputs(38)));
    layer0_outputs(8867) <= (inputs(26)) or (inputs(171));
    layer0_outputs(8868) <= inputs(121);
    layer0_outputs(8869) <= (inputs(224)) or (inputs(219));
    layer0_outputs(8870) <= inputs(148);
    layer0_outputs(8871) <= not(inputs(34)) or (inputs(185));
    layer0_outputs(8872) <= not((inputs(213)) or (inputs(174)));
    layer0_outputs(8873) <= not((inputs(186)) xor (inputs(7)));
    layer0_outputs(8874) <= not((inputs(42)) or (inputs(1)));
    layer0_outputs(8875) <= not((inputs(49)) and (inputs(240)));
    layer0_outputs(8876) <= inputs(55);
    layer0_outputs(8877) <= not(inputs(181));
    layer0_outputs(8878) <= (inputs(13)) and not (inputs(76));
    layer0_outputs(8879) <= not(inputs(185));
    layer0_outputs(8880) <= (inputs(239)) xor (inputs(41));
    layer0_outputs(8881) <= (inputs(230)) and not (inputs(243));
    layer0_outputs(8882) <= inputs(22);
    layer0_outputs(8883) <= (inputs(166)) or (inputs(2));
    layer0_outputs(8884) <= not(inputs(163));
    layer0_outputs(8885) <= (inputs(139)) and not (inputs(241));
    layer0_outputs(8886) <= not(inputs(104)) or (inputs(216));
    layer0_outputs(8887) <= inputs(25);
    layer0_outputs(8888) <= not(inputs(123)) or (inputs(98));
    layer0_outputs(8889) <= not(inputs(40)) or (inputs(236));
    layer0_outputs(8890) <= inputs(46);
    layer0_outputs(8891) <= not((inputs(53)) or (inputs(62)));
    layer0_outputs(8892) <= not((inputs(115)) xor (inputs(76)));
    layer0_outputs(8893) <= (inputs(54)) or (inputs(103));
    layer0_outputs(8894) <= not((inputs(74)) xor (inputs(23)));
    layer0_outputs(8895) <= not((inputs(97)) xor (inputs(170)));
    layer0_outputs(8896) <= (inputs(189)) and not (inputs(17));
    layer0_outputs(8897) <= not((inputs(59)) xor (inputs(3)));
    layer0_outputs(8898) <= inputs(146);
    layer0_outputs(8899) <= (inputs(214)) or (inputs(190));
    layer0_outputs(8900) <= not(inputs(94)) or (inputs(221));
    layer0_outputs(8901) <= (inputs(51)) and not (inputs(126));
    layer0_outputs(8902) <= (inputs(183)) and not (inputs(12));
    layer0_outputs(8903) <= not(inputs(70)) or (inputs(159));
    layer0_outputs(8904) <= (inputs(54)) or (inputs(78));
    layer0_outputs(8905) <= (inputs(107)) and not (inputs(143));
    layer0_outputs(8906) <= not(inputs(179)) or (inputs(125));
    layer0_outputs(8907) <= not(inputs(61));
    layer0_outputs(8908) <= (inputs(108)) and not (inputs(203));
    layer0_outputs(8909) <= (inputs(91)) and not (inputs(13));
    layer0_outputs(8910) <= not((inputs(17)) or (inputs(234)));
    layer0_outputs(8911) <= '0';
    layer0_outputs(8912) <= not((inputs(144)) xor (inputs(99)));
    layer0_outputs(8913) <= (inputs(233)) and not (inputs(85));
    layer0_outputs(8914) <= (inputs(15)) and not (inputs(214));
    layer0_outputs(8915) <= not(inputs(98));
    layer0_outputs(8916) <= inputs(47);
    layer0_outputs(8917) <= not((inputs(253)) or (inputs(30)));
    layer0_outputs(8918) <= (inputs(64)) or (inputs(77));
    layer0_outputs(8919) <= '0';
    layer0_outputs(8920) <= (inputs(237)) xor (inputs(4));
    layer0_outputs(8921) <= not(inputs(13));
    layer0_outputs(8922) <= (inputs(120)) xor (inputs(195));
    layer0_outputs(8923) <= not((inputs(72)) or (inputs(130)));
    layer0_outputs(8924) <= (inputs(140)) or (inputs(110));
    layer0_outputs(8925) <= not((inputs(182)) or (inputs(146)));
    layer0_outputs(8926) <= (inputs(52)) or (inputs(70));
    layer0_outputs(8927) <= '0';
    layer0_outputs(8928) <= (inputs(31)) and not (inputs(51));
    layer0_outputs(8929) <= inputs(9);
    layer0_outputs(8930) <= not((inputs(136)) or (inputs(104)));
    layer0_outputs(8931) <= not(inputs(120));
    layer0_outputs(8932) <= not(inputs(59)) or (inputs(206));
    layer0_outputs(8933) <= (inputs(137)) and not (inputs(36));
    layer0_outputs(8934) <= (inputs(42)) or (inputs(126));
    layer0_outputs(8935) <= not((inputs(126)) xor (inputs(108)));
    layer0_outputs(8936) <= not(inputs(161));
    layer0_outputs(8937) <= not(inputs(3));
    layer0_outputs(8938) <= not(inputs(166));
    layer0_outputs(8939) <= (inputs(160)) xor (inputs(129));
    layer0_outputs(8940) <= (inputs(169)) and not (inputs(97));
    layer0_outputs(8941) <= not((inputs(213)) or (inputs(88)));
    layer0_outputs(8942) <= (inputs(222)) xor (inputs(206));
    layer0_outputs(8943) <= not(inputs(36));
    layer0_outputs(8944) <= inputs(175);
    layer0_outputs(8945) <= not(inputs(211)) or (inputs(120));
    layer0_outputs(8946) <= not((inputs(95)) xor (inputs(192)));
    layer0_outputs(8947) <= not(inputs(197)) or (inputs(125));
    layer0_outputs(8948) <= not(inputs(230));
    layer0_outputs(8949) <= not((inputs(252)) or (inputs(115)));
    layer0_outputs(8950) <= not(inputs(178));
    layer0_outputs(8951) <= not(inputs(91)) or (inputs(178));
    layer0_outputs(8952) <= inputs(133);
    layer0_outputs(8953) <= not(inputs(54));
    layer0_outputs(8954) <= (inputs(49)) xor (inputs(247));
    layer0_outputs(8955) <= not(inputs(113));
    layer0_outputs(8956) <= not((inputs(115)) or (inputs(26)));
    layer0_outputs(8957) <= not(inputs(153)) or (inputs(3));
    layer0_outputs(8958) <= (inputs(51)) xor (inputs(73));
    layer0_outputs(8959) <= inputs(1);
    layer0_outputs(8960) <= inputs(147);
    layer0_outputs(8961) <= (inputs(59)) and not (inputs(236));
    layer0_outputs(8962) <= (inputs(74)) xor (inputs(43));
    layer0_outputs(8963) <= (inputs(220)) or (inputs(236));
    layer0_outputs(8964) <= (inputs(116)) and not (inputs(17));
    layer0_outputs(8965) <= not(inputs(54)) or (inputs(94));
    layer0_outputs(8966) <= not(inputs(116));
    layer0_outputs(8967) <= inputs(72);
    layer0_outputs(8968) <= (inputs(227)) and not (inputs(25));
    layer0_outputs(8969) <= not(inputs(211));
    layer0_outputs(8970) <= inputs(24);
    layer0_outputs(8971) <= (inputs(164)) xor (inputs(219));
    layer0_outputs(8972) <= (inputs(48)) xor (inputs(44));
    layer0_outputs(8973) <= not((inputs(202)) xor (inputs(145)));
    layer0_outputs(8974) <= inputs(230);
    layer0_outputs(8975) <= inputs(26);
    layer0_outputs(8976) <= not(inputs(98)) or (inputs(28));
    layer0_outputs(8977) <= inputs(214);
    layer0_outputs(8978) <= not(inputs(109));
    layer0_outputs(8979) <= not(inputs(15));
    layer0_outputs(8980) <= (inputs(216)) and (inputs(218));
    layer0_outputs(8981) <= not((inputs(8)) or (inputs(125)));
    layer0_outputs(8982) <= not((inputs(2)) or (inputs(12)));
    layer0_outputs(8983) <= (inputs(209)) or (inputs(223));
    layer0_outputs(8984) <= not(inputs(194));
    layer0_outputs(8985) <= not(inputs(145));
    layer0_outputs(8986) <= inputs(28);
    layer0_outputs(8987) <= not(inputs(255));
    layer0_outputs(8988) <= (inputs(86)) xor (inputs(35));
    layer0_outputs(8989) <= (inputs(243)) or (inputs(245));
    layer0_outputs(8990) <= not(inputs(80));
    layer0_outputs(8991) <= (inputs(202)) and (inputs(76));
    layer0_outputs(8992) <= (inputs(84)) and not (inputs(95));
    layer0_outputs(8993) <= (inputs(99)) or (inputs(174));
    layer0_outputs(8994) <= (inputs(91)) or (inputs(154));
    layer0_outputs(8995) <= (inputs(184)) or (inputs(200));
    layer0_outputs(8996) <= inputs(13);
    layer0_outputs(8997) <= not(inputs(71));
    layer0_outputs(8998) <= inputs(100);
    layer0_outputs(8999) <= (inputs(151)) or (inputs(228));
    layer0_outputs(9000) <= inputs(148);
    layer0_outputs(9001) <= inputs(130);
    layer0_outputs(9002) <= not((inputs(88)) and (inputs(87)));
    layer0_outputs(9003) <= (inputs(38)) and not (inputs(56));
    layer0_outputs(9004) <= not(inputs(246));
    layer0_outputs(9005) <= not(inputs(107)) or (inputs(103));
    layer0_outputs(9006) <= inputs(92);
    layer0_outputs(9007) <= not((inputs(188)) or (inputs(79)));
    layer0_outputs(9008) <= not((inputs(149)) xor (inputs(182)));
    layer0_outputs(9009) <= not(inputs(139));
    layer0_outputs(9010) <= not((inputs(154)) xor (inputs(207)));
    layer0_outputs(9011) <= not((inputs(124)) or (inputs(220)));
    layer0_outputs(9012) <= inputs(194);
    layer0_outputs(9013) <= (inputs(220)) and (inputs(219));
    layer0_outputs(9014) <= not((inputs(22)) xor (inputs(113)));
    layer0_outputs(9015) <= not((inputs(124)) xor (inputs(77)));
    layer0_outputs(9016) <= not(inputs(82));
    layer0_outputs(9017) <= not(inputs(14)) or (inputs(225));
    layer0_outputs(9018) <= not((inputs(68)) or (inputs(28)));
    layer0_outputs(9019) <= not((inputs(133)) xor (inputs(220)));
    layer0_outputs(9020) <= not((inputs(105)) xor (inputs(22)));
    layer0_outputs(9021) <= inputs(218);
    layer0_outputs(9022) <= inputs(214);
    layer0_outputs(9023) <= inputs(143);
    layer0_outputs(9024) <= not(inputs(116)) or (inputs(204));
    layer0_outputs(9025) <= not(inputs(107));
    layer0_outputs(9026) <= inputs(149);
    layer0_outputs(9027) <= (inputs(141)) or (inputs(140));
    layer0_outputs(9028) <= (inputs(192)) xor (inputs(215));
    layer0_outputs(9029) <= not((inputs(19)) or (inputs(72)));
    layer0_outputs(9030) <= not((inputs(214)) or (inputs(106)));
    layer0_outputs(9031) <= inputs(23);
    layer0_outputs(9032) <= not(inputs(104));
    layer0_outputs(9033) <= not(inputs(141));
    layer0_outputs(9034) <= inputs(160);
    layer0_outputs(9035) <= (inputs(96)) and (inputs(108));
    layer0_outputs(9036) <= not((inputs(26)) xor (inputs(173)));
    layer0_outputs(9037) <= not(inputs(68));
    layer0_outputs(9038) <= (inputs(61)) or (inputs(216));
    layer0_outputs(9039) <= not((inputs(226)) xor (inputs(118)));
    layer0_outputs(9040) <= (inputs(89)) and not (inputs(36));
    layer0_outputs(9041) <= not(inputs(118));
    layer0_outputs(9042) <= not((inputs(229)) or (inputs(172)));
    layer0_outputs(9043) <= (inputs(37)) xor (inputs(79));
    layer0_outputs(9044) <= not(inputs(108));
    layer0_outputs(9045) <= inputs(215);
    layer0_outputs(9046) <= not(inputs(55));
    layer0_outputs(9047) <= not((inputs(16)) or (inputs(105)));
    layer0_outputs(9048) <= (inputs(138)) and not (inputs(225));
    layer0_outputs(9049) <= inputs(113);
    layer0_outputs(9050) <= inputs(195);
    layer0_outputs(9051) <= not((inputs(189)) or (inputs(81)));
    layer0_outputs(9052) <= not(inputs(99)) or (inputs(127));
    layer0_outputs(9053) <= not(inputs(70));
    layer0_outputs(9054) <= not((inputs(149)) xor (inputs(167)));
    layer0_outputs(9055) <= not(inputs(138));
    layer0_outputs(9056) <= not(inputs(167)) or (inputs(185));
    layer0_outputs(9057) <= (inputs(122)) and not (inputs(209));
    layer0_outputs(9058) <= not(inputs(117)) or (inputs(189));
    layer0_outputs(9059) <= not((inputs(242)) or (inputs(37)));
    layer0_outputs(9060) <= not(inputs(174));
    layer0_outputs(9061) <= (inputs(145)) xor (inputs(190));
    layer0_outputs(9062) <= not((inputs(232)) xor (inputs(245)));
    layer0_outputs(9063) <= (inputs(173)) and not (inputs(32));
    layer0_outputs(9064) <= not((inputs(86)) or (inputs(176)));
    layer0_outputs(9065) <= not((inputs(28)) xor (inputs(61)));
    layer0_outputs(9066) <= not((inputs(199)) xor (inputs(180)));
    layer0_outputs(9067) <= (inputs(230)) and not (inputs(172));
    layer0_outputs(9068) <= not(inputs(228)) or (inputs(135));
    layer0_outputs(9069) <= inputs(175);
    layer0_outputs(9070) <= (inputs(21)) and not (inputs(148));
    layer0_outputs(9071) <= not((inputs(91)) or (inputs(255)));
    layer0_outputs(9072) <= not((inputs(152)) xor (inputs(119)));
    layer0_outputs(9073) <= inputs(213);
    layer0_outputs(9074) <= (inputs(42)) and not (inputs(234));
    layer0_outputs(9075) <= not((inputs(187)) xor (inputs(159)));
    layer0_outputs(9076) <= (inputs(84)) or (inputs(62));
    layer0_outputs(9077) <= (inputs(161)) or (inputs(202));
    layer0_outputs(9078) <= not((inputs(13)) or (inputs(88)));
    layer0_outputs(9079) <= not((inputs(191)) xor (inputs(97)));
    layer0_outputs(9080) <= not((inputs(196)) and (inputs(23)));
    layer0_outputs(9081) <= '1';
    layer0_outputs(9082) <= inputs(232);
    layer0_outputs(9083) <= inputs(185);
    layer0_outputs(9084) <= not(inputs(69)) or (inputs(58));
    layer0_outputs(9085) <= (inputs(163)) or (inputs(197));
    layer0_outputs(9086) <= not(inputs(47)) or (inputs(201));
    layer0_outputs(9087) <= (inputs(8)) or (inputs(150));
    layer0_outputs(9088) <= (inputs(163)) and not (inputs(254));
    layer0_outputs(9089) <= not(inputs(197));
    layer0_outputs(9090) <= (inputs(140)) and not (inputs(177));
    layer0_outputs(9091) <= not(inputs(122)) or (inputs(224));
    layer0_outputs(9092) <= not((inputs(94)) xor (inputs(107)));
    layer0_outputs(9093) <= (inputs(192)) and not (inputs(128));
    layer0_outputs(9094) <= not(inputs(155));
    layer0_outputs(9095) <= not(inputs(138)) or (inputs(146));
    layer0_outputs(9096) <= inputs(160);
    layer0_outputs(9097) <= (inputs(179)) xor (inputs(120));
    layer0_outputs(9098) <= not((inputs(104)) xor (inputs(152)));
    layer0_outputs(9099) <= not(inputs(184));
    layer0_outputs(9100) <= inputs(249);
    layer0_outputs(9101) <= inputs(233);
    layer0_outputs(9102) <= not(inputs(77));
    layer0_outputs(9103) <= not((inputs(236)) or (inputs(194)));
    layer0_outputs(9104) <= not(inputs(136)) or (inputs(205));
    layer0_outputs(9105) <= inputs(74);
    layer0_outputs(9106) <= (inputs(83)) and not (inputs(162));
    layer0_outputs(9107) <= (inputs(187)) xor (inputs(62));
    layer0_outputs(9108) <= not((inputs(246)) and (inputs(164)));
    layer0_outputs(9109) <= inputs(101);
    layer0_outputs(9110) <= (inputs(224)) or (inputs(33));
    layer0_outputs(9111) <= '1';
    layer0_outputs(9112) <= (inputs(205)) and not (inputs(191));
    layer0_outputs(9113) <= not(inputs(145)) or (inputs(63));
    layer0_outputs(9114) <= inputs(137);
    layer0_outputs(9115) <= (inputs(54)) or (inputs(65));
    layer0_outputs(9116) <= (inputs(135)) and not (inputs(48));
    layer0_outputs(9117) <= not((inputs(61)) xor (inputs(139)));
    layer0_outputs(9118) <= (inputs(167)) and not (inputs(93));
    layer0_outputs(9119) <= inputs(4);
    layer0_outputs(9120) <= not(inputs(89));
    layer0_outputs(9121) <= (inputs(213)) and not (inputs(18));
    layer0_outputs(9122) <= inputs(37);
    layer0_outputs(9123) <= (inputs(36)) and not (inputs(222));
    layer0_outputs(9124) <= not(inputs(173));
    layer0_outputs(9125) <= not(inputs(85)) or (inputs(78));
    layer0_outputs(9126) <= (inputs(87)) and not (inputs(220));
    layer0_outputs(9127) <= (inputs(169)) or (inputs(222));
    layer0_outputs(9128) <= (inputs(29)) and not (inputs(44));
    layer0_outputs(9129) <= not((inputs(17)) or (inputs(48)));
    layer0_outputs(9130) <= not(inputs(28));
    layer0_outputs(9131) <= not(inputs(212)) or (inputs(106));
    layer0_outputs(9132) <= (inputs(170)) and not (inputs(56));
    layer0_outputs(9133) <= not((inputs(232)) xor (inputs(168)));
    layer0_outputs(9134) <= not((inputs(174)) or (inputs(44)));
    layer0_outputs(9135) <= (inputs(76)) or (inputs(212));
    layer0_outputs(9136) <= inputs(216);
    layer0_outputs(9137) <= inputs(124);
    layer0_outputs(9138) <= (inputs(124)) xor (inputs(69));
    layer0_outputs(9139) <= not(inputs(23));
    layer0_outputs(9140) <= not((inputs(105)) xor (inputs(176)));
    layer0_outputs(9141) <= not((inputs(253)) or (inputs(130)));
    layer0_outputs(9142) <= (inputs(88)) xor (inputs(144));
    layer0_outputs(9143) <= not(inputs(172));
    layer0_outputs(9144) <= not(inputs(147));
    layer0_outputs(9145) <= inputs(117);
    layer0_outputs(9146) <= not(inputs(146)) or (inputs(97));
    layer0_outputs(9147) <= not((inputs(110)) or (inputs(38)));
    layer0_outputs(9148) <= not(inputs(221)) or (inputs(14));
    layer0_outputs(9149) <= inputs(144);
    layer0_outputs(9150) <= not(inputs(91)) or (inputs(131));
    layer0_outputs(9151) <= (inputs(145)) and (inputs(129));
    layer0_outputs(9152) <= not(inputs(146));
    layer0_outputs(9153) <= not(inputs(254)) or (inputs(47));
    layer0_outputs(9154) <= inputs(129);
    layer0_outputs(9155) <= inputs(70);
    layer0_outputs(9156) <= not(inputs(130)) or (inputs(243));
    layer0_outputs(9157) <= (inputs(0)) or (inputs(131));
    layer0_outputs(9158) <= (inputs(214)) or (inputs(13));
    layer0_outputs(9159) <= not(inputs(211)) or (inputs(76));
    layer0_outputs(9160) <= not((inputs(69)) or (inputs(38)));
    layer0_outputs(9161) <= (inputs(27)) and not (inputs(178));
    layer0_outputs(9162) <= not(inputs(204)) or (inputs(81));
    layer0_outputs(9163) <= not(inputs(45));
    layer0_outputs(9164) <= not(inputs(69));
    layer0_outputs(9165) <= not((inputs(175)) xor (inputs(19)));
    layer0_outputs(9166) <= inputs(215);
    layer0_outputs(9167) <= (inputs(47)) or (inputs(226));
    layer0_outputs(9168) <= (inputs(218)) and not (inputs(253));
    layer0_outputs(9169) <= (inputs(184)) and not (inputs(59));
    layer0_outputs(9170) <= not((inputs(164)) or (inputs(186)));
    layer0_outputs(9171) <= (inputs(136)) or (inputs(120));
    layer0_outputs(9172) <= (inputs(25)) xor (inputs(99));
    layer0_outputs(9173) <= '1';
    layer0_outputs(9174) <= not((inputs(253)) xor (inputs(14)));
    layer0_outputs(9175) <= inputs(73);
    layer0_outputs(9176) <= not(inputs(84)) or (inputs(195));
    layer0_outputs(9177) <= inputs(231);
    layer0_outputs(9178) <= (inputs(52)) and not (inputs(111));
    layer0_outputs(9179) <= inputs(25);
    layer0_outputs(9180) <= not((inputs(133)) xor (inputs(198)));
    layer0_outputs(9181) <= not(inputs(161));
    layer0_outputs(9182) <= (inputs(117)) or (inputs(206));
    layer0_outputs(9183) <= (inputs(18)) or (inputs(21));
    layer0_outputs(9184) <= not((inputs(254)) xor (inputs(67)));
    layer0_outputs(9185) <= not(inputs(197));
    layer0_outputs(9186) <= not((inputs(5)) xor (inputs(156)));
    layer0_outputs(9187) <= (inputs(206)) or (inputs(208));
    layer0_outputs(9188) <= (inputs(9)) and not (inputs(10));
    layer0_outputs(9189) <= (inputs(120)) and not (inputs(55));
    layer0_outputs(9190) <= (inputs(250)) and (inputs(61));
    layer0_outputs(9191) <= (inputs(113)) or (inputs(144));
    layer0_outputs(9192) <= inputs(218);
    layer0_outputs(9193) <= not(inputs(167)) or (inputs(240));
    layer0_outputs(9194) <= not((inputs(167)) xor (inputs(131)));
    layer0_outputs(9195) <= not(inputs(229));
    layer0_outputs(9196) <= (inputs(151)) and not (inputs(112));
    layer0_outputs(9197) <= not((inputs(66)) or (inputs(218)));
    layer0_outputs(9198) <= not(inputs(39));
    layer0_outputs(9199) <= not((inputs(101)) xor (inputs(59)));
    layer0_outputs(9200) <= not((inputs(134)) and (inputs(67)));
    layer0_outputs(9201) <= (inputs(11)) or (inputs(203));
    layer0_outputs(9202) <= (inputs(215)) and not (inputs(0));
    layer0_outputs(9203) <= inputs(217);
    layer0_outputs(9204) <= (inputs(155)) or (inputs(60));
    layer0_outputs(9205) <= not((inputs(20)) xor (inputs(62)));
    layer0_outputs(9206) <= not((inputs(212)) or (inputs(249)));
    layer0_outputs(9207) <= not(inputs(232)) or (inputs(19));
    layer0_outputs(9208) <= not(inputs(172)) or (inputs(30));
    layer0_outputs(9209) <= inputs(247);
    layer0_outputs(9210) <= not((inputs(42)) xor (inputs(229)));
    layer0_outputs(9211) <= not(inputs(38));
    layer0_outputs(9212) <= not((inputs(236)) xor (inputs(6)));
    layer0_outputs(9213) <= not((inputs(18)) or (inputs(255)));
    layer0_outputs(9214) <= not(inputs(31)) or (inputs(127));
    layer0_outputs(9215) <= not((inputs(98)) or (inputs(186)));
    layer0_outputs(9216) <= not(inputs(202));
    layer0_outputs(9217) <= (inputs(145)) or (inputs(105));
    layer0_outputs(9218) <= inputs(69);
    layer0_outputs(9219) <= not(inputs(24)) or (inputs(175));
    layer0_outputs(9220) <= not((inputs(34)) or (inputs(77)));
    layer0_outputs(9221) <= '0';
    layer0_outputs(9222) <= not((inputs(176)) or (inputs(231)));
    layer0_outputs(9223) <= not(inputs(182)) or (inputs(112));
    layer0_outputs(9224) <= not(inputs(203)) or (inputs(169));
    layer0_outputs(9225) <= not(inputs(145));
    layer0_outputs(9226) <= (inputs(110)) or (inputs(10));
    layer0_outputs(9227) <= inputs(100);
    layer0_outputs(9228) <= (inputs(190)) and not (inputs(201));
    layer0_outputs(9229) <= (inputs(249)) or (inputs(132));
    layer0_outputs(9230) <= not((inputs(229)) xor (inputs(0)));
    layer0_outputs(9231) <= not((inputs(34)) xor (inputs(253)));
    layer0_outputs(9232) <= not(inputs(182)) or (inputs(144));
    layer0_outputs(9233) <= inputs(39);
    layer0_outputs(9234) <= (inputs(48)) or (inputs(8));
    layer0_outputs(9235) <= not((inputs(37)) or (inputs(49)));
    layer0_outputs(9236) <= not((inputs(219)) xor (inputs(194)));
    layer0_outputs(9237) <= inputs(133);
    layer0_outputs(9238) <= not(inputs(22)) or (inputs(144));
    layer0_outputs(9239) <= not(inputs(50));
    layer0_outputs(9240) <= not(inputs(24)) or (inputs(187));
    layer0_outputs(9241) <= inputs(137);
    layer0_outputs(9242) <= not(inputs(47));
    layer0_outputs(9243) <= not(inputs(5)) or (inputs(83));
    layer0_outputs(9244) <= not(inputs(108));
    layer0_outputs(9245) <= not((inputs(126)) or (inputs(252)));
    layer0_outputs(9246) <= not((inputs(180)) xor (inputs(212)));
    layer0_outputs(9247) <= (inputs(113)) xor (inputs(87));
    layer0_outputs(9248) <= (inputs(86)) and not (inputs(94));
    layer0_outputs(9249) <= (inputs(47)) or (inputs(251));
    layer0_outputs(9250) <= not(inputs(42));
    layer0_outputs(9251) <= (inputs(32)) and (inputs(58));
    layer0_outputs(9252) <= inputs(169);
    layer0_outputs(9253) <= inputs(68);
    layer0_outputs(9254) <= not(inputs(19));
    layer0_outputs(9255) <= not((inputs(79)) or (inputs(57)));
    layer0_outputs(9256) <= not((inputs(242)) or (inputs(5)));
    layer0_outputs(9257) <= (inputs(119)) and not (inputs(32));
    layer0_outputs(9258) <= not(inputs(104));
    layer0_outputs(9259) <= not(inputs(71));
    layer0_outputs(9260) <= (inputs(175)) or (inputs(124));
    layer0_outputs(9261) <= (inputs(60)) and not (inputs(179));
    layer0_outputs(9262) <= not(inputs(115));
    layer0_outputs(9263) <= (inputs(135)) or (inputs(213));
    layer0_outputs(9264) <= inputs(126);
    layer0_outputs(9265) <= not((inputs(85)) xor (inputs(83)));
    layer0_outputs(9266) <= (inputs(34)) or (inputs(63));
    layer0_outputs(9267) <= not(inputs(238));
    layer0_outputs(9268) <= not(inputs(179));
    layer0_outputs(9269) <= not((inputs(34)) and (inputs(44)));
    layer0_outputs(9270) <= (inputs(145)) xor (inputs(131));
    layer0_outputs(9271) <= (inputs(200)) and not (inputs(54));
    layer0_outputs(9272) <= (inputs(245)) or (inputs(25));
    layer0_outputs(9273) <= (inputs(92)) and not (inputs(252));
    layer0_outputs(9274) <= not((inputs(227)) or (inputs(63)));
    layer0_outputs(9275) <= inputs(54);
    layer0_outputs(9276) <= (inputs(99)) or (inputs(254));
    layer0_outputs(9277) <= not((inputs(180)) xor (inputs(50)));
    layer0_outputs(9278) <= not((inputs(44)) xor (inputs(116)));
    layer0_outputs(9279) <= not(inputs(18));
    layer0_outputs(9280) <= (inputs(28)) and not (inputs(162));
    layer0_outputs(9281) <= inputs(6);
    layer0_outputs(9282) <= not((inputs(36)) xor (inputs(20)));
    layer0_outputs(9283) <= inputs(86);
    layer0_outputs(9284) <= (inputs(54)) and not (inputs(149));
    layer0_outputs(9285) <= not(inputs(171)) or (inputs(71));
    layer0_outputs(9286) <= inputs(212);
    layer0_outputs(9287) <= not(inputs(203));
    layer0_outputs(9288) <= not((inputs(7)) xor (inputs(33)));
    layer0_outputs(9289) <= not(inputs(107));
    layer0_outputs(9290) <= not((inputs(103)) or (inputs(242)));
    layer0_outputs(9291) <= (inputs(55)) or (inputs(97));
    layer0_outputs(9292) <= not((inputs(142)) or (inputs(111)));
    layer0_outputs(9293) <= not((inputs(174)) or (inputs(151)));
    layer0_outputs(9294) <= (inputs(138)) and not (inputs(224));
    layer0_outputs(9295) <= not(inputs(251)) or (inputs(234));
    layer0_outputs(9296) <= not((inputs(193)) or (inputs(239)));
    layer0_outputs(9297) <= not((inputs(184)) xor (inputs(217)));
    layer0_outputs(9298) <= inputs(215);
    layer0_outputs(9299) <= not((inputs(252)) or (inputs(237)));
    layer0_outputs(9300) <= not((inputs(216)) xor (inputs(186)));
    layer0_outputs(9301) <= not(inputs(203));
    layer0_outputs(9302) <= not(inputs(238));
    layer0_outputs(9303) <= (inputs(249)) and not (inputs(73));
    layer0_outputs(9304) <= (inputs(49)) or (inputs(53));
    layer0_outputs(9305) <= (inputs(121)) and not (inputs(32));
    layer0_outputs(9306) <= (inputs(123)) xor (inputs(156));
    layer0_outputs(9307) <= (inputs(178)) or (inputs(208));
    layer0_outputs(9308) <= not((inputs(3)) xor (inputs(124)));
    layer0_outputs(9309) <= not((inputs(33)) or (inputs(212)));
    layer0_outputs(9310) <= not((inputs(172)) or (inputs(20)));
    layer0_outputs(9311) <= not((inputs(107)) and (inputs(157)));
    layer0_outputs(9312) <= inputs(9);
    layer0_outputs(9313) <= not((inputs(44)) or (inputs(90)));
    layer0_outputs(9314) <= not((inputs(1)) or (inputs(203)));
    layer0_outputs(9315) <= (inputs(78)) xor (inputs(79));
    layer0_outputs(9316) <= not((inputs(248)) or (inputs(66)));
    layer0_outputs(9317) <= (inputs(138)) and not (inputs(120));
    layer0_outputs(9318) <= not((inputs(118)) or (inputs(204)));
    layer0_outputs(9319) <= (inputs(142)) or (inputs(195));
    layer0_outputs(9320) <= inputs(249);
    layer0_outputs(9321) <= not(inputs(190)) or (inputs(96));
    layer0_outputs(9322) <= (inputs(107)) or (inputs(70));
    layer0_outputs(9323) <= not(inputs(8)) or (inputs(210));
    layer0_outputs(9324) <= not((inputs(196)) or (inputs(14)));
    layer0_outputs(9325) <= (inputs(184)) and not (inputs(156));
    layer0_outputs(9326) <= not(inputs(74)) or (inputs(87));
    layer0_outputs(9327) <= (inputs(217)) or (inputs(211));
    layer0_outputs(9328) <= (inputs(28)) xor (inputs(72));
    layer0_outputs(9329) <= not((inputs(148)) or (inputs(116)));
    layer0_outputs(9330) <= not(inputs(24));
    layer0_outputs(9331) <= not(inputs(214));
    layer0_outputs(9332) <= not(inputs(204)) or (inputs(35));
    layer0_outputs(9333) <= inputs(29);
    layer0_outputs(9334) <= not(inputs(110));
    layer0_outputs(9335) <= (inputs(11)) and not (inputs(200));
    layer0_outputs(9336) <= not((inputs(30)) xor (inputs(34)));
    layer0_outputs(9337) <= (inputs(182)) and not (inputs(207));
    layer0_outputs(9338) <= not(inputs(76));
    layer0_outputs(9339) <= inputs(164);
    layer0_outputs(9340) <= not((inputs(178)) or (inputs(216)));
    layer0_outputs(9341) <= inputs(21);
    layer0_outputs(9342) <= (inputs(194)) xor (inputs(217));
    layer0_outputs(9343) <= not(inputs(190)) or (inputs(126));
    layer0_outputs(9344) <= not(inputs(25)) or (inputs(241));
    layer0_outputs(9345) <= not((inputs(40)) or (inputs(58)));
    layer0_outputs(9346) <= inputs(66);
    layer0_outputs(9347) <= not((inputs(206)) or (inputs(7)));
    layer0_outputs(9348) <= not((inputs(206)) or (inputs(90)));
    layer0_outputs(9349) <= not((inputs(159)) or (inputs(4)));
    layer0_outputs(9350) <= (inputs(143)) xor (inputs(136));
    layer0_outputs(9351) <= inputs(55);
    layer0_outputs(9352) <= (inputs(236)) xor (inputs(125));
    layer0_outputs(9353) <= (inputs(84)) and not (inputs(175));
    layer0_outputs(9354) <= not((inputs(183)) or (inputs(183)));
    layer0_outputs(9355) <= inputs(136);
    layer0_outputs(9356) <= not((inputs(75)) xor (inputs(146)));
    layer0_outputs(9357) <= (inputs(214)) and not (inputs(87));
    layer0_outputs(9358) <= inputs(78);
    layer0_outputs(9359) <= not(inputs(54)) or (inputs(156));
    layer0_outputs(9360) <= not(inputs(142));
    layer0_outputs(9361) <= (inputs(64)) or (inputs(151));
    layer0_outputs(9362) <= not((inputs(247)) or (inputs(41)));
    layer0_outputs(9363) <= not((inputs(61)) xor (inputs(104)));
    layer0_outputs(9364) <= not(inputs(156)) or (inputs(233));
    layer0_outputs(9365) <= not((inputs(96)) or (inputs(10)));
    layer0_outputs(9366) <= not(inputs(254));
    layer0_outputs(9367) <= not(inputs(154));
    layer0_outputs(9368) <= (inputs(17)) or (inputs(12));
    layer0_outputs(9369) <= not((inputs(251)) xor (inputs(171)));
    layer0_outputs(9370) <= inputs(13);
    layer0_outputs(9371) <= inputs(212);
    layer0_outputs(9372) <= (inputs(43)) xor (inputs(76));
    layer0_outputs(9373) <= not((inputs(102)) and (inputs(214)));
    layer0_outputs(9374) <= not(inputs(151)) or (inputs(94));
    layer0_outputs(9375) <= not(inputs(228)) or (inputs(5));
    layer0_outputs(9376) <= not(inputs(59));
    layer0_outputs(9377) <= (inputs(100)) and not (inputs(72));
    layer0_outputs(9378) <= inputs(230);
    layer0_outputs(9379) <= (inputs(232)) or (inputs(128));
    layer0_outputs(9380) <= not((inputs(27)) xor (inputs(9)));
    layer0_outputs(9381) <= not(inputs(141));
    layer0_outputs(9382) <= not(inputs(174)) or (inputs(41));
    layer0_outputs(9383) <= (inputs(150)) or (inputs(149));
    layer0_outputs(9384) <= (inputs(118)) or (inputs(93));
    layer0_outputs(9385) <= '0';
    layer0_outputs(9386) <= inputs(211);
    layer0_outputs(9387) <= (inputs(73)) and not (inputs(65));
    layer0_outputs(9388) <= not(inputs(236));
    layer0_outputs(9389) <= (inputs(47)) and not (inputs(152));
    layer0_outputs(9390) <= (inputs(16)) and not (inputs(242));
    layer0_outputs(9391) <= not(inputs(167)) or (inputs(176));
    layer0_outputs(9392) <= not(inputs(214)) or (inputs(217));
    layer0_outputs(9393) <= not((inputs(181)) xor (inputs(200)));
    layer0_outputs(9394) <= not(inputs(68)) or (inputs(134));
    layer0_outputs(9395) <= (inputs(241)) or (inputs(137));
    layer0_outputs(9396) <= not((inputs(231)) or (inputs(80)));
    layer0_outputs(9397) <= not((inputs(64)) or (inputs(209)));
    layer0_outputs(9398) <= (inputs(12)) and not (inputs(26));
    layer0_outputs(9399) <= (inputs(228)) xor (inputs(177));
    layer0_outputs(9400) <= not((inputs(106)) or (inputs(5)));
    layer0_outputs(9401) <= not((inputs(27)) xor (inputs(161)));
    layer0_outputs(9402) <= not((inputs(102)) or (inputs(105)));
    layer0_outputs(9403) <= not((inputs(20)) xor (inputs(187)));
    layer0_outputs(9404) <= not(inputs(232));
    layer0_outputs(9405) <= (inputs(56)) and not (inputs(12));
    layer0_outputs(9406) <= not(inputs(83));
    layer0_outputs(9407) <= (inputs(123)) and not (inputs(174));
    layer0_outputs(9408) <= not(inputs(21)) or (inputs(115));
    layer0_outputs(9409) <= inputs(207);
    layer0_outputs(9410) <= not((inputs(84)) or (inputs(19)));
    layer0_outputs(9411) <= '0';
    layer0_outputs(9412) <= not((inputs(247)) xor (inputs(216)));
    layer0_outputs(9413) <= not(inputs(92));
    layer0_outputs(9414) <= (inputs(202)) xor (inputs(160));
    layer0_outputs(9415) <= (inputs(23)) or (inputs(252));
    layer0_outputs(9416) <= (inputs(184)) and not (inputs(86));
    layer0_outputs(9417) <= not((inputs(204)) xor (inputs(135)));
    layer0_outputs(9418) <= not((inputs(250)) xor (inputs(36)));
    layer0_outputs(9419) <= not((inputs(125)) and (inputs(194)));
    layer0_outputs(9420) <= (inputs(72)) and not (inputs(3));
    layer0_outputs(9421) <= not(inputs(51));
    layer0_outputs(9422) <= not(inputs(252));
    layer0_outputs(9423) <= (inputs(225)) xor (inputs(173));
    layer0_outputs(9424) <= not((inputs(184)) or (inputs(96)));
    layer0_outputs(9425) <= (inputs(67)) or (inputs(106));
    layer0_outputs(9426) <= inputs(103);
    layer0_outputs(9427) <= not(inputs(117));
    layer0_outputs(9428) <= inputs(218);
    layer0_outputs(9429) <= not(inputs(11));
    layer0_outputs(9430) <= inputs(111);
    layer0_outputs(9431) <= (inputs(40)) or (inputs(193));
    layer0_outputs(9432) <= not(inputs(56)) or (inputs(160));
    layer0_outputs(9433) <= not(inputs(136)) or (inputs(30));
    layer0_outputs(9434) <= (inputs(211)) or (inputs(209));
    layer0_outputs(9435) <= (inputs(209)) xor (inputs(206));
    layer0_outputs(9436) <= inputs(230);
    layer0_outputs(9437) <= not(inputs(201));
    layer0_outputs(9438) <= (inputs(247)) xor (inputs(182));
    layer0_outputs(9439) <= not((inputs(198)) or (inputs(143)));
    layer0_outputs(9440) <= not((inputs(116)) xor (inputs(114)));
    layer0_outputs(9441) <= (inputs(97)) and (inputs(120));
    layer0_outputs(9442) <= not(inputs(132));
    layer0_outputs(9443) <= (inputs(210)) or (inputs(18));
    layer0_outputs(9444) <= not(inputs(238));
    layer0_outputs(9445) <= '1';
    layer0_outputs(9446) <= not((inputs(74)) xor (inputs(127)));
    layer0_outputs(9447) <= inputs(9);
    layer0_outputs(9448) <= (inputs(56)) or (inputs(228));
    layer0_outputs(9449) <= (inputs(172)) xor (inputs(196));
    layer0_outputs(9450) <= not(inputs(40));
    layer0_outputs(9451) <= not((inputs(251)) xor (inputs(219)));
    layer0_outputs(9452) <= not(inputs(143));
    layer0_outputs(9453) <= not(inputs(38)) or (inputs(34));
    layer0_outputs(9454) <= inputs(111);
    layer0_outputs(9455) <= not(inputs(113)) or (inputs(62));
    layer0_outputs(9456) <= (inputs(238)) or (inputs(62));
    layer0_outputs(9457) <= (inputs(204)) xor (inputs(121));
    layer0_outputs(9458) <= (inputs(231)) and not (inputs(251));
    layer0_outputs(9459) <= not((inputs(60)) xor (inputs(93)));
    layer0_outputs(9460) <= (inputs(238)) or (inputs(100));
    layer0_outputs(9461) <= not((inputs(30)) xor (inputs(254)));
    layer0_outputs(9462) <= not(inputs(75));
    layer0_outputs(9463) <= (inputs(152)) and not (inputs(10));
    layer0_outputs(9464) <= not(inputs(74));
    layer0_outputs(9465) <= not((inputs(194)) or (inputs(185)));
    layer0_outputs(9466) <= not(inputs(184));
    layer0_outputs(9467) <= (inputs(165)) xor (inputs(241));
    layer0_outputs(9468) <= (inputs(87)) xor (inputs(189));
    layer0_outputs(9469) <= (inputs(85)) and not (inputs(94));
    layer0_outputs(9470) <= (inputs(233)) or (inputs(101));
    layer0_outputs(9471) <= (inputs(180)) and not (inputs(112));
    layer0_outputs(9472) <= not(inputs(26)) or (inputs(200));
    layer0_outputs(9473) <= inputs(162);
    layer0_outputs(9474) <= not(inputs(176));
    layer0_outputs(9475) <= (inputs(55)) and not (inputs(48));
    layer0_outputs(9476) <= not((inputs(46)) xor (inputs(201)));
    layer0_outputs(9477) <= not((inputs(199)) xor (inputs(230)));
    layer0_outputs(9478) <= (inputs(247)) and not (inputs(127));
    layer0_outputs(9479) <= (inputs(216)) or (inputs(224));
    layer0_outputs(9480) <= (inputs(39)) xor (inputs(64));
    layer0_outputs(9481) <= (inputs(177)) xor (inputs(68));
    layer0_outputs(9482) <= (inputs(201)) or (inputs(207));
    layer0_outputs(9483) <= (inputs(227)) or (inputs(23));
    layer0_outputs(9484) <= not((inputs(117)) and (inputs(36)));
    layer0_outputs(9485) <= not((inputs(187)) xor (inputs(28)));
    layer0_outputs(9486) <= not(inputs(6));
    layer0_outputs(9487) <= not(inputs(37)) or (inputs(250));
    layer0_outputs(9488) <= not(inputs(114));
    layer0_outputs(9489) <= not((inputs(223)) xor (inputs(190)));
    layer0_outputs(9490) <= not(inputs(46));
    layer0_outputs(9491) <= not(inputs(194));
    layer0_outputs(9492) <= not((inputs(119)) or (inputs(22)));
    layer0_outputs(9493) <= not((inputs(38)) or (inputs(111)));
    layer0_outputs(9494) <= '1';
    layer0_outputs(9495) <= (inputs(133)) and not (inputs(239));
    layer0_outputs(9496) <= inputs(90);
    layer0_outputs(9497) <= inputs(196);
    layer0_outputs(9498) <= not((inputs(243)) or (inputs(208)));
    layer0_outputs(9499) <= not(inputs(39));
    layer0_outputs(9500) <= not(inputs(181));
    layer0_outputs(9501) <= not((inputs(168)) and (inputs(250)));
    layer0_outputs(9502) <= not((inputs(65)) or (inputs(13)));
    layer0_outputs(9503) <= not(inputs(2));
    layer0_outputs(9504) <= not(inputs(208)) or (inputs(253));
    layer0_outputs(9505) <= (inputs(39)) and not (inputs(251));
    layer0_outputs(9506) <= not((inputs(223)) or (inputs(215)));
    layer0_outputs(9507) <= (inputs(109)) and not (inputs(250));
    layer0_outputs(9508) <= not((inputs(212)) or (inputs(11)));
    layer0_outputs(9509) <= not((inputs(180)) and (inputs(252)));
    layer0_outputs(9510) <= not((inputs(88)) xor (inputs(62)));
    layer0_outputs(9511) <= (inputs(252)) or (inputs(69));
    layer0_outputs(9512) <= (inputs(59)) and not (inputs(239));
    layer0_outputs(9513) <= not((inputs(90)) xor (inputs(125)));
    layer0_outputs(9514) <= not(inputs(61));
    layer0_outputs(9515) <= not((inputs(56)) or (inputs(125)));
    layer0_outputs(9516) <= not(inputs(183));
    layer0_outputs(9517) <= (inputs(124)) and not (inputs(220));
    layer0_outputs(9518) <= '0';
    layer0_outputs(9519) <= not((inputs(190)) or (inputs(107)));
    layer0_outputs(9520) <= not((inputs(127)) or (inputs(206)));
    layer0_outputs(9521) <= not((inputs(171)) or (inputs(186)));
    layer0_outputs(9522) <= (inputs(79)) xor (inputs(222));
    layer0_outputs(9523) <= not(inputs(236));
    layer0_outputs(9524) <= not((inputs(228)) xor (inputs(183)));
    layer0_outputs(9525) <= not(inputs(63)) or (inputs(215));
    layer0_outputs(9526) <= inputs(65);
    layer0_outputs(9527) <= not(inputs(109));
    layer0_outputs(9528) <= (inputs(149)) and not (inputs(239));
    layer0_outputs(9529) <= (inputs(83)) and not (inputs(93));
    layer0_outputs(9530) <= (inputs(16)) xor (inputs(129));
    layer0_outputs(9531) <= inputs(56);
    layer0_outputs(9532) <= (inputs(39)) and not (inputs(0));
    layer0_outputs(9533) <= not((inputs(191)) xor (inputs(161)));
    layer0_outputs(9534) <= not((inputs(52)) xor (inputs(148)));
    layer0_outputs(9535) <= not((inputs(195)) xor (inputs(203)));
    layer0_outputs(9536) <= not((inputs(218)) or (inputs(156)));
    layer0_outputs(9537) <= inputs(146);
    layer0_outputs(9538) <= not(inputs(181)) or (inputs(171));
    layer0_outputs(9539) <= not(inputs(119));
    layer0_outputs(9540) <= (inputs(66)) and not (inputs(237));
    layer0_outputs(9541) <= not(inputs(177));
    layer0_outputs(9542) <= not(inputs(132)) or (inputs(220));
    layer0_outputs(9543) <= not(inputs(69));
    layer0_outputs(9544) <= (inputs(15)) or (inputs(65));
    layer0_outputs(9545) <= not((inputs(235)) xor (inputs(218)));
    layer0_outputs(9546) <= inputs(25);
    layer0_outputs(9547) <= (inputs(41)) or (inputs(57));
    layer0_outputs(9548) <= (inputs(158)) or (inputs(218));
    layer0_outputs(9549) <= inputs(216);
    layer0_outputs(9550) <= (inputs(174)) xor (inputs(21));
    layer0_outputs(9551) <= not(inputs(3));
    layer0_outputs(9552) <= (inputs(16)) or (inputs(36));
    layer0_outputs(9553) <= not((inputs(36)) and (inputs(34)));
    layer0_outputs(9554) <= not(inputs(59)) or (inputs(102));
    layer0_outputs(9555) <= not((inputs(98)) xor (inputs(186)));
    layer0_outputs(9556) <= not(inputs(166));
    layer0_outputs(9557) <= inputs(191);
    layer0_outputs(9558) <= inputs(35);
    layer0_outputs(9559) <= (inputs(97)) xor (inputs(149));
    layer0_outputs(9560) <= (inputs(249)) and not (inputs(77));
    layer0_outputs(9561) <= not(inputs(89));
    layer0_outputs(9562) <= not(inputs(252));
    layer0_outputs(9563) <= not(inputs(234));
    layer0_outputs(9564) <= (inputs(238)) or (inputs(165));
    layer0_outputs(9565) <= (inputs(74)) and not (inputs(204));
    layer0_outputs(9566) <= (inputs(169)) xor (inputs(150));
    layer0_outputs(9567) <= not(inputs(71));
    layer0_outputs(9568) <= not(inputs(60));
    layer0_outputs(9569) <= not((inputs(189)) or (inputs(154)));
    layer0_outputs(9570) <= not((inputs(198)) or (inputs(189)));
    layer0_outputs(9571) <= not((inputs(218)) xor (inputs(190)));
    layer0_outputs(9572) <= inputs(9);
    layer0_outputs(9573) <= not((inputs(174)) xor (inputs(236)));
    layer0_outputs(9574) <= (inputs(157)) xor (inputs(83));
    layer0_outputs(9575) <= (inputs(120)) and not (inputs(111));
    layer0_outputs(9576) <= (inputs(150)) or (inputs(211));
    layer0_outputs(9577) <= (inputs(128)) xor (inputs(158));
    layer0_outputs(9578) <= not(inputs(73));
    layer0_outputs(9579) <= not(inputs(192)) or (inputs(17));
    layer0_outputs(9580) <= (inputs(215)) and not (inputs(54));
    layer0_outputs(9581) <= not((inputs(101)) and (inputs(60)));
    layer0_outputs(9582) <= inputs(146);
    layer0_outputs(9583) <= not(inputs(163));
    layer0_outputs(9584) <= not(inputs(139));
    layer0_outputs(9585) <= not((inputs(219)) xor (inputs(211)));
    layer0_outputs(9586) <= not(inputs(10)) or (inputs(205));
    layer0_outputs(9587) <= (inputs(21)) and not (inputs(55));
    layer0_outputs(9588) <= (inputs(154)) or (inputs(168));
    layer0_outputs(9589) <= (inputs(202)) xor (inputs(121));
    layer0_outputs(9590) <= (inputs(71)) and (inputs(199));
    layer0_outputs(9591) <= not((inputs(109)) xor (inputs(219)));
    layer0_outputs(9592) <= not(inputs(223));
    layer0_outputs(9593) <= (inputs(7)) or (inputs(22));
    layer0_outputs(9594) <= not(inputs(160));
    layer0_outputs(9595) <= (inputs(44)) and not (inputs(250));
    layer0_outputs(9596) <= not((inputs(213)) or (inputs(205)));
    layer0_outputs(9597) <= not((inputs(91)) xor (inputs(60)));
    layer0_outputs(9598) <= not(inputs(14));
    layer0_outputs(9599) <= (inputs(254)) xor (inputs(95));
    layer0_outputs(9600) <= not(inputs(55));
    layer0_outputs(9601) <= not((inputs(183)) xor (inputs(184)));
    layer0_outputs(9602) <= (inputs(102)) xor (inputs(112));
    layer0_outputs(9603) <= (inputs(210)) or (inputs(186));
    layer0_outputs(9604) <= (inputs(221)) and not (inputs(18));
    layer0_outputs(9605) <= (inputs(216)) or (inputs(189));
    layer0_outputs(9606) <= inputs(179);
    layer0_outputs(9607) <= (inputs(23)) and not (inputs(222));
    layer0_outputs(9608) <= (inputs(182)) and not (inputs(83));
    layer0_outputs(9609) <= not(inputs(171));
    layer0_outputs(9610) <= inputs(124);
    layer0_outputs(9611) <= not(inputs(66));
    layer0_outputs(9612) <= not((inputs(40)) or (inputs(55)));
    layer0_outputs(9613) <= not(inputs(45));
    layer0_outputs(9614) <= (inputs(81)) or (inputs(246));
    layer0_outputs(9615) <= '0';
    layer0_outputs(9616) <= not(inputs(145)) or (inputs(239));
    layer0_outputs(9617) <= not(inputs(225));
    layer0_outputs(9618) <= inputs(160);
    layer0_outputs(9619) <= not(inputs(28));
    layer0_outputs(9620) <= inputs(65);
    layer0_outputs(9621) <= not(inputs(133)) or (inputs(125));
    layer0_outputs(9622) <= inputs(40);
    layer0_outputs(9623) <= (inputs(247)) and not (inputs(81));
    layer0_outputs(9624) <= (inputs(92)) and not (inputs(244));
    layer0_outputs(9625) <= (inputs(86)) or (inputs(251));
    layer0_outputs(9626) <= not(inputs(108)) or (inputs(243));
    layer0_outputs(9627) <= inputs(114);
    layer0_outputs(9628) <= not((inputs(47)) or (inputs(251)));
    layer0_outputs(9629) <= not((inputs(117)) xor (inputs(232)));
    layer0_outputs(9630) <= inputs(128);
    layer0_outputs(9631) <= not(inputs(127));
    layer0_outputs(9632) <= not(inputs(193));
    layer0_outputs(9633) <= (inputs(61)) and not (inputs(255));
    layer0_outputs(9634) <= inputs(38);
    layer0_outputs(9635) <= not(inputs(198));
    layer0_outputs(9636) <= not(inputs(163));
    layer0_outputs(9637) <= not(inputs(94));
    layer0_outputs(9638) <= not(inputs(79)) or (inputs(236));
    layer0_outputs(9639) <= (inputs(42)) xor (inputs(75));
    layer0_outputs(9640) <= (inputs(80)) or (inputs(50));
    layer0_outputs(9641) <= (inputs(178)) xor (inputs(198));
    layer0_outputs(9642) <= (inputs(90)) and not (inputs(128));
    layer0_outputs(9643) <= not((inputs(171)) or (inputs(112)));
    layer0_outputs(9644) <= inputs(78);
    layer0_outputs(9645) <= not(inputs(118));
    layer0_outputs(9646) <= not((inputs(12)) or (inputs(224)));
    layer0_outputs(9647) <= not(inputs(219)) or (inputs(147));
    layer0_outputs(9648) <= not((inputs(68)) or (inputs(15)));
    layer0_outputs(9649) <= not(inputs(138)) or (inputs(111));
    layer0_outputs(9650) <= (inputs(221)) xor (inputs(248));
    layer0_outputs(9651) <= inputs(100);
    layer0_outputs(9652) <= not(inputs(70)) or (inputs(223));
    layer0_outputs(9653) <= not(inputs(40));
    layer0_outputs(9654) <= not((inputs(19)) or (inputs(56)));
    layer0_outputs(9655) <= (inputs(235)) or (inputs(252));
    layer0_outputs(9656) <= inputs(180);
    layer0_outputs(9657) <= not((inputs(186)) xor (inputs(105)));
    layer0_outputs(9658) <= (inputs(237)) xor (inputs(90));
    layer0_outputs(9659) <= not(inputs(229)) or (inputs(42));
    layer0_outputs(9660) <= not((inputs(137)) xor (inputs(189)));
    layer0_outputs(9661) <= not((inputs(80)) xor (inputs(91)));
    layer0_outputs(9662) <= inputs(36);
    layer0_outputs(9663) <= (inputs(204)) and not (inputs(152));
    layer0_outputs(9664) <= not((inputs(109)) or (inputs(85)));
    layer0_outputs(9665) <= inputs(210);
    layer0_outputs(9666) <= not(inputs(179)) or (inputs(130));
    layer0_outputs(9667) <= (inputs(194)) or (inputs(3));
    layer0_outputs(9668) <= not((inputs(56)) and (inputs(30)));
    layer0_outputs(9669) <= not(inputs(20)) or (inputs(207));
    layer0_outputs(9670) <= '0';
    layer0_outputs(9671) <= not(inputs(114));
    layer0_outputs(9672) <= not((inputs(96)) or (inputs(96)));
    layer0_outputs(9673) <= not((inputs(123)) or (inputs(63)));
    layer0_outputs(9674) <= (inputs(162)) or (inputs(108));
    layer0_outputs(9675) <= not((inputs(112)) or (inputs(124)));
    layer0_outputs(9676) <= not((inputs(130)) xor (inputs(103)));
    layer0_outputs(9677) <= '1';
    layer0_outputs(9678) <= (inputs(70)) and not (inputs(163));
    layer0_outputs(9679) <= (inputs(93)) and not (inputs(208));
    layer0_outputs(9680) <= inputs(246);
    layer0_outputs(9681) <= inputs(104);
    layer0_outputs(9682) <= not(inputs(216)) or (inputs(126));
    layer0_outputs(9683) <= not((inputs(49)) or (inputs(167)));
    layer0_outputs(9684) <= (inputs(212)) or (inputs(148));
    layer0_outputs(9685) <= not(inputs(34));
    layer0_outputs(9686) <= not((inputs(137)) xor (inputs(170)));
    layer0_outputs(9687) <= (inputs(50)) and not (inputs(1));
    layer0_outputs(9688) <= not(inputs(90)) or (inputs(55));
    layer0_outputs(9689) <= (inputs(235)) xor (inputs(193));
    layer0_outputs(9690) <= not(inputs(12)) or (inputs(232));
    layer0_outputs(9691) <= (inputs(190)) and not (inputs(168));
    layer0_outputs(9692) <= not((inputs(171)) or (inputs(188)));
    layer0_outputs(9693) <= inputs(152);
    layer0_outputs(9694) <= inputs(248);
    layer0_outputs(9695) <= not(inputs(60));
    layer0_outputs(9696) <= inputs(85);
    layer0_outputs(9697) <= (inputs(85)) and not (inputs(2));
    layer0_outputs(9698) <= inputs(155);
    layer0_outputs(9699) <= not(inputs(199)) or (inputs(95));
    layer0_outputs(9700) <= (inputs(94)) or (inputs(248));
    layer0_outputs(9701) <= (inputs(88)) and (inputs(142));
    layer0_outputs(9702) <= not((inputs(157)) xor (inputs(4)));
    layer0_outputs(9703) <= not(inputs(167));
    layer0_outputs(9704) <= not((inputs(139)) xor (inputs(4)));
    layer0_outputs(9705) <= inputs(73);
    layer0_outputs(9706) <= not(inputs(115));
    layer0_outputs(9707) <= inputs(240);
    layer0_outputs(9708) <= (inputs(16)) and not (inputs(18));
    layer0_outputs(9709) <= not(inputs(25));
    layer0_outputs(9710) <= not(inputs(135)) or (inputs(143));
    layer0_outputs(9711) <= not((inputs(50)) or (inputs(235)));
    layer0_outputs(9712) <= (inputs(80)) and not (inputs(72));
    layer0_outputs(9713) <= (inputs(87)) and not (inputs(179));
    layer0_outputs(9714) <= not(inputs(226));
    layer0_outputs(9715) <= '1';
    layer0_outputs(9716) <= inputs(134);
    layer0_outputs(9717) <= not((inputs(140)) xor (inputs(94)));
    layer0_outputs(9718) <= inputs(234);
    layer0_outputs(9719) <= inputs(227);
    layer0_outputs(9720) <= (inputs(165)) xor (inputs(237));
    layer0_outputs(9721) <= not(inputs(223));
    layer0_outputs(9722) <= (inputs(22)) or (inputs(188));
    layer0_outputs(9723) <= (inputs(99)) xor (inputs(53));
    layer0_outputs(9724) <= not((inputs(196)) and (inputs(235)));
    layer0_outputs(9725) <= not(inputs(118)) or (inputs(237));
    layer0_outputs(9726) <= inputs(8);
    layer0_outputs(9727) <= not(inputs(211));
    layer0_outputs(9728) <= (inputs(107)) xor (inputs(59));
    layer0_outputs(9729) <= (inputs(117)) and not (inputs(93));
    layer0_outputs(9730) <= (inputs(100)) xor (inputs(102));
    layer0_outputs(9731) <= not((inputs(247)) or (inputs(208)));
    layer0_outputs(9732) <= (inputs(184)) or (inputs(190));
    layer0_outputs(9733) <= (inputs(106)) or (inputs(116));
    layer0_outputs(9734) <= not(inputs(122));
    layer0_outputs(9735) <= not((inputs(207)) xor (inputs(17)));
    layer0_outputs(9736) <= (inputs(212)) or (inputs(196));
    layer0_outputs(9737) <= not(inputs(164));
    layer0_outputs(9738) <= (inputs(57)) and not (inputs(77));
    layer0_outputs(9739) <= not((inputs(123)) xor (inputs(238)));
    layer0_outputs(9740) <= not((inputs(38)) and (inputs(122)));
    layer0_outputs(9741) <= not(inputs(123)) or (inputs(6));
    layer0_outputs(9742) <= (inputs(227)) and not (inputs(49));
    layer0_outputs(9743) <= not((inputs(113)) xor (inputs(118)));
    layer0_outputs(9744) <= not((inputs(134)) xor (inputs(117)));
    layer0_outputs(9745) <= not((inputs(243)) or (inputs(167)));
    layer0_outputs(9746) <= inputs(89);
    layer0_outputs(9747) <= not(inputs(12)) or (inputs(153));
    layer0_outputs(9748) <= (inputs(160)) or (inputs(97));
    layer0_outputs(9749) <= not(inputs(59)) or (inputs(2));
    layer0_outputs(9750) <= (inputs(242)) or (inputs(170));
    layer0_outputs(9751) <= (inputs(237)) and not (inputs(127));
    layer0_outputs(9752) <= not(inputs(58));
    layer0_outputs(9753) <= inputs(178);
    layer0_outputs(9754) <= inputs(52);
    layer0_outputs(9755) <= not(inputs(207)) or (inputs(205));
    layer0_outputs(9756) <= not((inputs(119)) and (inputs(180)));
    layer0_outputs(9757) <= (inputs(142)) or (inputs(144));
    layer0_outputs(9758) <= not(inputs(87));
    layer0_outputs(9759) <= not((inputs(255)) or (inputs(167)));
    layer0_outputs(9760) <= inputs(99);
    layer0_outputs(9761) <= inputs(144);
    layer0_outputs(9762) <= (inputs(191)) or (inputs(202));
    layer0_outputs(9763) <= (inputs(53)) or (inputs(5));
    layer0_outputs(9764) <= (inputs(201)) and not (inputs(47));
    layer0_outputs(9765) <= not(inputs(176));
    layer0_outputs(9766) <= not(inputs(22));
    layer0_outputs(9767) <= inputs(90);
    layer0_outputs(9768) <= (inputs(70)) xor (inputs(106));
    layer0_outputs(9769) <= inputs(95);
    layer0_outputs(9770) <= (inputs(201)) xor (inputs(214));
    layer0_outputs(9771) <= (inputs(61)) and not (inputs(124));
    layer0_outputs(9772) <= not((inputs(25)) xor (inputs(193)));
    layer0_outputs(9773) <= not(inputs(151)) or (inputs(145));
    layer0_outputs(9774) <= (inputs(142)) or (inputs(227));
    layer0_outputs(9775) <= inputs(126);
    layer0_outputs(9776) <= inputs(84);
    layer0_outputs(9777) <= not(inputs(54));
    layer0_outputs(9778) <= not((inputs(220)) xor (inputs(217)));
    layer0_outputs(9779) <= (inputs(245)) and (inputs(163));
    layer0_outputs(9780) <= not(inputs(122)) or (inputs(255));
    layer0_outputs(9781) <= not((inputs(88)) or (inputs(22)));
    layer0_outputs(9782) <= not(inputs(229));
    layer0_outputs(9783) <= inputs(212);
    layer0_outputs(9784) <= inputs(37);
    layer0_outputs(9785) <= not(inputs(197)) or (inputs(51));
    layer0_outputs(9786) <= (inputs(222)) or (inputs(136));
    layer0_outputs(9787) <= (inputs(167)) and not (inputs(118));
    layer0_outputs(9788) <= '0';
    layer0_outputs(9789) <= (inputs(84)) and not (inputs(160));
    layer0_outputs(9790) <= not(inputs(229)) or (inputs(6));
    layer0_outputs(9791) <= (inputs(182)) and not (inputs(208));
    layer0_outputs(9792) <= not(inputs(177));
    layer0_outputs(9793) <= not((inputs(154)) and (inputs(192)));
    layer0_outputs(9794) <= not(inputs(248)) or (inputs(41));
    layer0_outputs(9795) <= not((inputs(43)) xor (inputs(62)));
    layer0_outputs(9796) <= (inputs(79)) and not (inputs(240));
    layer0_outputs(9797) <= not((inputs(49)) or (inputs(121)));
    layer0_outputs(9798) <= inputs(198);
    layer0_outputs(9799) <= inputs(231);
    layer0_outputs(9800) <= not((inputs(216)) xor (inputs(184)));
    layer0_outputs(9801) <= (inputs(209)) or (inputs(218));
    layer0_outputs(9802) <= not((inputs(192)) xor (inputs(13)));
    layer0_outputs(9803) <= not(inputs(216));
    layer0_outputs(9804) <= inputs(184);
    layer0_outputs(9805) <= not((inputs(33)) or (inputs(61)));
    layer0_outputs(9806) <= not(inputs(82));
    layer0_outputs(9807) <= not(inputs(48));
    layer0_outputs(9808) <= (inputs(53)) and not (inputs(224));
    layer0_outputs(9809) <= (inputs(147)) and not (inputs(206));
    layer0_outputs(9810) <= not(inputs(16)) or (inputs(185));
    layer0_outputs(9811) <= (inputs(125)) or (inputs(126));
    layer0_outputs(9812) <= not((inputs(143)) xor (inputs(165)));
    layer0_outputs(9813) <= (inputs(168)) or (inputs(147));
    layer0_outputs(9814) <= not(inputs(132));
    layer0_outputs(9815) <= inputs(30);
    layer0_outputs(9816) <= not((inputs(196)) xor (inputs(47)));
    layer0_outputs(9817) <= inputs(92);
    layer0_outputs(9818) <= not(inputs(155));
    layer0_outputs(9819) <= not(inputs(29)) or (inputs(82));
    layer0_outputs(9820) <= not((inputs(15)) or (inputs(83)));
    layer0_outputs(9821) <= (inputs(54)) or (inputs(92));
    layer0_outputs(9822) <= (inputs(52)) and not (inputs(141));
    layer0_outputs(9823) <= (inputs(228)) and not (inputs(104));
    layer0_outputs(9824) <= not(inputs(96)) or (inputs(112));
    layer0_outputs(9825) <= not((inputs(171)) or (inputs(222)));
    layer0_outputs(9826) <= not((inputs(41)) or (inputs(199)));
    layer0_outputs(9827) <= inputs(62);
    layer0_outputs(9828) <= not((inputs(197)) or (inputs(176)));
    layer0_outputs(9829) <= (inputs(240)) or (inputs(77));
    layer0_outputs(9830) <= (inputs(47)) or (inputs(99));
    layer0_outputs(9831) <= (inputs(72)) and (inputs(9));
    layer0_outputs(9832) <= not((inputs(175)) or (inputs(140)));
    layer0_outputs(9833) <= inputs(20);
    layer0_outputs(9834) <= not(inputs(139));
    layer0_outputs(9835) <= inputs(104);
    layer0_outputs(9836) <= not(inputs(94));
    layer0_outputs(9837) <= not(inputs(183));
    layer0_outputs(9838) <= '0';
    layer0_outputs(9839) <= inputs(86);
    layer0_outputs(9840) <= not(inputs(214)) or (inputs(46));
    layer0_outputs(9841) <= inputs(103);
    layer0_outputs(9842) <= not(inputs(181));
    layer0_outputs(9843) <= not((inputs(147)) or (inputs(186)));
    layer0_outputs(9844) <= (inputs(200)) and not (inputs(62));
    layer0_outputs(9845) <= not(inputs(231)) or (inputs(156));
    layer0_outputs(9846) <= not(inputs(249));
    layer0_outputs(9847) <= not(inputs(57));
    layer0_outputs(9848) <= not(inputs(230));
    layer0_outputs(9849) <= not((inputs(58)) xor (inputs(217)));
    layer0_outputs(9850) <= (inputs(24)) or (inputs(163));
    layer0_outputs(9851) <= (inputs(168)) xor (inputs(99));
    layer0_outputs(9852) <= inputs(88);
    layer0_outputs(9853) <= (inputs(167)) xor (inputs(134));
    layer0_outputs(9854) <= (inputs(250)) xor (inputs(51));
    layer0_outputs(9855) <= (inputs(134)) and not (inputs(115));
    layer0_outputs(9856) <= not((inputs(47)) or (inputs(155)));
    layer0_outputs(9857) <= (inputs(25)) or (inputs(35));
    layer0_outputs(9858) <= not((inputs(38)) or (inputs(92)));
    layer0_outputs(9859) <= (inputs(223)) or (inputs(96));
    layer0_outputs(9860) <= (inputs(215)) and (inputs(41));
    layer0_outputs(9861) <= not((inputs(102)) and (inputs(103)));
    layer0_outputs(9862) <= (inputs(117)) and not (inputs(39));
    layer0_outputs(9863) <= (inputs(213)) or (inputs(199));
    layer0_outputs(9864) <= inputs(9);
    layer0_outputs(9865) <= not(inputs(91)) or (inputs(23));
    layer0_outputs(9866) <= inputs(84);
    layer0_outputs(9867) <= (inputs(8)) and not (inputs(114));
    layer0_outputs(9868) <= (inputs(108)) xor (inputs(116));
    layer0_outputs(9869) <= not(inputs(105)) or (inputs(240));
    layer0_outputs(9870) <= inputs(248);
    layer0_outputs(9871) <= not(inputs(22));
    layer0_outputs(9872) <= inputs(216);
    layer0_outputs(9873) <= inputs(114);
    layer0_outputs(9874) <= (inputs(25)) or (inputs(97));
    layer0_outputs(9875) <= inputs(144);
    layer0_outputs(9876) <= (inputs(235)) xor (inputs(179));
    layer0_outputs(9877) <= (inputs(106)) or (inputs(12));
    layer0_outputs(9878) <= not(inputs(159)) or (inputs(48));
    layer0_outputs(9879) <= not(inputs(120));
    layer0_outputs(9880) <= not((inputs(56)) xor (inputs(101)));
    layer0_outputs(9881) <= not(inputs(72)) or (inputs(195));
    layer0_outputs(9882) <= not(inputs(178));
    layer0_outputs(9883) <= (inputs(19)) and not (inputs(136));
    layer0_outputs(9884) <= (inputs(118)) xor (inputs(116));
    layer0_outputs(9885) <= not((inputs(2)) xor (inputs(227)));
    layer0_outputs(9886) <= not(inputs(188)) or (inputs(97));
    layer0_outputs(9887) <= (inputs(132)) xor (inputs(21));
    layer0_outputs(9888) <= not(inputs(70)) or (inputs(0));
    layer0_outputs(9889) <= not(inputs(148));
    layer0_outputs(9890) <= not(inputs(68)) or (inputs(1));
    layer0_outputs(9891) <= '1';
    layer0_outputs(9892) <= not((inputs(128)) xor (inputs(226)));
    layer0_outputs(9893) <= inputs(213);
    layer0_outputs(9894) <= not((inputs(100)) xor (inputs(85)));
    layer0_outputs(9895) <= inputs(35);
    layer0_outputs(9896) <= not(inputs(26)) or (inputs(224));
    layer0_outputs(9897) <= not(inputs(28)) or (inputs(241));
    layer0_outputs(9898) <= not(inputs(24));
    layer0_outputs(9899) <= (inputs(48)) or (inputs(167));
    layer0_outputs(9900) <= not(inputs(82));
    layer0_outputs(9901) <= not(inputs(123));
    layer0_outputs(9902) <= not((inputs(49)) or (inputs(2)));
    layer0_outputs(9903) <= inputs(60);
    layer0_outputs(9904) <= (inputs(42)) and not (inputs(33));
    layer0_outputs(9905) <= (inputs(241)) or (inputs(124));
    layer0_outputs(9906) <= not(inputs(39));
    layer0_outputs(9907) <= inputs(111);
    layer0_outputs(9908) <= not((inputs(114)) xor (inputs(104)));
    layer0_outputs(9909) <= (inputs(198)) xor (inputs(185));
    layer0_outputs(9910) <= not((inputs(57)) or (inputs(127)));
    layer0_outputs(9911) <= not((inputs(242)) xor (inputs(254)));
    layer0_outputs(9912) <= inputs(189);
    layer0_outputs(9913) <= inputs(227);
    layer0_outputs(9914) <= '1';
    layer0_outputs(9915) <= not(inputs(240)) or (inputs(132));
    layer0_outputs(9916) <= inputs(229);
    layer0_outputs(9917) <= (inputs(224)) xor (inputs(247));
    layer0_outputs(9918) <= (inputs(31)) xor (inputs(145));
    layer0_outputs(9919) <= not(inputs(84));
    layer0_outputs(9920) <= not(inputs(93));
    layer0_outputs(9921) <= inputs(128);
    layer0_outputs(9922) <= not((inputs(121)) or (inputs(103)));
    layer0_outputs(9923) <= (inputs(107)) and not (inputs(227));
    layer0_outputs(9924) <= (inputs(27)) xor (inputs(131));
    layer0_outputs(9925) <= not(inputs(171));
    layer0_outputs(9926) <= (inputs(157)) and not (inputs(65));
    layer0_outputs(9927) <= (inputs(129)) or (inputs(189));
    layer0_outputs(9928) <= (inputs(155)) or (inputs(63));
    layer0_outputs(9929) <= '1';
    layer0_outputs(9930) <= not(inputs(205)) or (inputs(6));
    layer0_outputs(9931) <= not((inputs(119)) and (inputs(246)));
    layer0_outputs(9932) <= (inputs(216)) and not (inputs(94));
    layer0_outputs(9933) <= not(inputs(78));
    layer0_outputs(9934) <= not(inputs(19));
    layer0_outputs(9935) <= (inputs(29)) or (inputs(109));
    layer0_outputs(9936) <= inputs(214);
    layer0_outputs(9937) <= not(inputs(105)) or (inputs(203));
    layer0_outputs(9938) <= inputs(142);
    layer0_outputs(9939) <= not(inputs(116)) or (inputs(61));
    layer0_outputs(9940) <= (inputs(153)) or (inputs(163));
    layer0_outputs(9941) <= (inputs(122)) and (inputs(5));
    layer0_outputs(9942) <= (inputs(105)) xor (inputs(1));
    layer0_outputs(9943) <= not(inputs(243)) or (inputs(131));
    layer0_outputs(9944) <= (inputs(250)) or (inputs(191));
    layer0_outputs(9945) <= (inputs(54)) and not (inputs(162));
    layer0_outputs(9946) <= not((inputs(184)) or (inputs(226)));
    layer0_outputs(9947) <= not(inputs(95));
    layer0_outputs(9948) <= not(inputs(188));
    layer0_outputs(9949) <= not((inputs(53)) and (inputs(242)));
    layer0_outputs(9950) <= '1';
    layer0_outputs(9951) <= (inputs(194)) xor (inputs(236));
    layer0_outputs(9952) <= (inputs(127)) xor (inputs(141));
    layer0_outputs(9953) <= (inputs(62)) xor (inputs(74));
    layer0_outputs(9954) <= not((inputs(240)) or (inputs(193)));
    layer0_outputs(9955) <= (inputs(15)) or (inputs(83));
    layer0_outputs(9956) <= not((inputs(108)) or (inputs(21)));
    layer0_outputs(9957) <= inputs(128);
    layer0_outputs(9958) <= (inputs(195)) xor (inputs(162));
    layer0_outputs(9959) <= (inputs(24)) xor (inputs(27));
    layer0_outputs(9960) <= not(inputs(219)) or (inputs(87));
    layer0_outputs(9961) <= (inputs(199)) and not (inputs(78));
    layer0_outputs(9962) <= not(inputs(20)) or (inputs(206));
    layer0_outputs(9963) <= not(inputs(56));
    layer0_outputs(9964) <= (inputs(23)) or (inputs(56));
    layer0_outputs(9965) <= (inputs(109)) xor (inputs(177));
    layer0_outputs(9966) <= not(inputs(102)) or (inputs(140));
    layer0_outputs(9967) <= not((inputs(98)) or (inputs(115)));
    layer0_outputs(9968) <= (inputs(228)) and not (inputs(88));
    layer0_outputs(9969) <= (inputs(177)) or (inputs(145));
    layer0_outputs(9970) <= (inputs(173)) and not (inputs(60));
    layer0_outputs(9971) <= not(inputs(114));
    layer0_outputs(9972) <= (inputs(229)) and not (inputs(54));
    layer0_outputs(9973) <= inputs(100);
    layer0_outputs(9974) <= not(inputs(102));
    layer0_outputs(9975) <= (inputs(83)) or (inputs(171));
    layer0_outputs(9976) <= (inputs(115)) and not (inputs(17));
    layer0_outputs(9977) <= not((inputs(132)) xor (inputs(86)));
    layer0_outputs(9978) <= not(inputs(241));
    layer0_outputs(9979) <= not(inputs(52)) or (inputs(179));
    layer0_outputs(9980) <= (inputs(54)) and not (inputs(108));
    layer0_outputs(9981) <= (inputs(178)) and (inputs(109));
    layer0_outputs(9982) <= (inputs(185)) and not (inputs(17));
    layer0_outputs(9983) <= inputs(215);
    layer0_outputs(9984) <= (inputs(16)) or (inputs(94));
    layer0_outputs(9985) <= not((inputs(49)) xor (inputs(206)));
    layer0_outputs(9986) <= not(inputs(84));
    layer0_outputs(9987) <= inputs(82);
    layer0_outputs(9988) <= (inputs(198)) and (inputs(198));
    layer0_outputs(9989) <= not(inputs(217));
    layer0_outputs(9990) <= inputs(201);
    layer0_outputs(9991) <= not(inputs(68));
    layer0_outputs(9992) <= inputs(227);
    layer0_outputs(9993) <= not((inputs(247)) or (inputs(208)));
    layer0_outputs(9994) <= not(inputs(235)) or (inputs(93));
    layer0_outputs(9995) <= (inputs(187)) or (inputs(208));
    layer0_outputs(9996) <= not(inputs(172)) or (inputs(207));
    layer0_outputs(9997) <= '0';
    layer0_outputs(9998) <= (inputs(95)) and not (inputs(243));
    layer0_outputs(9999) <= not(inputs(6)) or (inputs(29));
    layer0_outputs(10000) <= not(inputs(241)) or (inputs(130));
    layer0_outputs(10001) <= not(inputs(138)) or (inputs(221));
    layer0_outputs(10002) <= not(inputs(225));
    layer0_outputs(10003) <= not(inputs(89)) or (inputs(126));
    layer0_outputs(10004) <= inputs(235);
    layer0_outputs(10005) <= inputs(166);
    layer0_outputs(10006) <= not((inputs(96)) or (inputs(146)));
    layer0_outputs(10007) <= not((inputs(189)) and (inputs(144)));
    layer0_outputs(10008) <= inputs(195);
    layer0_outputs(10009) <= not(inputs(231));
    layer0_outputs(10010) <= not(inputs(218)) or (inputs(46));
    layer0_outputs(10011) <= inputs(47);
    layer0_outputs(10012) <= not((inputs(195)) xor (inputs(79)));
    layer0_outputs(10013) <= inputs(71);
    layer0_outputs(10014) <= not((inputs(178)) xor (inputs(92)));
    layer0_outputs(10015) <= (inputs(58)) and not (inputs(166));
    layer0_outputs(10016) <= not((inputs(194)) xor (inputs(80)));
    layer0_outputs(10017) <= not((inputs(205)) or (inputs(246)));
    layer0_outputs(10018) <= inputs(117);
    layer0_outputs(10019) <= not(inputs(36));
    layer0_outputs(10020) <= not(inputs(117));
    layer0_outputs(10021) <= not(inputs(115)) or (inputs(214));
    layer0_outputs(10022) <= (inputs(191)) xor (inputs(17));
    layer0_outputs(10023) <= (inputs(80)) or (inputs(179));
    layer0_outputs(10024) <= inputs(129);
    layer0_outputs(10025) <= not((inputs(202)) or (inputs(159)));
    layer0_outputs(10026) <= not(inputs(234));
    layer0_outputs(10027) <= inputs(167);
    layer0_outputs(10028) <= not((inputs(240)) or (inputs(223)));
    layer0_outputs(10029) <= (inputs(135)) and not (inputs(143));
    layer0_outputs(10030) <= not((inputs(11)) or (inputs(112)));
    layer0_outputs(10031) <= inputs(210);
    layer0_outputs(10032) <= not(inputs(119));
    layer0_outputs(10033) <= not((inputs(249)) or (inputs(216)));
    layer0_outputs(10034) <= not((inputs(49)) or (inputs(54)));
    layer0_outputs(10035) <= (inputs(38)) and (inputs(17));
    layer0_outputs(10036) <= inputs(198);
    layer0_outputs(10037) <= not(inputs(123));
    layer0_outputs(10038) <= not((inputs(210)) xor (inputs(222)));
    layer0_outputs(10039) <= not(inputs(205)) or (inputs(111));
    layer0_outputs(10040) <= inputs(180);
    layer0_outputs(10041) <= (inputs(81)) and (inputs(251));
    layer0_outputs(10042) <= not(inputs(241));
    layer0_outputs(10043) <= not(inputs(182)) or (inputs(28));
    layer0_outputs(10044) <= inputs(161);
    layer0_outputs(10045) <= not(inputs(196));
    layer0_outputs(10046) <= (inputs(80)) or (inputs(159));
    layer0_outputs(10047) <= inputs(8);
    layer0_outputs(10048) <= inputs(231);
    layer0_outputs(10049) <= inputs(22);
    layer0_outputs(10050) <= inputs(153);
    layer0_outputs(10051) <= inputs(250);
    layer0_outputs(10052) <= not((inputs(176)) and (inputs(178)));
    layer0_outputs(10053) <= not((inputs(16)) or (inputs(73)));
    layer0_outputs(10054) <= not((inputs(169)) xor (inputs(172)));
    layer0_outputs(10055) <= not(inputs(148));
    layer0_outputs(10056) <= not(inputs(181)) or (inputs(34));
    layer0_outputs(10057) <= not(inputs(203));
    layer0_outputs(10058) <= inputs(187);
    layer0_outputs(10059) <= inputs(7);
    layer0_outputs(10060) <= not((inputs(204)) and (inputs(134)));
    layer0_outputs(10061) <= inputs(212);
    layer0_outputs(10062) <= inputs(239);
    layer0_outputs(10063) <= (inputs(53)) and not (inputs(231));
    layer0_outputs(10064) <= not(inputs(87));
    layer0_outputs(10065) <= not((inputs(165)) or (inputs(224)));
    layer0_outputs(10066) <= not(inputs(168)) or (inputs(189));
    layer0_outputs(10067) <= (inputs(3)) xor (inputs(95));
    layer0_outputs(10068) <= inputs(49);
    layer0_outputs(10069) <= not(inputs(177));
    layer0_outputs(10070) <= (inputs(41)) or (inputs(136));
    layer0_outputs(10071) <= (inputs(149)) and not (inputs(236));
    layer0_outputs(10072) <= not((inputs(94)) xor (inputs(12)));
    layer0_outputs(10073) <= (inputs(235)) and not (inputs(238));
    layer0_outputs(10074) <= inputs(130);
    layer0_outputs(10075) <= not(inputs(104));
    layer0_outputs(10076) <= not((inputs(108)) xor (inputs(36)));
    layer0_outputs(10077) <= not(inputs(249)) or (inputs(136));
    layer0_outputs(10078) <= not(inputs(114));
    layer0_outputs(10079) <= not(inputs(196));
    layer0_outputs(10080) <= inputs(253);
    layer0_outputs(10081) <= (inputs(142)) xor (inputs(246));
    layer0_outputs(10082) <= (inputs(129)) xor (inputs(151));
    layer0_outputs(10083) <= (inputs(189)) or (inputs(221));
    layer0_outputs(10084) <= not(inputs(57)) or (inputs(206));
    layer0_outputs(10085) <= (inputs(38)) and not (inputs(114));
    layer0_outputs(10086) <= (inputs(55)) xor (inputs(85));
    layer0_outputs(10087) <= not(inputs(122)) or (inputs(225));
    layer0_outputs(10088) <= not(inputs(154)) or (inputs(112));
    layer0_outputs(10089) <= inputs(7);
    layer0_outputs(10090) <= (inputs(217)) and not (inputs(162));
    layer0_outputs(10091) <= (inputs(132)) xor (inputs(140));
    layer0_outputs(10092) <= not((inputs(128)) xor (inputs(172)));
    layer0_outputs(10093) <= inputs(233);
    layer0_outputs(10094) <= (inputs(63)) or (inputs(87));
    layer0_outputs(10095) <= (inputs(176)) xor (inputs(214));
    layer0_outputs(10096) <= (inputs(97)) xor (inputs(71));
    layer0_outputs(10097) <= not(inputs(75)) or (inputs(252));
    layer0_outputs(10098) <= (inputs(107)) xor (inputs(143));
    layer0_outputs(10099) <= not(inputs(159)) or (inputs(82));
    layer0_outputs(10100) <= not(inputs(192)) or (inputs(29));
    layer0_outputs(10101) <= inputs(3);
    layer0_outputs(10102) <= not((inputs(181)) or (inputs(11)));
    layer0_outputs(10103) <= not(inputs(231));
    layer0_outputs(10104) <= inputs(134);
    layer0_outputs(10105) <= not(inputs(139));
    layer0_outputs(10106) <= not((inputs(87)) or (inputs(202)));
    layer0_outputs(10107) <= (inputs(252)) or (inputs(185));
    layer0_outputs(10108) <= not((inputs(116)) xor (inputs(35)));
    layer0_outputs(10109) <= not(inputs(43));
    layer0_outputs(10110) <= inputs(127);
    layer0_outputs(10111) <= inputs(166);
    layer0_outputs(10112) <= not(inputs(104)) or (inputs(202));
    layer0_outputs(10113) <= not((inputs(222)) or (inputs(163)));
    layer0_outputs(10114) <= (inputs(245)) or (inputs(38));
    layer0_outputs(10115) <= not(inputs(89)) or (inputs(242));
    layer0_outputs(10116) <= not((inputs(20)) xor (inputs(33)));
    layer0_outputs(10117) <= (inputs(107)) and (inputs(27));
    layer0_outputs(10118) <= not((inputs(160)) or (inputs(23)));
    layer0_outputs(10119) <= not(inputs(95));
    layer0_outputs(10120) <= not(inputs(209));
    layer0_outputs(10121) <= not((inputs(193)) xor (inputs(83)));
    layer0_outputs(10122) <= not((inputs(244)) or (inputs(101)));
    layer0_outputs(10123) <= (inputs(58)) and not (inputs(13));
    layer0_outputs(10124) <= not(inputs(101)) or (inputs(2));
    layer0_outputs(10125) <= not(inputs(185)) or (inputs(1));
    layer0_outputs(10126) <= not(inputs(126));
    layer0_outputs(10127) <= not((inputs(165)) and (inputs(197)));
    layer0_outputs(10128) <= inputs(8);
    layer0_outputs(10129) <= not((inputs(71)) and (inputs(46)));
    layer0_outputs(10130) <= not((inputs(28)) xor (inputs(45)));
    layer0_outputs(10131) <= not(inputs(127)) or (inputs(142));
    layer0_outputs(10132) <= (inputs(252)) xor (inputs(60));
    layer0_outputs(10133) <= (inputs(60)) or (inputs(162));
    layer0_outputs(10134) <= inputs(105);
    layer0_outputs(10135) <= (inputs(79)) or (inputs(53));
    layer0_outputs(10136) <= (inputs(65)) and (inputs(100));
    layer0_outputs(10137) <= not((inputs(71)) and (inputs(198)));
    layer0_outputs(10138) <= not(inputs(19));
    layer0_outputs(10139) <= not((inputs(184)) xor (inputs(231)));
    layer0_outputs(10140) <= not((inputs(88)) xor (inputs(130)));
    layer0_outputs(10141) <= not(inputs(22));
    layer0_outputs(10142) <= not((inputs(162)) xor (inputs(192)));
    layer0_outputs(10143) <= not(inputs(215));
    layer0_outputs(10144) <= not(inputs(139));
    layer0_outputs(10145) <= not(inputs(59));
    layer0_outputs(10146) <= not(inputs(103));
    layer0_outputs(10147) <= '1';
    layer0_outputs(10148) <= (inputs(123)) and not (inputs(208));
    layer0_outputs(10149) <= inputs(137);
    layer0_outputs(10150) <= (inputs(89)) and (inputs(66));
    layer0_outputs(10151) <= (inputs(178)) or (inputs(36));
    layer0_outputs(10152) <= not(inputs(115));
    layer0_outputs(10153) <= (inputs(87)) xor (inputs(130));
    layer0_outputs(10154) <= (inputs(201)) and not (inputs(127));
    layer0_outputs(10155) <= (inputs(151)) or (inputs(245));
    layer0_outputs(10156) <= inputs(200);
    layer0_outputs(10157) <= not((inputs(58)) xor (inputs(39)));
    layer0_outputs(10158) <= not(inputs(148)) or (inputs(96));
    layer0_outputs(10159) <= inputs(140);
    layer0_outputs(10160) <= not(inputs(55));
    layer0_outputs(10161) <= (inputs(90)) xor (inputs(137));
    layer0_outputs(10162) <= inputs(22);
    layer0_outputs(10163) <= (inputs(84)) xor (inputs(55));
    layer0_outputs(10164) <= not(inputs(1)) or (inputs(4));
    layer0_outputs(10165) <= (inputs(28)) and not (inputs(146));
    layer0_outputs(10166) <= (inputs(128)) or (inputs(148));
    layer0_outputs(10167) <= inputs(7);
    layer0_outputs(10168) <= inputs(199);
    layer0_outputs(10169) <= (inputs(238)) and not (inputs(235));
    layer0_outputs(10170) <= (inputs(237)) or (inputs(248));
    layer0_outputs(10171) <= not(inputs(163));
    layer0_outputs(10172) <= (inputs(146)) or (inputs(255));
    layer0_outputs(10173) <= '1';
    layer0_outputs(10174) <= not(inputs(25));
    layer0_outputs(10175) <= not(inputs(84));
    layer0_outputs(10176) <= not((inputs(221)) or (inputs(169)));
    layer0_outputs(10177) <= (inputs(98)) and not (inputs(225));
    layer0_outputs(10178) <= inputs(41);
    layer0_outputs(10179) <= inputs(114);
    layer0_outputs(10180) <= inputs(239);
    layer0_outputs(10181) <= not((inputs(209)) xor (inputs(159)));
    layer0_outputs(10182) <= '1';
    layer0_outputs(10183) <= not((inputs(142)) or (inputs(218)));
    layer0_outputs(10184) <= not(inputs(249));
    layer0_outputs(10185) <= (inputs(92)) xor (inputs(3));
    layer0_outputs(10186) <= (inputs(100)) or (inputs(202));
    layer0_outputs(10187) <= (inputs(15)) xor (inputs(95));
    layer0_outputs(10188) <= (inputs(100)) and not (inputs(1));
    layer0_outputs(10189) <= (inputs(17)) or (inputs(241));
    layer0_outputs(10190) <= (inputs(229)) or (inputs(191));
    layer0_outputs(10191) <= (inputs(246)) or (inputs(31));
    layer0_outputs(10192) <= not(inputs(125)) or (inputs(32));
    layer0_outputs(10193) <= not((inputs(62)) or (inputs(156)));
    layer0_outputs(10194) <= not(inputs(8)) or (inputs(83));
    layer0_outputs(10195) <= inputs(133);
    layer0_outputs(10196) <= not(inputs(88)) or (inputs(110));
    layer0_outputs(10197) <= not(inputs(104));
    layer0_outputs(10198) <= (inputs(157)) or (inputs(206));
    layer0_outputs(10199) <= not(inputs(165));
    layer0_outputs(10200) <= (inputs(97)) xor (inputs(5));
    layer0_outputs(10201) <= not(inputs(243)) or (inputs(128));
    layer0_outputs(10202) <= not(inputs(59));
    layer0_outputs(10203) <= (inputs(221)) or (inputs(219));
    layer0_outputs(10204) <= not(inputs(222));
    layer0_outputs(10205) <= not(inputs(89)) or (inputs(204));
    layer0_outputs(10206) <= not((inputs(79)) or (inputs(95)));
    layer0_outputs(10207) <= inputs(116);
    layer0_outputs(10208) <= not((inputs(166)) or (inputs(141)));
    layer0_outputs(10209) <= not(inputs(30));
    layer0_outputs(10210) <= inputs(37);
    layer0_outputs(10211) <= inputs(232);
    layer0_outputs(10212) <= not(inputs(56)) or (inputs(15));
    layer0_outputs(10213) <= not((inputs(197)) and (inputs(209)));
    layer0_outputs(10214) <= inputs(177);
    layer0_outputs(10215) <= not((inputs(84)) xor (inputs(158)));
    layer0_outputs(10216) <= not(inputs(170)) or (inputs(204));
    layer0_outputs(10217) <= inputs(195);
    layer0_outputs(10218) <= inputs(40);
    layer0_outputs(10219) <= not((inputs(72)) xor (inputs(115)));
    layer0_outputs(10220) <= inputs(58);
    layer0_outputs(10221) <= (inputs(229)) xor (inputs(149));
    layer0_outputs(10222) <= not(inputs(116)) or (inputs(10));
    layer0_outputs(10223) <= not((inputs(79)) and (inputs(255)));
    layer0_outputs(10224) <= (inputs(77)) and not (inputs(243));
    layer0_outputs(10225) <= (inputs(179)) or (inputs(196));
    layer0_outputs(10226) <= (inputs(193)) or (inputs(186));
    layer0_outputs(10227) <= (inputs(116)) xor (inputs(146));
    layer0_outputs(10228) <= not((inputs(35)) xor (inputs(37)));
    layer0_outputs(10229) <= (inputs(151)) xor (inputs(132));
    layer0_outputs(10230) <= (inputs(57)) and not (inputs(39));
    layer0_outputs(10231) <= (inputs(119)) and not (inputs(191));
    layer0_outputs(10232) <= not((inputs(15)) xor (inputs(83)));
    layer0_outputs(10233) <= not(inputs(233));
    layer0_outputs(10234) <= (inputs(219)) and (inputs(173));
    layer0_outputs(10235) <= not((inputs(169)) or (inputs(11)));
    layer0_outputs(10236) <= (inputs(29)) xor (inputs(74));
    layer0_outputs(10237) <= not((inputs(252)) or (inputs(85)));
    layer0_outputs(10238) <= inputs(158);
    layer0_outputs(10239) <= inputs(65);
    outputs(0) <= not((layer0_outputs(8250)) xor (layer0_outputs(6404)));
    outputs(1) <= layer0_outputs(4407);
    outputs(2) <= (layer0_outputs(5885)) and not (layer0_outputs(5011));
    outputs(3) <= (layer0_outputs(4910)) and not (layer0_outputs(3786));
    outputs(4) <= (layer0_outputs(1383)) and not (layer0_outputs(7592));
    outputs(5) <= not((layer0_outputs(2992)) xor (layer0_outputs(9170)));
    outputs(6) <= (layer0_outputs(660)) or (layer0_outputs(7491));
    outputs(7) <= layer0_outputs(5218);
    outputs(8) <= (layer0_outputs(7369)) or (layer0_outputs(888));
    outputs(9) <= (layer0_outputs(130)) and not (layer0_outputs(5134));
    outputs(10) <= (layer0_outputs(286)) and not (layer0_outputs(8272));
    outputs(11) <= (layer0_outputs(8365)) and not (layer0_outputs(7020));
    outputs(12) <= (layer0_outputs(2245)) and not (layer0_outputs(7783));
    outputs(13) <= layer0_outputs(5568);
    outputs(14) <= (layer0_outputs(7765)) and (layer0_outputs(184));
    outputs(15) <= (layer0_outputs(8221)) and not (layer0_outputs(487));
    outputs(16) <= not(layer0_outputs(5388));
    outputs(17) <= layer0_outputs(4383);
    outputs(18) <= not((layer0_outputs(8483)) xor (layer0_outputs(547)));
    outputs(19) <= not(layer0_outputs(7612)) or (layer0_outputs(8028));
    outputs(20) <= (layer0_outputs(4520)) xor (layer0_outputs(3145));
    outputs(21) <= layer0_outputs(4239);
    outputs(22) <= not(layer0_outputs(4557));
    outputs(23) <= not(layer0_outputs(3071));
    outputs(24) <= (layer0_outputs(8770)) and (layer0_outputs(2599));
    outputs(25) <= not(layer0_outputs(9717));
    outputs(26) <= layer0_outputs(8336);
    outputs(27) <= not(layer0_outputs(9574));
    outputs(28) <= not(layer0_outputs(5576));
    outputs(29) <= not((layer0_outputs(1466)) xor (layer0_outputs(7389)));
    outputs(30) <= not(layer0_outputs(10012)) or (layer0_outputs(9209));
    outputs(31) <= (layer0_outputs(7233)) and not (layer0_outputs(2635));
    outputs(32) <= (layer0_outputs(5120)) and (layer0_outputs(1014));
    outputs(33) <= (layer0_outputs(10032)) and (layer0_outputs(9459));
    outputs(34) <= (layer0_outputs(5655)) xor (layer0_outputs(2040));
    outputs(35) <= not((layer0_outputs(1976)) or (layer0_outputs(9110)));
    outputs(36) <= layer0_outputs(3647);
    outputs(37) <= (layer0_outputs(7555)) xor (layer0_outputs(4998));
    outputs(38) <= not(layer0_outputs(3406));
    outputs(39) <= (layer0_outputs(9556)) and (layer0_outputs(3620));
    outputs(40) <= layer0_outputs(8961);
    outputs(41) <= (layer0_outputs(7005)) xor (layer0_outputs(4620));
    outputs(42) <= not(layer0_outputs(2764));
    outputs(43) <= not(layer0_outputs(2453)) or (layer0_outputs(2337));
    outputs(44) <= layer0_outputs(3255);
    outputs(45) <= layer0_outputs(1873);
    outputs(46) <= not(layer0_outputs(2236));
    outputs(47) <= not(layer0_outputs(3277));
    outputs(48) <= layer0_outputs(47);
    outputs(49) <= (layer0_outputs(10026)) xor (layer0_outputs(275));
    outputs(50) <= not(layer0_outputs(8792));
    outputs(51) <= (layer0_outputs(5902)) xor (layer0_outputs(76));
    outputs(52) <= (layer0_outputs(4043)) or (layer0_outputs(6752));
    outputs(53) <= layer0_outputs(1949);
    outputs(54) <= not(layer0_outputs(8326));
    outputs(55) <= not(layer0_outputs(6982));
    outputs(56) <= layer0_outputs(4220);
    outputs(57) <= (layer0_outputs(1388)) and (layer0_outputs(5160));
    outputs(58) <= layer0_outputs(4132);
    outputs(59) <= not(layer0_outputs(9360));
    outputs(60) <= not((layer0_outputs(8040)) or (layer0_outputs(7791)));
    outputs(61) <= layer0_outputs(1815);
    outputs(62) <= layer0_outputs(5430);
    outputs(63) <= (layer0_outputs(5339)) or (layer0_outputs(3967));
    outputs(64) <= not(layer0_outputs(1603));
    outputs(65) <= layer0_outputs(3078);
    outputs(66) <= not(layer0_outputs(8900));
    outputs(67) <= layer0_outputs(3427);
    outputs(68) <= not((layer0_outputs(3424)) xor (layer0_outputs(1840)));
    outputs(69) <= layer0_outputs(3701);
    outputs(70) <= (layer0_outputs(9487)) and (layer0_outputs(4471));
    outputs(71) <= (layer0_outputs(8814)) xor (layer0_outputs(8818));
    outputs(72) <= (layer0_outputs(10116)) and not (layer0_outputs(7999));
    outputs(73) <= not(layer0_outputs(5188));
    outputs(74) <= layer0_outputs(2685);
    outputs(75) <= layer0_outputs(8335);
    outputs(76) <= (layer0_outputs(1610)) or (layer0_outputs(5297));
    outputs(77) <= not(layer0_outputs(3302));
    outputs(78) <= not(layer0_outputs(2716));
    outputs(79) <= (layer0_outputs(5095)) and not (layer0_outputs(2603));
    outputs(80) <= not(layer0_outputs(5648));
    outputs(81) <= not(layer0_outputs(4927)) or (layer0_outputs(6248));
    outputs(82) <= layer0_outputs(7565);
    outputs(83) <= not(layer0_outputs(7394)) or (layer0_outputs(277));
    outputs(84) <= not(layer0_outputs(139));
    outputs(85) <= (layer0_outputs(9221)) xor (layer0_outputs(3915));
    outputs(86) <= not((layer0_outputs(8443)) and (layer0_outputs(465)));
    outputs(87) <= not(layer0_outputs(2153));
    outputs(88) <= layer0_outputs(6581);
    outputs(89) <= not(layer0_outputs(4814)) or (layer0_outputs(7298));
    outputs(90) <= not((layer0_outputs(5613)) xor (layer0_outputs(3103)));
    outputs(91) <= layer0_outputs(2423);
    outputs(92) <= (layer0_outputs(4607)) and not (layer0_outputs(2795));
    outputs(93) <= not(layer0_outputs(977)) or (layer0_outputs(1154));
    outputs(94) <= not((layer0_outputs(8239)) or (layer0_outputs(2075)));
    outputs(95) <= (layer0_outputs(6251)) and not (layer0_outputs(3594));
    outputs(96) <= not(layer0_outputs(3637));
    outputs(97) <= not(layer0_outputs(7172));
    outputs(98) <= layer0_outputs(6992);
    outputs(99) <= (layer0_outputs(10028)) and not (layer0_outputs(830));
    outputs(100) <= (layer0_outputs(667)) or (layer0_outputs(7460));
    outputs(101) <= not((layer0_outputs(5486)) and (layer0_outputs(5707)));
    outputs(102) <= not(layer0_outputs(8482));
    outputs(103) <= not((layer0_outputs(6618)) xor (layer0_outputs(2733)));
    outputs(104) <= not((layer0_outputs(4359)) xor (layer0_outputs(5166)));
    outputs(105) <= (layer0_outputs(5272)) or (layer0_outputs(6870));
    outputs(106) <= not(layer0_outputs(3236));
    outputs(107) <= (layer0_outputs(1195)) and not (layer0_outputs(1241));
    outputs(108) <= (layer0_outputs(9069)) xor (layer0_outputs(6127));
    outputs(109) <= (layer0_outputs(5012)) xor (layer0_outputs(7474));
    outputs(110) <= (layer0_outputs(6)) and not (layer0_outputs(8339));
    outputs(111) <= not(layer0_outputs(6684));
    outputs(112) <= (layer0_outputs(6077)) or (layer0_outputs(5198));
    outputs(113) <= not(layer0_outputs(9749));
    outputs(114) <= layer0_outputs(4148);
    outputs(115) <= (layer0_outputs(9482)) xor (layer0_outputs(4989));
    outputs(116) <= layer0_outputs(8120);
    outputs(117) <= not(layer0_outputs(9117));
    outputs(118) <= not(layer0_outputs(6723));
    outputs(119) <= (layer0_outputs(4199)) xor (layer0_outputs(5151));
    outputs(120) <= layer0_outputs(6533);
    outputs(121) <= (layer0_outputs(9609)) xor (layer0_outputs(9060));
    outputs(122) <= not(layer0_outputs(8467));
    outputs(123) <= not(layer0_outputs(6527));
    outputs(124) <= not(layer0_outputs(201)) or (layer0_outputs(3404));
    outputs(125) <= not(layer0_outputs(6179));
    outputs(126) <= not((layer0_outputs(718)) or (layer0_outputs(3204)));
    outputs(127) <= not(layer0_outputs(6407));
    outputs(128) <= layer0_outputs(1535);
    outputs(129) <= (layer0_outputs(5588)) and not (layer0_outputs(4453));
    outputs(130) <= (layer0_outputs(4681)) and not (layer0_outputs(8007));
    outputs(131) <= (layer0_outputs(8177)) or (layer0_outputs(1122));
    outputs(132) <= not((layer0_outputs(4774)) xor (layer0_outputs(2332)));
    outputs(133) <= (layer0_outputs(3)) xor (layer0_outputs(6576));
    outputs(134) <= (layer0_outputs(5113)) and (layer0_outputs(524));
    outputs(135) <= not((layer0_outputs(10137)) and (layer0_outputs(1057)));
    outputs(136) <= (layer0_outputs(3766)) xor (layer0_outputs(5515));
    outputs(137) <= (layer0_outputs(8808)) xor (layer0_outputs(8744));
    outputs(138) <= not(layer0_outputs(8920));
    outputs(139) <= layer0_outputs(9736);
    outputs(140) <= (layer0_outputs(7899)) xor (layer0_outputs(9291));
    outputs(141) <= (layer0_outputs(6895)) and not (layer0_outputs(9608));
    outputs(142) <= not((layer0_outputs(3019)) xor (layer0_outputs(6830)));
    outputs(143) <= not(layer0_outputs(4195));
    outputs(144) <= not(layer0_outputs(100));
    outputs(145) <= (layer0_outputs(8508)) and not (layer0_outputs(7827));
    outputs(146) <= (layer0_outputs(8849)) or (layer0_outputs(3870));
    outputs(147) <= not((layer0_outputs(2970)) and (layer0_outputs(9360)));
    outputs(148) <= not(layer0_outputs(8407));
    outputs(149) <= layer0_outputs(5829);
    outputs(150) <= (layer0_outputs(7778)) xor (layer0_outputs(1930));
    outputs(151) <= not(layer0_outputs(5636));
    outputs(152) <= (layer0_outputs(5292)) and not (layer0_outputs(4299));
    outputs(153) <= not((layer0_outputs(1346)) xor (layer0_outputs(7660)));
    outputs(154) <= not(layer0_outputs(5256)) or (layer0_outputs(3496));
    outputs(155) <= layer0_outputs(3286);
    outputs(156) <= not((layer0_outputs(9109)) xor (layer0_outputs(6728)));
    outputs(157) <= layer0_outputs(7408);
    outputs(158) <= not(layer0_outputs(8607)) or (layer0_outputs(7571));
    outputs(159) <= not((layer0_outputs(5889)) or (layer0_outputs(8367)));
    outputs(160) <= not((layer0_outputs(7455)) xor (layer0_outputs(3937)));
    outputs(161) <= layer0_outputs(2230);
    outputs(162) <= not(layer0_outputs(3570));
    outputs(163) <= (layer0_outputs(4033)) xor (layer0_outputs(964));
    outputs(164) <= not(layer0_outputs(637)) or (layer0_outputs(6014));
    outputs(165) <= layer0_outputs(2494);
    outputs(166) <= (layer0_outputs(658)) and not (layer0_outputs(7401));
    outputs(167) <= layer0_outputs(3384);
    outputs(168) <= not(layer0_outputs(2023));
    outputs(169) <= layer0_outputs(4403);
    outputs(170) <= layer0_outputs(8347);
    outputs(171) <= not((layer0_outputs(3387)) or (layer0_outputs(8246)));
    outputs(172) <= not(layer0_outputs(9297));
    outputs(173) <= layer0_outputs(8498);
    outputs(174) <= layer0_outputs(4932);
    outputs(175) <= not(layer0_outputs(1886));
    outputs(176) <= not(layer0_outputs(5867));
    outputs(177) <= not(layer0_outputs(10108));
    outputs(178) <= not((layer0_outputs(3907)) xor (layer0_outputs(8175)));
    outputs(179) <= not(layer0_outputs(6289));
    outputs(180) <= layer0_outputs(8357);
    outputs(181) <= not(layer0_outputs(1933)) or (layer0_outputs(5685));
    outputs(182) <= not(layer0_outputs(633));
    outputs(183) <= not(layer0_outputs(3962));
    outputs(184) <= (layer0_outputs(7005)) and not (layer0_outputs(5690));
    outputs(185) <= layer0_outputs(990);
    outputs(186) <= layer0_outputs(8492);
    outputs(187) <= not(layer0_outputs(6737));
    outputs(188) <= not((layer0_outputs(6415)) xor (layer0_outputs(9726)));
    outputs(189) <= not(layer0_outputs(148)) or (layer0_outputs(5719));
    outputs(190) <= not(layer0_outputs(5039));
    outputs(191) <= layer0_outputs(1773);
    outputs(192) <= (layer0_outputs(9159)) xor (layer0_outputs(8588));
    outputs(193) <= (layer0_outputs(5467)) and not (layer0_outputs(3096));
    outputs(194) <= not(layer0_outputs(5838));
    outputs(195) <= not((layer0_outputs(2715)) and (layer0_outputs(7461)));
    outputs(196) <= (layer0_outputs(5032)) and not (layer0_outputs(4719));
    outputs(197) <= (layer0_outputs(2604)) and (layer0_outputs(30));
    outputs(198) <= not((layer0_outputs(5411)) or (layer0_outputs(3781)));
    outputs(199) <= (layer0_outputs(4805)) xor (layer0_outputs(5939));
    outputs(200) <= (layer0_outputs(1100)) or (layer0_outputs(2306));
    outputs(201) <= not(layer0_outputs(1482));
    outputs(202) <= (layer0_outputs(9503)) and (layer0_outputs(7634));
    outputs(203) <= not((layer0_outputs(6657)) xor (layer0_outputs(9596)));
    outputs(204) <= not(layer0_outputs(2526)) or (layer0_outputs(9656));
    outputs(205) <= (layer0_outputs(9278)) xor (layer0_outputs(8308));
    outputs(206) <= (layer0_outputs(901)) xor (layer0_outputs(6913));
    outputs(207) <= layer0_outputs(1755);
    outputs(208) <= not(layer0_outputs(5648));
    outputs(209) <= (layer0_outputs(5047)) xor (layer0_outputs(995));
    outputs(210) <= not(layer0_outputs(8789));
    outputs(211) <= (layer0_outputs(4392)) and not (layer0_outputs(5324));
    outputs(212) <= (layer0_outputs(6589)) and not (layer0_outputs(4955));
    outputs(213) <= layer0_outputs(8163);
    outputs(214) <= not((layer0_outputs(1155)) xor (layer0_outputs(7155)));
    outputs(215) <= not((layer0_outputs(7174)) xor (layer0_outputs(7537)));
    outputs(216) <= (layer0_outputs(1103)) and (layer0_outputs(5286));
    outputs(217) <= layer0_outputs(9592);
    outputs(218) <= (layer0_outputs(3804)) xor (layer0_outputs(4715));
    outputs(219) <= (layer0_outputs(2468)) and not (layer0_outputs(4072));
    outputs(220) <= (layer0_outputs(73)) or (layer0_outputs(2385));
    outputs(221) <= layer0_outputs(3584);
    outputs(222) <= not((layer0_outputs(6871)) xor (layer0_outputs(269)));
    outputs(223) <= not(layer0_outputs(10063));
    outputs(224) <= not(layer0_outputs(9171));
    outputs(225) <= layer0_outputs(873);
    outputs(226) <= not(layer0_outputs(3609));
    outputs(227) <= (layer0_outputs(6993)) xor (layer0_outputs(3092));
    outputs(228) <= layer0_outputs(6245);
    outputs(229) <= (layer0_outputs(5232)) and not (layer0_outputs(8147));
    outputs(230) <= layer0_outputs(6652);
    outputs(231) <= (layer0_outputs(7451)) and not (layer0_outputs(2510));
    outputs(232) <= not(layer0_outputs(207)) or (layer0_outputs(9998));
    outputs(233) <= not(layer0_outputs(2508));
    outputs(234) <= layer0_outputs(5190);
    outputs(235) <= not(layer0_outputs(9337)) or (layer0_outputs(9952));
    outputs(236) <= layer0_outputs(3064);
    outputs(237) <= layer0_outputs(2728);
    outputs(238) <= not((layer0_outputs(1761)) and (layer0_outputs(6914)));
    outputs(239) <= not(layer0_outputs(2027));
    outputs(240) <= not(layer0_outputs(7589));
    outputs(241) <= not((layer0_outputs(5765)) xor (layer0_outputs(4500)));
    outputs(242) <= not(layer0_outputs(4297));
    outputs(243) <= layer0_outputs(2702);
    outputs(244) <= not(layer0_outputs(8985));
    outputs(245) <= layer0_outputs(2845);
    outputs(246) <= not((layer0_outputs(6832)) and (layer0_outputs(2149)));
    outputs(247) <= layer0_outputs(3670);
    outputs(248) <= not((layer0_outputs(8188)) xor (layer0_outputs(5159)));
    outputs(249) <= layer0_outputs(3775);
    outputs(250) <= not((layer0_outputs(6959)) xor (layer0_outputs(5381)));
    outputs(251) <= (layer0_outputs(3739)) and not (layer0_outputs(5059));
    outputs(252) <= (layer0_outputs(1807)) and not (layer0_outputs(4323));
    outputs(253) <= not(layer0_outputs(5216));
    outputs(254) <= not((layer0_outputs(8560)) or (layer0_outputs(5308)));
    outputs(255) <= not(layer0_outputs(4543)) or (layer0_outputs(5101));
    outputs(256) <= not(layer0_outputs(3239)) or (layer0_outputs(4208));
    outputs(257) <= not(layer0_outputs(5271));
    outputs(258) <= not(layer0_outputs(8138));
    outputs(259) <= layer0_outputs(9769);
    outputs(260) <= (layer0_outputs(7055)) and (layer0_outputs(1288));
    outputs(261) <= not(layer0_outputs(1798));
    outputs(262) <= not((layer0_outputs(1912)) or (layer0_outputs(1742)));
    outputs(263) <= layer0_outputs(3053);
    outputs(264) <= (layer0_outputs(5514)) and not (layer0_outputs(8942));
    outputs(265) <= (layer0_outputs(2503)) and not (layer0_outputs(3727));
    outputs(266) <= not(layer0_outputs(2670)) or (layer0_outputs(9981));
    outputs(267) <= not(layer0_outputs(3876)) or (layer0_outputs(3372));
    outputs(268) <= not((layer0_outputs(8640)) and (layer0_outputs(3715)));
    outputs(269) <= not(layer0_outputs(7886));
    outputs(270) <= not((layer0_outputs(927)) xor (layer0_outputs(7111)));
    outputs(271) <= not((layer0_outputs(7794)) and (layer0_outputs(9308)));
    outputs(272) <= (layer0_outputs(4644)) or (layer0_outputs(2504));
    outputs(273) <= (layer0_outputs(5222)) and (layer0_outputs(1703));
    outputs(274) <= layer0_outputs(8189);
    outputs(275) <= not((layer0_outputs(567)) xor (layer0_outputs(4650)));
    outputs(276) <= not((layer0_outputs(8348)) xor (layer0_outputs(2241)));
    outputs(277) <= layer0_outputs(9742);
    outputs(278) <= not(layer0_outputs(6954)) or (layer0_outputs(3792));
    outputs(279) <= not(layer0_outputs(1585));
    outputs(280) <= not(layer0_outputs(6020));
    outputs(281) <= not((layer0_outputs(5509)) xor (layer0_outputs(379)));
    outputs(282) <= not(layer0_outputs(6179)) or (layer0_outputs(7917));
    outputs(283) <= not(layer0_outputs(7717));
    outputs(284) <= (layer0_outputs(8763)) or (layer0_outputs(8893));
    outputs(285) <= not(layer0_outputs(2668));
    outputs(286) <= layer0_outputs(7296);
    outputs(287) <= (layer0_outputs(8172)) and (layer0_outputs(3007));
    outputs(288) <= (layer0_outputs(8363)) and not (layer0_outputs(2096));
    outputs(289) <= (layer0_outputs(860)) and not (layer0_outputs(7364));
    outputs(290) <= not(layer0_outputs(5240));
    outputs(291) <= (layer0_outputs(3728)) and not (layer0_outputs(3352));
    outputs(292) <= not((layer0_outputs(3413)) and (layer0_outputs(3187)));
    outputs(293) <= not((layer0_outputs(9628)) xor (layer0_outputs(9551)));
    outputs(294) <= not((layer0_outputs(10006)) xor (layer0_outputs(10195)));
    outputs(295) <= not(layer0_outputs(5798)) or (layer0_outputs(895));
    outputs(296) <= not(layer0_outputs(8574));
    outputs(297) <= (layer0_outputs(5842)) and not (layer0_outputs(1870));
    outputs(298) <= not(layer0_outputs(4386));
    outputs(299) <= layer0_outputs(8529);
    outputs(300) <= (layer0_outputs(3136)) and not (layer0_outputs(5059));
    outputs(301) <= (layer0_outputs(7296)) and (layer0_outputs(9321));
    outputs(302) <= (layer0_outputs(790)) or (layer0_outputs(6652));
    outputs(303) <= not(layer0_outputs(6257));
    outputs(304) <= not(layer0_outputs(4693)) or (layer0_outputs(7743));
    outputs(305) <= (layer0_outputs(7257)) xor (layer0_outputs(6146));
    outputs(306) <= layer0_outputs(6157);
    outputs(307) <= not(layer0_outputs(6737));
    outputs(308) <= layer0_outputs(6802);
    outputs(309) <= layer0_outputs(9809);
    outputs(310) <= layer0_outputs(1854);
    outputs(311) <= (layer0_outputs(5620)) and (layer0_outputs(3214));
    outputs(312) <= not(layer0_outputs(4088));
    outputs(313) <= (layer0_outputs(9683)) and not (layer0_outputs(2413));
    outputs(314) <= layer0_outputs(7566);
    outputs(315) <= (layer0_outputs(6571)) and (layer0_outputs(6958));
    outputs(316) <= not(layer0_outputs(6915));
    outputs(317) <= not(layer0_outputs(5985)) or (layer0_outputs(3190));
    outputs(318) <= not(layer0_outputs(7717));
    outputs(319) <= not(layer0_outputs(3882)) or (layer0_outputs(6206));
    outputs(320) <= (layer0_outputs(5776)) and (layer0_outputs(1838));
    outputs(321) <= layer0_outputs(1572);
    outputs(322) <= not(layer0_outputs(707));
    outputs(323) <= not(layer0_outputs(7503));
    outputs(324) <= not(layer0_outputs(3578));
    outputs(325) <= not(layer0_outputs(6336));
    outputs(326) <= layer0_outputs(2513);
    outputs(327) <= (layer0_outputs(8700)) and (layer0_outputs(6109));
    outputs(328) <= not((layer0_outputs(8523)) xor (layer0_outputs(7105)));
    outputs(329) <= layer0_outputs(25);
    outputs(330) <= not(layer0_outputs(6017));
    outputs(331) <= not((layer0_outputs(6705)) xor (layer0_outputs(7480)));
    outputs(332) <= not(layer0_outputs(8900));
    outputs(333) <= layer0_outputs(4167);
    outputs(334) <= not((layer0_outputs(8716)) xor (layer0_outputs(368)));
    outputs(335) <= not(layer0_outputs(9932));
    outputs(336) <= not(layer0_outputs(4319)) or (layer0_outputs(5364));
    outputs(337) <= (layer0_outputs(1844)) and not (layer0_outputs(7853));
    outputs(338) <= not((layer0_outputs(3283)) xor (layer0_outputs(8446)));
    outputs(339) <= not(layer0_outputs(2812));
    outputs(340) <= (layer0_outputs(774)) xor (layer0_outputs(1849));
    outputs(341) <= not((layer0_outputs(3403)) xor (layer0_outputs(8062)));
    outputs(342) <= not(layer0_outputs(10055));
    outputs(343) <= not(layer0_outputs(7405)) or (layer0_outputs(1068));
    outputs(344) <= (layer0_outputs(6446)) xor (layer0_outputs(8131));
    outputs(345) <= (layer0_outputs(9898)) or (layer0_outputs(9634));
    outputs(346) <= not((layer0_outputs(9904)) xor (layer0_outputs(3540)));
    outputs(347) <= not((layer0_outputs(1634)) xor (layer0_outputs(7104)));
    outputs(348) <= layer0_outputs(9734);
    outputs(349) <= not(layer0_outputs(4184)) or (layer0_outputs(1564));
    outputs(350) <= not(layer0_outputs(1578));
    outputs(351) <= (layer0_outputs(2955)) xor (layer0_outputs(7231));
    outputs(352) <= layer0_outputs(524);
    outputs(353) <= layer0_outputs(7206);
    outputs(354) <= layer0_outputs(7951);
    outputs(355) <= layer0_outputs(6910);
    outputs(356) <= not((layer0_outputs(8348)) or (layer0_outputs(5597)));
    outputs(357) <= not(layer0_outputs(2923));
    outputs(358) <= not(layer0_outputs(9370));
    outputs(359) <= (layer0_outputs(2689)) and not (layer0_outputs(1254));
    outputs(360) <= not((layer0_outputs(2181)) and (layer0_outputs(8)));
    outputs(361) <= not(layer0_outputs(7236));
    outputs(362) <= layer0_outputs(8961);
    outputs(363) <= (layer0_outputs(8911)) xor (layer0_outputs(4));
    outputs(364) <= not(layer0_outputs(9877)) or (layer0_outputs(307));
    outputs(365) <= not((layer0_outputs(7008)) or (layer0_outputs(1865)));
    outputs(366) <= (layer0_outputs(2692)) xor (layer0_outputs(1611));
    outputs(367) <= not((layer0_outputs(1867)) or (layer0_outputs(9815)));
    outputs(368) <= (layer0_outputs(5504)) or (layer0_outputs(3767));
    outputs(369) <= layer0_outputs(2604);
    outputs(370) <= not(layer0_outputs(3391));
    outputs(371) <= (layer0_outputs(8200)) and not (layer0_outputs(1808));
    outputs(372) <= not(layer0_outputs(3762));
    outputs(373) <= not(layer0_outputs(3424)) or (layer0_outputs(4492));
    outputs(374) <= layer0_outputs(8142);
    outputs(375) <= layer0_outputs(1803);
    outputs(376) <= layer0_outputs(4287);
    outputs(377) <= (layer0_outputs(2300)) and not (layer0_outputs(7922));
    outputs(378) <= not(layer0_outputs(6457));
    outputs(379) <= (layer0_outputs(775)) or (layer0_outputs(295));
    outputs(380) <= (layer0_outputs(8257)) and not (layer0_outputs(3418));
    outputs(381) <= not(layer0_outputs(2204));
    outputs(382) <= (layer0_outputs(4121)) and not (layer0_outputs(3921));
    outputs(383) <= (layer0_outputs(2988)) and not (layer0_outputs(7731));
    outputs(384) <= not((layer0_outputs(1001)) xor (layer0_outputs(2904)));
    outputs(385) <= layer0_outputs(2657);
    outputs(386) <= (layer0_outputs(3945)) or (layer0_outputs(3677));
    outputs(387) <= layer0_outputs(8842);
    outputs(388) <= not(layer0_outputs(2089)) or (layer0_outputs(3945));
    outputs(389) <= not((layer0_outputs(4895)) xor (layer0_outputs(1719)));
    outputs(390) <= (layer0_outputs(8992)) xor (layer0_outputs(5655));
    outputs(391) <= (layer0_outputs(1879)) or (layer0_outputs(5710));
    outputs(392) <= layer0_outputs(5457);
    outputs(393) <= not(layer0_outputs(7287));
    outputs(394) <= not((layer0_outputs(2875)) xor (layer0_outputs(7719)));
    outputs(395) <= (layer0_outputs(2529)) or (layer0_outputs(7542));
    outputs(396) <= not(layer0_outputs(10076)) or (layer0_outputs(323));
    outputs(397) <= not(layer0_outputs(3001)) or (layer0_outputs(3901));
    outputs(398) <= layer0_outputs(1244);
    outputs(399) <= layer0_outputs(3253);
    outputs(400) <= layer0_outputs(4527);
    outputs(401) <= not((layer0_outputs(1214)) xor (layer0_outputs(6989)));
    outputs(402) <= not((layer0_outputs(6170)) xor (layer0_outputs(8001)));
    outputs(403) <= layer0_outputs(2500);
    outputs(404) <= not((layer0_outputs(1029)) xor (layer0_outputs(837)));
    outputs(405) <= not((layer0_outputs(8468)) xor (layer0_outputs(2456)));
    outputs(406) <= not((layer0_outputs(434)) xor (layer0_outputs(1553)));
    outputs(407) <= (layer0_outputs(9506)) xor (layer0_outputs(6942));
    outputs(408) <= (layer0_outputs(7932)) and not (layer0_outputs(6667));
    outputs(409) <= (layer0_outputs(7980)) xor (layer0_outputs(1268));
    outputs(410) <= not(layer0_outputs(7778));
    outputs(411) <= (layer0_outputs(2104)) xor (layer0_outputs(787));
    outputs(412) <= layer0_outputs(5934);
    outputs(413) <= not(layer0_outputs(7227));
    outputs(414) <= (layer0_outputs(5149)) or (layer0_outputs(7407));
    outputs(415) <= not(layer0_outputs(217)) or (layer0_outputs(7567));
    outputs(416) <= not((layer0_outputs(8370)) xor (layer0_outputs(1293)));
    outputs(417) <= not(layer0_outputs(4326)) or (layer0_outputs(1891));
    outputs(418) <= layer0_outputs(851);
    outputs(419) <= layer0_outputs(4899);
    outputs(420) <= layer0_outputs(2732);
    outputs(421) <= layer0_outputs(5261);
    outputs(422) <= not((layer0_outputs(1608)) xor (layer0_outputs(10079)));
    outputs(423) <= layer0_outputs(2038);
    outputs(424) <= not((layer0_outputs(347)) xor (layer0_outputs(4010)));
    outputs(425) <= not((layer0_outputs(5838)) or (layer0_outputs(5681)));
    outputs(426) <= (layer0_outputs(2582)) xor (layer0_outputs(5492));
    outputs(427) <= not(layer0_outputs(9446));
    outputs(428) <= (layer0_outputs(9212)) and not (layer0_outputs(3537));
    outputs(429) <= not(layer0_outputs(4604)) or (layer0_outputs(4641));
    outputs(430) <= not(layer0_outputs(1468)) or (layer0_outputs(361));
    outputs(431) <= not(layer0_outputs(1082));
    outputs(432) <= not(layer0_outputs(3815)) or (layer0_outputs(3176));
    outputs(433) <= not(layer0_outputs(6335));
    outputs(434) <= layer0_outputs(8962);
    outputs(435) <= not(layer0_outputs(7050));
    outputs(436) <= not((layer0_outputs(9042)) or (layer0_outputs(10091)));
    outputs(437) <= (layer0_outputs(8427)) or (layer0_outputs(7465));
    outputs(438) <= not(layer0_outputs(3840));
    outputs(439) <= not(layer0_outputs(10089)) or (layer0_outputs(5767));
    outputs(440) <= not(layer0_outputs(5931));
    outputs(441) <= not((layer0_outputs(8367)) xor (layer0_outputs(2601)));
    outputs(442) <= not((layer0_outputs(8396)) and (layer0_outputs(755)));
    outputs(443) <= not(layer0_outputs(28));
    outputs(444) <= layer0_outputs(9436);
    outputs(445) <= not((layer0_outputs(3435)) xor (layer0_outputs(9974)));
    outputs(446) <= (layer0_outputs(9180)) or (layer0_outputs(3857));
    outputs(447) <= not(layer0_outputs(9868));
    outputs(448) <= (layer0_outputs(2039)) and (layer0_outputs(2536));
    outputs(449) <= not((layer0_outputs(6503)) and (layer0_outputs(8521)));
    outputs(450) <= not(layer0_outputs(3570));
    outputs(451) <= layer0_outputs(582);
    outputs(452) <= layer0_outputs(6771);
    outputs(453) <= not(layer0_outputs(1804)) or (layer0_outputs(4525));
    outputs(454) <= not(layer0_outputs(2625)) or (layer0_outputs(841));
    outputs(455) <= not(layer0_outputs(8782));
    outputs(456) <= not(layer0_outputs(3928));
    outputs(457) <= not((layer0_outputs(7590)) xor (layer0_outputs(2905)));
    outputs(458) <= not(layer0_outputs(3342)) or (layer0_outputs(2070));
    outputs(459) <= (layer0_outputs(2110)) and not (layer0_outputs(5545));
    outputs(460) <= layer0_outputs(4141);
    outputs(461) <= not(layer0_outputs(1271));
    outputs(462) <= (layer0_outputs(6718)) and (layer0_outputs(4932));
    outputs(463) <= layer0_outputs(1514);
    outputs(464) <= not((layer0_outputs(6395)) xor (layer0_outputs(10031)));
    outputs(465) <= (layer0_outputs(5537)) and not (layer0_outputs(5295));
    outputs(466) <= (layer0_outputs(5189)) xor (layer0_outputs(1604));
    outputs(467) <= not(layer0_outputs(1597));
    outputs(468) <= not(layer0_outputs(8895)) or (layer0_outputs(5249));
    outputs(469) <= (layer0_outputs(5449)) or (layer0_outputs(4417));
    outputs(470) <= not((layer0_outputs(3749)) xor (layer0_outputs(9656)));
    outputs(471) <= (layer0_outputs(3487)) or (layer0_outputs(4953));
    outputs(472) <= not(layer0_outputs(7349));
    outputs(473) <= not(layer0_outputs(2664)) or (layer0_outputs(4156));
    outputs(474) <= not(layer0_outputs(4222)) or (layer0_outputs(1653));
    outputs(475) <= not(layer0_outputs(5197)) or (layer0_outputs(7427));
    outputs(476) <= not(layer0_outputs(7406));
    outputs(477) <= not(layer0_outputs(6546));
    outputs(478) <= not((layer0_outputs(5933)) xor (layer0_outputs(1671)));
    outputs(479) <= not((layer0_outputs(2873)) or (layer0_outputs(7785)));
    outputs(480) <= layer0_outputs(6460);
    outputs(481) <= not(layer0_outputs(9068)) or (layer0_outputs(2986));
    outputs(482) <= not((layer0_outputs(6891)) and (layer0_outputs(1743)));
    outputs(483) <= (layer0_outputs(7974)) and not (layer0_outputs(6165));
    outputs(484) <= (layer0_outputs(9556)) and (layer0_outputs(825));
    outputs(485) <= not((layer0_outputs(785)) xor (layer0_outputs(4363)));
    outputs(486) <= not((layer0_outputs(488)) or (layer0_outputs(74)));
    outputs(487) <= (layer0_outputs(10220)) xor (layer0_outputs(9540));
    outputs(488) <= (layer0_outputs(8862)) and not (layer0_outputs(5671));
    outputs(489) <= not((layer0_outputs(4939)) xor (layer0_outputs(8767)));
    outputs(490) <= layer0_outputs(5102);
    outputs(491) <= not(layer0_outputs(7940)) or (layer0_outputs(2555));
    outputs(492) <= not(layer0_outputs(5756));
    outputs(493) <= not(layer0_outputs(5977));
    outputs(494) <= layer0_outputs(5984);
    outputs(495) <= not((layer0_outputs(7722)) or (layer0_outputs(291)));
    outputs(496) <= layer0_outputs(9315);
    outputs(497) <= not(layer0_outputs(7077));
    outputs(498) <= not(layer0_outputs(6044));
    outputs(499) <= layer0_outputs(6195);
    outputs(500) <= not((layer0_outputs(1876)) and (layer0_outputs(7745)));
    outputs(501) <= not((layer0_outputs(6782)) xor (layer0_outputs(2302)));
    outputs(502) <= not((layer0_outputs(5187)) and (layer0_outputs(7766)));
    outputs(503) <= layer0_outputs(6802);
    outputs(504) <= not(layer0_outputs(9225));
    outputs(505) <= (layer0_outputs(8376)) and not (layer0_outputs(7102));
    outputs(506) <= (layer0_outputs(4483)) and (layer0_outputs(3492));
    outputs(507) <= not(layer0_outputs(4210));
    outputs(508) <= layer0_outputs(7064);
    outputs(509) <= (layer0_outputs(7319)) and not (layer0_outputs(937));
    outputs(510) <= not(layer0_outputs(4631));
    outputs(511) <= (layer0_outputs(144)) or (layer0_outputs(391));
    outputs(512) <= (layer0_outputs(294)) and (layer0_outputs(9077));
    outputs(513) <= not(layer0_outputs(2822));
    outputs(514) <= (layer0_outputs(1852)) or (layer0_outputs(490));
    outputs(515) <= not((layer0_outputs(2078)) xor (layer0_outputs(6656)));
    outputs(516) <= not(layer0_outputs(1253));
    outputs(517) <= layer0_outputs(7983);
    outputs(518) <= not((layer0_outputs(6159)) xor (layer0_outputs(7704)));
    outputs(519) <= layer0_outputs(5743);
    outputs(520) <= (layer0_outputs(2557)) and not (layer0_outputs(5563));
    outputs(521) <= not(layer0_outputs(4419));
    outputs(522) <= not((layer0_outputs(4231)) xor (layer0_outputs(6713)));
    outputs(523) <= (layer0_outputs(6221)) and not (layer0_outputs(10145));
    outputs(524) <= not((layer0_outputs(2452)) xor (layer0_outputs(1957)));
    outputs(525) <= not(layer0_outputs(7662));
    outputs(526) <= not(layer0_outputs(3408));
    outputs(527) <= layer0_outputs(7566);
    outputs(528) <= not((layer0_outputs(1134)) and (layer0_outputs(8766)));
    outputs(529) <= (layer0_outputs(10110)) or (layer0_outputs(8395));
    outputs(530) <= not(layer0_outputs(305));
    outputs(531) <= (layer0_outputs(2908)) or (layer0_outputs(2179));
    outputs(532) <= layer0_outputs(5982);
    outputs(533) <= (layer0_outputs(3195)) or (layer0_outputs(6818));
    outputs(534) <= not((layer0_outputs(2730)) and (layer0_outputs(9265)));
    outputs(535) <= not(layer0_outputs(7793));
    outputs(536) <= (layer0_outputs(1306)) or (layer0_outputs(9530));
    outputs(537) <= not(layer0_outputs(10142));
    outputs(538) <= not((layer0_outputs(844)) and (layer0_outputs(9513)));
    outputs(539) <= not((layer0_outputs(7095)) and (layer0_outputs(1394)));
    outputs(540) <= not((layer0_outputs(3464)) and (layer0_outputs(2467)));
    outputs(541) <= (layer0_outputs(3763)) and not (layer0_outputs(9542));
    outputs(542) <= layer0_outputs(9430);
    outputs(543) <= not((layer0_outputs(915)) or (layer0_outputs(7922)));
    outputs(544) <= not(layer0_outputs(1107));
    outputs(545) <= layer0_outputs(9694);
    outputs(546) <= not(layer0_outputs(6753));
    outputs(547) <= not(layer0_outputs(922));
    outputs(548) <= not(layer0_outputs(2013));
    outputs(549) <= not(layer0_outputs(9713));
    outputs(550) <= not(layer0_outputs(2276)) or (layer0_outputs(9916));
    outputs(551) <= not(layer0_outputs(4968));
    outputs(552) <= not(layer0_outputs(7469));
    outputs(553) <= not(layer0_outputs(8945));
    outputs(554) <= not(layer0_outputs(7776));
    outputs(555) <= not(layer0_outputs(9108));
    outputs(556) <= (layer0_outputs(4219)) xor (layer0_outputs(4746));
    outputs(557) <= (layer0_outputs(3084)) or (layer0_outputs(2232));
    outputs(558) <= not(layer0_outputs(8539));
    outputs(559) <= not((layer0_outputs(528)) xor (layer0_outputs(2037)));
    outputs(560) <= not(layer0_outputs(9330)) or (layer0_outputs(1626));
    outputs(561) <= not(layer0_outputs(9092));
    outputs(562) <= not(layer0_outputs(8314));
    outputs(563) <= (layer0_outputs(6413)) or (layer0_outputs(10236));
    outputs(564) <= not(layer0_outputs(3460));
    outputs(565) <= (layer0_outputs(2763)) and not (layer0_outputs(7701));
    outputs(566) <= layer0_outputs(5501);
    outputs(567) <= layer0_outputs(4206);
    outputs(568) <= layer0_outputs(5908);
    outputs(569) <= layer0_outputs(4900);
    outputs(570) <= layer0_outputs(6430);
    outputs(571) <= not(layer0_outputs(4548)) or (layer0_outputs(6449));
    outputs(572) <= not(layer0_outputs(704));
    outputs(573) <= layer0_outputs(88);
    outputs(574) <= (layer0_outputs(3636)) and not (layer0_outputs(1498));
    outputs(575) <= not((layer0_outputs(5015)) or (layer0_outputs(1814)));
    outputs(576) <= (layer0_outputs(8721)) xor (layer0_outputs(3380));
    outputs(577) <= not(layer0_outputs(1309));
    outputs(578) <= not((layer0_outputs(1252)) and (layer0_outputs(6660)));
    outputs(579) <= not(layer0_outputs(4684));
    outputs(580) <= not(layer0_outputs(1906));
    outputs(581) <= (layer0_outputs(3335)) and not (layer0_outputs(2587));
    outputs(582) <= layer0_outputs(9981);
    outputs(583) <= not((layer0_outputs(1410)) or (layer0_outputs(7767)));
    outputs(584) <= not((layer0_outputs(8923)) xor (layer0_outputs(10181)));
    outputs(585) <= not((layer0_outputs(1622)) xor (layer0_outputs(5295)));
    outputs(586) <= not(layer0_outputs(1422)) or (layer0_outputs(7328));
    outputs(587) <= (layer0_outputs(2336)) and not (layer0_outputs(912));
    outputs(588) <= not(layer0_outputs(7295));
    outputs(589) <= not(layer0_outputs(231)) or (layer0_outputs(4961));
    outputs(590) <= layer0_outputs(6294);
    outputs(591) <= layer0_outputs(3710);
    outputs(592) <= (layer0_outputs(9218)) and not (layer0_outputs(1224));
    outputs(593) <= (layer0_outputs(2994)) and not (layer0_outputs(8190));
    outputs(594) <= (layer0_outputs(5607)) and not (layer0_outputs(2731));
    outputs(595) <= layer0_outputs(6874);
    outputs(596) <= layer0_outputs(5044);
    outputs(597) <= layer0_outputs(7495);
    outputs(598) <= not(layer0_outputs(8147));
    outputs(599) <= (layer0_outputs(4212)) xor (layer0_outputs(3719));
    outputs(600) <= not(layer0_outputs(9005)) or (layer0_outputs(8498));
    outputs(601) <= not(layer0_outputs(9782));
    outputs(602) <= not((layer0_outputs(6180)) xor (layer0_outputs(3414)));
    outputs(603) <= (layer0_outputs(954)) and (layer0_outputs(6236));
    outputs(604) <= not((layer0_outputs(9140)) xor (layer0_outputs(4540)));
    outputs(605) <= (layer0_outputs(7430)) and (layer0_outputs(1810));
    outputs(606) <= layer0_outputs(13);
    outputs(607) <= not(layer0_outputs(4398)) or (layer0_outputs(4131));
    outputs(608) <= not(layer0_outputs(7598));
    outputs(609) <= not((layer0_outputs(7564)) xor (layer0_outputs(62)));
    outputs(610) <= not(layer0_outputs(6539)) or (layer0_outputs(6127));
    outputs(611) <= not((layer0_outputs(1642)) and (layer0_outputs(1101)));
    outputs(612) <= not((layer0_outputs(5940)) or (layer0_outputs(7286)));
    outputs(613) <= layer0_outputs(6948);
    outputs(614) <= (layer0_outputs(9495)) xor (layer0_outputs(4346));
    outputs(615) <= (layer0_outputs(279)) xor (layer0_outputs(4085));
    outputs(616) <= (layer0_outputs(3351)) and not (layer0_outputs(9868));
    outputs(617) <= layer0_outputs(3769);
    outputs(618) <= not(layer0_outputs(8694));
    outputs(619) <= (layer0_outputs(2959)) xor (layer0_outputs(9792));
    outputs(620) <= (layer0_outputs(3319)) xor (layer0_outputs(6042));
    outputs(621) <= not(layer0_outputs(2791));
    outputs(622) <= not(layer0_outputs(10212));
    outputs(623) <= not(layer0_outputs(9144)) or (layer0_outputs(4834));
    outputs(624) <= not((layer0_outputs(6250)) or (layer0_outputs(9294)));
    outputs(625) <= layer0_outputs(132);
    outputs(626) <= not(layer0_outputs(3446));
    outputs(627) <= not((layer0_outputs(4864)) xor (layer0_outputs(3200)));
    outputs(628) <= (layer0_outputs(5824)) xor (layer0_outputs(5702));
    outputs(629) <= not((layer0_outputs(4852)) and (layer0_outputs(7729)));
    outputs(630) <= (layer0_outputs(980)) xor (layer0_outputs(7520));
    outputs(631) <= layer0_outputs(9388);
    outputs(632) <= not(layer0_outputs(8935));
    outputs(633) <= (layer0_outputs(3281)) or (layer0_outputs(9957));
    outputs(634) <= not(layer0_outputs(2349));
    outputs(635) <= (layer0_outputs(5739)) and not (layer0_outputs(2884));
    outputs(636) <= (layer0_outputs(8366)) and not (layer0_outputs(7385));
    outputs(637) <= not(layer0_outputs(6308));
    outputs(638) <= layer0_outputs(1652);
    outputs(639) <= not(layer0_outputs(1941));
    outputs(640) <= (layer0_outputs(1624)) and (layer0_outputs(6579));
    outputs(641) <= layer0_outputs(7491);
    outputs(642) <= not(layer0_outputs(8963)) or (layer0_outputs(6516));
    outputs(643) <= not(layer0_outputs(9125)) or (layer0_outputs(10234));
    outputs(644) <= not((layer0_outputs(7045)) xor (layer0_outputs(4737)));
    outputs(645) <= not((layer0_outputs(7140)) xor (layer0_outputs(2032)));
    outputs(646) <= layer0_outputs(2768);
    outputs(647) <= not(layer0_outputs(8616));
    outputs(648) <= not(layer0_outputs(8328));
    outputs(649) <= (layer0_outputs(9302)) and (layer0_outputs(4089));
    outputs(650) <= (layer0_outputs(4699)) and (layer0_outputs(8988));
    outputs(651) <= (layer0_outputs(4254)) xor (layer0_outputs(5172));
    outputs(652) <= (layer0_outputs(7956)) or (layer0_outputs(8025));
    outputs(653) <= layer0_outputs(5595);
    outputs(654) <= not(layer0_outputs(8299)) or (layer0_outputs(501));
    outputs(655) <= (layer0_outputs(4371)) and not (layer0_outputs(9692));
    outputs(656) <= (layer0_outputs(3663)) and (layer0_outputs(1277));
    outputs(657) <= not((layer0_outputs(8088)) and (layer0_outputs(2638)));
    outputs(658) <= not(layer0_outputs(6777));
    outputs(659) <= (layer0_outputs(8861)) and (layer0_outputs(8280));
    outputs(660) <= not(layer0_outputs(9058));
    outputs(661) <= not((layer0_outputs(1339)) xor (layer0_outputs(473)));
    outputs(662) <= (layer0_outputs(3047)) xor (layer0_outputs(6103));
    outputs(663) <= not((layer0_outputs(1271)) or (layer0_outputs(8307)));
    outputs(664) <= (layer0_outputs(7125)) and (layer0_outputs(5472));
    outputs(665) <= layer0_outputs(1433);
    outputs(666) <= not(layer0_outputs(3057));
    outputs(667) <= not((layer0_outputs(2704)) and (layer0_outputs(6052)));
    outputs(668) <= (layer0_outputs(1201)) and not (layer0_outputs(1889));
    outputs(669) <= not(layer0_outputs(6525));
    outputs(670) <= not(layer0_outputs(6949)) or (layer0_outputs(4225));
    outputs(671) <= (layer0_outputs(7433)) and not (layer0_outputs(749));
    outputs(672) <= not(layer0_outputs(97));
    outputs(673) <= layer0_outputs(9420);
    outputs(674) <= not((layer0_outputs(4879)) and (layer0_outputs(2277)));
    outputs(675) <= not(layer0_outputs(8026));
    outputs(676) <= layer0_outputs(3764);
    outputs(677) <= layer0_outputs(763);
    outputs(678) <= not(layer0_outputs(8948)) or (layer0_outputs(1509));
    outputs(679) <= not(layer0_outputs(6592)) or (layer0_outputs(5752));
    outputs(680) <= not(layer0_outputs(2675));
    outputs(681) <= layer0_outputs(4715);
    outputs(682) <= layer0_outputs(8090);
    outputs(683) <= layer0_outputs(5687);
    outputs(684) <= not(layer0_outputs(10175)) or (layer0_outputs(10204));
    outputs(685) <= layer0_outputs(8085);
    outputs(686) <= (layer0_outputs(4363)) and (layer0_outputs(5307));
    outputs(687) <= (layer0_outputs(2342)) xor (layer0_outputs(9925));
    outputs(688) <= not(layer0_outputs(1022));
    outputs(689) <= (layer0_outputs(4565)) xor (layer0_outputs(8580));
    outputs(690) <= layer0_outputs(6718);
    outputs(691) <= not(layer0_outputs(8350));
    outputs(692) <= not((layer0_outputs(7015)) xor (layer0_outputs(1373)));
    outputs(693) <= not(layer0_outputs(4414)) or (layer0_outputs(3958));
    outputs(694) <= not(layer0_outputs(1118));
    outputs(695) <= not((layer0_outputs(8481)) xor (layer0_outputs(8497)));
    outputs(696) <= (layer0_outputs(4435)) or (layer0_outputs(1400));
    outputs(697) <= not((layer0_outputs(6923)) xor (layer0_outputs(9259)));
    outputs(698) <= not(layer0_outputs(9033));
    outputs(699) <= not(layer0_outputs(3068));
    outputs(700) <= not(layer0_outputs(278));
    outputs(701) <= not(layer0_outputs(8379));
    outputs(702) <= layer0_outputs(8787);
    outputs(703) <= not(layer0_outputs(4295));
    outputs(704) <= not((layer0_outputs(8591)) xor (layer0_outputs(1789)));
    outputs(705) <= (layer0_outputs(3805)) or (layer0_outputs(9149));
    outputs(706) <= (layer0_outputs(4856)) xor (layer0_outputs(8569));
    outputs(707) <= (layer0_outputs(7906)) xor (layer0_outputs(9184));
    outputs(708) <= not(layer0_outputs(2428));
    outputs(709) <= (layer0_outputs(7591)) and not (layer0_outputs(2829));
    outputs(710) <= layer0_outputs(416);
    outputs(711) <= not((layer0_outputs(4128)) xor (layer0_outputs(4397)));
    outputs(712) <= (layer0_outputs(7392)) xor (layer0_outputs(7415));
    outputs(713) <= (layer0_outputs(3339)) xor (layer0_outputs(10113));
    outputs(714) <= (layer0_outputs(1413)) xor (layer0_outputs(2524));
    outputs(715) <= not(layer0_outputs(8134));
    outputs(716) <= not((layer0_outputs(6774)) xor (layer0_outputs(9168)));
    outputs(717) <= not(layer0_outputs(8550));
    outputs(718) <= (layer0_outputs(2352)) xor (layer0_outputs(4720));
    outputs(719) <= layer0_outputs(2301);
    outputs(720) <= (layer0_outputs(4083)) and not (layer0_outputs(5526));
    outputs(721) <= layer0_outputs(4606);
    outputs(722) <= layer0_outputs(7672);
    outputs(723) <= (layer0_outputs(1560)) or (layer0_outputs(5989));
    outputs(724) <= not(layer0_outputs(9910));
    outputs(725) <= not(layer0_outputs(2176));
    outputs(726) <= layer0_outputs(8938);
    outputs(727) <= layer0_outputs(7240);
    outputs(728) <= (layer0_outputs(7543)) and (layer0_outputs(8549));
    outputs(729) <= layer0_outputs(3754);
    outputs(730) <= (layer0_outputs(9824)) and (layer0_outputs(8569));
    outputs(731) <= layer0_outputs(7597);
    outputs(732) <= not((layer0_outputs(9114)) xor (layer0_outputs(6653)));
    outputs(733) <= (layer0_outputs(2142)) and not (layer0_outputs(6615));
    outputs(734) <= (layer0_outputs(1763)) or (layer0_outputs(608));
    outputs(735) <= layer0_outputs(893);
    outputs(736) <= not(layer0_outputs(1841));
    outputs(737) <= layer0_outputs(2596);
    outputs(738) <= layer0_outputs(2036);
    outputs(739) <= not(layer0_outputs(972));
    outputs(740) <= (layer0_outputs(5569)) and not (layer0_outputs(8487));
    outputs(741) <= not(layer0_outputs(9594));
    outputs(742) <= not(layer0_outputs(1953));
    outputs(743) <= not(layer0_outputs(1875));
    outputs(744) <= (layer0_outputs(4145)) and not (layer0_outputs(2602));
    outputs(745) <= layer0_outputs(9490);
    outputs(746) <= not(layer0_outputs(6339));
    outputs(747) <= not((layer0_outputs(6282)) xor (layer0_outputs(6166)));
    outputs(748) <= layer0_outputs(4302);
    outputs(749) <= not(layer0_outputs(3645));
    outputs(750) <= not((layer0_outputs(1011)) xor (layer0_outputs(1416)));
    outputs(751) <= not(layer0_outputs(6530)) or (layer0_outputs(6843));
    outputs(752) <= (layer0_outputs(2838)) and (layer0_outputs(5300));
    outputs(753) <= not(layer0_outputs(2196));
    outputs(754) <= not((layer0_outputs(7751)) and (layer0_outputs(312)));
    outputs(755) <= layer0_outputs(5990);
    outputs(756) <= (layer0_outputs(8594)) and (layer0_outputs(2074));
    outputs(757) <= (layer0_outputs(5342)) and not (layer0_outputs(5840));
    outputs(758) <= not(layer0_outputs(2098)) or (layer0_outputs(2643));
    outputs(759) <= (layer0_outputs(10178)) or (layer0_outputs(7103));
    outputs(760) <= (layer0_outputs(1490)) and (layer0_outputs(7993));
    outputs(761) <= not(layer0_outputs(4835)) or (layer0_outputs(5617));
    outputs(762) <= not(layer0_outputs(6491));
    outputs(763) <= (layer0_outputs(6221)) xor (layer0_outputs(1915));
    outputs(764) <= layer0_outputs(9559);
    outputs(765) <= not(layer0_outputs(4710)) or (layer0_outputs(3902));
    outputs(766) <= not(layer0_outputs(7383));
    outputs(767) <= (layer0_outputs(5105)) xor (layer0_outputs(9834));
    outputs(768) <= (layer0_outputs(2317)) and not (layer0_outputs(1002));
    outputs(769) <= not(layer0_outputs(6477));
    outputs(770) <= (layer0_outputs(6039)) and not (layer0_outputs(8733));
    outputs(771) <= layer0_outputs(1297);
    outputs(772) <= (layer0_outputs(4432)) xor (layer0_outputs(1908));
    outputs(773) <= layer0_outputs(1207);
    outputs(774) <= layer0_outputs(136);
    outputs(775) <= not((layer0_outputs(2442)) xor (layer0_outputs(3402)));
    outputs(776) <= not((layer0_outputs(1715)) xor (layer0_outputs(5697)));
    outputs(777) <= not(layer0_outputs(4311));
    outputs(778) <= (layer0_outputs(7074)) xor (layer0_outputs(4279));
    outputs(779) <= (layer0_outputs(1877)) and not (layer0_outputs(8984));
    outputs(780) <= not((layer0_outputs(9722)) xor (layer0_outputs(10071)));
    outputs(781) <= (layer0_outputs(9969)) or (layer0_outputs(9610));
    outputs(782) <= (layer0_outputs(3195)) xor (layer0_outputs(8980));
    outputs(783) <= not(layer0_outputs(3154));
    outputs(784) <= not(layer0_outputs(7675));
    outputs(785) <= not((layer0_outputs(5536)) or (layer0_outputs(465)));
    outputs(786) <= (layer0_outputs(577)) and (layer0_outputs(9758));
    outputs(787) <= not(layer0_outputs(2117));
    outputs(788) <= layer0_outputs(2894);
    outputs(789) <= (layer0_outputs(452)) and not (layer0_outputs(3995));
    outputs(790) <= layer0_outputs(9417);
    outputs(791) <= not((layer0_outputs(8511)) xor (layer0_outputs(2734)));
    outputs(792) <= not(layer0_outputs(8491));
    outputs(793) <= (layer0_outputs(4247)) and (layer0_outputs(9734));
    outputs(794) <= not(layer0_outputs(4051));
    outputs(795) <= (layer0_outputs(9902)) and not (layer0_outputs(7608));
    outputs(796) <= not(layer0_outputs(2430));
    outputs(797) <= layer0_outputs(1700);
    outputs(798) <= (layer0_outputs(2469)) xor (layer0_outputs(4594));
    outputs(799) <= not((layer0_outputs(5339)) xor (layer0_outputs(8296)));
    outputs(800) <= (layer0_outputs(8038)) xor (layer0_outputs(3693));
    outputs(801) <= (layer0_outputs(1298)) and not (layer0_outputs(9587));
    outputs(802) <= layer0_outputs(3194);
    outputs(803) <= (layer0_outputs(6622)) xor (layer0_outputs(3545));
    outputs(804) <= (layer0_outputs(4875)) and (layer0_outputs(7989));
    outputs(805) <= not(layer0_outputs(1417));
    outputs(806) <= layer0_outputs(1475);
    outputs(807) <= not((layer0_outputs(2703)) and (layer0_outputs(6615)));
    outputs(808) <= (layer0_outputs(6707)) xor (layer0_outputs(3268));
    outputs(809) <= not(layer0_outputs(4273));
    outputs(810) <= not(layer0_outputs(7412));
    outputs(811) <= layer0_outputs(9953);
    outputs(812) <= layer0_outputs(6478);
    outputs(813) <= not(layer0_outputs(4040));
    outputs(814) <= layer0_outputs(1264);
    outputs(815) <= (layer0_outputs(4563)) and not (layer0_outputs(5019));
    outputs(816) <= (layer0_outputs(7455)) xor (layer0_outputs(566));
    outputs(817) <= not((layer0_outputs(5230)) or (layer0_outputs(6232)));
    outputs(818) <= not(layer0_outputs(227));
    outputs(819) <= (layer0_outputs(9223)) and not (layer0_outputs(8385));
    outputs(820) <= not((layer0_outputs(2940)) and (layer0_outputs(2956)));
    outputs(821) <= (layer0_outputs(7690)) xor (layer0_outputs(1618));
    outputs(822) <= not(layer0_outputs(7552));
    outputs(823) <= (layer0_outputs(968)) and (layer0_outputs(4271));
    outputs(824) <= layer0_outputs(2915);
    outputs(825) <= (layer0_outputs(1157)) and (layer0_outputs(8413));
    outputs(826) <= (layer0_outputs(7709)) and not (layer0_outputs(3891));
    outputs(827) <= (layer0_outputs(4421)) and not (layer0_outputs(1594));
    outputs(828) <= (layer0_outputs(5238)) and not (layer0_outputs(2227));
    outputs(829) <= not((layer0_outputs(1811)) xor (layer0_outputs(618)));
    outputs(830) <= not(layer0_outputs(7970));
    outputs(831) <= (layer0_outputs(208)) xor (layer0_outputs(6131));
    outputs(832) <= layer0_outputs(5693);
    outputs(833) <= not((layer0_outputs(2314)) and (layer0_outputs(9558)));
    outputs(834) <= not(layer0_outputs(9515)) or (layer0_outputs(7071));
    outputs(835) <= layer0_outputs(4591);
    outputs(836) <= (layer0_outputs(5299)) xor (layer0_outputs(1914));
    outputs(837) <= (layer0_outputs(8194)) or (layer0_outputs(2925));
    outputs(838) <= (layer0_outputs(7197)) and (layer0_outputs(7575));
    outputs(839) <= not(layer0_outputs(3560));
    outputs(840) <= not(layer0_outputs(2132));
    outputs(841) <= (layer0_outputs(9321)) and not (layer0_outputs(8799));
    outputs(842) <= (layer0_outputs(4507)) and not (layer0_outputs(5092));
    outputs(843) <= (layer0_outputs(10164)) xor (layer0_outputs(568));
    outputs(844) <= not(layer0_outputs(2106));
    outputs(845) <= not(layer0_outputs(3326));
    outputs(846) <= not(layer0_outputs(5079)) or (layer0_outputs(7336));
    outputs(847) <= not(layer0_outputs(1638));
    outputs(848) <= (layer0_outputs(8301)) xor (layer0_outputs(4868));
    outputs(849) <= layer0_outputs(3818);
    outputs(850) <= not((layer0_outputs(241)) or (layer0_outputs(8567)));
    outputs(851) <= layer0_outputs(3499);
    outputs(852) <= (layer0_outputs(6610)) xor (layer0_outputs(9622));
    outputs(853) <= layer0_outputs(7539);
    outputs(854) <= (layer0_outputs(7150)) and not (layer0_outputs(3533));
    outputs(855) <= not((layer0_outputs(9786)) or (layer0_outputs(1031)));
    outputs(856) <= (layer0_outputs(9379)) xor (layer0_outputs(8600));
    outputs(857) <= not(layer0_outputs(3032));
    outputs(858) <= not(layer0_outputs(9836));
    outputs(859) <= not((layer0_outputs(275)) or (layer0_outputs(3947)));
    outputs(860) <= not(layer0_outputs(2876));
    outputs(861) <= not(layer0_outputs(5513));
    outputs(862) <= not(layer0_outputs(1285)) or (layer0_outputs(4073));
    outputs(863) <= not((layer0_outputs(1225)) or (layer0_outputs(7128)));
    outputs(864) <= not(layer0_outputs(2488));
    outputs(865) <= (layer0_outputs(2507)) and not (layer0_outputs(8126));
    outputs(866) <= (layer0_outputs(1168)) and (layer0_outputs(4335));
    outputs(867) <= layer0_outputs(3322);
    outputs(868) <= not(layer0_outputs(1262));
    outputs(869) <= not(layer0_outputs(4154));
    outputs(870) <= (layer0_outputs(5097)) xor (layer0_outputs(8875));
    outputs(871) <= not((layer0_outputs(2499)) xor (layer0_outputs(6388)));
    outputs(872) <= layer0_outputs(7352);
    outputs(873) <= not(layer0_outputs(8588));
    outputs(874) <= (layer0_outputs(5758)) xor (layer0_outputs(467));
    outputs(875) <= layer0_outputs(2120);
    outputs(876) <= not(layer0_outputs(4722));
    outputs(877) <= layer0_outputs(1402);
    outputs(878) <= (layer0_outputs(8620)) xor (layer0_outputs(5900));
    outputs(879) <= layer0_outputs(5176);
    outputs(880) <= not(layer0_outputs(2673)) or (layer0_outputs(8861));
    outputs(881) <= not((layer0_outputs(7959)) xor (layer0_outputs(3746)));
    outputs(882) <= not((layer0_outputs(2236)) xor (layer0_outputs(878)));
    outputs(883) <= not(layer0_outputs(7895));
    outputs(884) <= not((layer0_outputs(380)) or (layer0_outputs(4835)));
    outputs(885) <= not(layer0_outputs(9524));
    outputs(886) <= not((layer0_outputs(7748)) and (layer0_outputs(8285)));
    outputs(887) <= (layer0_outputs(1098)) or (layer0_outputs(869));
    outputs(888) <= not((layer0_outputs(819)) or (layer0_outputs(2620)));
    outputs(889) <= not((layer0_outputs(6497)) xor (layer0_outputs(7028)));
    outputs(890) <= not(layer0_outputs(8421)) or (layer0_outputs(2678));
    outputs(891) <= (layer0_outputs(1601)) and not (layer0_outputs(610));
    outputs(892) <= not((layer0_outputs(6316)) xor (layer0_outputs(8623)));
    outputs(893) <= not(layer0_outputs(10149));
    outputs(894) <= (layer0_outputs(5984)) and not (layer0_outputs(4923));
    outputs(895) <= (layer0_outputs(10075)) and not (layer0_outputs(6919));
    outputs(896) <= layer0_outputs(5670);
    outputs(897) <= layer0_outputs(7846);
    outputs(898) <= (layer0_outputs(6371)) xor (layer0_outputs(8225));
    outputs(899) <= not(layer0_outputs(2084)) or (layer0_outputs(3769));
    outputs(900) <= (layer0_outputs(2471)) and not (layer0_outputs(5570));
    outputs(901) <= layer0_outputs(5122);
    outputs(902) <= not((layer0_outputs(5063)) or (layer0_outputs(3702)));
    outputs(903) <= not(layer0_outputs(5028)) or (layer0_outputs(1208));
    outputs(904) <= layer0_outputs(1746);
    outputs(905) <= layer0_outputs(3481);
    outputs(906) <= not(layer0_outputs(3662));
    outputs(907) <= layer0_outputs(3266);
    outputs(908) <= (layer0_outputs(10115)) xor (layer0_outputs(8578));
    outputs(909) <= not(layer0_outputs(6315));
    outputs(910) <= layer0_outputs(8687);
    outputs(911) <= layer0_outputs(7803);
    outputs(912) <= not(layer0_outputs(317)) or (layer0_outputs(4044));
    outputs(913) <= (layer0_outputs(7412)) xor (layer0_outputs(178));
    outputs(914) <= (layer0_outputs(1242)) and not (layer0_outputs(5385));
    outputs(915) <= not(layer0_outputs(6907));
    outputs(916) <= layer0_outputs(3775);
    outputs(917) <= not(layer0_outputs(7477)) or (layer0_outputs(4055));
    outputs(918) <= layer0_outputs(894);
    outputs(919) <= not(layer0_outputs(3724)) or (layer0_outputs(7992));
    outputs(920) <= layer0_outputs(3393);
    outputs(921) <= layer0_outputs(10003);
    outputs(922) <= not((layer0_outputs(2240)) xor (layer0_outputs(10051)));
    outputs(923) <= not(layer0_outputs(7873));
    outputs(924) <= not(layer0_outputs(1108));
    outputs(925) <= not((layer0_outputs(1421)) xor (layer0_outputs(7159)));
    outputs(926) <= layer0_outputs(2405);
    outputs(927) <= not(layer0_outputs(2234));
    outputs(928) <= not((layer0_outputs(287)) xor (layer0_outputs(6337)));
    outputs(929) <= not((layer0_outputs(984)) or (layer0_outputs(5765)));
    outputs(930) <= not(layer0_outputs(1922));
    outputs(931) <= layer0_outputs(5741);
    outputs(932) <= layer0_outputs(10081);
    outputs(933) <= (layer0_outputs(5501)) xor (layer0_outputs(7677));
    outputs(934) <= (layer0_outputs(4350)) xor (layer0_outputs(8424));
    outputs(935) <= not(layer0_outputs(9899));
    outputs(936) <= (layer0_outputs(4730)) or (layer0_outputs(3264));
    outputs(937) <= (layer0_outputs(7025)) and not (layer0_outputs(7686));
    outputs(938) <= not((layer0_outputs(109)) xor (layer0_outputs(9561)));
    outputs(939) <= layer0_outputs(1491);
    outputs(940) <= not((layer0_outputs(4500)) or (layer0_outputs(1712)));
    outputs(941) <= layer0_outputs(6081);
    outputs(942) <= (layer0_outputs(413)) and (layer0_outputs(4801));
    outputs(943) <= layer0_outputs(1572);
    outputs(944) <= (layer0_outputs(7312)) and not (layer0_outputs(910));
    outputs(945) <= not(layer0_outputs(4097));
    outputs(946) <= not((layer0_outputs(792)) and (layer0_outputs(5953)));
    outputs(947) <= layer0_outputs(790);
    outputs(948) <= not(layer0_outputs(637));
    outputs(949) <= not((layer0_outputs(2001)) or (layer0_outputs(8816)));
    outputs(950) <= not(layer0_outputs(7886));
    outputs(951) <= (layer0_outputs(419)) xor (layer0_outputs(5103));
    outputs(952) <= (layer0_outputs(7852)) and not (layer0_outputs(3541));
    outputs(953) <= (layer0_outputs(5737)) xor (layer0_outputs(7222));
    outputs(954) <= (layer0_outputs(8470)) xor (layer0_outputs(3851));
    outputs(955) <= not(layer0_outputs(7343));
    outputs(956) <= (layer0_outputs(764)) or (layer0_outputs(6132));
    outputs(957) <= not(layer0_outputs(4176)) or (layer0_outputs(3529));
    outputs(958) <= not(layer0_outputs(7344));
    outputs(959) <= not((layer0_outputs(4553)) xor (layer0_outputs(3002)));
    outputs(960) <= not((layer0_outputs(10119)) and (layer0_outputs(520)));
    outputs(961) <= not(layer0_outputs(9280));
    outputs(962) <= not(layer0_outputs(5015));
    outputs(963) <= not((layer0_outputs(5986)) or (layer0_outputs(7834)));
    outputs(964) <= not(layer0_outputs(5681));
    outputs(965) <= not(layer0_outputs(2418));
    outputs(966) <= not(layer0_outputs(1664));
    outputs(967) <= (layer0_outputs(7322)) and (layer0_outputs(2946));
    outputs(968) <= not(layer0_outputs(2853));
    outputs(969) <= not(layer0_outputs(4572));
    outputs(970) <= layer0_outputs(2320);
    outputs(971) <= layer0_outputs(1844);
    outputs(972) <= not((layer0_outputs(8631)) or (layer0_outputs(2294)));
    outputs(973) <= layer0_outputs(7587);
    outputs(974) <= not(layer0_outputs(1296)) or (layer0_outputs(3616));
    outputs(975) <= layer0_outputs(4138);
    outputs(976) <= layer0_outputs(4551);
    outputs(977) <= not((layer0_outputs(7771)) xor (layer0_outputs(6197)));
    outputs(978) <= layer0_outputs(660);
    outputs(979) <= (layer0_outputs(76)) xor (layer0_outputs(8515));
    outputs(980) <= not(layer0_outputs(8197));
    outputs(981) <= not((layer0_outputs(6690)) or (layer0_outputs(9036)));
    outputs(982) <= not(layer0_outputs(7143));
    outputs(983) <= not((layer0_outputs(8541)) and (layer0_outputs(2564)));
    outputs(984) <= layer0_outputs(7149);
    outputs(985) <= not(layer0_outputs(3249));
    outputs(986) <= not(layer0_outputs(4357)) or (layer0_outputs(7414));
    outputs(987) <= layer0_outputs(2975);
    outputs(988) <= layer0_outputs(2297);
    outputs(989) <= not(layer0_outputs(10069)) or (layer0_outputs(7103));
    outputs(990) <= not(layer0_outputs(1667));
    outputs(991) <= not((layer0_outputs(8738)) or (layer0_outputs(6842)));
    outputs(992) <= layer0_outputs(4445);
    outputs(993) <= not(layer0_outputs(1104));
    outputs(994) <= (layer0_outputs(1376)) and not (layer0_outputs(7511));
    outputs(995) <= layer0_outputs(4958);
    outputs(996) <= not(layer0_outputs(3808)) or (layer0_outputs(6376));
    outputs(997) <= not(layer0_outputs(3903));
    outputs(998) <= (layer0_outputs(4944)) and not (layer0_outputs(6156));
    outputs(999) <= not((layer0_outputs(8107)) xor (layer0_outputs(8539)));
    outputs(1000) <= not(layer0_outputs(6655));
    outputs(1001) <= not(layer0_outputs(4358));
    outputs(1002) <= layer0_outputs(6549);
    outputs(1003) <= (layer0_outputs(9233)) xor (layer0_outputs(5453));
    outputs(1004) <= (layer0_outputs(214)) and not (layer0_outputs(1367));
    outputs(1005) <= (layer0_outputs(9121)) or (layer0_outputs(9100));
    outputs(1006) <= layer0_outputs(4550);
    outputs(1007) <= not((layer0_outputs(6907)) or (layer0_outputs(1341)));
    outputs(1008) <= not((layer0_outputs(1422)) or (layer0_outputs(7806)));
    outputs(1009) <= not(layer0_outputs(534)) or (layer0_outputs(706));
    outputs(1010) <= not(layer0_outputs(2606));
    outputs(1011) <= not(layer0_outputs(3228));
    outputs(1012) <= not(layer0_outputs(7786));
    outputs(1013) <= not(layer0_outputs(838)) or (layer0_outputs(7536));
    outputs(1014) <= not((layer0_outputs(3918)) xor (layer0_outputs(4869)));
    outputs(1015) <= (layer0_outputs(4121)) and not (layer0_outputs(4993));
    outputs(1016) <= (layer0_outputs(6292)) or (layer0_outputs(3953));
    outputs(1017) <= not((layer0_outputs(2497)) xor (layer0_outputs(3442)));
    outputs(1018) <= (layer0_outputs(8795)) or (layer0_outputs(1969));
    outputs(1019) <= (layer0_outputs(27)) and (layer0_outputs(8352));
    outputs(1020) <= layer0_outputs(1423);
    outputs(1021) <= layer0_outputs(8747);
    outputs(1022) <= (layer0_outputs(4393)) and not (layer0_outputs(3216));
    outputs(1023) <= layer0_outputs(1145);
    outputs(1024) <= (layer0_outputs(6700)) and not (layer0_outputs(6826));
    outputs(1025) <= layer0_outputs(814);
    outputs(1026) <= not((layer0_outputs(8216)) xor (layer0_outputs(8183)));
    outputs(1027) <= not((layer0_outputs(7826)) xor (layer0_outputs(9664)));
    outputs(1028) <= (layer0_outputs(2785)) xor (layer0_outputs(6333));
    outputs(1029) <= layer0_outputs(3967);
    outputs(1030) <= not((layer0_outputs(8258)) or (layer0_outputs(2246)));
    outputs(1031) <= (layer0_outputs(4664)) and not (layer0_outputs(7129));
    outputs(1032) <= (layer0_outputs(7376)) and not (layer0_outputs(8043));
    outputs(1033) <= (layer0_outputs(9971)) and not (layer0_outputs(9927));
    outputs(1034) <= (layer0_outputs(2772)) and (layer0_outputs(1055));
    outputs(1035) <= (layer0_outputs(4754)) and (layer0_outputs(2170));
    outputs(1036) <= not(layer0_outputs(439));
    outputs(1037) <= (layer0_outputs(8713)) and not (layer0_outputs(3542));
    outputs(1038) <= not((layer0_outputs(7986)) or (layer0_outputs(10044)));
    outputs(1039) <= (layer0_outputs(2934)) and not (layer0_outputs(7816));
    outputs(1040) <= layer0_outputs(9297);
    outputs(1041) <= not((layer0_outputs(8159)) or (layer0_outputs(2995)));
    outputs(1042) <= not(layer0_outputs(8471));
    outputs(1043) <= (layer0_outputs(9557)) and not (layer0_outputs(7164));
    outputs(1044) <= (layer0_outputs(7807)) and (layer0_outputs(1631));
    outputs(1045) <= (layer0_outputs(1146)) and (layer0_outputs(5661));
    outputs(1046) <= not(layer0_outputs(7712));
    outputs(1047) <= layer0_outputs(34);
    outputs(1048) <= not((layer0_outputs(2740)) xor (layer0_outputs(187)));
    outputs(1049) <= (layer0_outputs(6399)) xor (layer0_outputs(9699));
    outputs(1050) <= (layer0_outputs(8617)) and (layer0_outputs(6475));
    outputs(1051) <= layer0_outputs(263);
    outputs(1052) <= (layer0_outputs(9565)) and not (layer0_outputs(6848));
    outputs(1053) <= (layer0_outputs(5963)) xor (layer0_outputs(7919));
    outputs(1054) <= not(layer0_outputs(7331));
    outputs(1055) <= layer0_outputs(9246);
    outputs(1056) <= not((layer0_outputs(4411)) xor (layer0_outputs(5045)));
    outputs(1057) <= (layer0_outputs(9956)) and not (layer0_outputs(3812));
    outputs(1058) <= not((layer0_outputs(1617)) xor (layer0_outputs(2195)));
    outputs(1059) <= (layer0_outputs(2837)) and (layer0_outputs(6504));
    outputs(1060) <= (layer0_outputs(1476)) and (layer0_outputs(6580));
    outputs(1061) <= not(layer0_outputs(2015));
    outputs(1062) <= (layer0_outputs(7359)) and (layer0_outputs(1228));
    outputs(1063) <= (layer0_outputs(7564)) and not (layer0_outputs(10223));
    outputs(1064) <= (layer0_outputs(1328)) and not (layer0_outputs(9587));
    outputs(1065) <= (layer0_outputs(6503)) and not (layer0_outputs(5207));
    outputs(1066) <= not((layer0_outputs(1192)) or (layer0_outputs(4779)));
    outputs(1067) <= (layer0_outputs(676)) and not (layer0_outputs(10066));
    outputs(1068) <= (layer0_outputs(5391)) and not (layer0_outputs(7035));
    outputs(1069) <= (layer0_outputs(796)) xor (layer0_outputs(784));
    outputs(1070) <= (layer0_outputs(3154)) and not (layer0_outputs(8788));
    outputs(1071) <= not(layer0_outputs(4393));
    outputs(1072) <= not((layer0_outputs(517)) xor (layer0_outputs(2696)));
    outputs(1073) <= layer0_outputs(9398);
    outputs(1074) <= not(layer0_outputs(8095));
    outputs(1075) <= not((layer0_outputs(4255)) or (layer0_outputs(835)));
    outputs(1076) <= not(layer0_outputs(1916));
    outputs(1077) <= (layer0_outputs(10090)) and (layer0_outputs(9717));
    outputs(1078) <= (layer0_outputs(1649)) and not (layer0_outputs(6731));
    outputs(1079) <= layer0_outputs(2756);
    outputs(1080) <= not(layer0_outputs(2292));
    outputs(1081) <= not(layer0_outputs(4908)) or (layer0_outputs(5712));
    outputs(1082) <= (layer0_outputs(9765)) and (layer0_outputs(6695));
    outputs(1083) <= not((layer0_outputs(2476)) xor (layer0_outputs(1273)));
    outputs(1084) <= not((layer0_outputs(862)) or (layer0_outputs(4213)));
    outputs(1085) <= (layer0_outputs(9727)) and not (layer0_outputs(1078));
    outputs(1086) <= layer0_outputs(8968);
    outputs(1087) <= (layer0_outputs(9488)) and (layer0_outputs(8291));
    outputs(1088) <= (layer0_outputs(2089)) and (layer0_outputs(1880));
    outputs(1089) <= not((layer0_outputs(4967)) or (layer0_outputs(9895)));
    outputs(1090) <= not((layer0_outputs(5515)) xor (layer0_outputs(7684)));
    outputs(1091) <= (layer0_outputs(5899)) xor (layer0_outputs(6867));
    outputs(1092) <= (layer0_outputs(2231)) and not (layer0_outputs(5830));
    outputs(1093) <= (layer0_outputs(7938)) and not (layer0_outputs(10161));
    outputs(1094) <= not(layer0_outputs(2113));
    outputs(1095) <= (layer0_outputs(171)) xor (layer0_outputs(4427));
    outputs(1096) <= layer0_outputs(2507);
    outputs(1097) <= not((layer0_outputs(8372)) xor (layer0_outputs(7523)));
    outputs(1098) <= not((layer0_outputs(8336)) or (layer0_outputs(4855)));
    outputs(1099) <= layer0_outputs(7083);
    outputs(1100) <= layer0_outputs(6537);
    outputs(1101) <= not((layer0_outputs(266)) or (layer0_outputs(8137)));
    outputs(1102) <= (layer0_outputs(6668)) and not (layer0_outputs(1706));
    outputs(1103) <= (layer0_outputs(1220)) xor (layer0_outputs(1272));
    outputs(1104) <= not((layer0_outputs(4369)) or (layer0_outputs(7769)));
    outputs(1105) <= (layer0_outputs(5114)) and not (layer0_outputs(6431));
    outputs(1106) <= not((layer0_outputs(9473)) or (layer0_outputs(7355)));
    outputs(1107) <= (layer0_outputs(6785)) and (layer0_outputs(6933));
    outputs(1108) <= not((layer0_outputs(1980)) or (layer0_outputs(304)));
    outputs(1109) <= not((layer0_outputs(1984)) xor (layer0_outputs(6663)));
    outputs(1110) <= (layer0_outputs(5138)) xor (layer0_outputs(462));
    outputs(1111) <= not((layer0_outputs(2)) xor (layer0_outputs(7520)));
    outputs(1112) <= layer0_outputs(7796);
    outputs(1113) <= (layer0_outputs(6523)) and (layer0_outputs(7410));
    outputs(1114) <= layer0_outputs(2676);
    outputs(1115) <= not((layer0_outputs(9424)) xor (layer0_outputs(3982)));
    outputs(1116) <= not((layer0_outputs(538)) xor (layer0_outputs(8010)));
    outputs(1117) <= (layer0_outputs(6808)) and not (layer0_outputs(2835));
    outputs(1118) <= (layer0_outputs(2234)) and (layer0_outputs(2014));
    outputs(1119) <= (layer0_outputs(2250)) xor (layer0_outputs(7026));
    outputs(1120) <= (layer0_outputs(4086)) and not (layer0_outputs(3140));
    outputs(1121) <= not((layer0_outputs(4973)) xor (layer0_outputs(2834)));
    outputs(1122) <= (layer0_outputs(4598)) xor (layer0_outputs(535));
    outputs(1123) <= not((layer0_outputs(2750)) xor (layer0_outputs(4168)));
    outputs(1124) <= not((layer0_outputs(6640)) and (layer0_outputs(8548)));
    outputs(1125) <= layer0_outputs(8168);
    outputs(1126) <= not((layer0_outputs(2330)) or (layer0_outputs(10198)));
    outputs(1127) <= layer0_outputs(1735);
    outputs(1128) <= not((layer0_outputs(9363)) xor (layer0_outputs(3273)));
    outputs(1129) <= (layer0_outputs(8139)) and not (layer0_outputs(5817));
    outputs(1130) <= layer0_outputs(4568);
    outputs(1131) <= not((layer0_outputs(8130)) or (layer0_outputs(9194)));
    outputs(1132) <= not((layer0_outputs(8803)) or (layer0_outputs(2434)));
    outputs(1133) <= (layer0_outputs(288)) and (layer0_outputs(5935));
    outputs(1134) <= (layer0_outputs(7323)) xor (layer0_outputs(9713));
    outputs(1135) <= (layer0_outputs(7320)) xor (layer0_outputs(1630));
    outputs(1136) <= layer0_outputs(4036);
    outputs(1137) <= (layer0_outputs(161)) and (layer0_outputs(173));
    outputs(1138) <= not((layer0_outputs(2690)) xor (layer0_outputs(1842)));
    outputs(1139) <= (layer0_outputs(8735)) xor (layer0_outputs(6401));
    outputs(1140) <= not((layer0_outputs(2327)) or (layer0_outputs(4755)));
    outputs(1141) <= (layer0_outputs(2912)) and (layer0_outputs(1092));
    outputs(1142) <= (layer0_outputs(3833)) and not (layer0_outputs(1214));
    outputs(1143) <= layer0_outputs(7693);
    outputs(1144) <= (layer0_outputs(2821)) and (layer0_outputs(4356));
    outputs(1145) <= not((layer0_outputs(628)) xor (layer0_outputs(2600)));
    outputs(1146) <= (layer0_outputs(5351)) xor (layer0_outputs(8801));
    outputs(1147) <= (layer0_outputs(5791)) and (layer0_outputs(8728));
    outputs(1148) <= not((layer0_outputs(9975)) xor (layer0_outputs(5669)));
    outputs(1149) <= (layer0_outputs(9287)) xor (layer0_outputs(1715));
    outputs(1150) <= not(layer0_outputs(1625));
    outputs(1151) <= not((layer0_outputs(9912)) xor (layer0_outputs(5713)));
    outputs(1152) <= (layer0_outputs(119)) and (layer0_outputs(8048));
    outputs(1153) <= (layer0_outputs(574)) and (layer0_outputs(6720));
    outputs(1154) <= (layer0_outputs(2566)) and not (layer0_outputs(10196));
    outputs(1155) <= (layer0_outputs(10191)) and not (layer0_outputs(663));
    outputs(1156) <= not(layer0_outputs(3324));
    outputs(1157) <= not((layer0_outputs(8475)) xor (layer0_outputs(4880)));
    outputs(1158) <= layer0_outputs(10152);
    outputs(1159) <= not(layer0_outputs(3222));
    outputs(1160) <= not((layer0_outputs(3592)) xor (layer0_outputs(4125)));
    outputs(1161) <= (layer0_outputs(1260)) and (layer0_outputs(6974));
    outputs(1162) <= (layer0_outputs(8374)) xor (layer0_outputs(3875));
    outputs(1163) <= (layer0_outputs(9740)) or (layer0_outputs(1405));
    outputs(1164) <= not((layer0_outputs(8812)) or (layer0_outputs(5584)));
    outputs(1165) <= layer0_outputs(6415);
    outputs(1166) <= (layer0_outputs(640)) xor (layer0_outputs(8818));
    outputs(1167) <= (layer0_outputs(7955)) and not (layer0_outputs(8159));
    outputs(1168) <= not(layer0_outputs(4384));
    outputs(1169) <= not(layer0_outputs(3100));
    outputs(1170) <= (layer0_outputs(5773)) and not (layer0_outputs(515));
    outputs(1171) <= not((layer0_outputs(4314)) xor (layer0_outputs(8598)));
    outputs(1172) <= (layer0_outputs(597)) and (layer0_outputs(3345));
    outputs(1173) <= (layer0_outputs(8871)) and not (layer0_outputs(9922));
    outputs(1174) <= not(layer0_outputs(9161));
    outputs(1175) <= (layer0_outputs(738)) and not (layer0_outputs(10236));
    outputs(1176) <= (layer0_outputs(9983)) and (layer0_outputs(3529));
    outputs(1177) <= not(layer0_outputs(1281));
    outputs(1178) <= not((layer0_outputs(2140)) xor (layer0_outputs(1492)));
    outputs(1179) <= not((layer0_outputs(6184)) or (layer0_outputs(8252)));
    outputs(1180) <= (layer0_outputs(9035)) and not (layer0_outputs(7774));
    outputs(1181) <= not(layer0_outputs(7816));
    outputs(1182) <= (layer0_outputs(857)) and not (layer0_outputs(3085));
    outputs(1183) <= (layer0_outputs(3720)) xor (layer0_outputs(10221));
    outputs(1184) <= (layer0_outputs(1023)) and not (layer0_outputs(7997));
    outputs(1185) <= (layer0_outputs(9493)) and not (layer0_outputs(10179));
    outputs(1186) <= (layer0_outputs(2779)) and (layer0_outputs(9690));
    outputs(1187) <= not(layer0_outputs(2703));
    outputs(1188) <= '0';
    outputs(1189) <= (layer0_outputs(9819)) xor (layer0_outputs(987));
    outputs(1190) <= layer0_outputs(7350);
    outputs(1191) <= (layer0_outputs(7626)) and not (layer0_outputs(1813));
    outputs(1192) <= (layer0_outputs(662)) and (layer0_outputs(4748));
    outputs(1193) <= (layer0_outputs(5114)) and (layer0_outputs(8291));
    outputs(1194) <= layer0_outputs(9072);
    outputs(1195) <= (layer0_outputs(9328)) and (layer0_outputs(8036));
    outputs(1196) <= layer0_outputs(7030);
    outputs(1197) <= not((layer0_outputs(2175)) xor (layer0_outputs(9414)));
    outputs(1198) <= (layer0_outputs(9748)) xor (layer0_outputs(8554));
    outputs(1199) <= (layer0_outputs(929)) and not (layer0_outputs(5920));
    outputs(1200) <= not(layer0_outputs(678));
    outputs(1201) <= not(layer0_outputs(6613));
    outputs(1202) <= layer0_outputs(4054);
    outputs(1203) <= (layer0_outputs(2390)) and not (layer0_outputs(8685));
    outputs(1204) <= not((layer0_outputs(9876)) xor (layer0_outputs(7024)));
    outputs(1205) <= not((layer0_outputs(4871)) xor (layer0_outputs(44)));
    outputs(1206) <= not(layer0_outputs(9196));
    outputs(1207) <= (layer0_outputs(8339)) xor (layer0_outputs(587));
    outputs(1208) <= (layer0_outputs(2445)) and not (layer0_outputs(9921));
    outputs(1209) <= (layer0_outputs(8135)) and not (layer0_outputs(114));
    outputs(1210) <= not(layer0_outputs(8656));
    outputs(1211) <= layer0_outputs(4296);
    outputs(1212) <= not(layer0_outputs(4937));
    outputs(1213) <= (layer0_outputs(9986)) and not (layer0_outputs(3606));
    outputs(1214) <= not(layer0_outputs(7476));
    outputs(1215) <= not(layer0_outputs(9458));
    outputs(1216) <= not(layer0_outputs(7759));
    outputs(1217) <= (layer0_outputs(589)) and (layer0_outputs(3174));
    outputs(1218) <= not((layer0_outputs(146)) or (layer0_outputs(7115)));
    outputs(1219) <= not((layer0_outputs(4076)) or (layer0_outputs(8503)));
    outputs(1220) <= (layer0_outputs(2457)) and not (layer0_outputs(5223));
    outputs(1221) <= (layer0_outputs(7532)) and (layer0_outputs(9489));
    outputs(1222) <= (layer0_outputs(7459)) and not (layer0_outputs(5942));
    outputs(1223) <= layer0_outputs(2335);
    outputs(1224) <= not(layer0_outputs(6764));
    outputs(1225) <= not((layer0_outputs(3554)) xor (layer0_outputs(6646)));
    outputs(1226) <= '0';
    outputs(1227) <= not((layer0_outputs(3904)) or (layer0_outputs(6647)));
    outputs(1228) <= not((layer0_outputs(6018)) or (layer0_outputs(9026)));
    outputs(1229) <= (layer0_outputs(6174)) and not (layer0_outputs(10064));
    outputs(1230) <= not((layer0_outputs(6722)) or (layer0_outputs(3208)));
    outputs(1231) <= (layer0_outputs(6795)) xor (layer0_outputs(5929));
    outputs(1232) <= (layer0_outputs(7225)) and not (layer0_outputs(1670));
    outputs(1233) <= not(layer0_outputs(8676));
    outputs(1234) <= not((layer0_outputs(2109)) or (layer0_outputs(7762)));
    outputs(1235) <= not(layer0_outputs(5762));
    outputs(1236) <= (layer0_outputs(10092)) and not (layer0_outputs(5473));
    outputs(1237) <= not((layer0_outputs(7689)) or (layer0_outputs(8597)));
    outputs(1238) <= (layer0_outputs(5720)) and not (layer0_outputs(7151));
    outputs(1239) <= not((layer0_outputs(6996)) xor (layer0_outputs(6445)));
    outputs(1240) <= (layer0_outputs(4443)) and not (layer0_outputs(8380));
    outputs(1241) <= layer0_outputs(2428);
    outputs(1242) <= not(layer0_outputs(2005));
    outputs(1243) <= layer0_outputs(7250);
    outputs(1244) <= (layer0_outputs(7154)) xor (layer0_outputs(8023));
    outputs(1245) <= layer0_outputs(6834);
    outputs(1246) <= '0';
    outputs(1247) <= (layer0_outputs(7333)) and (layer0_outputs(9979));
    outputs(1248) <= not(layer0_outputs(5955));
    outputs(1249) <= layer0_outputs(813);
    outputs(1250) <= not((layer0_outputs(5707)) or (layer0_outputs(1418)));
    outputs(1251) <= (layer0_outputs(9589)) xor (layer0_outputs(6183));
    outputs(1252) <= layer0_outputs(6866);
    outputs(1253) <= not(layer0_outputs(3572));
    outputs(1254) <= (layer0_outputs(1729)) and not (layer0_outputs(7248));
    outputs(1255) <= (layer0_outputs(7943)) and not (layer0_outputs(9540));
    outputs(1256) <= (layer0_outputs(6202)) and (layer0_outputs(2218));
    outputs(1257) <= layer0_outputs(4820);
    outputs(1258) <= (layer0_outputs(1495)) and (layer0_outputs(3470));
    outputs(1259) <= not(layer0_outputs(1806));
    outputs(1260) <= (layer0_outputs(2248)) and not (layer0_outputs(2327));
    outputs(1261) <= not((layer0_outputs(3031)) xor (layer0_outputs(4346)));
    outputs(1262) <= not((layer0_outputs(2778)) or (layer0_outputs(2583)));
    outputs(1263) <= not(layer0_outputs(720));
    outputs(1264) <= (layer0_outputs(6345)) xor (layer0_outputs(9398));
    outputs(1265) <= (layer0_outputs(8306)) xor (layer0_outputs(9935));
    outputs(1266) <= (layer0_outputs(8350)) and not (layer0_outputs(1237));
    outputs(1267) <= (layer0_outputs(4627)) and not (layer0_outputs(9849));
    outputs(1268) <= not((layer0_outputs(6592)) xor (layer0_outputs(5570)));
    outputs(1269) <= (layer0_outputs(1533)) and (layer0_outputs(4530));
    outputs(1270) <= (layer0_outputs(5512)) xor (layer0_outputs(911));
    outputs(1271) <= not(layer0_outputs(10157));
    outputs(1272) <= layer0_outputs(8123);
    outputs(1273) <= not((layer0_outputs(5989)) or (layer0_outputs(652)));
    outputs(1274) <= not(layer0_outputs(5289));
    outputs(1275) <= (layer0_outputs(3944)) and not (layer0_outputs(8638));
    outputs(1276) <= not(layer0_outputs(7129)) or (layer0_outputs(957));
    outputs(1277) <= not((layer0_outputs(5728)) xor (layer0_outputs(9491)));
    outputs(1278) <= not((layer0_outputs(6284)) or (layer0_outputs(6151)));
    outputs(1279) <= not((layer0_outputs(2287)) or (layer0_outputs(8408)));
    outputs(1280) <= not((layer0_outputs(3173)) xor (layer0_outputs(9522)));
    outputs(1281) <= (layer0_outputs(727)) xor (layer0_outputs(4154));
    outputs(1282) <= layer0_outputs(1077);
    outputs(1283) <= (layer0_outputs(3391)) xor (layer0_outputs(1032));
    outputs(1284) <= (layer0_outputs(1821)) and not (layer0_outputs(6675));
    outputs(1285) <= (layer0_outputs(794)) xor (layer0_outputs(3087));
    outputs(1286) <= not(layer0_outputs(5871));
    outputs(1287) <= (layer0_outputs(2659)) and (layer0_outputs(8118));
    outputs(1288) <= not(layer0_outputs(7023));
    outputs(1289) <= not((layer0_outputs(2365)) xor (layer0_outputs(5992)));
    outputs(1290) <= not(layer0_outputs(4061));
    outputs(1291) <= (layer0_outputs(6254)) xor (layer0_outputs(5864));
    outputs(1292) <= not(layer0_outputs(4371));
    outputs(1293) <= not((layer0_outputs(2052)) xor (layer0_outputs(4905)));
    outputs(1294) <= not(layer0_outputs(8826));
    outputs(1295) <= not((layer0_outputs(9049)) or (layer0_outputs(2874)));
    outputs(1296) <= not(layer0_outputs(2437));
    outputs(1297) <= (layer0_outputs(6064)) and (layer0_outputs(4442));
    outputs(1298) <= layer0_outputs(7716);
    outputs(1299) <= (layer0_outputs(2196)) and (layer0_outputs(3644));
    outputs(1300) <= (layer0_outputs(6678)) and not (layer0_outputs(4401));
    outputs(1301) <= (layer0_outputs(9165)) xor (layer0_outputs(725));
    outputs(1302) <= (layer0_outputs(8814)) and not (layer0_outputs(9272));
    outputs(1303) <= not(layer0_outputs(8611));
    outputs(1304) <= (layer0_outputs(3303)) and not (layer0_outputs(1958));
    outputs(1305) <= not((layer0_outputs(740)) xor (layer0_outputs(6442)));
    outputs(1306) <= (layer0_outputs(5110)) and not (layer0_outputs(6331));
    outputs(1307) <= not(layer0_outputs(9546));
    outputs(1308) <= (layer0_outputs(7199)) and not (layer0_outputs(8693));
    outputs(1309) <= not((layer0_outputs(5897)) xor (layer0_outputs(5208)));
    outputs(1310) <= layer0_outputs(4517);
    outputs(1311) <= not((layer0_outputs(302)) or (layer0_outputs(6587)));
    outputs(1312) <= (layer0_outputs(8346)) xor (layer0_outputs(8459));
    outputs(1313) <= (layer0_outputs(1612)) xor (layer0_outputs(5892));
    outputs(1314) <= (layer0_outputs(722)) and not (layer0_outputs(9258));
    outputs(1315) <= (layer0_outputs(9344)) and (layer0_outputs(1687));
    outputs(1316) <= layer0_outputs(4969);
    outputs(1317) <= not((layer0_outputs(5355)) xor (layer0_outputs(7037)));
    outputs(1318) <= not((layer0_outputs(8798)) or (layer0_outputs(5173)));
    outputs(1319) <= (layer0_outputs(7238)) xor (layer0_outputs(2119));
    outputs(1320) <= (layer0_outputs(2770)) and (layer0_outputs(9421));
    outputs(1321) <= (layer0_outputs(606)) xor (layer0_outputs(3075));
    outputs(1322) <= (layer0_outputs(1726)) and (layer0_outputs(10079));
    outputs(1323) <= (layer0_outputs(3097)) and (layer0_outputs(8289));
    outputs(1324) <= layer0_outputs(8981);
    outputs(1325) <= (layer0_outputs(10133)) xor (layer0_outputs(1350));
    outputs(1326) <= (layer0_outputs(981)) xor (layer0_outputs(8678));
    outputs(1327) <= layer0_outputs(1656);
    outputs(1328) <= (layer0_outputs(1137)) xor (layer0_outputs(3146));
    outputs(1329) <= layer0_outputs(8306);
    outputs(1330) <= (layer0_outputs(6629)) xor (layer0_outputs(2564));
    outputs(1331) <= (layer0_outputs(5345)) and not (layer0_outputs(4674));
    outputs(1332) <= (layer0_outputs(6883)) and not (layer0_outputs(8610));
    outputs(1333) <= layer0_outputs(731);
    outputs(1334) <= not((layer0_outputs(6625)) or (layer0_outputs(8357)));
    outputs(1335) <= (layer0_outputs(2744)) and (layer0_outputs(4534));
    outputs(1336) <= layer0_outputs(6858);
    outputs(1337) <= (layer0_outputs(4588)) and (layer0_outputs(337));
    outputs(1338) <= (layer0_outputs(2714)) and (layer0_outputs(5414));
    outputs(1339) <= layer0_outputs(8271);
    outputs(1340) <= (layer0_outputs(1619)) xor (layer0_outputs(1343));
    outputs(1341) <= not((layer0_outputs(2565)) xor (layer0_outputs(6412)));
    outputs(1342) <= not((layer0_outputs(434)) xor (layer0_outputs(5076)));
    outputs(1343) <= layer0_outputs(7704);
    outputs(1344) <= (layer0_outputs(4166)) xor (layer0_outputs(7901));
    outputs(1345) <= (layer0_outputs(228)) xor (layer0_outputs(1109));
    outputs(1346) <= (layer0_outputs(7475)) and not (layer0_outputs(3516));
    outputs(1347) <= not((layer0_outputs(3664)) or (layer0_outputs(5478)));
    outputs(1348) <= (layer0_outputs(2991)) and (layer0_outputs(4447));
    outputs(1349) <= (layer0_outputs(1930)) and not (layer0_outputs(6387));
    outputs(1350) <= not(layer0_outputs(6163));
    outputs(1351) <= (layer0_outputs(1000)) xor (layer0_outputs(4274));
    outputs(1352) <= not((layer0_outputs(1057)) and (layer0_outputs(8669)));
    outputs(1353) <= (layer0_outputs(3653)) xor (layer0_outputs(9259));
    outputs(1354) <= not(layer0_outputs(1188));
    outputs(1355) <= (layer0_outputs(5254)) and not (layer0_outputs(4041));
    outputs(1356) <= (layer0_outputs(9215)) and not (layer0_outputs(7136));
    outputs(1357) <= (layer0_outputs(3716)) and not (layer0_outputs(946));
    outputs(1358) <= layer0_outputs(9768);
    outputs(1359) <= (layer0_outputs(9024)) xor (layer0_outputs(4422));
    outputs(1360) <= not((layer0_outputs(5103)) xor (layer0_outputs(4416)));
    outputs(1361) <= layer0_outputs(1964);
    outputs(1362) <= not((layer0_outputs(4173)) xor (layer0_outputs(1356)));
    outputs(1363) <= (layer0_outputs(4970)) xor (layer0_outputs(9864));
    outputs(1364) <= (layer0_outputs(7299)) and not (layer0_outputs(1054));
    outputs(1365) <= not((layer0_outputs(4309)) or (layer0_outputs(7600)));
    outputs(1366) <= not((layer0_outputs(6540)) or (layer0_outputs(7931)));
    outputs(1367) <= (layer0_outputs(2716)) xor (layer0_outputs(5860));
    outputs(1368) <= (layer0_outputs(8204)) and not (layer0_outputs(8255));
    outputs(1369) <= layer0_outputs(6899);
    outputs(1370) <= (layer0_outputs(7541)) and not (layer0_outputs(5776));
    outputs(1371) <= (layer0_outputs(10070)) xor (layer0_outputs(3037));
    outputs(1372) <= not((layer0_outputs(2983)) or (layer0_outputs(1499)));
    outputs(1373) <= (layer0_outputs(6071)) xor (layer0_outputs(113));
    outputs(1374) <= not(layer0_outputs(7974));
    outputs(1375) <= (layer0_outputs(9534)) and not (layer0_outputs(7485));
    outputs(1376) <= layer0_outputs(6900);
    outputs(1377) <= '0';
    outputs(1378) <= (layer0_outputs(9118)) and not (layer0_outputs(4975));
    outputs(1379) <= layer0_outputs(3301);
    outputs(1380) <= (layer0_outputs(9397)) and not (layer0_outputs(1565));
    outputs(1381) <= not(layer0_outputs(575));
    outputs(1382) <= layer0_outputs(3979);
    outputs(1383) <= (layer0_outputs(7641)) or (layer0_outputs(3556));
    outputs(1384) <= (layer0_outputs(2711)) xor (layer0_outputs(2164));
    outputs(1385) <= (layer0_outputs(6474)) and not (layer0_outputs(10167));
    outputs(1386) <= (layer0_outputs(9241)) and not (layer0_outputs(390));
    outputs(1387) <= layer0_outputs(3472);
    outputs(1388) <= (layer0_outputs(2740)) and (layer0_outputs(3165));
    outputs(1389) <= (layer0_outputs(2896)) and (layer0_outputs(3421));
    outputs(1390) <= (layer0_outputs(3815)) and not (layer0_outputs(7456));
    outputs(1391) <= (layer0_outputs(6507)) and not (layer0_outputs(6231));
    outputs(1392) <= (layer0_outputs(8837)) and not (layer0_outputs(1326));
    outputs(1393) <= (layer0_outputs(2652)) and (layer0_outputs(9030));
    outputs(1394) <= (layer0_outputs(6801)) and (layer0_outputs(6260));
    outputs(1395) <= (layer0_outputs(1623)) and (layer0_outputs(8504));
    outputs(1396) <= layer0_outputs(4866);
    outputs(1397) <= not(layer0_outputs(6254));
    outputs(1398) <= (layer0_outputs(6593)) and not (layer0_outputs(8896));
    outputs(1399) <= layer0_outputs(1005);
    outputs(1400) <= (layer0_outputs(2622)) xor (layer0_outputs(9578));
    outputs(1401) <= (layer0_outputs(5206)) and not (layer0_outputs(3904));
    outputs(1402) <= (layer0_outputs(5453)) and not (layer0_outputs(5247));
    outputs(1403) <= layer0_outputs(8174);
    outputs(1404) <= not((layer0_outputs(342)) xor (layer0_outputs(6773)));
    outputs(1405) <= not((layer0_outputs(7804)) xor (layer0_outputs(5487)));
    outputs(1406) <= not((layer0_outputs(1120)) or (layer0_outputs(8219)));
    outputs(1407) <= (layer0_outputs(7630)) xor (layer0_outputs(6015));
    outputs(1408) <= (layer0_outputs(4075)) xor (layer0_outputs(7484));
    outputs(1409) <= (layer0_outputs(9832)) and not (layer0_outputs(2937));
    outputs(1410) <= not((layer0_outputs(7663)) xor (layer0_outputs(9111)));
    outputs(1411) <= (layer0_outputs(3810)) xor (layer0_outputs(3394));
    outputs(1412) <= not(layer0_outputs(3652));
    outputs(1413) <= (layer0_outputs(1449)) and (layer0_outputs(2402));
    outputs(1414) <= layer0_outputs(6776);
    outputs(1415) <= (layer0_outputs(10029)) and not (layer0_outputs(7187));
    outputs(1416) <= (layer0_outputs(9500)) and not (layer0_outputs(2311));
    outputs(1417) <= (layer0_outputs(7051)) xor (layer0_outputs(1880));
    outputs(1418) <= (layer0_outputs(9247)) and not (layer0_outputs(3686));
    outputs(1419) <= (layer0_outputs(1272)) and (layer0_outputs(2021));
    outputs(1420) <= (layer0_outputs(3902)) and (layer0_outputs(5987));
    outputs(1421) <= layer0_outputs(6411);
    outputs(1422) <= not((layer0_outputs(2328)) xor (layer0_outputs(1862)));
    outputs(1423) <= (layer0_outputs(5572)) and not (layer0_outputs(3256));
    outputs(1424) <= (layer0_outputs(213)) and not (layer0_outputs(8625));
    outputs(1425) <= (layer0_outputs(7560)) and not (layer0_outputs(2902));
    outputs(1426) <= (layer0_outputs(3331)) and not (layer0_outputs(5330));
    outputs(1427) <= (layer0_outputs(9040)) and not (layer0_outputs(5260));
    outputs(1428) <= not((layer0_outputs(7828)) or (layer0_outputs(6489)));
    outputs(1429) <= (layer0_outputs(2333)) and not (layer0_outputs(3742));
    outputs(1430) <= (layer0_outputs(5758)) xor (layer0_outputs(1089));
    outputs(1431) <= (layer0_outputs(3495)) and not (layer0_outputs(160));
    outputs(1432) <= not(layer0_outputs(9857));
    outputs(1433) <= (layer0_outputs(7863)) and not (layer0_outputs(4972));
    outputs(1434) <= layer0_outputs(919);
    outputs(1435) <= layer0_outputs(9870);
    outputs(1436) <= (layer0_outputs(2773)) xor (layer0_outputs(1683));
    outputs(1437) <= (layer0_outputs(4428)) xor (layer0_outputs(5193));
    outputs(1438) <= (layer0_outputs(3153)) and not (layer0_outputs(9187));
    outputs(1439) <= not((layer0_outputs(9454)) or (layer0_outputs(939)));
    outputs(1440) <= (layer0_outputs(8384)) and not (layer0_outputs(2108));
    outputs(1441) <= not((layer0_outputs(5980)) or (layer0_outputs(8176)));
    outputs(1442) <= (layer0_outputs(2235)) xor (layer0_outputs(3471));
    outputs(1443) <= (layer0_outputs(3525)) and not (layer0_outputs(2077));
    outputs(1444) <= not((layer0_outputs(6153)) xor (layer0_outputs(6274)));
    outputs(1445) <= layer0_outputs(2212);
    outputs(1446) <= (layer0_outputs(9334)) and not (layer0_outputs(10151));
    outputs(1447) <= (layer0_outputs(1269)) xor (layer0_outputs(7844));
    outputs(1448) <= not((layer0_outputs(9958)) or (layer0_outputs(9107)));
    outputs(1449) <= (layer0_outputs(8474)) and (layer0_outputs(6591));
    outputs(1450) <= not((layer0_outputs(1336)) xor (layer0_outputs(8049)));
    outputs(1451) <= layer0_outputs(7309);
    outputs(1452) <= layer0_outputs(3925);
    outputs(1453) <= (layer0_outputs(5148)) and (layer0_outputs(6197));
    outputs(1454) <= (layer0_outputs(563)) and not (layer0_outputs(4342));
    outputs(1455) <= not(layer0_outputs(9054));
    outputs(1456) <= not((layer0_outputs(9182)) or (layer0_outputs(1085)));
    outputs(1457) <= (layer0_outputs(283)) and not (layer0_outputs(189));
    outputs(1458) <= layer0_outputs(3226);
    outputs(1459) <= not((layer0_outputs(5128)) xor (layer0_outputs(1752)));
    outputs(1460) <= not(layer0_outputs(8522));
    outputs(1461) <= not((layer0_outputs(7702)) xor (layer0_outputs(1236)));
    outputs(1462) <= (layer0_outputs(3484)) and (layer0_outputs(5787));
    outputs(1463) <= (layer0_outputs(6601)) and not (layer0_outputs(6123));
    outputs(1464) <= not((layer0_outputs(4592)) xor (layer0_outputs(7496)));
    outputs(1465) <= not((layer0_outputs(4583)) or (layer0_outputs(439)));
    outputs(1466) <= not((layer0_outputs(5887)) xor (layer0_outputs(1950)));
    outputs(1467) <= (layer0_outputs(8712)) xor (layer0_outputs(6543));
    outputs(1468) <= (layer0_outputs(6982)) and (layer0_outputs(5336));
    outputs(1469) <= layer0_outputs(4267);
    outputs(1470) <= (layer0_outputs(5337)) xor (layer0_outputs(2055));
    outputs(1471) <= not((layer0_outputs(9515)) xor (layer0_outputs(4676)));
    outputs(1472) <= '0';
    outputs(1473) <= (layer0_outputs(3930)) and not (layer0_outputs(834));
    outputs(1474) <= layer0_outputs(7339);
    outputs(1475) <= not((layer0_outputs(7960)) xor (layer0_outputs(9605)));
    outputs(1476) <= (layer0_outputs(8518)) and not (layer0_outputs(6037));
    outputs(1477) <= not(layer0_outputs(4983));
    outputs(1478) <= layer0_outputs(1358);
    outputs(1479) <= (layer0_outputs(9440)) and not (layer0_outputs(7478));
    outputs(1480) <= (layer0_outputs(9344)) xor (layer0_outputs(9142));
    outputs(1481) <= (layer0_outputs(10009)) and not (layer0_outputs(1676));
    outputs(1482) <= (layer0_outputs(6576)) and not (layer0_outputs(6120));
    outputs(1483) <= layer0_outputs(6749);
    outputs(1484) <= (layer0_outputs(6423)) and not (layer0_outputs(7263));
    outputs(1485) <= (layer0_outputs(827)) and not (layer0_outputs(6135));
    outputs(1486) <= not((layer0_outputs(1133)) or (layer0_outputs(9618)));
    outputs(1487) <= (layer0_outputs(960)) xor (layer0_outputs(8315));
    outputs(1488) <= (layer0_outputs(5243)) and not (layer0_outputs(3011));
    outputs(1489) <= (layer0_outputs(5371)) and (layer0_outputs(5433));
    outputs(1490) <= layer0_outputs(5183);
    outputs(1491) <= not((layer0_outputs(1375)) or (layer0_outputs(6401)));
    outputs(1492) <= (layer0_outputs(5841)) xor (layer0_outputs(2465));
    outputs(1493) <= not((layer0_outputs(2433)) xor (layer0_outputs(8840)));
    outputs(1494) <= not((layer0_outputs(7955)) xor (layer0_outputs(8929)));
    outputs(1495) <= (layer0_outputs(6092)) and (layer0_outputs(2312));
    outputs(1496) <= (layer0_outputs(1906)) and not (layer0_outputs(7643));
    outputs(1497) <= not((layer0_outputs(3989)) xor (layer0_outputs(5627)));
    outputs(1498) <= (layer0_outputs(1723)) xor (layer0_outputs(1313));
    outputs(1499) <= (layer0_outputs(9956)) and (layer0_outputs(5481));
    outputs(1500) <= not((layer0_outputs(135)) and (layer0_outputs(9784)));
    outputs(1501) <= not((layer0_outputs(3753)) xor (layer0_outputs(2830)));
    outputs(1502) <= (layer0_outputs(8793)) xor (layer0_outputs(5242));
    outputs(1503) <= (layer0_outputs(6828)) and not (layer0_outputs(5862));
    outputs(1504) <= (layer0_outputs(4353)) and not (layer0_outputs(1010));
    outputs(1505) <= not((layer0_outputs(2099)) or (layer0_outputs(5654)));
    outputs(1506) <= not((layer0_outputs(6607)) or (layer0_outputs(782)));
    outputs(1507) <= not(layer0_outputs(4710));
    outputs(1508) <= not((layer0_outputs(2595)) or (layer0_outputs(190)));
    outputs(1509) <= not((layer0_outputs(9449)) xor (layer0_outputs(1558)));
    outputs(1510) <= (layer0_outputs(4513)) and (layer0_outputs(9401));
    outputs(1511) <= (layer0_outputs(3605)) xor (layer0_outputs(1292));
    outputs(1512) <= (layer0_outputs(2011)) and not (layer0_outputs(8511));
    outputs(1513) <= (layer0_outputs(5608)) and (layer0_outputs(9490));
    outputs(1514) <= (layer0_outputs(9704)) and (layer0_outputs(9747));
    outputs(1515) <= (layer0_outputs(7399)) xor (layer0_outputs(5056));
    outputs(1516) <= not((layer0_outputs(9678)) xor (layer0_outputs(7109)));
    outputs(1517) <= (layer0_outputs(4200)) xor (layer0_outputs(3965));
    outputs(1518) <= not((layer0_outputs(5049)) or (layer0_outputs(3544)));
    outputs(1519) <= (layer0_outputs(2842)) and not (layer0_outputs(142));
    outputs(1520) <= (layer0_outputs(4134)) and (layer0_outputs(8447));
    outputs(1521) <= (layer0_outputs(4053)) and (layer0_outputs(2710));
    outputs(1522) <= layer0_outputs(6258);
    outputs(1523) <= (layer0_outputs(4437)) xor (layer0_outputs(1633));
    outputs(1524) <= '0';
    outputs(1525) <= not((layer0_outputs(4406)) or (layer0_outputs(9304)));
    outputs(1526) <= not((layer0_outputs(1878)) xor (layer0_outputs(1642)));
    outputs(1527) <= not((layer0_outputs(5586)) xor (layer0_outputs(5394)));
    outputs(1528) <= layer0_outputs(1793);
    outputs(1529) <= (layer0_outputs(7260)) and (layer0_outputs(1009));
    outputs(1530) <= not((layer0_outputs(6983)) xor (layer0_outputs(146)));
    outputs(1531) <= (layer0_outputs(6274)) xor (layer0_outputs(5967));
    outputs(1532) <= not((layer0_outputs(7614)) or (layer0_outputs(483)));
    outputs(1533) <= not((layer0_outputs(292)) or (layer0_outputs(5625)));
    outputs(1534) <= (layer0_outputs(1251)) xor (layer0_outputs(5654));
    outputs(1535) <= (layer0_outputs(7110)) and not (layer0_outputs(4990));
    outputs(1536) <= not(layer0_outputs(8081));
    outputs(1537) <= not((layer0_outputs(9234)) or (layer0_outputs(6101)));
    outputs(1538) <= (layer0_outputs(5021)) xor (layer0_outputs(2237));
    outputs(1539) <= (layer0_outputs(8652)) and (layer0_outputs(1074));
    outputs(1540) <= (layer0_outputs(81)) and not (layer0_outputs(6450));
    outputs(1541) <= (layer0_outputs(7811)) xor (layer0_outputs(3129));
    outputs(1542) <= not((layer0_outputs(643)) or (layer0_outputs(6289)));
    outputs(1543) <= (layer0_outputs(2045)) and not (layer0_outputs(323));
    outputs(1544) <= not(layer0_outputs(3432));
    outputs(1545) <= (layer0_outputs(2309)) and not (layer0_outputs(7930));
    outputs(1546) <= not((layer0_outputs(9465)) xor (layer0_outputs(4656)));
    outputs(1547) <= not((layer0_outputs(2441)) or (layer0_outputs(144)));
    outputs(1548) <= (layer0_outputs(7673)) xor (layer0_outputs(3778));
    outputs(1549) <= (layer0_outputs(7658)) and (layer0_outputs(7756));
    outputs(1550) <= (layer0_outputs(1639)) and (layer0_outputs(9805));
    outputs(1551) <= (layer0_outputs(3124)) xor (layer0_outputs(2642));
    outputs(1552) <= layer0_outputs(6024);
    outputs(1553) <= not((layer0_outputs(2420)) or (layer0_outputs(178)));
    outputs(1554) <= not(layer0_outputs(861));
    outputs(1555) <= (layer0_outputs(8124)) xor (layer0_outputs(8371));
    outputs(1556) <= (layer0_outputs(7391)) xor (layer0_outputs(2137));
    outputs(1557) <= (layer0_outputs(8913)) xor (layer0_outputs(9383));
    outputs(1558) <= (layer0_outputs(1014)) xor (layer0_outputs(8094));
    outputs(1559) <= layer0_outputs(2044);
    outputs(1560) <= not((layer0_outputs(2140)) xor (layer0_outputs(3305)));
    outputs(1561) <= (layer0_outputs(9305)) and not (layer0_outputs(2980));
    outputs(1562) <= not(layer0_outputs(4145));
    outputs(1563) <= not((layer0_outputs(6797)) xor (layer0_outputs(553)));
    outputs(1564) <= not((layer0_outputs(2426)) xor (layer0_outputs(298)));
    outputs(1565) <= not((layer0_outputs(8887)) xor (layer0_outputs(4582)));
    outputs(1566) <= '0';
    outputs(1567) <= not((layer0_outputs(965)) or (layer0_outputs(9862)));
    outputs(1568) <= not((layer0_outputs(2190)) or (layer0_outputs(1791)));
    outputs(1569) <= not((layer0_outputs(9368)) or (layer0_outputs(5175)));
    outputs(1570) <= (layer0_outputs(4964)) and not (layer0_outputs(7450));
    outputs(1571) <= not((layer0_outputs(9002)) and (layer0_outputs(1223)));
    outputs(1572) <= layer0_outputs(3265);
    outputs(1573) <= (layer0_outputs(3906)) and not (layer0_outputs(5399));
    outputs(1574) <= not((layer0_outputs(2609)) or (layer0_outputs(2920)));
    outputs(1575) <= (layer0_outputs(3360)) and (layer0_outputs(7338));
    outputs(1576) <= not((layer0_outputs(8068)) xor (layer0_outputs(333)));
    outputs(1577) <= not((layer0_outputs(5502)) xor (layer0_outputs(3102)));
    outputs(1578) <= (layer0_outputs(1979)) and (layer0_outputs(3158));
    outputs(1579) <= (layer0_outputs(5671)) xor (layer0_outputs(560));
    outputs(1580) <= not((layer0_outputs(9011)) xor (layer0_outputs(6582)));
    outputs(1581) <= not((layer0_outputs(4065)) xor (layer0_outputs(53)));
    outputs(1582) <= not((layer0_outputs(8832)) xor (layer0_outputs(10031)));
    outputs(1583) <= (layer0_outputs(4690)) and (layer0_outputs(4891));
    outputs(1584) <= not(layer0_outputs(237));
    outputs(1585) <= not(layer0_outputs(6085));
    outputs(1586) <= not((layer0_outputs(3116)) or (layer0_outputs(10214)));
    outputs(1587) <= (layer0_outputs(679)) xor (layer0_outputs(4038));
    outputs(1588) <= '0';
    outputs(1589) <= not((layer0_outputs(5663)) xor (layer0_outputs(110)));
    outputs(1590) <= (layer0_outputs(2880)) and not (layer0_outputs(1974));
    outputs(1591) <= (layer0_outputs(1825)) and not (layer0_outputs(5815));
    outputs(1592) <= (layer0_outputs(4195)) and not (layer0_outputs(5467));
    outputs(1593) <= layer0_outputs(9959);
    outputs(1594) <= (layer0_outputs(8206)) xor (layer0_outputs(8375));
    outputs(1595) <= (layer0_outputs(5791)) xor (layer0_outputs(8376));
    outputs(1596) <= (layer0_outputs(9642)) and not (layer0_outputs(5087));
    outputs(1597) <= not((layer0_outputs(5739)) xor (layer0_outputs(1548)));
    outputs(1598) <= (layer0_outputs(5304)) and (layer0_outputs(7863));
    outputs(1599) <= (layer0_outputs(8116)) or (layer0_outputs(10153));
    outputs(1600) <= (layer0_outputs(5206)) and not (layer0_outputs(7572));
    outputs(1601) <= not((layer0_outputs(5766)) or (layer0_outputs(3371)));
    outputs(1602) <= (layer0_outputs(2870)) and (layer0_outputs(9767));
    outputs(1603) <= (layer0_outputs(3261)) xor (layer0_outputs(1189));
    outputs(1604) <= (layer0_outputs(7316)) xor (layer0_outputs(5450));
    outputs(1605) <= not(layer0_outputs(4012));
    outputs(1606) <= (layer0_outputs(7468)) and not (layer0_outputs(8834));
    outputs(1607) <= (layer0_outputs(3330)) and (layer0_outputs(4117));
    outputs(1608) <= (layer0_outputs(10166)) xor (layer0_outputs(7384));
    outputs(1609) <= not((layer0_outputs(2759)) or (layer0_outputs(8580)));
    outputs(1610) <= (layer0_outputs(4180)) xor (layer0_outputs(6035));
    outputs(1611) <= not(layer0_outputs(8669));
    outputs(1612) <= (layer0_outputs(9604)) and not (layer0_outputs(9112));
    outputs(1613) <= (layer0_outputs(6751)) and not (layer0_outputs(367));
    outputs(1614) <= (layer0_outputs(6821)) and not (layer0_outputs(313));
    outputs(1615) <= layer0_outputs(4717);
    outputs(1616) <= (layer0_outputs(2215)) and not (layer0_outputs(6861));
    outputs(1617) <= not(layer0_outputs(5135));
    outputs(1618) <= (layer0_outputs(2479)) and not (layer0_outputs(9187));
    outputs(1619) <= (layer0_outputs(3777)) xor (layer0_outputs(1915));
    outputs(1620) <= (layer0_outputs(7257)) and not (layer0_outputs(9105));
    outputs(1621) <= '0';
    outputs(1622) <= (layer0_outputs(5488)) xor (layer0_outputs(4842));
    outputs(1623) <= (layer0_outputs(2212)) and not (layer0_outputs(268));
    outputs(1624) <= (layer0_outputs(1446)) and (layer0_outputs(6451));
    outputs(1625) <= not((layer0_outputs(7173)) or (layer0_outputs(1324)));
    outputs(1626) <= (layer0_outputs(1250)) xor (layer0_outputs(4265));
    outputs(1627) <= (layer0_outputs(5534)) xor (layer0_outputs(6400));
    outputs(1628) <= (layer0_outputs(10193)) and not (layer0_outputs(5422));
    outputs(1629) <= (layer0_outputs(6099)) and not (layer0_outputs(9745));
    outputs(1630) <= (layer0_outputs(7176)) xor (layer0_outputs(8951));
    outputs(1631) <= not((layer0_outputs(2199)) or (layer0_outputs(10091)));
    outputs(1632) <= (layer0_outputs(1998)) and not (layer0_outputs(5058));
    outputs(1633) <= not(layer0_outputs(3796));
    outputs(1634) <= not((layer0_outputs(5546)) xor (layer0_outputs(3849)));
    outputs(1635) <= layer0_outputs(1358);
    outputs(1636) <= not((layer0_outputs(3580)) or (layer0_outputs(7987)));
    outputs(1637) <= (layer0_outputs(562)) and (layer0_outputs(1084));
    outputs(1638) <= not((layer0_outputs(7091)) or (layer0_outputs(7866)));
    outputs(1639) <= (layer0_outputs(4397)) and not (layer0_outputs(6710));
    outputs(1640) <= layer0_outputs(9856);
    outputs(1641) <= (layer0_outputs(7774)) and (layer0_outputs(1284));
    outputs(1642) <= (layer0_outputs(6554)) and (layer0_outputs(3009));
    outputs(1643) <= layer0_outputs(3823);
    outputs(1644) <= (layer0_outputs(733)) and not (layer0_outputs(1916));
    outputs(1645) <= not(layer0_outputs(6075));
    outputs(1646) <= not((layer0_outputs(2121)) xor (layer0_outputs(10129)));
    outputs(1647) <= (layer0_outputs(8522)) xor (layer0_outputs(2886));
    outputs(1648) <= (layer0_outputs(7086)) and not (layer0_outputs(5162));
    outputs(1649) <= not(layer0_outputs(2894));
    outputs(1650) <= not(layer0_outputs(309));
    outputs(1651) <= not(layer0_outputs(6769));
    outputs(1652) <= not(layer0_outputs(4869));
    outputs(1653) <= layer0_outputs(3056);
    outputs(1654) <= (layer0_outputs(6459)) and (layer0_outputs(5656));
    outputs(1655) <= not((layer0_outputs(8121)) xor (layer0_outputs(9262)));
    outputs(1656) <= not((layer0_outputs(2155)) or (layer0_outputs(9644)));
    outputs(1657) <= not((layer0_outputs(8774)) xor (layer0_outputs(9882)));
    outputs(1658) <= not((layer0_outputs(2816)) xor (layer0_outputs(3345)));
    outputs(1659) <= layer0_outputs(9834);
    outputs(1660) <= (layer0_outputs(3783)) xor (layer0_outputs(7401));
    outputs(1661) <= (layer0_outputs(3338)) and not (layer0_outputs(8135));
    outputs(1662) <= (layer0_outputs(6148)) and (layer0_outputs(436));
    outputs(1663) <= layer0_outputs(4630);
    outputs(1664) <= not((layer0_outputs(303)) xor (layer0_outputs(4609)));
    outputs(1665) <= (layer0_outputs(6302)) xor (layer0_outputs(5916));
    outputs(1666) <= not((layer0_outputs(7319)) or (layer0_outputs(5627)));
    outputs(1667) <= (layer0_outputs(1845)) and not (layer0_outputs(8704));
    outputs(1668) <= layer0_outputs(9477);
    outputs(1669) <= (layer0_outputs(9942)) and not (layer0_outputs(4321));
    outputs(1670) <= (layer0_outputs(9509)) and not (layer0_outputs(4498));
    outputs(1671) <= (layer0_outputs(3639)) and (layer0_outputs(6065));
    outputs(1672) <= (layer0_outputs(813)) and not (layer0_outputs(169));
    outputs(1673) <= not((layer0_outputs(2455)) xor (layer0_outputs(3765)));
    outputs(1674) <= (layer0_outputs(4909)) xor (layer0_outputs(8111));
    outputs(1675) <= (layer0_outputs(134)) xor (layer0_outputs(2278));
    outputs(1676) <= (layer0_outputs(9772)) and not (layer0_outputs(651));
    outputs(1677) <= (layer0_outputs(7487)) and not (layer0_outputs(9917));
    outputs(1678) <= (layer0_outputs(4793)) xor (layer0_outputs(4822));
    outputs(1679) <= (layer0_outputs(2373)) xor (layer0_outputs(4046));
    outputs(1680) <= (layer0_outputs(4217)) and not (layer0_outputs(8416));
    outputs(1681) <= (layer0_outputs(5424)) xor (layer0_outputs(9281));
    outputs(1682) <= (layer0_outputs(7982)) xor (layer0_outputs(1069));
    outputs(1683) <= (layer0_outputs(3547)) and (layer0_outputs(5234));
    outputs(1684) <= (layer0_outputs(2840)) and (layer0_outputs(3294));
    outputs(1685) <= not(layer0_outputs(6071));
    outputs(1686) <= not((layer0_outputs(1383)) xor (layer0_outputs(1224)));
    outputs(1687) <= not(layer0_outputs(9020));
    outputs(1688) <= (layer0_outputs(5971)) and not (layer0_outputs(4712));
    outputs(1689) <= not((layer0_outputs(7278)) or (layer0_outputs(4583)));
    outputs(1690) <= (layer0_outputs(3819)) and (layer0_outputs(5507));
    outputs(1691) <= layer0_outputs(7043);
    outputs(1692) <= not((layer0_outputs(702)) or (layer0_outputs(8865)));
    outputs(1693) <= not((layer0_outputs(7907)) or (layer0_outputs(2109)));
    outputs(1694) <= layer0_outputs(3505);
    outputs(1695) <= (layer0_outputs(4137)) xor (layer0_outputs(3148));
    outputs(1696) <= not((layer0_outputs(3874)) xor (layer0_outputs(1722)));
    outputs(1697) <= layer0_outputs(6306);
    outputs(1698) <= not((layer0_outputs(7315)) xor (layer0_outputs(5036)));
    outputs(1699) <= (layer0_outputs(8020)) and not (layer0_outputs(8882));
    outputs(1700) <= layer0_outputs(5793);
    outputs(1701) <= layer0_outputs(1545);
    outputs(1702) <= (layer0_outputs(9292)) and (layer0_outputs(8956));
    outputs(1703) <= not(layer0_outputs(1989)) or (layer0_outputs(6442));
    outputs(1704) <= (layer0_outputs(4223)) xor (layer0_outputs(10176));
    outputs(1705) <= (layer0_outputs(3836)) xor (layer0_outputs(8744));
    outputs(1706) <= (layer0_outputs(7308)) and (layer0_outputs(62));
    outputs(1707) <= not(layer0_outputs(6619));
    outputs(1708) <= (layer0_outputs(9152)) and (layer0_outputs(4686));
    outputs(1709) <= not((layer0_outputs(7622)) xor (layer0_outputs(9403)));
    outputs(1710) <= not(layer0_outputs(1757));
    outputs(1711) <= not(layer0_outputs(1563));
    outputs(1712) <= layer0_outputs(4131);
    outputs(1713) <= (layer0_outputs(7481)) and not (layer0_outputs(1062));
    outputs(1714) <= (layer0_outputs(4478)) and not (layer0_outputs(944));
    outputs(1715) <= not(layer0_outputs(6505));
    outputs(1716) <= not((layer0_outputs(1776)) and (layer0_outputs(1096)));
    outputs(1717) <= layer0_outputs(5701);
    outputs(1718) <= layer0_outputs(7132);
    outputs(1719) <= (layer0_outputs(8286)) and not (layer0_outputs(10159));
    outputs(1720) <= (layer0_outputs(4277)) and not (layer0_outputs(8029));
    outputs(1721) <= (layer0_outputs(5923)) and not (layer0_outputs(1978));
    outputs(1722) <= (layer0_outputs(3484)) and not (layer0_outputs(2919));
    outputs(1723) <= (layer0_outputs(8559)) and not (layer0_outputs(6860));
    outputs(1724) <= (layer0_outputs(5140)) and (layer0_outputs(6070));
    outputs(1725) <= layer0_outputs(1210);
    outputs(1726) <= (layer0_outputs(3421)) and not (layer0_outputs(2399));
    outputs(1727) <= not((layer0_outputs(8607)) xor (layer0_outputs(5665)));
    outputs(1728) <= (layer0_outputs(3138)) and not (layer0_outputs(9431));
    outputs(1729) <= layer0_outputs(891);
    outputs(1730) <= not(layer0_outputs(2057));
    outputs(1731) <= (layer0_outputs(7848)) and (layer0_outputs(9277));
    outputs(1732) <= not(layer0_outputs(9937));
    outputs(1733) <= (layer0_outputs(910)) and (layer0_outputs(5771));
    outputs(1734) <= not(layer0_outputs(3083));
    outputs(1735) <= (layer0_outputs(4270)) xor (layer0_outputs(615));
    outputs(1736) <= not((layer0_outputs(5001)) or (layer0_outputs(2701)));
    outputs(1737) <= (layer0_outputs(6433)) and (layer0_outputs(3916));
    outputs(1738) <= (layer0_outputs(8453)) and not (layer0_outputs(8542));
    outputs(1739) <= (layer0_outputs(1787)) and not (layer0_outputs(4574));
    outputs(1740) <= (layer0_outputs(8112)) xor (layer0_outputs(8237));
    outputs(1741) <= (layer0_outputs(7533)) and not (layer0_outputs(7025));
    outputs(1742) <= not(layer0_outputs(986));
    outputs(1743) <= (layer0_outputs(7417)) and not (layer0_outputs(1118));
    outputs(1744) <= (layer0_outputs(4585)) xor (layer0_outputs(832));
    outputs(1745) <= not((layer0_outputs(9864)) xor (layer0_outputs(6369)));
    outputs(1746) <= not(layer0_outputs(7754));
    outputs(1747) <= (layer0_outputs(5356)) xor (layer0_outputs(9489));
    outputs(1748) <= (layer0_outputs(7551)) and not (layer0_outputs(5231));
    outputs(1749) <= layer0_outputs(9327);
    outputs(1750) <= not((layer0_outputs(8162)) xor (layer0_outputs(3349)));
    outputs(1751) <= not((layer0_outputs(8723)) and (layer0_outputs(4306)));
    outputs(1752) <= (layer0_outputs(6165)) and (layer0_outputs(5783));
    outputs(1753) <= (layer0_outputs(3520)) xor (layer0_outputs(9120));
    outputs(1754) <= not((layer0_outputs(9049)) xor (layer0_outputs(4742)));
    outputs(1755) <= layer0_outputs(4070);
    outputs(1756) <= not((layer0_outputs(2997)) xor (layer0_outputs(4750)));
    outputs(1757) <= not((layer0_outputs(2803)) or (layer0_outputs(10024)));
    outputs(1758) <= layer0_outputs(5196);
    outputs(1759) <= not(layer0_outputs(9066));
    outputs(1760) <= not((layer0_outputs(6313)) or (layer0_outputs(2755)));
    outputs(1761) <= not((layer0_outputs(226)) xor (layer0_outputs(21)));
    outputs(1762) <= (layer0_outputs(5073)) and (layer0_outputs(7479));
    outputs(1763) <= not((layer0_outputs(4762)) xor (layer0_outputs(2028)));
    outputs(1764) <= not((layer0_outputs(8556)) xor (layer0_outputs(4825)));
    outputs(1765) <= layer0_outputs(4969);
    outputs(1766) <= (layer0_outputs(838)) and not (layer0_outputs(3566));
    outputs(1767) <= (layer0_outputs(1742)) and not (layer0_outputs(9438));
    outputs(1768) <= layer0_outputs(4067);
    outputs(1769) <= (layer0_outputs(5540)) and not (layer0_outputs(4637));
    outputs(1770) <= not(layer0_outputs(5468));
    outputs(1771) <= (layer0_outputs(5789)) and not (layer0_outputs(442));
    outputs(1772) <= (layer0_outputs(2511)) xor (layer0_outputs(3060));
    outputs(1773) <= layer0_outputs(9322);
    outputs(1774) <= (layer0_outputs(1861)) and not (layer0_outputs(7050));
    outputs(1775) <= not(layer0_outputs(1474));
    outputs(1776) <= (layer0_outputs(1456)) and not (layer0_outputs(2746));
    outputs(1777) <= not((layer0_outputs(5635)) xor (layer0_outputs(3658)));
    outputs(1778) <= not((layer0_outputs(9065)) xor (layer0_outputs(9920)));
    outputs(1779) <= layer0_outputs(3896);
    outputs(1780) <= not(layer0_outputs(2985));
    outputs(1781) <= (layer0_outputs(9261)) xor (layer0_outputs(9011));
    outputs(1782) <= (layer0_outputs(6612)) and not (layer0_outputs(9965));
    outputs(1783) <= not((layer0_outputs(5965)) xor (layer0_outputs(6261)));
    outputs(1784) <= (layer0_outputs(4284)) and not (layer0_outputs(3164));
    outputs(1785) <= (layer0_outputs(3270)) and not (layer0_outputs(8337));
    outputs(1786) <= (layer0_outputs(8698)) and not (layer0_outputs(1990));
    outputs(1787) <= (layer0_outputs(4811)) and not (layer0_outputs(4275));
    outputs(1788) <= not((layer0_outputs(9087)) xor (layer0_outputs(3793)));
    outputs(1789) <= (layer0_outputs(10235)) and (layer0_outputs(2188));
    outputs(1790) <= (layer0_outputs(9521)) and not (layer0_outputs(10128));
    outputs(1791) <= layer0_outputs(6986);
    outputs(1792) <= not((layer0_outputs(10162)) or (layer0_outputs(8894)));
    outputs(1793) <= (layer0_outputs(2353)) xor (layer0_outputs(6632));
    outputs(1794) <= not((layer0_outputs(4102)) xor (layer0_outputs(222)));
    outputs(1795) <= not((layer0_outputs(319)) xor (layer0_outputs(7686)));
    outputs(1796) <= not(layer0_outputs(3494));
    outputs(1797) <= not(layer0_outputs(9874));
    outputs(1798) <= not(layer0_outputs(4698));
    outputs(1799) <= (layer0_outputs(299)) and not (layer0_outputs(4460));
    outputs(1800) <= not((layer0_outputs(3475)) or (layer0_outputs(3880)));
    outputs(1801) <= (layer0_outputs(3742)) and not (layer0_outputs(1385));
    outputs(1802) <= layer0_outputs(9566);
    outputs(1803) <= (layer0_outputs(5668)) and not (layer0_outputs(3636));
    outputs(1804) <= (layer0_outputs(933)) and not (layer0_outputs(10110));
    outputs(1805) <= not((layer0_outputs(5544)) xor (layer0_outputs(6894)));
    outputs(1806) <= (layer0_outputs(9794)) xor (layer0_outputs(1513));
    outputs(1807) <= (layer0_outputs(1036)) and (layer0_outputs(6920));
    outputs(1808) <= (layer0_outputs(7420)) xor (layer0_outputs(9113));
    outputs(1809) <= (layer0_outputs(9451)) and not (layer0_outputs(5504));
    outputs(1810) <= (layer0_outputs(10130)) and (layer0_outputs(8233));
    outputs(1811) <= (layer0_outputs(1536)) xor (layer0_outputs(8914));
    outputs(1812) <= (layer0_outputs(5935)) xor (layer0_outputs(5452));
    outputs(1813) <= not((layer0_outputs(2161)) xor (layer0_outputs(5902)));
    outputs(1814) <= layer0_outputs(4773);
    outputs(1815) <= layer0_outputs(804);
    outputs(1816) <= not(layer0_outputs(5111));
    outputs(1817) <= not((layer0_outputs(1852)) xor (layer0_outputs(2221)));
    outputs(1818) <= (layer0_outputs(8695)) and (layer0_outputs(8666));
    outputs(1819) <= (layer0_outputs(1152)) xor (layer0_outputs(3678));
    outputs(1820) <= not(layer0_outputs(5096));
    outputs(1821) <= not((layer0_outputs(2679)) or (layer0_outputs(2383)));
    outputs(1822) <= (layer0_outputs(9642)) and not (layer0_outputs(7908));
    outputs(1823) <= (layer0_outputs(6381)) xor (layer0_outputs(7107));
    outputs(1824) <= not((layer0_outputs(8262)) xor (layer0_outputs(9135)));
    outputs(1825) <= (layer0_outputs(2741)) and (layer0_outputs(3290));
    outputs(1826) <= not(layer0_outputs(8849));
    outputs(1827) <= not((layer0_outputs(3398)) xor (layer0_outputs(2130)));
    outputs(1828) <= (layer0_outputs(7637)) and not (layer0_outputs(956));
    outputs(1829) <= (layer0_outputs(3964)) and not (layer0_outputs(2450));
    outputs(1830) <= '0';
    outputs(1831) <= not((layer0_outputs(2799)) or (layer0_outputs(7628)));
    outputs(1832) <= (layer0_outputs(1831)) and not (layer0_outputs(9458));
    outputs(1833) <= layer0_outputs(3543);
    outputs(1834) <= (layer0_outputs(2567)) xor (layer0_outputs(6320));
    outputs(1835) <= not((layer0_outputs(7854)) or (layer0_outputs(757)));
    outputs(1836) <= (layer0_outputs(3851)) and not (layer0_outputs(2886));
    outputs(1837) <= layer0_outputs(7182);
    outputs(1838) <= not((layer0_outputs(2857)) xor (layer0_outputs(4136)));
    outputs(1839) <= layer0_outputs(2334);
    outputs(1840) <= layer0_outputs(3050);
    outputs(1841) <= not(layer0_outputs(7160));
    outputs(1842) <= (layer0_outputs(3814)) and not (layer0_outputs(987));
    outputs(1843) <= (layer0_outputs(3333)) and not (layer0_outputs(305));
    outputs(1844) <= (layer0_outputs(3557)) and not (layer0_outputs(5173));
    outputs(1845) <= (layer0_outputs(5691)) xor (layer0_outputs(5106));
    outputs(1846) <= (layer0_outputs(7425)) xor (layer0_outputs(5861));
    outputs(1847) <= not((layer0_outputs(6016)) xor (layer0_outputs(5787)));
    outputs(1848) <= not((layer0_outputs(7849)) or (layer0_outputs(1283)));
    outputs(1849) <= (layer0_outputs(447)) and not (layer0_outputs(4432));
    outputs(1850) <= (layer0_outputs(1311)) and (layer0_outputs(8345));
    outputs(1851) <= (layer0_outputs(9818)) and not (layer0_outputs(442));
    outputs(1852) <= (layer0_outputs(4966)) and (layer0_outputs(7272));
    outputs(1853) <= layer0_outputs(6984);
    outputs(1854) <= not(layer0_outputs(5410));
    outputs(1855) <= (layer0_outputs(1673)) xor (layer0_outputs(4667));
    outputs(1856) <= (layer0_outputs(9220)) and not (layer0_outputs(211));
    outputs(1857) <= layer0_outputs(3731);
    outputs(1858) <= (layer0_outputs(914)) and not (layer0_outputs(8392));
    outputs(1859) <= (layer0_outputs(2475)) xor (layer0_outputs(1965));
    outputs(1860) <= (layer0_outputs(9007)) and not (layer0_outputs(2945));
    outputs(1861) <= not((layer0_outputs(4489)) xor (layer0_outputs(5065)));
    outputs(1862) <= (layer0_outputs(2119)) xor (layer0_outputs(4968));
    outputs(1863) <= (layer0_outputs(1554)) and not (layer0_outputs(2739));
    outputs(1864) <= not((layer0_outputs(181)) xor (layer0_outputs(9347)));
    outputs(1865) <= (layer0_outputs(4508)) and not (layer0_outputs(3383));
    outputs(1866) <= (layer0_outputs(8444)) and (layer0_outputs(7623));
    outputs(1867) <= layer0_outputs(1769);
    outputs(1868) <= layer0_outputs(2019);
    outputs(1869) <= not((layer0_outputs(7380)) xor (layer0_outputs(6488)));
    outputs(1870) <= not((layer0_outputs(4266)) or (layer0_outputs(9000)));
    outputs(1871) <= (layer0_outputs(8741)) and (layer0_outputs(550));
    outputs(1872) <= (layer0_outputs(6152)) and not (layer0_outputs(7963));
    outputs(1873) <= layer0_outputs(8126);
    outputs(1874) <= not(layer0_outputs(5182));
    outputs(1875) <= not((layer0_outputs(7801)) or (layer0_outputs(6426)));
    outputs(1876) <= not((layer0_outputs(1231)) xor (layer0_outputs(8490)));
    outputs(1877) <= layer0_outputs(5723);
    outputs(1878) <= (layer0_outputs(2170)) and not (layer0_outputs(1650));
    outputs(1879) <= (layer0_outputs(2069)) and not (layer0_outputs(1115));
    outputs(1880) <= not((layer0_outputs(1387)) xor (layer0_outputs(7168)));
    outputs(1881) <= layer0_outputs(8532);
    outputs(1882) <= not((layer0_outputs(37)) xor (layer0_outputs(2284)));
    outputs(1883) <= not((layer0_outputs(8846)) xor (layer0_outputs(9791)));
    outputs(1884) <= (layer0_outputs(1020)) and (layer0_outputs(7027));
    outputs(1885) <= not((layer0_outputs(1290)) or (layer0_outputs(5797)));
    outputs(1886) <= not((layer0_outputs(1539)) or (layer0_outputs(5249)));
    outputs(1887) <= layer0_outputs(6779);
    outputs(1888) <= (layer0_outputs(4317)) and not (layer0_outputs(5843));
    outputs(1889) <= layer0_outputs(8009);
    outputs(1890) <= (layer0_outputs(177)) and not (layer0_outputs(6352));
    outputs(1891) <= layer0_outputs(4963);
    outputs(1892) <= (layer0_outputs(8516)) and not (layer0_outputs(3297));
    outputs(1893) <= not(layer0_outputs(4155));
    outputs(1894) <= not(layer0_outputs(8885));
    outputs(1895) <= (layer0_outputs(1960)) and (layer0_outputs(7503));
    outputs(1896) <= not((layer0_outputs(4468)) xor (layer0_outputs(7910)));
    outputs(1897) <= not((layer0_outputs(3187)) xor (layer0_outputs(4223)));
    outputs(1898) <= not((layer0_outputs(2864)) xor (layer0_outputs(603)));
    outputs(1899) <= (layer0_outputs(8844)) and not (layer0_outputs(3359));
    outputs(1900) <= (layer0_outputs(5262)) xor (layer0_outputs(7209));
    outputs(1901) <= (layer0_outputs(2753)) and not (layer0_outputs(1237));
    outputs(1902) <= not((layer0_outputs(5470)) xor (layer0_outputs(5039)));
    outputs(1903) <= (layer0_outputs(10005)) xor (layer0_outputs(6299));
    outputs(1904) <= (layer0_outputs(2085)) and not (layer0_outputs(6597));
    outputs(1905) <= not((layer0_outputs(7820)) xor (layer0_outputs(4764)));
    outputs(1906) <= (layer0_outputs(1779)) and not (layer0_outputs(967));
    outputs(1907) <= (layer0_outputs(4110)) and (layer0_outputs(3961));
    outputs(1908) <= not((layer0_outputs(2500)) xor (layer0_outputs(9781)));
    outputs(1909) <= (layer0_outputs(4435)) and not (layer0_outputs(1063));
    outputs(1910) <= not(layer0_outputs(7548));
    outputs(1911) <= not((layer0_outputs(1965)) or (layer0_outputs(8316)));
    outputs(1912) <= layer0_outputs(2636);
    outputs(1913) <= (layer0_outputs(2414)) and not (layer0_outputs(2790));
    outputs(1914) <= (layer0_outputs(5516)) xor (layer0_outputs(3723));
    outputs(1915) <= '0';
    outputs(1916) <= not(layer0_outputs(8867));
    outputs(1917) <= not(layer0_outputs(9728));
    outputs(1918) <= (layer0_outputs(7770)) and (layer0_outputs(9496));
    outputs(1919) <= (layer0_outputs(7341)) and (layer0_outputs(3631));
    outputs(1920) <= (layer0_outputs(3)) and (layer0_outputs(9139));
    outputs(1921) <= layer0_outputs(3480);
    outputs(1922) <= not(layer0_outputs(1391));
    outputs(1923) <= layer0_outputs(7972);
    outputs(1924) <= (layer0_outputs(3149)) and not (layer0_outputs(3105));
    outputs(1925) <= not((layer0_outputs(7747)) or (layer0_outputs(3217)));
    outputs(1926) <= (layer0_outputs(1680)) xor (layer0_outputs(7619));
    outputs(1927) <= not((layer0_outputs(9866)) xor (layer0_outputs(10046)));
    outputs(1928) <= (layer0_outputs(5034)) and (layer0_outputs(6013));
    outputs(1929) <= layer0_outputs(8030);
    outputs(1930) <= layer0_outputs(1685);
    outputs(1931) <= (layer0_outputs(8320)) xor (layer0_outputs(2763));
    outputs(1932) <= (layer0_outputs(2341)) and not (layer0_outputs(9700));
    outputs(1933) <= layer0_outputs(3180);
    outputs(1934) <= (layer0_outputs(9014)) and (layer0_outputs(5146));
    outputs(1935) <= not((layer0_outputs(7391)) or (layer0_outputs(9908)));
    outputs(1936) <= not(layer0_outputs(5482));
    outputs(1937) <= not((layer0_outputs(2504)) xor (layer0_outputs(2672)));
    outputs(1938) <= (layer0_outputs(988)) and (layer0_outputs(4345));
    outputs(1939) <= (layer0_outputs(4849)) and not (layer0_outputs(2249));
    outputs(1940) <= (layer0_outputs(6623)) and not (layer0_outputs(5631));
    outputs(1941) <= not((layer0_outputs(6076)) or (layer0_outputs(1255)));
    outputs(1942) <= not(layer0_outputs(6195));
    outputs(1943) <= not((layer0_outputs(822)) xor (layer0_outputs(7281)));
    outputs(1944) <= (layer0_outputs(3206)) or (layer0_outputs(6041));
    outputs(1945) <= (layer0_outputs(6806)) and (layer0_outputs(8226));
    outputs(1946) <= (layer0_outputs(4799)) and not (layer0_outputs(9667));
    outputs(1947) <= layer0_outputs(8254);
    outputs(1948) <= '0';
    outputs(1949) <= not((layer0_outputs(625)) xor (layer0_outputs(8660)));
    outputs(1950) <= (layer0_outputs(3618)) xor (layer0_outputs(4863));
    outputs(1951) <= (layer0_outputs(7262)) xor (layer0_outputs(3703));
    outputs(1952) <= not((layer0_outputs(8866)) or (layer0_outputs(9552)));
    outputs(1953) <= layer0_outputs(5100);
    outputs(1954) <= layer0_outputs(3726);
    outputs(1955) <= layer0_outputs(9463);
    outputs(1956) <= (layer0_outputs(4878)) and not (layer0_outputs(4112));
    outputs(1957) <= not(layer0_outputs(1532));
    outputs(1958) <= (layer0_outputs(3051)) xor (layer0_outputs(5237));
    outputs(1959) <= not((layer0_outputs(4506)) or (layer0_outputs(874)));
    outputs(1960) <= not((layer0_outputs(8340)) or (layer0_outputs(9404)));
    outputs(1961) <= (layer0_outputs(2948)) and not (layer0_outputs(7940));
    outputs(1962) <= (layer0_outputs(8926)) xor (layer0_outputs(6082));
    outputs(1963) <= (layer0_outputs(1547)) and not (layer0_outputs(7885));
    outputs(1964) <= (layer0_outputs(3579)) xor (layer0_outputs(5592));
    outputs(1965) <= not((layer0_outputs(2353)) xor (layer0_outputs(10195)));
    outputs(1966) <= layer0_outputs(4686);
    outputs(1967) <= (layer0_outputs(6280)) and (layer0_outputs(2953));
    outputs(1968) <= not(layer0_outputs(4465)) or (layer0_outputs(3596));
    outputs(1969) <= (layer0_outputs(276)) and not (layer0_outputs(7647));
    outputs(1970) <= not(layer0_outputs(8534));
    outputs(1971) <= (layer0_outputs(2880)) and not (layer0_outputs(6608));
    outputs(1972) <= not(layer0_outputs(9812)) or (layer0_outputs(5285));
    outputs(1973) <= not(layer0_outputs(9978));
    outputs(1974) <= (layer0_outputs(2111)) and not (layer0_outputs(2102));
    outputs(1975) <= (layer0_outputs(3099)) and not (layer0_outputs(5429));
    outputs(1976) <= '0';
    outputs(1977) <= (layer0_outputs(7898)) xor (layer0_outputs(3357));
    outputs(1978) <= (layer0_outputs(7961)) and (layer0_outputs(9841));
    outputs(1979) <= (layer0_outputs(8434)) xor (layer0_outputs(6329));
    outputs(1980) <= not((layer0_outputs(3182)) or (layer0_outputs(9756)));
    outputs(1981) <= (layer0_outputs(8472)) and not (layer0_outputs(2382));
    outputs(1982) <= not((layer0_outputs(9745)) or (layer0_outputs(4477)));
    outputs(1983) <= (layer0_outputs(5914)) and not (layer0_outputs(8313));
    outputs(1984) <= (layer0_outputs(9094)) and not (layer0_outputs(883));
    outputs(1985) <= (layer0_outputs(6045)) and not (layer0_outputs(3561));
    outputs(1986) <= layer0_outputs(1398);
    outputs(1987) <= (layer0_outputs(8369)) and not (layer0_outputs(5224));
    outputs(1988) <= not(layer0_outputs(5));
    outputs(1989) <= not(layer0_outputs(9174));
    outputs(1990) <= not((layer0_outputs(2173)) or (layer0_outputs(8057)));
    outputs(1991) <= not((layer0_outputs(6532)) xor (layer0_outputs(1165)));
    outputs(1992) <= layer0_outputs(4724);
    outputs(1993) <= (layer0_outputs(2947)) and not (layer0_outputs(4637));
    outputs(1994) <= (layer0_outputs(3608)) and not (layer0_outputs(9062));
    outputs(1995) <= not((layer0_outputs(1340)) or (layer0_outputs(9753)));
    outputs(1996) <= (layer0_outputs(5252)) xor (layer0_outputs(2603));
    outputs(1997) <= (layer0_outputs(6298)) and (layer0_outputs(6999));
    outputs(1998) <= '0';
    outputs(1999) <= (layer0_outputs(1389)) and (layer0_outputs(5479));
    outputs(2000) <= (layer0_outputs(2063)) xor (layer0_outputs(8636));
    outputs(2001) <= not((layer0_outputs(3556)) xor (layer0_outputs(7282)));
    outputs(2002) <= (layer0_outputs(7001)) xor (layer0_outputs(8141));
    outputs(2003) <= (layer0_outputs(1303)) and (layer0_outputs(8734));
    outputs(2004) <= not((layer0_outputs(3369)) or (layer0_outputs(4474)));
    outputs(2005) <= not((layer0_outputs(1632)) xor (layer0_outputs(8001)));
    outputs(2006) <= not((layer0_outputs(9163)) xor (layer0_outputs(4643)));
    outputs(2007) <= not((layer0_outputs(5558)) or (layer0_outputs(8251)));
    outputs(2008) <= not((layer0_outputs(617)) or (layer0_outputs(7144)));
    outputs(2009) <= (layer0_outputs(6840)) and not (layer0_outputs(7984));
    outputs(2010) <= not((layer0_outputs(8757)) or (layer0_outputs(7782)));
    outputs(2011) <= not(layer0_outputs(2629));
    outputs(2012) <= (layer0_outputs(7046)) and (layer0_outputs(474));
    outputs(2013) <= (layer0_outputs(6367)) and not (layer0_outputs(5057));
    outputs(2014) <= (layer0_outputs(46)) xor (layer0_outputs(2483));
    outputs(2015) <= (layer0_outputs(2781)) and (layer0_outputs(4313));
    outputs(2016) <= (layer0_outputs(9844)) xor (layer0_outputs(8562));
    outputs(2017) <= not((layer0_outputs(8657)) xor (layer0_outputs(8240)));
    outputs(2018) <= (layer0_outputs(3835)) and not (layer0_outputs(5069));
    outputs(2019) <= (layer0_outputs(9807)) and not (layer0_outputs(3081));
    outputs(2020) <= (layer0_outputs(6964)) and not (layer0_outputs(3393));
    outputs(2021) <= (layer0_outputs(6869)) and not (layer0_outputs(3501));
    outputs(2022) <= not((layer0_outputs(7191)) or (layer0_outputs(8458)));
    outputs(2023) <= (layer0_outputs(4976)) and not (layer0_outputs(4330));
    outputs(2024) <= (layer0_outputs(8090)) and not (layer0_outputs(5526));
    outputs(2025) <= (layer0_outputs(1569)) and not (layer0_outputs(6919));
    outputs(2026) <= (layer0_outputs(6872)) and (layer0_outputs(9855));
    outputs(2027) <= '0';
    outputs(2028) <= (layer0_outputs(9873)) and not (layer0_outputs(4462));
    outputs(2029) <= not((layer0_outputs(4546)) xor (layer0_outputs(5429)));
    outputs(2030) <= (layer0_outputs(2258)) and not (layer0_outputs(1551));
    outputs(2031) <= layer0_outputs(2270);
    outputs(2032) <= (layer0_outputs(5657)) and not (layer0_outputs(712));
    outputs(2033) <= not((layer0_outputs(6203)) xor (layer0_outputs(6293)));
    outputs(2034) <= (layer0_outputs(4096)) and not (layer0_outputs(9715));
    outputs(2035) <= not((layer0_outputs(2859)) or (layer0_outputs(9230)));
    outputs(2036) <= (layer0_outputs(8504)) and not (layer0_outputs(5026));
    outputs(2037) <= (layer0_outputs(5890)) and not (layer0_outputs(2840));
    outputs(2038) <= (layer0_outputs(2268)) and not (layer0_outputs(4460));
    outputs(2039) <= not((layer0_outputs(210)) or (layer0_outputs(2914)));
    outputs(2040) <= (layer0_outputs(6921)) xor (layer0_outputs(6182));
    outputs(2041) <= (layer0_outputs(6091)) and (layer0_outputs(3043));
    outputs(2042) <= layer0_outputs(6259);
    outputs(2043) <= not(layer0_outputs(824));
    outputs(2044) <= layer0_outputs(2552);
    outputs(2045) <= layer0_outputs(8428);
    outputs(2046) <= layer0_outputs(2494);
    outputs(2047) <= (layer0_outputs(8356)) and (layer0_outputs(2489));
    outputs(2048) <= not(layer0_outputs(9426));
    outputs(2049) <= not((layer0_outputs(9582)) xor (layer0_outputs(185)));
    outputs(2050) <= not(layer0_outputs(7448));
    outputs(2051) <= (layer0_outputs(2666)) and not (layer0_outputs(2346));
    outputs(2052) <= layer0_outputs(5497);
    outputs(2053) <= not(layer0_outputs(7706)) or (layer0_outputs(7335));
    outputs(2054) <= not(layer0_outputs(3651));
    outputs(2055) <= not(layer0_outputs(2551)) or (layer0_outputs(8183));
    outputs(2056) <= (layer0_outputs(9208)) or (layer0_outputs(7068));
    outputs(2057) <= layer0_outputs(5002);
    outputs(2058) <= not(layer0_outputs(2550)) or (layer0_outputs(4901));
    outputs(2059) <= layer0_outputs(10040);
    outputs(2060) <= not(layer0_outputs(884));
    outputs(2061) <= not(layer0_outputs(9591));
    outputs(2062) <= (layer0_outputs(8933)) xor (layer0_outputs(1843));
    outputs(2063) <= not((layer0_outputs(4299)) or (layer0_outputs(2979)));
    outputs(2064) <= not(layer0_outputs(7573));
    outputs(2065) <= layer0_outputs(2082);
    outputs(2066) <= layer0_outputs(1539);
    outputs(2067) <= layer0_outputs(7973);
    outputs(2068) <= not((layer0_outputs(7157)) and (layer0_outputs(734)));
    outputs(2069) <= not((layer0_outputs(9712)) xor (layer0_outputs(5203)));
    outputs(2070) <= not(layer0_outputs(7835));
    outputs(2071) <= not(layer0_outputs(2868));
    outputs(2072) <= not(layer0_outputs(5762));
    outputs(2073) <= not(layer0_outputs(932));
    outputs(2074) <= (layer0_outputs(7942)) or (layer0_outputs(5703));
    outputs(2075) <= layer0_outputs(8966);
    outputs(2076) <= layer0_outputs(9743);
    outputs(2077) <= (layer0_outputs(1917)) and not (layer0_outputs(8952));
    outputs(2078) <= (layer0_outputs(384)) and not (layer0_outputs(7692));
    outputs(2079) <= not((layer0_outputs(9313)) xor (layer0_outputs(8012)));
    outputs(2080) <= not(layer0_outputs(6220));
    outputs(2081) <= not((layer0_outputs(8105)) xor (layer0_outputs(7033)));
    outputs(2082) <= layer0_outputs(3368);
    outputs(2083) <= (layer0_outputs(9850)) or (layer0_outputs(7862));
    outputs(2084) <= (layer0_outputs(6447)) xor (layer0_outputs(9826));
    outputs(2085) <= not((layer0_outputs(3817)) xor (layer0_outputs(6712)));
    outputs(2086) <= layer0_outputs(1136);
    outputs(2087) <= layer0_outputs(788);
    outputs(2088) <= (layer0_outputs(5228)) or (layer0_outputs(9968));
    outputs(2089) <= layer0_outputs(8920);
    outputs(2090) <= not(layer0_outputs(5035));
    outputs(2091) <= not((layer0_outputs(7818)) xor (layer0_outputs(5673)));
    outputs(2092) <= not(layer0_outputs(5807));
    outputs(2093) <= not(layer0_outputs(9326));
    outputs(2094) <= not(layer0_outputs(6480)) or (layer0_outputs(6006));
    outputs(2095) <= not(layer0_outputs(5635));
    outputs(2096) <= layer0_outputs(2213);
    outputs(2097) <= layer0_outputs(9961);
    outputs(2098) <= not((layer0_outputs(4539)) xor (layer0_outputs(1264)));
    outputs(2099) <= not(layer0_outputs(7339)) or (layer0_outputs(8942));
    outputs(2100) <= not((layer0_outputs(2127)) xor (layer0_outputs(1149)));
    outputs(2101) <= layer0_outputs(4437);
    outputs(2102) <= (layer0_outputs(9650)) and not (layer0_outputs(7161));
    outputs(2103) <= (layer0_outputs(8005)) xor (layer0_outputs(1493));
    outputs(2104) <= (layer0_outputs(770)) and not (layer0_outputs(5958));
    outputs(2105) <= (layer0_outputs(5121)) xor (layer0_outputs(5373));
    outputs(2106) <= layer0_outputs(905);
    outputs(2107) <= not(layer0_outputs(6508));
    outputs(2108) <= not(layer0_outputs(6034));
    outputs(2109) <= layer0_outputs(5915);
    outputs(2110) <= layer0_outputs(5632);
    outputs(2111) <= not((layer0_outputs(2535)) xor (layer0_outputs(413)));
    outputs(2112) <= (layer0_outputs(8079)) or (layer0_outputs(7349));
    outputs(2113) <= not((layer0_outputs(10188)) or (layer0_outputs(2026)));
    outputs(2114) <= (layer0_outputs(1774)) xor (layer0_outputs(2346));
    outputs(2115) <= not(layer0_outputs(5539));
    outputs(2116) <= (layer0_outputs(722)) xor (layer0_outputs(9803));
    outputs(2117) <= layer0_outputs(6987);
    outputs(2118) <= not(layer0_outputs(6638));
    outputs(2119) <= (layer0_outputs(638)) xor (layer0_outputs(8516));
    outputs(2120) <= layer0_outputs(8182);
    outputs(2121) <= layer0_outputs(9589);
    outputs(2122) <= not(layer0_outputs(7872));
    outputs(2123) <= layer0_outputs(3573);
    outputs(2124) <= (layer0_outputs(902)) or (layer0_outputs(1050));
    outputs(2125) <= not((layer0_outputs(6595)) xor (layer0_outputs(4999)));
    outputs(2126) <= not(layer0_outputs(7580));
    outputs(2127) <= not(layer0_outputs(2131)) or (layer0_outputs(6557));
    outputs(2128) <= layer0_outputs(2362);
    outputs(2129) <= not(layer0_outputs(8310)) or (layer0_outputs(2887));
    outputs(2130) <= not(layer0_outputs(5552)) or (layer0_outputs(6732));
    outputs(2131) <= not(layer0_outputs(2858));
    outputs(2132) <= layer0_outputs(8622);
    outputs(2133) <= not((layer0_outputs(2275)) and (layer0_outputs(9231)));
    outputs(2134) <= not(layer0_outputs(2859));
    outputs(2135) <= (layer0_outputs(3032)) xor (layer0_outputs(8802));
    outputs(2136) <= not((layer0_outputs(2049)) and (layer0_outputs(5194)));
    outputs(2137) <= layer0_outputs(6201);
    outputs(2138) <= layer0_outputs(8851);
    outputs(2139) <= not(layer0_outputs(3838)) or (layer0_outputs(3561));
    outputs(2140) <= layer0_outputs(4300);
    outputs(2141) <= (layer0_outputs(1724)) or (layer0_outputs(1395));
    outputs(2142) <= (layer0_outputs(4270)) xor (layer0_outputs(3671));
    outputs(2143) <= (layer0_outputs(3271)) xor (layer0_outputs(9987));
    outputs(2144) <= not(layer0_outputs(381));
    outputs(2145) <= not(layer0_outputs(12)) or (layer0_outputs(713));
    outputs(2146) <= layer0_outputs(5977);
    outputs(2147) <= not(layer0_outputs(6512)) or (layer0_outputs(4776));
    outputs(2148) <= not(layer0_outputs(7727));
    outputs(2149) <= layer0_outputs(4916);
    outputs(2150) <= not(layer0_outputs(5315)) or (layer0_outputs(4007));
    outputs(2151) <= not(layer0_outputs(2445)) or (layer0_outputs(4795));
    outputs(2152) <= not(layer0_outputs(9803)) or (layer0_outputs(3144));
    outputs(2153) <= not(layer0_outputs(4216)) or (layer0_outputs(5602));
    outputs(2154) <= layer0_outputs(8342);
    outputs(2155) <= (layer0_outputs(3219)) and not (layer0_outputs(5988));
    outputs(2156) <= not(layer0_outputs(8205));
    outputs(2157) <= (layer0_outputs(1442)) or (layer0_outputs(9104));
    outputs(2158) <= not(layer0_outputs(6486)) or (layer0_outputs(502));
    outputs(2159) <= layer0_outputs(855);
    outputs(2160) <= (layer0_outputs(8230)) xor (layer0_outputs(5580));
    outputs(2161) <= not(layer0_outputs(8430));
    outputs(2162) <= layer0_outputs(7260);
    outputs(2163) <= not(layer0_outputs(1037));
    outputs(2164) <= not(layer0_outputs(395));
    outputs(2165) <= not(layer0_outputs(4729));
    outputs(2166) <= layer0_outputs(7210);
    outputs(2167) <= not(layer0_outputs(5474)) or (layer0_outputs(2756));
    outputs(2168) <= (layer0_outputs(7106)) xor (layer0_outputs(234));
    outputs(2169) <= not(layer0_outputs(9697));
    outputs(2170) <= not((layer0_outputs(5272)) and (layer0_outputs(321)));
    outputs(2171) <= not(layer0_outputs(726));
    outputs(2172) <= layer0_outputs(10156);
    outputs(2173) <= not(layer0_outputs(8503));
    outputs(2174) <= layer0_outputs(2927);
    outputs(2175) <= (layer0_outputs(2982)) and not (layer0_outputs(7830));
    outputs(2176) <= not((layer0_outputs(2399)) xor (layer0_outputs(7730)));
    outputs(2177) <= not(layer0_outputs(3024));
    outputs(2178) <= not(layer0_outputs(4629));
    outputs(2179) <= layer0_outputs(8584);
    outputs(2180) <= not(layer0_outputs(6544));
    outputs(2181) <= not((layer0_outputs(876)) and (layer0_outputs(4370)));
    outputs(2182) <= not(layer0_outputs(9364)) or (layer0_outputs(9853));
    outputs(2183) <= layer0_outputs(4320);
    outputs(2184) <= (layer0_outputs(3246)) or (layer0_outputs(718));
    outputs(2185) <= layer0_outputs(7466);
    outputs(2186) <= not(layer0_outputs(2046)) or (layer0_outputs(9132));
    outputs(2187) <= layer0_outputs(3212);
    outputs(2188) <= (layer0_outputs(5853)) and not (layer0_outputs(3750));
    outputs(2189) <= not(layer0_outputs(7582));
    outputs(2190) <= (layer0_outputs(1239)) xor (layer0_outputs(9722));
    outputs(2191) <= (layer0_outputs(682)) xor (layer0_outputs(4200));
    outputs(2192) <= not(layer0_outputs(6760)) or (layer0_outputs(1275));
    outputs(2193) <= not(layer0_outputs(2342));
    outputs(2194) <= not(layer0_outputs(2483));
    outputs(2195) <= not(layer0_outputs(3162));
    outputs(2196) <= (layer0_outputs(3738)) or (layer0_outputs(10180));
    outputs(2197) <= not((layer0_outputs(5726)) and (layer0_outputs(5774)));
    outputs(2198) <= not(layer0_outputs(4980));
    outputs(2199) <= not(layer0_outputs(2542)) or (layer0_outputs(7753));
    outputs(2200) <= not(layer0_outputs(6774));
    outputs(2201) <= not(layer0_outputs(2375));
    outputs(2202) <= not(layer0_outputs(9830));
    outputs(2203) <= layer0_outputs(4829);
    outputs(2204) <= not(layer0_outputs(9841));
    outputs(2205) <= not((layer0_outputs(1426)) and (layer0_outputs(6295)));
    outputs(2206) <= not(layer0_outputs(9678));
    outputs(2207) <= not((layer0_outputs(6940)) and (layer0_outputs(3872)));
    outputs(2208) <= not(layer0_outputs(5361));
    outputs(2209) <= not(layer0_outputs(7636));
    outputs(2210) <= (layer0_outputs(6359)) xor (layer0_outputs(8700));
    outputs(2211) <= layer0_outputs(1747);
    outputs(2212) <= not(layer0_outputs(9133));
    outputs(2213) <= not(layer0_outputs(457));
    outputs(2214) <= layer0_outputs(8983);
    outputs(2215) <= not((layer0_outputs(4921)) and (layer0_outputs(3356)));
    outputs(2216) <= not(layer0_outputs(33));
    outputs(2217) <= not(layer0_outputs(5148));
    outputs(2218) <= (layer0_outputs(6920)) xor (layer0_outputs(9191));
    outputs(2219) <= (layer0_outputs(6803)) or (layer0_outputs(4192));
    outputs(2220) <= not(layer0_outputs(1010)) or (layer0_outputs(4286));
    outputs(2221) <= (layer0_outputs(9739)) and not (layer0_outputs(7276));
    outputs(2222) <= not(layer0_outputs(5549));
    outputs(2223) <= (layer0_outputs(8192)) xor (layer0_outputs(8852));
    outputs(2224) <= not(layer0_outputs(9627));
    outputs(2225) <= not((layer0_outputs(7372)) xor (layer0_outputs(10045)));
    outputs(2226) <= not(layer0_outputs(4399)) or (layer0_outputs(1417));
    outputs(2227) <= layer0_outputs(9684);
    outputs(2228) <= layer0_outputs(162);
    outputs(2229) <= (layer0_outputs(3539)) and not (layer0_outputs(4352));
    outputs(2230) <= (layer0_outputs(3130)) or (layer0_outputs(5505));
    outputs(2231) <= not((layer0_outputs(10129)) xor (layer0_outputs(3309)));
    outputs(2232) <= layer0_outputs(5185);
    outputs(2233) <= not(layer0_outputs(8552)) or (layer0_outputs(1779));
    outputs(2234) <= layer0_outputs(5486);
    outputs(2235) <= not(layer0_outputs(7780));
    outputs(2236) <= not((layer0_outputs(1090)) and (layer0_outputs(3279)));
    outputs(2237) <= not((layer0_outputs(2782)) xor (layer0_outputs(6077)));
    outputs(2238) <= not((layer0_outputs(565)) and (layer0_outputs(7139)));
    outputs(2239) <= layer0_outputs(4954);
    outputs(2240) <= (layer0_outputs(3774)) and not (layer0_outputs(2090));
    outputs(2241) <= (layer0_outputs(2879)) or (layer0_outputs(6858));
    outputs(2242) <= not(layer0_outputs(6390));
    outputs(2243) <= (layer0_outputs(5170)) and not (layer0_outputs(3209));
    outputs(2244) <= layer0_outputs(1169);
    outputs(2245) <= not(layer0_outputs(4642)) or (layer0_outputs(6248));
    outputs(2246) <= not(layer0_outputs(900));
    outputs(2247) <= not(layer0_outputs(804)) or (layer0_outputs(9134));
    outputs(2248) <= (layer0_outputs(6134)) or (layer0_outputs(527));
    outputs(2249) <= (layer0_outputs(3095)) and (layer0_outputs(10219));
    outputs(2250) <= not((layer0_outputs(1030)) xor (layer0_outputs(7979)));
    outputs(2251) <= not(layer0_outputs(2939));
    outputs(2252) <= not(layer0_outputs(530));
    outputs(2253) <= not((layer0_outputs(7504)) and (layer0_outputs(204)));
    outputs(2254) <= layer0_outputs(8122);
    outputs(2255) <= not(layer0_outputs(3259));
    outputs(2256) <= not(layer0_outputs(5220));
    outputs(2257) <= layer0_outputs(407);
    outputs(2258) <= (layer0_outputs(7072)) xor (layer0_outputs(7786));
    outputs(2259) <= layer0_outputs(4575);
    outputs(2260) <= (layer0_outputs(9013)) or (layer0_outputs(5143));
    outputs(2261) <= (layer0_outputs(5448)) and (layer0_outputs(7524));
    outputs(2262) <= not(layer0_outputs(2282));
    outputs(2263) <= layer0_outputs(60);
    outputs(2264) <= not(layer0_outputs(3467));
    outputs(2265) <= (layer0_outputs(5308)) xor (layer0_outputs(549));
    outputs(2266) <= (layer0_outputs(7354)) xor (layer0_outputs(5942));
    outputs(2267) <= not(layer0_outputs(7748));
    outputs(2268) <= not((layer0_outputs(5754)) and (layer0_outputs(17)));
    outputs(2269) <= layer0_outputs(7281);
    outputs(2270) <= (layer0_outputs(4014)) and (layer0_outputs(7554));
    outputs(2271) <= (layer0_outputs(4224)) xor (layer0_outputs(1186));
    outputs(2272) <= not((layer0_outputs(7347)) or (layer0_outputs(118)));
    outputs(2273) <= layer0_outputs(8678);
    outputs(2274) <= not(layer0_outputs(5859));
    outputs(2275) <= (layer0_outputs(8373)) and not (layer0_outputs(4951));
    outputs(2276) <= not(layer0_outputs(9189));
    outputs(2277) <= not((layer0_outputs(2139)) xor (layer0_outputs(4615)));
    outputs(2278) <= layer0_outputs(1139);
    outputs(2279) <= not(layer0_outputs(9724)) or (layer0_outputs(370));
    outputs(2280) <= (layer0_outputs(8829)) xor (layer0_outputs(6361));
    outputs(2281) <= not(layer0_outputs(9223)) or (layer0_outputs(1299));
    outputs(2282) <= layer0_outputs(8613);
    outputs(2283) <= not(layer0_outputs(2997));
    outputs(2284) <= not(layer0_outputs(4071));
    outputs(2285) <= not(layer0_outputs(532));
    outputs(2286) <= not(layer0_outputs(3527));
    outputs(2287) <= (layer0_outputs(240)) and not (layer0_outputs(6232));
    outputs(2288) <= layer0_outputs(5067);
    outputs(2289) <= not((layer0_outputs(10043)) and (layer0_outputs(7779)));
    outputs(2290) <= not(layer0_outputs(2398));
    outputs(2291) <= (layer0_outputs(8497)) xor (layer0_outputs(4561));
    outputs(2292) <= layer0_outputs(1925);
    outputs(2293) <= not(layer0_outputs(5713));
    outputs(2294) <= not(layer0_outputs(9828));
    outputs(2295) <= layer0_outputs(8730);
    outputs(2296) <= not(layer0_outputs(9721)) or (layer0_outputs(9965));
    outputs(2297) <= not(layer0_outputs(8820));
    outputs(2298) <= layer0_outputs(3827);
    outputs(2299) <= (layer0_outputs(5716)) xor (layer0_outputs(6468));
    outputs(2300) <= not(layer0_outputs(10016)) or (layer0_outputs(6992));
    outputs(2301) <= not(layer0_outputs(3044)) or (layer0_outputs(3679));
    outputs(2302) <= (layer0_outputs(1647)) and not (layer0_outputs(8755));
    outputs(2303) <= not(layer0_outputs(9283)) or (layer0_outputs(858));
    outputs(2304) <= layer0_outputs(4391);
    outputs(2305) <= not((layer0_outputs(7311)) or (layer0_outputs(7534)));
    outputs(2306) <= layer0_outputs(5672);
    outputs(2307) <= (layer0_outputs(9900)) and not (layer0_outputs(5551));
    outputs(2308) <= (layer0_outputs(3897)) and not (layer0_outputs(10015));
    outputs(2309) <= not((layer0_outputs(6449)) xor (layer0_outputs(6437)));
    outputs(2310) <= layer0_outputs(880);
    outputs(2311) <= (layer0_outputs(6130)) and not (layer0_outputs(4045));
    outputs(2312) <= (layer0_outputs(9881)) and not (layer0_outputs(194));
    outputs(2313) <= not((layer0_outputs(5071)) and (layer0_outputs(3052)));
    outputs(2314) <= not(layer0_outputs(5485));
    outputs(2315) <= not(layer0_outputs(5229)) or (layer0_outputs(8866));
    outputs(2316) <= not(layer0_outputs(3838)) or (layer0_outputs(8188));
    outputs(2317) <= not(layer0_outputs(2806));
    outputs(2318) <= layer0_outputs(4829);
    outputs(2319) <= not(layer0_outputs(1279));
    outputs(2320) <= layer0_outputs(9262);
    outputs(2321) <= (layer0_outputs(1871)) xor (layer0_outputs(9037));
    outputs(2322) <= layer0_outputs(2747);
    outputs(2323) <= (layer0_outputs(761)) and not (layer0_outputs(4757));
    outputs(2324) <= not((layer0_outputs(621)) or (layer0_outputs(1218)));
    outputs(2325) <= not(layer0_outputs(8056)) or (layer0_outputs(5297));
    outputs(2326) <= not(layer0_outputs(4848));
    outputs(2327) <= not(layer0_outputs(233));
    outputs(2328) <= not((layer0_outputs(4033)) or (layer0_outputs(6554)));
    outputs(2329) <= not(layer0_outputs(3541)) or (layer0_outputs(4306));
    outputs(2330) <= not((layer0_outputs(3162)) or (layer0_outputs(8152)));
    outputs(2331) <= not(layer0_outputs(3872)) or (layer0_outputs(3669));
    outputs(2332) <= not(layer0_outputs(7528));
    outputs(2333) <= layer0_outputs(7934);
    outputs(2334) <= not((layer0_outputs(7473)) or (layer0_outputs(2287)));
    outputs(2335) <= not(layer0_outputs(4709)) or (layer0_outputs(1637));
    outputs(2336) <= layer0_outputs(3248);
    outputs(2337) <= (layer0_outputs(3307)) xor (layer0_outputs(336));
    outputs(2338) <= not((layer0_outputs(7142)) or (layer0_outputs(531)));
    outputs(2339) <= not(layer0_outputs(1265));
    outputs(2340) <= layer0_outputs(3897);
    outputs(2341) <= layer0_outputs(7512);
    outputs(2342) <= not((layer0_outputs(2949)) xor (layer0_outputs(1263)));
    outputs(2343) <= not((layer0_outputs(5204)) or (layer0_outputs(6569)));
    outputs(2344) <= layer0_outputs(1707);
    outputs(2345) <= layer0_outputs(1105);
    outputs(2346) <= (layer0_outputs(8841)) or (layer0_outputs(8599));
    outputs(2347) <= layer0_outputs(1145);
    outputs(2348) <= not((layer0_outputs(5821)) or (layer0_outputs(9080)));
    outputs(2349) <= not(layer0_outputs(9759));
    outputs(2350) <= layer0_outputs(5400);
    outputs(2351) <= not((layer0_outputs(3550)) and (layer0_outputs(4545)));
    outputs(2352) <= not(layer0_outputs(699));
    outputs(2353) <= layer0_outputs(8099);
    outputs(2354) <= not((layer0_outputs(6620)) and (layer0_outputs(3896)));
    outputs(2355) <= not(layer0_outputs(5814));
    outputs(2356) <= layer0_outputs(6144);
    outputs(2357) <= not(layer0_outputs(6346)) or (layer0_outputs(4691));
    outputs(2358) <= layer0_outputs(573);
    outputs(2359) <= layer0_outputs(7162);
    outputs(2360) <= layer0_outputs(623);
    outputs(2361) <= (layer0_outputs(5806)) and (layer0_outputs(9780));
    outputs(2362) <= (layer0_outputs(9511)) xor (layer0_outputs(9229));
    outputs(2363) <= (layer0_outputs(1476)) or (layer0_outputs(7361));
    outputs(2364) <= layer0_outputs(7464);
    outputs(2365) <= (layer0_outputs(5312)) and not (layer0_outputs(1432));
    outputs(2366) <= layer0_outputs(7202);
    outputs(2367) <= (layer0_outputs(10077)) and not (layer0_outputs(3134));
    outputs(2368) <= (layer0_outputs(5109)) and not (layer0_outputs(8916));
    outputs(2369) <= layer0_outputs(7466);
    outputs(2370) <= not((layer0_outputs(5364)) xor (layer0_outputs(1277)));
    outputs(2371) <= not((layer0_outputs(5852)) xor (layer0_outputs(2694)));
    outputs(2372) <= layer0_outputs(7290);
    outputs(2373) <= not(layer0_outputs(4019));
    outputs(2374) <= layer0_outputs(1769);
    outputs(2375) <= not(layer0_outputs(6788));
    outputs(2376) <= (layer0_outputs(4927)) and (layer0_outputs(4028));
    outputs(2377) <= (layer0_outputs(4281)) and not (layer0_outputs(7941));
    outputs(2378) <= (layer0_outputs(5865)) or (layer0_outputs(1934));
    outputs(2379) <= not((layer0_outputs(6865)) xor (layer0_outputs(10232)));
    outputs(2380) <= (layer0_outputs(10226)) and (layer0_outputs(9127));
    outputs(2381) <= (layer0_outputs(859)) xor (layer0_outputs(478));
    outputs(2382) <= layer0_outputs(8475);
    outputs(2383) <= (layer0_outputs(6017)) and not (layer0_outputs(9910));
    outputs(2384) <= not(layer0_outputs(6253));
    outputs(2385) <= not(layer0_outputs(4077)) or (layer0_outputs(6822));
    outputs(2386) <= (layer0_outputs(2518)) xor (layer0_outputs(492));
    outputs(2387) <= not(layer0_outputs(8947));
    outputs(2388) <= layer0_outputs(8523);
    outputs(2389) <= layer0_outputs(1164);
    outputs(2390) <= (layer0_outputs(8323)) xor (layer0_outputs(2274));
    outputs(2391) <= (layer0_outputs(1591)) or (layer0_outputs(1112));
    outputs(2392) <= (layer0_outputs(7365)) and not (layer0_outputs(7082));
    outputs(2393) <= not((layer0_outputs(6772)) and (layer0_outputs(5456)));
    outputs(2394) <= (layer0_outputs(4444)) xor (layer0_outputs(593));
    outputs(2395) <= layer0_outputs(5645);
    outputs(2396) <= layer0_outputs(6877);
    outputs(2397) <= not((layer0_outputs(3956)) or (layer0_outputs(2951)));
    outputs(2398) <= not(layer0_outputs(1184));
    outputs(2399) <= (layer0_outputs(5806)) and not (layer0_outputs(8310));
    outputs(2400) <= not(layer0_outputs(7042)) or (layer0_outputs(6447));
    outputs(2401) <= not(layer0_outputs(925));
    outputs(2402) <= not((layer0_outputs(932)) or (layer0_outputs(7824)));
    outputs(2403) <= not(layer0_outputs(6993)) or (layer0_outputs(8555));
    outputs(2404) <= not((layer0_outputs(4496)) xor (layer0_outputs(4515)));
    outputs(2405) <= not((layer0_outputs(1052)) and (layer0_outputs(6909)));
    outputs(2406) <= not(layer0_outputs(3403));
    outputs(2407) <= layer0_outputs(935);
    outputs(2408) <= not((layer0_outputs(1536)) xor (layer0_outputs(5379)));
    outputs(2409) <= layer0_outputs(8705);
    outputs(2410) <= not((layer0_outputs(4019)) xor (layer0_outputs(9784)));
    outputs(2411) <= (layer0_outputs(7444)) and (layer0_outputs(9706));
    outputs(2412) <= (layer0_outputs(2501)) and not (layer0_outputs(5900));
    outputs(2413) <= not((layer0_outputs(1314)) xor (layer0_outputs(1606)));
    outputs(2414) <= not((layer0_outputs(7721)) or (layer0_outputs(7762)));
    outputs(2415) <= not((layer0_outputs(7301)) or (layer0_outputs(8996)));
    outputs(2416) <= not(layer0_outputs(10227)) or (layer0_outputs(44));
    outputs(2417) <= not(layer0_outputs(2590));
    outputs(2418) <= (layer0_outputs(6675)) and not (layer0_outputs(4867));
    outputs(2419) <= not((layer0_outputs(3188)) and (layer0_outputs(3487)));
    outputs(2420) <= not((layer0_outputs(4650)) xor (layer0_outputs(5921)));
    outputs(2421) <= (layer0_outputs(3887)) or (layer0_outputs(9853));
    outputs(2422) <= not(layer0_outputs(8964));
    outputs(2423) <= not((layer0_outputs(7807)) or (layer0_outputs(7340)));
    outputs(2424) <= layer0_outputs(8416);
    outputs(2425) <= not((layer0_outputs(8222)) xor (layer0_outputs(42)));
    outputs(2426) <= (layer0_outputs(3298)) xor (layer0_outputs(4262));
    outputs(2427) <= not(layer0_outputs(5718));
    outputs(2428) <= (layer0_outputs(744)) and not (layer0_outputs(8538));
    outputs(2429) <= not(layer0_outputs(3924));
    outputs(2430) <= layer0_outputs(9971);
    outputs(2431) <= (layer0_outputs(158)) and not (layer0_outputs(1914));
    outputs(2432) <= layer0_outputs(8902);
    outputs(2433) <= not((layer0_outputs(3943)) or (layer0_outputs(490)));
    outputs(2434) <= not((layer0_outputs(7478)) and (layer0_outputs(6606)));
    outputs(2435) <= not(layer0_outputs(998));
    outputs(2436) <= not(layer0_outputs(4280)) or (layer0_outputs(7954));
    outputs(2437) <= not((layer0_outputs(7791)) xor (layer0_outputs(1985)));
    outputs(2438) <= not(layer0_outputs(975));
    outputs(2439) <= not(layer0_outputs(2739));
    outputs(2440) <= (layer0_outputs(9913)) or (layer0_outputs(6281));
    outputs(2441) <= layer0_outputs(6124);
    outputs(2442) <= not(layer0_outputs(3131)) or (layer0_outputs(4304));
    outputs(2443) <= not((layer0_outputs(5263)) or (layer0_outputs(3940)));
    outputs(2444) <= not((layer0_outputs(4670)) or (layer0_outputs(9209)));
    outputs(2445) <= not(layer0_outputs(9103));
    outputs(2446) <= not(layer0_outputs(9426));
    outputs(2447) <= not(layer0_outputs(7635)) or (layer0_outputs(6953));
    outputs(2448) <= (layer0_outputs(9077)) and not (layer0_outputs(9389));
    outputs(2449) <= not((layer0_outputs(8137)) and (layer0_outputs(4523)));
    outputs(2450) <= (layer0_outputs(7505)) xor (layer0_outputs(3462));
    outputs(2451) <= not(layer0_outputs(2198)) or (layer0_outputs(5740));
    outputs(2452) <= not(layer0_outputs(3614)) or (layer0_outputs(8280));
    outputs(2453) <= not((layer0_outputs(3555)) xor (layer0_outputs(2070)));
    outputs(2454) <= not((layer0_outputs(1196)) or (layer0_outputs(1157)));
    outputs(2455) <= not(layer0_outputs(7248)) or (layer0_outputs(1070));
    outputs(2456) <= not(layer0_outputs(8098)) or (layer0_outputs(6944));
    outputs(2457) <= not(layer0_outputs(7952));
    outputs(2458) <= (layer0_outputs(8775)) and (layer0_outputs(8663));
    outputs(2459) <= not(layer0_outputs(5896));
    outputs(2460) <= (layer0_outputs(2588)) and not (layer0_outputs(3033));
    outputs(2461) <= (layer0_outputs(5749)) and not (layer0_outputs(8646));
    outputs(2462) <= layer0_outputs(935);
    outputs(2463) <= not(layer0_outputs(8273)) or (layer0_outputs(4798));
    outputs(2464) <= not(layer0_outputs(4665));
    outputs(2465) <= not(layer0_outputs(2889));
    outputs(2466) <= (layer0_outputs(5583)) xor (layer0_outputs(5352));
    outputs(2467) <= layer0_outputs(297);
    outputs(2468) <= layer0_outputs(1173);
    outputs(2469) <= not(layer0_outputs(8039)) or (layer0_outputs(4780));
    outputs(2470) <= not(layer0_outputs(5895)) or (layer0_outputs(3597));
    outputs(2471) <= layer0_outputs(1701);
    outputs(2472) <= (layer0_outputs(1782)) xor (layer0_outputs(5746));
    outputs(2473) <= not((layer0_outputs(8699)) or (layer0_outputs(5101)));
    outputs(2474) <= (layer0_outputs(4404)) or (layer0_outputs(9742));
    outputs(2475) <= not(layer0_outputs(5245));
    outputs(2476) <= layer0_outputs(7913);
    outputs(2477) <= not((layer0_outputs(2682)) and (layer0_outputs(1926)));
    outputs(2478) <= layer0_outputs(2004);
    outputs(2479) <= (layer0_outputs(86)) and (layer0_outputs(2438));
    outputs(2480) <= layer0_outputs(9922);
    outputs(2481) <= layer0_outputs(6285);
    outputs(2482) <= (layer0_outputs(9078)) and not (layer0_outputs(6959));
    outputs(2483) <= layer0_outputs(9443);
    outputs(2484) <= not((layer0_outputs(115)) xor (layer0_outputs(4022)));
    outputs(2485) <= not(layer0_outputs(8764));
    outputs(2486) <= layer0_outputs(7207);
    outputs(2487) <= layer0_outputs(894);
    outputs(2488) <= (layer0_outputs(7253)) and not (layer0_outputs(4967));
    outputs(2489) <= layer0_outputs(418);
    outputs(2490) <= not(layer0_outputs(6301));
    outputs(2491) <= not(layer0_outputs(7117)) or (layer0_outputs(9566));
    outputs(2492) <= layer0_outputs(691);
    outputs(2493) <= (layer0_outputs(3015)) or (layer0_outputs(9649));
    outputs(2494) <= layer0_outputs(8785);
    outputs(2495) <= not(layer0_outputs(857)) or (layer0_outputs(8854));
    outputs(2496) <= (layer0_outputs(2397)) xor (layer0_outputs(5210));
    outputs(2497) <= not((layer0_outputs(3361)) xor (layer0_outputs(3207)));
    outputs(2498) <= layer0_outputs(491);
    outputs(2499) <= (layer0_outputs(6080)) and (layer0_outputs(5510));
    outputs(2500) <= (layer0_outputs(6304)) or (layer0_outputs(5244));
    outputs(2501) <= not(layer0_outputs(3577)) or (layer0_outputs(2145));
    outputs(2502) <= (layer0_outputs(1509)) xor (layer0_outputs(10084));
    outputs(2503) <= (layer0_outputs(5270)) xor (layer0_outputs(10191));
    outputs(2504) <= not(layer0_outputs(4973));
    outputs(2505) <= layer0_outputs(5233);
    outputs(2506) <= layer0_outputs(3166);
    outputs(2507) <= not(layer0_outputs(9946));
    outputs(2508) <= not(layer0_outputs(5848));
    outputs(2509) <= not((layer0_outputs(9499)) and (layer0_outputs(9387)));
    outputs(2510) <= (layer0_outputs(1772)) and not (layer0_outputs(10143));
    outputs(2511) <= not((layer0_outputs(3868)) xor (layer0_outputs(9723)));
    outputs(2512) <= layer0_outputs(7382);
    outputs(2513) <= layer0_outputs(497);
    outputs(2514) <= not((layer0_outputs(9949)) and (layer0_outputs(8076)));
    outputs(2515) <= not(layer0_outputs(1265));
    outputs(2516) <= layer0_outputs(2001);
    outputs(2517) <= layer0_outputs(4242);
    outputs(2518) <= not((layer0_outputs(1067)) xor (layer0_outputs(8133)));
    outputs(2519) <= not(layer0_outputs(9733));
    outputs(2520) <= (layer0_outputs(6674)) xor (layer0_outputs(6003));
    outputs(2521) <= not(layer0_outputs(3108));
    outputs(2522) <= not(layer0_outputs(9524));
    outputs(2523) <= not(layer0_outputs(342));
    outputs(2524) <= (layer0_outputs(8855)) and not (layer0_outputs(5082));
    outputs(2525) <= layer0_outputs(5938);
    outputs(2526) <= not(layer0_outputs(3853));
    outputs(2527) <= (layer0_outputs(5810)) and (layer0_outputs(5449));
    outputs(2528) <= not(layer0_outputs(5848)) or (layer0_outputs(1917));
    outputs(2529) <= layer0_outputs(1293);
    outputs(2530) <= (layer0_outputs(4782)) xor (layer0_outputs(6181));
    outputs(2531) <= layer0_outputs(526);
    outputs(2532) <= not((layer0_outputs(3142)) xor (layer0_outputs(6451)));
    outputs(2533) <= not((layer0_outputs(8397)) and (layer0_outputs(5689)));
    outputs(2534) <= layer0_outputs(4765);
    outputs(2535) <= layer0_outputs(3122);
    outputs(2536) <= layer0_outputs(440);
    outputs(2537) <= not(layer0_outputs(3389));
    outputs(2538) <= not((layer0_outputs(3423)) xor (layer0_outputs(8228)));
    outputs(2539) <= not(layer0_outputs(8878));
    outputs(2540) <= (layer0_outputs(8727)) xor (layer0_outputs(7403));
    outputs(2541) <= not(layer0_outputs(2555));
    outputs(2542) <= (layer0_outputs(8810)) or (layer0_outputs(426));
    outputs(2543) <= (layer0_outputs(3226)) xor (layer0_outputs(4060));
    outputs(2544) <= not(layer0_outputs(1304)) or (layer0_outputs(10184));
    outputs(2545) <= (layer0_outputs(8918)) xor (layer0_outputs(9266));
    outputs(2546) <= not((layer0_outputs(8668)) xor (layer0_outputs(1796)));
    outputs(2547) <= layer0_outputs(7599);
    outputs(2548) <= not(layer0_outputs(7522));
    outputs(2549) <= not(layer0_outputs(6709));
    outputs(2550) <= (layer0_outputs(5239)) and not (layer0_outputs(6193));
    outputs(2551) <= (layer0_outputs(9969)) and not (layer0_outputs(7841));
    outputs(2552) <= not(layer0_outputs(1718));
    outputs(2553) <= (layer0_outputs(6848)) xor (layer0_outputs(5872));
    outputs(2554) <= not((layer0_outputs(2815)) xor (layer0_outputs(9346)));
    outputs(2555) <= not((layer0_outputs(9602)) and (layer0_outputs(7404)));
    outputs(2556) <= '1';
    outputs(2557) <= not((layer0_outputs(4574)) and (layer0_outputs(6174)));
    outputs(2558) <= layer0_outputs(5199);
    outputs(2559) <= not((layer0_outputs(4175)) xor (layer0_outputs(8627)));
    outputs(2560) <= layer0_outputs(3109);
    outputs(2561) <= not((layer0_outputs(5406)) or (layer0_outputs(1386)));
    outputs(2562) <= (layer0_outputs(1869)) and not (layer0_outputs(5555));
    outputs(2563) <= (layer0_outputs(4579)) or (layer0_outputs(7198));
    outputs(2564) <= not(layer0_outputs(2370)) or (layer0_outputs(3302));
    outputs(2565) <= not((layer0_outputs(7902)) xor (layer0_outputs(7828)));
    outputs(2566) <= layer0_outputs(1207);
    outputs(2567) <= (layer0_outputs(6285)) and (layer0_outputs(9854));
    outputs(2568) <= not(layer0_outputs(3064));
    outputs(2569) <= not(layer0_outputs(5572)) or (layer0_outputs(8930));
    outputs(2570) <= not((layer0_outputs(7655)) xor (layer0_outputs(4084)));
    outputs(2571) <= (layer0_outputs(8531)) and not (layer0_outputs(132));
    outputs(2572) <= (layer0_outputs(3845)) and not (layer0_outputs(9938));
    outputs(2573) <= layer0_outputs(8454);
    outputs(2574) <= not(layer0_outputs(6067));
    outputs(2575) <= (layer0_outputs(8019)) and not (layer0_outputs(2585));
    outputs(2576) <= layer0_outputs(8650);
    outputs(2577) <= not((layer0_outputs(8157)) and (layer0_outputs(2944)));
    outputs(2578) <= not(layer0_outputs(4405));
    outputs(2579) <= (layer0_outputs(9091)) and not (layer0_outputs(2896));
    outputs(2580) <= layer0_outputs(9380);
    outputs(2581) <= (layer0_outputs(4081)) xor (layer0_outputs(4257));
    outputs(2582) <= not(layer0_outputs(3621)) or (layer0_outputs(4586));
    outputs(2583) <= layer0_outputs(8915);
    outputs(2584) <= (layer0_outputs(6318)) or (layer0_outputs(9306));
    outputs(2585) <= layer0_outputs(8609);
    outputs(2586) <= not(layer0_outputs(5496));
    outputs(2587) <= (layer0_outputs(6793)) or (layer0_outputs(2075));
    outputs(2588) <= (layer0_outputs(1373)) or (layer0_outputs(7380));
    outputs(2589) <= not((layer0_outputs(2439)) xor (layer0_outputs(1190)));
    outputs(2590) <= not(layer0_outputs(5035)) or (layer0_outputs(8342));
    outputs(2591) <= (layer0_outputs(1462)) or (layer0_outputs(1112));
    outputs(2592) <= not(layer0_outputs(7031)) or (layer0_outputs(9394));
    outputs(2593) <= (layer0_outputs(5447)) or (layer0_outputs(1525));
    outputs(2594) <= layer0_outputs(5454);
    outputs(2595) <= layer0_outputs(6145);
    outputs(2596) <= not(layer0_outputs(5994));
    outputs(2597) <= layer0_outputs(5948);
    outputs(2598) <= not(layer0_outputs(2899)) or (layer0_outputs(8122));
    outputs(2599) <= not((layer0_outputs(2867)) and (layer0_outputs(2607)));
    outputs(2600) <= not((layer0_outputs(3797)) and (layer0_outputs(3994)));
    outputs(2601) <= not((layer0_outputs(5561)) and (layer0_outputs(2293)));
    outputs(2602) <= not((layer0_outputs(2546)) or (layer0_outputs(284)));
    outputs(2603) <= not(layer0_outputs(8452));
    outputs(2604) <= not(layer0_outputs(9476)) or (layer0_outputs(9893));
    outputs(2605) <= layer0_outputs(104);
    outputs(2606) <= not((layer0_outputs(4862)) xor (layer0_outputs(6613)));
    outputs(2607) <= not((layer0_outputs(7768)) and (layer0_outputs(9840)));
    outputs(2608) <= not((layer0_outputs(9874)) xor (layer0_outputs(1669)));
    outputs(2609) <= (layer0_outputs(1745)) and (layer0_outputs(9311));
    outputs(2610) <= (layer0_outputs(8673)) or (layer0_outputs(4947));
    outputs(2611) <= (layer0_outputs(5971)) and (layer0_outputs(1884));
    outputs(2612) <= not(layer0_outputs(5320));
    outputs(2613) <= not(layer0_outputs(4713));
    outputs(2614) <= not(layer0_outputs(8461));
    outputs(2615) <= (layer0_outputs(942)) or (layer0_outputs(9958));
    outputs(2616) <= not(layer0_outputs(3601));
    outputs(2617) <= not(layer0_outputs(720));
    outputs(2618) <= not((layer0_outputs(1003)) or (layer0_outputs(10042)));
    outputs(2619) <= layer0_outputs(6711);
    outputs(2620) <= not((layer0_outputs(4977)) xor (layer0_outputs(9218)));
    outputs(2621) <= not(layer0_outputs(842)) or (layer0_outputs(6714));
    outputs(2622) <= not(layer0_outputs(8762)) or (layer0_outputs(4189));
    outputs(2623) <= not((layer0_outputs(9413)) and (layer0_outputs(4408)));
    outputs(2624) <= (layer0_outputs(6755)) and not (layer0_outputs(2038));
    outputs(2625) <= not(layer0_outputs(9828));
    outputs(2626) <= (layer0_outputs(9643)) and not (layer0_outputs(9231));
    outputs(2627) <= (layer0_outputs(3343)) and not (layer0_outputs(6787));
    outputs(2628) <= (layer0_outputs(5578)) xor (layer0_outputs(2068));
    outputs(2629) <= not((layer0_outputs(9092)) and (layer0_outputs(7107)));
    outputs(2630) <= layer0_outputs(222);
    outputs(2631) <= layer0_outputs(683);
    outputs(2632) <= layer0_outputs(7967);
    outputs(2633) <= not(layer0_outputs(5863)) or (layer0_outputs(2240));
    outputs(2634) <= not(layer0_outputs(3789));
    outputs(2635) <= not(layer0_outputs(624));
    outputs(2636) <= not(layer0_outputs(6733));
    outputs(2637) <= not((layer0_outputs(8429)) or (layer0_outputs(7543)));
    outputs(2638) <= not(layer0_outputs(9194)) or (layer0_outputs(9972));
    outputs(2639) <= not((layer0_outputs(7147)) and (layer0_outputs(4787)));
    outputs(2640) <= not(layer0_outputs(7414));
    outputs(2641) <= not(layer0_outputs(8948)) or (layer0_outputs(5070));
    outputs(2642) <= not(layer0_outputs(10065));
    outputs(2643) <= layer0_outputs(3723);
    outputs(2644) <= (layer0_outputs(1400)) xor (layer0_outputs(346));
    outputs(2645) <= layer0_outputs(1024);
    outputs(2646) <= (layer0_outputs(3611)) and not (layer0_outputs(9595));
    outputs(2647) <= not((layer0_outputs(4327)) or (layer0_outputs(9565)));
    outputs(2648) <= layer0_outputs(10215);
    outputs(2649) <= not((layer0_outputs(4630)) xor (layer0_outputs(6098)));
    outputs(2650) <= (layer0_outputs(6935)) and not (layer0_outputs(4165));
    outputs(2651) <= layer0_outputs(6372);
    outputs(2652) <= layer0_outputs(8801);
    outputs(2653) <= (layer0_outputs(1256)) and (layer0_outputs(6089));
    outputs(2654) <= (layer0_outputs(6634)) and (layer0_outputs(5957));
    outputs(2655) <= (layer0_outputs(6648)) or (layer0_outputs(7495));
    outputs(2656) <= (layer0_outputs(2592)) and not (layer0_outputs(4632));
    outputs(2657) <= layer0_outputs(2569);
    outputs(2658) <= (layer0_outputs(182)) xor (layer0_outputs(9055));
    outputs(2659) <= (layer0_outputs(1188)) xor (layer0_outputs(4219));
    outputs(2660) <= not(layer0_outputs(2104)) or (layer0_outputs(443));
    outputs(2661) <= (layer0_outputs(5746)) and not (layer0_outputs(2053));
    outputs(2662) <= not(layer0_outputs(2260)) or (layer0_outputs(1860));
    outputs(2663) <= not(layer0_outputs(2205));
    outputs(2664) <= not(layer0_outputs(80));
    outputs(2665) <= layer0_outputs(3519);
    outputs(2666) <= not(layer0_outputs(5098));
    outputs(2667) <= (layer0_outputs(8121)) xor (layer0_outputs(3053));
    outputs(2668) <= (layer0_outputs(4006)) xor (layer0_outputs(2665));
    outputs(2669) <= not(layer0_outputs(9001)) or (layer0_outputs(6326));
    outputs(2670) <= not(layer0_outputs(522));
    outputs(2671) <= (layer0_outputs(5419)) and (layer0_outputs(8619));
    outputs(2672) <= not(layer0_outputs(9884));
    outputs(2673) <= not((layer0_outputs(6777)) xor (layer0_outputs(5833)));
    outputs(2674) <= (layer0_outputs(6917)) xor (layer0_outputs(877));
    outputs(2675) <= layer0_outputs(7467);
    outputs(2676) <= layer0_outputs(9263);
    outputs(2677) <= (layer0_outputs(7203)) or (layer0_outputs(2626));
    outputs(2678) <= not((layer0_outputs(6991)) or (layer0_outputs(3549)));
    outputs(2679) <= not((layer0_outputs(2205)) and (layer0_outputs(5669)));
    outputs(2680) <= layer0_outputs(4188);
    outputs(2681) <= (layer0_outputs(6213)) xor (layer0_outputs(7542));
    outputs(2682) <= not(layer0_outputs(921)) or (layer0_outputs(3676));
    outputs(2683) <= layer0_outputs(940);
    outputs(2684) <= (layer0_outputs(3015)) xor (layer0_outputs(3431));
    outputs(2685) <= not(layer0_outputs(7995)) or (layer0_outputs(6026));
    outputs(2686) <= not(layer0_outputs(9257)) or (layer0_outputs(8378));
    outputs(2687) <= not((layer0_outputs(3127)) or (layer0_outputs(2466)));
    outputs(2688) <= layer0_outputs(8544);
    outputs(2689) <= not(layer0_outputs(2686));
    outputs(2690) <= not(layer0_outputs(2647));
    outputs(2691) <= not(layer0_outputs(5361));
    outputs(2692) <= (layer0_outputs(7708)) xor (layer0_outputs(2474));
    outputs(2693) <= not(layer0_outputs(7089)) or (layer0_outputs(5866));
    outputs(2694) <= not(layer0_outputs(6673)) or (layer0_outputs(7862));
    outputs(2695) <= not(layer0_outputs(4380)) or (layer0_outputs(8186));
    outputs(2696) <= not(layer0_outputs(5077)) or (layer0_outputs(6317));
    outputs(2697) <= (layer0_outputs(6824)) xor (layer0_outputs(4208));
    outputs(2698) <= layer0_outputs(1723);
    outputs(2699) <= layer0_outputs(7390);
    outputs(2700) <= not(layer0_outputs(1802));
    outputs(2701) <= not((layer0_outputs(675)) xor (layer0_outputs(7054)));
    outputs(2702) <= not(layer0_outputs(6932));
    outputs(2703) <= layer0_outputs(8438);
    outputs(2704) <= not(layer0_outputs(6239)) or (layer0_outputs(1187));
    outputs(2705) <= not((layer0_outputs(9560)) or (layer0_outputs(2864)));
    outputs(2706) <= not(layer0_outputs(5941)) or (layer0_outputs(1038));
    outputs(2707) <= not((layer0_outputs(848)) and (layer0_outputs(7038)));
    outputs(2708) <= not(layer0_outputs(1877));
    outputs(2709) <= (layer0_outputs(8981)) xor (layer0_outputs(8751));
    outputs(2710) <= layer0_outputs(5911);
    outputs(2711) <= not((layer0_outputs(9837)) or (layer0_outputs(6276)));
    outputs(2712) <= not((layer0_outputs(246)) xor (layer0_outputs(3094)));
    outputs(2713) <= not(layer0_outputs(3398)) or (layer0_outputs(1872));
    outputs(2714) <= (layer0_outputs(482)) or (layer0_outputs(5451));
    outputs(2715) <= not(layer0_outputs(2271));
    outputs(2716) <= (layer0_outputs(3305)) or (layer0_outputs(1038));
    outputs(2717) <= not(layer0_outputs(9076));
    outputs(2718) <= not((layer0_outputs(9625)) and (layer0_outputs(6988)));
    outputs(2719) <= layer0_outputs(3217);
    outputs(2720) <= not(layer0_outputs(4589));
    outputs(2721) <= not(layer0_outputs(7073));
    outputs(2722) <= layer0_outputs(8709);
    outputs(2723) <= (layer0_outputs(1890)) and (layer0_outputs(81));
    outputs(2724) <= not(layer0_outputs(3936)) or (layer0_outputs(7629));
    outputs(2725) <= not((layer0_outputs(1171)) and (layer0_outputs(9985)));
    outputs(2726) <= not((layer0_outputs(10231)) and (layer0_outputs(3179)));
    outputs(2727) <= (layer0_outputs(6145)) and not (layer0_outputs(2271));
    outputs(2728) <= not((layer0_outputs(649)) xor (layer0_outputs(6349)));
    outputs(2729) <= layer0_outputs(9967);
    outputs(2730) <= not((layer0_outputs(516)) and (layer0_outputs(4265)));
    outputs(2731) <= layer0_outputs(6021);
    outputs(2732) <= not((layer0_outputs(3923)) xor (layer0_outputs(3456)));
    outputs(2733) <= not((layer0_outputs(112)) xor (layer0_outputs(7964)));
    outputs(2734) <= not(layer0_outputs(4064));
    outputs(2735) <= (layer0_outputs(4360)) xor (layer0_outputs(2883));
    outputs(2736) <= layer0_outputs(3666);
    outputs(2737) <= not((layer0_outputs(5711)) or (layer0_outputs(8726)));
    outputs(2738) <= (layer0_outputs(5601)) and (layer0_outputs(9865));
    outputs(2739) <= (layer0_outputs(3858)) and not (layer0_outputs(4376));
    outputs(2740) <= not(layer0_outputs(3434)) or (layer0_outputs(392));
    outputs(2741) <= layer0_outputs(2556);
    outputs(2742) <= not(layer0_outputs(4318));
    outputs(2743) <= layer0_outputs(2443);
    outputs(2744) <= not(layer0_outputs(9666));
    outputs(2745) <= not((layer0_outputs(6393)) xor (layer0_outputs(8409)));
    outputs(2746) <= not((layer0_outputs(1803)) xor (layer0_outputs(8672)));
    outputs(2747) <= layer0_outputs(4651);
    outputs(2748) <= not((layer0_outputs(9624)) xor (layer0_outputs(4678)));
    outputs(2749) <= not(layer0_outputs(1740));
    outputs(2750) <= (layer0_outputs(7665)) and not (layer0_outputs(2148));
    outputs(2751) <= layer0_outputs(2257);
    outputs(2752) <= not((layer0_outputs(3859)) and (layer0_outputs(10100)));
    outputs(2753) <= not((layer0_outputs(6520)) xor (layer0_outputs(9268)));
    outputs(2754) <= not((layer0_outputs(6841)) and (layer0_outputs(3955)));
    outputs(2755) <= (layer0_outputs(4343)) xor (layer0_outputs(4162));
    outputs(2756) <= (layer0_outputs(10022)) and (layer0_outputs(2419));
    outputs(2757) <= not(layer0_outputs(4338));
    outputs(2758) <= not(layer0_outputs(2724));
    outputs(2759) <= not(layer0_outputs(6386)) or (layer0_outputs(4401));
    outputs(2760) <= layer0_outputs(9908);
    outputs(2761) <= not((layer0_outputs(7822)) and (layer0_outputs(2587)));
    outputs(2762) <= not(layer0_outputs(9746)) or (layer0_outputs(4258));
    outputs(2763) <= not((layer0_outputs(1333)) and (layer0_outputs(6107)));
    outputs(2764) <= layer0_outputs(7978);
    outputs(2765) <= (layer0_outputs(7171)) and (layer0_outputs(6555));
    outputs(2766) <= not(layer0_outputs(8998));
    outputs(2767) <= layer0_outputs(7510);
    outputs(2768) <= not((layer0_outputs(66)) xor (layer0_outputs(254)));
    outputs(2769) <= (layer0_outputs(8398)) and not (layer0_outputs(2602));
    outputs(2770) <= layer0_outputs(5832);
    outputs(2771) <= (layer0_outputs(4018)) and not (layer0_outputs(7105));
    outputs(2772) <= not((layer0_outputs(1150)) or (layer0_outputs(4513)));
    outputs(2773) <= layer0_outputs(5260);
    outputs(2774) <= (layer0_outputs(7761)) xor (layer0_outputs(7037));
    outputs(2775) <= layer0_outputs(2822);
    outputs(2776) <= not(layer0_outputs(5928)) or (layer0_outputs(6404));
    outputs(2777) <= not((layer0_outputs(5107)) xor (layer0_outputs(9875)));
    outputs(2778) <= not(layer0_outputs(5023)) or (layer0_outputs(4777));
    outputs(2779) <= (layer0_outputs(1190)) xor (layer0_outputs(5763));
    outputs(2780) <= not(layer0_outputs(3959)) or (layer0_outputs(9564));
    outputs(2781) <= not(layer0_outputs(9617)) or (layer0_outputs(343));
    outputs(2782) <= layer0_outputs(2545);
    outputs(2783) <= (layer0_outputs(4771)) and not (layer0_outputs(3444));
    outputs(2784) <= (layer0_outputs(5731)) or (layer0_outputs(8037));
    outputs(2785) <= layer0_outputs(2376);
    outputs(2786) <= (layer0_outputs(5812)) xor (layer0_outputs(1174));
    outputs(2787) <= not(layer0_outputs(1693));
    outputs(2788) <= not(layer0_outputs(6733));
    outputs(2789) <= layer0_outputs(8536);
    outputs(2790) <= layer0_outputs(6271);
    outputs(2791) <= not((layer0_outputs(7494)) or (layer0_outputs(3453)));
    outputs(2792) <= layer0_outputs(10054);
    outputs(2793) <= (layer0_outputs(4308)) or (layer0_outputs(479));
    outputs(2794) <= (layer0_outputs(9557)) or (layer0_outputs(10020));
    outputs(2795) <= not(layer0_outputs(4503));
    outputs(2796) <= not((layer0_outputs(821)) xor (layer0_outputs(7958)));
    outputs(2797) <= layer0_outputs(2956);
    outputs(2798) <= layer0_outputs(8341);
    outputs(2799) <= (layer0_outputs(8887)) and not (layer0_outputs(6854));
    outputs(2800) <= (layer0_outputs(7131)) or (layer0_outputs(4936));
    outputs(2801) <= (layer0_outputs(4548)) and not (layer0_outputs(8813));
    outputs(2802) <= not((layer0_outputs(1471)) xor (layer0_outputs(6923)));
    outputs(2803) <= layer0_outputs(556);
    outputs(2804) <= layer0_outputs(1973);
    outputs(2805) <= layer0_outputs(6830);
    outputs(2806) <= layer0_outputs(9641);
    outputs(2807) <= not((layer0_outputs(1559)) or (layer0_outputs(3523)));
    outputs(2808) <= (layer0_outputs(5863)) xor (layer0_outputs(4141));
    outputs(2809) <= not((layer0_outputs(1227)) or (layer0_outputs(9516)));
    outputs(2810) <= not(layer0_outputs(2634));
    outputs(2811) <= not(layer0_outputs(9227));
    outputs(2812) <= layer0_outputs(1166);
    outputs(2813) <= not(layer0_outputs(2856)) or (layer0_outputs(2289));
    outputs(2814) <= (layer0_outputs(4122)) xor (layer0_outputs(5871));
    outputs(2815) <= layer0_outputs(3825);
    outputs(2816) <= (layer0_outputs(424)) and (layer0_outputs(7632));
    outputs(2817) <= not((layer0_outputs(7514)) or (layer0_outputs(8585)));
    outputs(2818) <= (layer0_outputs(7096)) xor (layer0_outputs(3272));
    outputs(2819) <= layer0_outputs(444);
    outputs(2820) <= not(layer0_outputs(7212)) or (layer0_outputs(8067));
    outputs(2821) <= not((layer0_outputs(5708)) and (layer0_outputs(10000)));
    outputs(2822) <= (layer0_outputs(7512)) and not (layer0_outputs(4757));
    outputs(2823) <= not(layer0_outputs(507)) or (layer0_outputs(3396));
    outputs(2824) <= layer0_outputs(4982);
    outputs(2825) <= not(layer0_outputs(5533)) or (layer0_outputs(4976));
    outputs(2826) <= layer0_outputs(3137);
    outputs(2827) <= (layer0_outputs(4422)) xor (layer0_outputs(8811));
    outputs(2828) <= (layer0_outputs(3294)) and not (layer0_outputs(1026));
    outputs(2829) <= not(layer0_outputs(9735));
    outputs(2830) <= (layer0_outputs(7262)) and not (layer0_outputs(1557));
    outputs(2831) <= layer0_outputs(7332);
    outputs(2832) <= layer0_outputs(8710);
    outputs(2833) <= not(layer0_outputs(3764)) or (layer0_outputs(3243));
    outputs(2834) <= layer0_outputs(7755);
    outputs(2835) <= not(layer0_outputs(3538));
    outputs(2836) <= not((layer0_outputs(8626)) and (layer0_outputs(3132)));
    outputs(2837) <= (layer0_outputs(5662)) and (layer0_outputs(10124));
    outputs(2838) <= not(layer0_outputs(196));
    outputs(2839) <= not(layer0_outputs(7909));
    outputs(2840) <= not(layer0_outputs(9274));
    outputs(2841) <= layer0_outputs(1691);
    outputs(2842) <= not(layer0_outputs(9681));
    outputs(2843) <= not((layer0_outputs(10177)) or (layer0_outputs(7654)));
    outputs(2844) <= not((layer0_outputs(6154)) and (layer0_outputs(2372)));
    outputs(2845) <= layer0_outputs(7832);
    outputs(2846) <= layer0_outputs(8730);
    outputs(2847) <= (layer0_outputs(5522)) and not (layer0_outputs(5485));
    outputs(2848) <= not((layer0_outputs(4911)) or (layer0_outputs(7419)));
    outputs(2849) <= layer0_outputs(6537);
    outputs(2850) <= not((layer0_outputs(9486)) xor (layer0_outputs(377)));
    outputs(2851) <= (layer0_outputs(3816)) or (layer0_outputs(2633));
    outputs(2852) <= layer0_outputs(9823);
    outputs(2853) <= (layer0_outputs(5845)) and (layer0_outputs(2680));
    outputs(2854) <= (layer0_outputs(8823)) and (layer0_outputs(6143));
    outputs(2855) <= not((layer0_outputs(5819)) and (layer0_outputs(3172)));
    outputs(2856) <= layer0_outputs(58);
    outputs(2857) <= not(layer0_outputs(470));
    outputs(2858) <= (layer0_outputs(2789)) and (layer0_outputs(3911));
    outputs(2859) <= not(layer0_outputs(9131));
    outputs(2860) <= not(layer0_outputs(123)) or (layer0_outputs(1730));
    outputs(2861) <= not((layer0_outputs(4351)) xor (layer0_outputs(1668)));
    outputs(2862) <= (layer0_outputs(10174)) xor (layer0_outputs(7220));
    outputs(2863) <= not(layer0_outputs(10024));
    outputs(2864) <= not(layer0_outputs(1887)) or (layer0_outputs(324));
    outputs(2865) <= not((layer0_outputs(3445)) and (layer0_outputs(6129)));
    outputs(2866) <= (layer0_outputs(5753)) or (layer0_outputs(3708));
    outputs(2867) <= (layer0_outputs(6651)) or (layer0_outputs(487));
    outputs(2868) <= not(layer0_outputs(2560));
    outputs(2869) <= (layer0_outputs(1183)) xor (layer0_outputs(2969));
    outputs(2870) <= not(layer0_outputs(9453)) or (layer0_outputs(1076));
    outputs(2871) <= layer0_outputs(3343);
    outputs(2872) <= not((layer0_outputs(5219)) and (layer0_outputs(7551)));
    outputs(2873) <= layer0_outputs(7918);
    outputs(2874) <= not(layer0_outputs(5966)) or (layer0_outputs(7307));
    outputs(2875) <= (layer0_outputs(7688)) xor (layer0_outputs(5348));
    outputs(2876) <= not((layer0_outputs(5587)) xor (layer0_outputs(70)));
    outputs(2877) <= not((layer0_outputs(854)) and (layer0_outputs(3530)));
    outputs(2878) <= (layer0_outputs(2233)) xor (layer0_outputs(2158));
    outputs(2879) <= not(layer0_outputs(5227)) or (layer0_outputs(8477));
    outputs(2880) <= not(layer0_outputs(4632));
    outputs(2881) <= layer0_outputs(7993);
    outputs(2882) <= not(layer0_outputs(10134)) or (layer0_outputs(1538));
    outputs(2883) <= not(layer0_outputs(6738));
    outputs(2884) <= layer0_outputs(7252);
    outputs(2885) <= not(layer0_outputs(359)) or (layer0_outputs(3088));
    outputs(2886) <= not(layer0_outputs(7372)) or (layer0_outputs(3202));
    outputs(2887) <= not(layer0_outputs(54)) or (layer0_outputs(6794));
    outputs(2888) <= layer0_outputs(3986);
    outputs(2889) <= not(layer0_outputs(1978));
    outputs(2890) <= layer0_outputs(2978);
    outputs(2891) <= not(layer0_outputs(9299));
    outputs(2892) <= (layer0_outputs(538)) and (layer0_outputs(6584));
    outputs(2893) <= not((layer0_outputs(4828)) xor (layer0_outputs(10233)));
    outputs(2894) <= layer0_outputs(903);
    outputs(2895) <= not(layer0_outputs(4812)) or (layer0_outputs(5748));
    outputs(2896) <= not(layer0_outputs(5803)) or (layer0_outputs(7880));
    outputs(2897) <= not((layer0_outputs(6972)) xor (layer0_outputs(7211)));
    outputs(2898) <= not(layer0_outputs(9573));
    outputs(2899) <= not((layer0_outputs(5445)) or (layer0_outputs(3314)));
    outputs(2900) <= not(layer0_outputs(8273)) or (layer0_outputs(1783));
    outputs(2901) <= not(layer0_outputs(4687));
    outputs(2902) <= not(layer0_outputs(3785));
    outputs(2903) <= not((layer0_outputs(6941)) or (layer0_outputs(7211)));
    outputs(2904) <= layer0_outputs(3968);
    outputs(2905) <= not((layer0_outputs(5781)) or (layer0_outputs(5603)));
    outputs(2906) <= layer0_outputs(4506);
    outputs(2907) <= layer0_outputs(6859);
    outputs(2908) <= not(layer0_outputs(477));
    outputs(2909) <= not(layer0_outputs(6548));
    outputs(2910) <= not(layer0_outputs(10139));
    outputs(2911) <= not(layer0_outputs(302)) or (layer0_outputs(8202));
    outputs(2912) <= not(layer0_outputs(6918));
    outputs(2913) <= (layer0_outputs(8230)) or (layer0_outputs(1677));
    outputs(2914) <= not(layer0_outputs(8564)) or (layer0_outputs(279));
    outputs(2915) <= not(layer0_outputs(8873));
    outputs(2916) <= layer0_outputs(2181);
    outputs(2917) <= (layer0_outputs(9255)) xor (layer0_outputs(9250));
    outputs(2918) <= not(layer0_outputs(3107));
    outputs(2919) <= (layer0_outputs(3687)) xor (layer0_outputs(10007));
    outputs(2920) <= not(layer0_outputs(2994));
    outputs(2921) <= not(layer0_outputs(7167));
    outputs(2922) <= not((layer0_outputs(9181)) and (layer0_outputs(6635)));
    outputs(2923) <= (layer0_outputs(7166)) or (layer0_outputs(10180));
    outputs(2924) <= not(layer0_outputs(6084));
    outputs(2925) <= not((layer0_outputs(8457)) xor (layer0_outputs(4177)));
    outputs(2926) <= layer0_outputs(8050);
    outputs(2927) <= not((layer0_outputs(6383)) and (layer0_outputs(8249)));
    outputs(2928) <= (layer0_outputs(257)) and not (layer0_outputs(9303));
    outputs(2929) <= (layer0_outputs(2034)) xor (layer0_outputs(4897));
    outputs(2930) <= (layer0_outputs(4716)) and not (layer0_outputs(7611));
    outputs(2931) <= layer0_outputs(8256);
    outputs(2932) <= not(layer0_outputs(8893));
    outputs(2933) <= (layer0_outputs(1359)) or (layer0_outputs(1576));
    outputs(2934) <= not((layer0_outputs(6650)) xor (layer0_outputs(7413)));
    outputs(2935) <= '1';
    outputs(2936) <= layer0_outputs(3416);
    outputs(2937) <= not(layer0_outputs(1761)) or (layer0_outputs(663));
    outputs(2938) <= not(layer0_outputs(8590));
    outputs(2939) <= not(layer0_outputs(653)) or (layer0_outputs(7547));
    outputs(2940) <= (layer0_outputs(9943)) xor (layer0_outputs(4206));
    outputs(2941) <= layer0_outputs(3319);
    outputs(2942) <= (layer0_outputs(2029)) xor (layer0_outputs(1588));
    outputs(2943) <= not(layer0_outputs(373));
    outputs(2944) <= not((layer0_outputs(1620)) and (layer0_outputs(1479)));
    outputs(2945) <= (layer0_outputs(9961)) or (layer0_outputs(4085));
    outputs(2946) <= layer0_outputs(9169);
    outputs(2947) <= layer0_outputs(7934);
    outputs(2948) <= not((layer0_outputs(7293)) or (layer0_outputs(9237)));
    outputs(2949) <= not((layer0_outputs(9830)) or (layer0_outputs(6092)));
    outputs(2950) <= layer0_outputs(5465);
    outputs(2951) <= not(layer0_outputs(10052)) or (layer0_outputs(1500));
    outputs(2952) <= layer0_outputs(2403);
    outputs(2953) <= not(layer0_outputs(7579));
    outputs(2954) <= layer0_outputs(996);
    outputs(2955) <= (layer0_outputs(3562)) xor (layer0_outputs(2846));
    outputs(2956) <= layer0_outputs(5753);
    outputs(2957) <= not((layer0_outputs(536)) xor (layer0_outputs(1835)));
    outputs(2958) <= layer0_outputs(9012);
    outputs(2959) <= (layer0_outputs(1008)) and not (layer0_outputs(9771));
    outputs(2960) <= not((layer0_outputs(4226)) or (layer0_outputs(3126)));
    outputs(2961) <= (layer0_outputs(9406)) and (layer0_outputs(5714));
    outputs(2962) <= not((layer0_outputs(5358)) xor (layer0_outputs(4137)));
    outputs(2963) <= not(layer0_outputs(5331)) or (layer0_outputs(9673));
    outputs(2964) <= not(layer0_outputs(4679)) or (layer0_outputs(1529));
    outputs(2965) <= not(layer0_outputs(6229)) or (layer0_outputs(4810));
    outputs(2966) <= layer0_outputs(5953);
    outputs(2967) <= layer0_outputs(9606);
    outputs(2968) <= (layer0_outputs(4420)) or (layer0_outputs(1099));
    outputs(2969) <= (layer0_outputs(8970)) xor (layer0_outputs(1520));
    outputs(2970) <= not((layer0_outputs(1295)) or (layer0_outputs(3783)));
    outputs(2971) <= not((layer0_outputs(7996)) and (layer0_outputs(3067)));
    outputs(2972) <= layer0_outputs(7284);
    outputs(2973) <= not(layer0_outputs(2006));
    outputs(2974) <= (layer0_outputs(5061)) or (layer0_outputs(8449));
    outputs(2975) <= not((layer0_outputs(6314)) xor (layer0_outputs(6397)));
    outputs(2976) <= (layer0_outputs(6735)) and not (layer0_outputs(2048));
    outputs(2977) <= not((layer0_outputs(4903)) and (layer0_outputs(7235)));
    outputs(2978) <= not(layer0_outputs(2220));
    outputs(2979) <= not(layer0_outputs(8149));
    outputs(2980) <= layer0_outputs(803);
    outputs(2981) <= not((layer0_outputs(2026)) and (layer0_outputs(1718)));
    outputs(2982) <= not((layer0_outputs(8586)) xor (layer0_outputs(892)));
    outputs(2983) <= (layer0_outputs(2849)) and not (layer0_outputs(382));
    outputs(2984) <= (layer0_outputs(1077)) and (layer0_outputs(8260));
    outputs(2985) <= (layer0_outputs(9705)) xor (layer0_outputs(4669));
    outputs(2986) <= (layer0_outputs(224)) xor (layer0_outputs(544));
    outputs(2987) <= layer0_outputs(5251);
    outputs(2988) <= not(layer0_outputs(630));
    outputs(2989) <= not((layer0_outputs(4070)) and (layer0_outputs(2198)));
    outputs(2990) <= (layer0_outputs(10095)) and (layer0_outputs(1141));
    outputs(2991) <= not((layer0_outputs(1218)) or (layer0_outputs(6847)));
    outputs(2992) <= not(layer0_outputs(1340));
    outputs(2993) <= layer0_outputs(2141);
    outputs(2994) <= not(layer0_outputs(5683));
    outputs(2995) <= not(layer0_outputs(1278)) or (layer0_outputs(6832));
    outputs(2996) <= (layer0_outputs(7916)) and not (layer0_outputs(9923));
    outputs(2997) <= not((layer0_outputs(8377)) and (layer0_outputs(3167)));
    outputs(2998) <= not((layer0_outputs(9708)) or (layer0_outputs(8527)));
    outputs(2999) <= (layer0_outputs(8578)) or (layer0_outputs(6030));
    outputs(3000) <= not(layer0_outputs(6569));
    outputs(3001) <= (layer0_outputs(4239)) and (layer0_outputs(7912));
    outputs(3002) <= layer0_outputs(6171);
    outputs(3003) <= not(layer0_outputs(6381));
    outputs(3004) <= (layer0_outputs(7518)) and (layer0_outputs(2094));
    outputs(3005) <= (layer0_outputs(592)) and not (layer0_outputs(9954));
    outputs(3006) <= not(layer0_outputs(7236));
    outputs(3007) <= not((layer0_outputs(7765)) and (layer0_outputs(9994)));
    outputs(3008) <= not(layer0_outputs(1988));
    outputs(3009) <= layer0_outputs(1713);
    outputs(3010) <= layer0_outputs(4237);
    outputs(3011) <= (layer0_outputs(5261)) and not (layer0_outputs(6403));
    outputs(3012) <= not(layer0_outputs(9444));
    outputs(3013) <= not((layer0_outputs(4147)) and (layer0_outputs(7657)));
    outputs(3014) <= not(layer0_outputs(6934));
    outputs(3015) <= (layer0_outputs(5593)) xor (layer0_outputs(1688));
    outputs(3016) <= (layer0_outputs(2508)) and not (layer0_outputs(820));
    outputs(3017) <= layer0_outputs(9865);
    outputs(3018) <= not((layer0_outputs(9345)) xor (layer0_outputs(795)));
    outputs(3019) <= not((layer0_outputs(3729)) and (layer0_outputs(2379)));
    outputs(3020) <= not((layer0_outputs(7299)) xor (layer0_outputs(6725)));
    outputs(3021) <= not(layer0_outputs(8809));
    outputs(3022) <= (layer0_outputs(8453)) or (layer0_outputs(9205));
    outputs(3023) <= (layer0_outputs(9671)) and (layer0_outputs(7732));
    outputs(3024) <= (layer0_outputs(252)) or (layer0_outputs(5822));
    outputs(3025) <= not(layer0_outputs(2095)) or (layer0_outputs(7590));
    outputs(3026) <= layer0_outputs(9130);
    outputs(3027) <= layer0_outputs(5159);
    outputs(3028) <= not(layer0_outputs(2962));
    outputs(3029) <= not(layer0_outputs(2112)) or (layer0_outputs(2447));
    outputs(3030) <= (layer0_outputs(92)) or (layer0_outputs(4860));
    outputs(3031) <= (layer0_outputs(8167)) and not (layer0_outputs(9680));
    outputs(3032) <= not(layer0_outputs(8403));
    outputs(3033) <= (layer0_outputs(775)) or (layer0_outputs(4479));
    outputs(3034) <= not(layer0_outputs(618));
    outputs(3035) <= not((layer0_outputs(1223)) and (layer0_outputs(2360)));
    outputs(3036) <= not(layer0_outputs(2803)) or (layer0_outputs(6745));
    outputs(3037) <= not(layer0_outputs(7883));
    outputs(3038) <= not(layer0_outputs(1419));
    outputs(3039) <= (layer0_outputs(3170)) and not (layer0_outputs(9816));
    outputs(3040) <= not((layer0_outputs(10096)) or (layer0_outputs(2629)));
    outputs(3041) <= not(layer0_outputs(8309));
    outputs(3042) <= not(layer0_outputs(6336)) or (layer0_outputs(3596));
    outputs(3043) <= not((layer0_outputs(2044)) xor (layer0_outputs(6850)));
    outputs(3044) <= not(layer0_outputs(8328)) or (layer0_outputs(7656));
    outputs(3045) <= not(layer0_outputs(8407)) or (layer0_outputs(7800));
    outputs(3046) <= not(layer0_outputs(1780));
    outputs(3047) <= not((layer0_outputs(7409)) or (layer0_outputs(7990)));
    outputs(3048) <= (layer0_outputs(1042)) and not (layer0_outputs(2645));
    outputs(3049) <= not(layer0_outputs(9800));
    outputs(3050) <= not(layer0_outputs(5983));
    outputs(3051) <= layer0_outputs(2771);
    outputs(3052) <= layer0_outputs(533);
    outputs(3053) <= layer0_outputs(7873);
    outputs(3054) <= not((layer0_outputs(3068)) xor (layer0_outputs(7739)));
    outputs(3055) <= not(layer0_outputs(1131)) or (layer0_outputs(8759));
    outputs(3056) <= layer0_outputs(8940);
    outputs(3057) <= not(layer0_outputs(8831)) or (layer0_outputs(1644));
    outputs(3058) <= (layer0_outputs(9078)) or (layer0_outputs(1940));
    outputs(3059) <= (layer0_outputs(5201)) and not (layer0_outputs(7409));
    outputs(3060) <= (layer0_outputs(3844)) or (layer0_outputs(4240));
    outputs(3061) <= not((layer0_outputs(7327)) xor (layer0_outputs(7855)));
    outputs(3062) <= not(layer0_outputs(6280)) or (layer0_outputs(7222));
    outputs(3063) <= not(layer0_outputs(2711));
    outputs(3064) <= not((layer0_outputs(6024)) xor (layer0_outputs(6321)));
    outputs(3065) <= layer0_outputs(2185);
    outputs(3066) <= (layer0_outputs(4199)) xor (layer0_outputs(3438));
    outputs(3067) <= not((layer0_outputs(2334)) and (layer0_outputs(2670)));
    outputs(3068) <= not(layer0_outputs(735));
    outputs(3069) <= layer0_outputs(5343);
    outputs(3070) <= (layer0_outputs(116)) and not (layer0_outputs(3684));
    outputs(3071) <= (layer0_outputs(756)) xor (layer0_outputs(2532));
    outputs(3072) <= not(layer0_outputs(3434));
    outputs(3073) <= not(layer0_outputs(8204));
    outputs(3074) <= layer0_outputs(9359);
    outputs(3075) <= (layer0_outputs(8842)) and not (layer0_outputs(325));
    outputs(3076) <= (layer0_outputs(3213)) xor (layer0_outputs(7423));
    outputs(3077) <= not((layer0_outputs(9067)) xor (layer0_outputs(4220)));
    outputs(3078) <= not(layer0_outputs(8734));
    outputs(3079) <= layer0_outputs(6297);
    outputs(3080) <= not(layer0_outputs(1045));
    outputs(3081) <= (layer0_outputs(4266)) and not (layer0_outputs(7086));
    outputs(3082) <= (layer0_outputs(6339)) xor (layer0_outputs(471));
    outputs(3083) <= layer0_outputs(3745);
    outputs(3084) <= (layer0_outputs(875)) and not (layer0_outputs(8405));
    outputs(3085) <= not(layer0_outputs(823));
    outputs(3086) <= (layer0_outputs(2200)) and (layer0_outputs(10154));
    outputs(3087) <= not((layer0_outputs(4804)) or (layer0_outputs(3748)));
    outputs(3088) <= (layer0_outputs(4477)) and not (layer0_outputs(6599));
    outputs(3089) <= not((layer0_outputs(1842)) xor (layer0_outputs(9630)));
    outputs(3090) <= not((layer0_outputs(2343)) or (layer0_outputs(1824)));
    outputs(3091) <= not((layer0_outputs(2722)) xor (layer0_outputs(9673)));
    outputs(3092) <= not(layer0_outputs(4303));
    outputs(3093) <= layer0_outputs(3624);
    outputs(3094) <= not(layer0_outputs(2157));
    outputs(3095) <= not(layer0_outputs(1182));
    outputs(3096) <= layer0_outputs(8007);
    outputs(3097) <= not(layer0_outputs(9250));
    outputs(3098) <= (layer0_outputs(3758)) and (layer0_outputs(2409));
    outputs(3099) <= not(layer0_outputs(3984));
    outputs(3100) <= not((layer0_outputs(3746)) or (layer0_outputs(6641)));
    outputs(3101) <= not((layer0_outputs(981)) or (layer0_outputs(4230)));
    outputs(3102) <= (layer0_outputs(6530)) and not (layer0_outputs(1113));
    outputs(3103) <= layer0_outputs(8419);
    outputs(3104) <= (layer0_outputs(3341)) xor (layer0_outputs(3814));
    outputs(3105) <= not((layer0_outputs(689)) or (layer0_outputs(2868)));
    outputs(3106) <= not((layer0_outputs(4160)) and (layer0_outputs(6650)));
    outputs(3107) <= (layer0_outputs(5009)) and (layer0_outputs(3448));
    outputs(3108) <= layer0_outputs(474);
    outputs(3109) <= not((layer0_outputs(3074)) and (layer0_outputs(4705)));
    outputs(3110) <= not(layer0_outputs(537));
    outputs(3111) <= layer0_outputs(6278);
    outputs(3112) <= layer0_outputs(8667);
    outputs(3113) <= layer0_outputs(5698);
    outputs(3114) <= not((layer0_outputs(6172)) and (layer0_outputs(6102)));
    outputs(3115) <= not((layer0_outputs(7007)) xor (layer0_outputs(2644)));
    outputs(3116) <= (layer0_outputs(8070)) and not (layer0_outputs(2583));
    outputs(3117) <= not(layer0_outputs(2060));
    outputs(3118) <= (layer0_outputs(10220)) and not (layer0_outputs(8672));
    outputs(3119) <= (layer0_outputs(7766)) xor (layer0_outputs(6590));
    outputs(3120) <= (layer0_outputs(771)) and not (layer0_outputs(7046));
    outputs(3121) <= not(layer0_outputs(7653));
    outputs(3122) <= not((layer0_outputs(188)) xor (layer0_outputs(9984)));
    outputs(3123) <= not(layer0_outputs(4036));
    outputs(3124) <= not((layer0_outputs(4436)) or (layer0_outputs(6633)));
    outputs(3125) <= not(layer0_outputs(4802)) or (layer0_outputs(4053));
    outputs(3126) <= layer0_outputs(3536);
    outputs(3127) <= (layer0_outputs(626)) and (layer0_outputs(6616));
    outputs(3128) <= not((layer0_outputs(7698)) and (layer0_outputs(1425)));
    outputs(3129) <= layer0_outputs(656);
    outputs(3130) <= not((layer0_outputs(9689)) xor (layer0_outputs(2610)));
    outputs(3131) <= (layer0_outputs(4600)) and not (layer0_outputs(5387));
    outputs(3132) <= (layer0_outputs(8213)) and not (layer0_outputs(5520));
    outputs(3133) <= (layer0_outputs(8169)) and not (layer0_outputs(7141));
    outputs(3134) <= not((layer0_outputs(6900)) xor (layer0_outputs(2460)));
    outputs(3135) <= not(layer0_outputs(4893));
    outputs(3136) <= (layer0_outputs(9156)) and not (layer0_outputs(4943));
    outputs(3137) <= not((layer0_outputs(6191)) or (layer0_outputs(764)));
    outputs(3138) <= layer0_outputs(10011);
    outputs(3139) <= not(layer0_outputs(3906));
    outputs(3140) <= not((layer0_outputs(86)) or (layer0_outputs(8940)));
    outputs(3141) <= layer0_outputs(9024);
    outputs(3142) <= not((layer0_outputs(248)) xor (layer0_outputs(1757)));
    outputs(3143) <= not((layer0_outputs(8930)) or (layer0_outputs(149)));
    outputs(3144) <= (layer0_outputs(2913)) and not (layer0_outputs(7000));
    outputs(3145) <= (layer0_outputs(5258)) and not (layer0_outputs(5911));
    outputs(3146) <= (layer0_outputs(6456)) and not (layer0_outputs(825));
    outputs(3147) <= layer0_outputs(3013);
    outputs(3148) <= layer0_outputs(7914);
    outputs(3149) <= (layer0_outputs(6487)) xor (layer0_outputs(9491));
    outputs(3150) <= not((layer0_outputs(367)) and (layer0_outputs(28)));
    outputs(3151) <= layer0_outputs(9894);
    outputs(3152) <= not(layer0_outputs(1725));
    outputs(3153) <= layer0_outputs(6389);
    outputs(3154) <= (layer0_outputs(403)) and not (layer0_outputs(9402));
    outputs(3155) <= not(layer0_outputs(4580)) or (layer0_outputs(266));
    outputs(3156) <= not((layer0_outputs(10141)) xor (layer0_outputs(7756)));
    outputs(3157) <= not((layer0_outputs(9504)) and (layer0_outputs(9208)));
    outputs(3158) <= (layer0_outputs(5331)) xor (layer0_outputs(9434));
    outputs(3159) <= not(layer0_outputs(9346));
    outputs(3160) <= (layer0_outputs(5761)) or (layer0_outputs(1602));
    outputs(3161) <= not(layer0_outputs(8636));
    outputs(3162) <= not((layer0_outputs(1567)) xor (layer0_outputs(7469)));
    outputs(3163) <= not(layer0_outputs(8500));
    outputs(3164) <= (layer0_outputs(174)) xor (layer0_outputs(8797));
    outputs(3165) <= layer0_outputs(5267);
    outputs(3166) <= (layer0_outputs(9571)) xor (layer0_outputs(10183));
    outputs(3167) <= not(layer0_outputs(3599));
    outputs(3168) <= not(layer0_outputs(8016)) or (layer0_outputs(1516));
    outputs(3169) <= (layer0_outputs(3791)) xor (layer0_outputs(5833));
    outputs(3170) <= not((layer0_outputs(450)) and (layer0_outputs(4226)));
    outputs(3171) <= (layer0_outputs(786)) and not (layer0_outputs(2357));
    outputs(3172) <= not((layer0_outputs(1702)) or (layer0_outputs(8680)));
    outputs(3173) <= layer0_outputs(3734);
    outputs(3174) <= (layer0_outputs(5682)) xor (layer0_outputs(3597));
    outputs(3175) <= not(layer0_outputs(2636));
    outputs(3176) <= (layer0_outputs(10014)) and (layer0_outputs(9380));
    outputs(3177) <= layer0_outputs(759);
    outputs(3178) <= (layer0_outputs(7911)) xor (layer0_outputs(4258));
    outputs(3179) <= (layer0_outputs(2489)) and not (layer0_outputs(2172));
    outputs(3180) <= not(layer0_outputs(8265));
    outputs(3181) <= not(layer0_outputs(7306));
    outputs(3182) <= not((layer0_outputs(8426)) xor (layer0_outputs(4772)));
    outputs(3183) <= layer0_outputs(1907);
    outputs(3184) <= (layer0_outputs(7483)) and not (layer0_outputs(3019));
    outputs(3185) <= (layer0_outputs(7454)) and not (layer0_outputs(862));
    outputs(3186) <= not((layer0_outputs(1257)) xor (layer0_outputs(2254)));
    outputs(3187) <= not(layer0_outputs(8369)) or (layer0_outputs(6162));
    outputs(3188) <= (layer0_outputs(4987)) and (layer0_outputs(9777));
    outputs(3189) <= not((layer0_outputs(1990)) or (layer0_outputs(9770)));
    outputs(3190) <= layer0_outputs(3629);
    outputs(3191) <= not(layer0_outputs(8795));
    outputs(3192) <= (layer0_outputs(6283)) xor (layer0_outputs(4795));
    outputs(3193) <= (layer0_outputs(1679)) and (layer0_outputs(3136));
    outputs(3194) <= not(layer0_outputs(4974));
    outputs(3195) <= (layer0_outputs(10067)) xor (layer0_outputs(6235));
    outputs(3196) <= not(layer0_outputs(2363));
    outputs(3197) <= (layer0_outputs(8989)) and not (layer0_outputs(3518));
    outputs(3198) <= (layer0_outputs(3359)) xor (layer0_outputs(9984));
    outputs(3199) <= (layer0_outputs(6714)) xor (layer0_outputs(10146));
    outputs(3200) <= not((layer0_outputs(8467)) or (layer0_outputs(6564)));
    outputs(3201) <= not(layer0_outputs(5108));
    outputs(3202) <= (layer0_outputs(6525)) or (layer0_outputs(937));
    outputs(3203) <= layer0_outputs(2675);
    outputs(3204) <= not(layer0_outputs(2619)) or (layer0_outputs(7145));
    outputs(3205) <= (layer0_outputs(7725)) xor (layer0_outputs(1686));
    outputs(3206) <= not(layer0_outputs(4328));
    outputs(3207) <= layer0_outputs(8706);
    outputs(3208) <= not(layer0_outputs(9243));
    outputs(3209) <= (layer0_outputs(348)) xor (layer0_outputs(3700));
    outputs(3210) <= (layer0_outputs(10002)) xor (layer0_outputs(10165));
    outputs(3211) <= layer0_outputs(1956);
    outputs(3212) <= layer0_outputs(6173);
    outputs(3213) <= (layer0_outputs(876)) and not (layer0_outputs(4391));
    outputs(3214) <= layer0_outputs(9777);
    outputs(3215) <= (layer0_outputs(737)) and (layer0_outputs(2296));
    outputs(3216) <= layer0_outputs(9995);
    outputs(3217) <= not((layer0_outputs(514)) and (layer0_outputs(8817)));
    outputs(3218) <= layer0_outputs(2758);
    outputs(3219) <= not(layer0_outputs(6057)) or (layer0_outputs(6727));
    outputs(3220) <= layer0_outputs(2674);
    outputs(3221) <= not(layer0_outputs(2336));
    outputs(3222) <= not(layer0_outputs(2304));
    outputs(3223) <= (layer0_outputs(5247)) and not (layer0_outputs(1465));
    outputs(3224) <= not(layer0_outputs(2128)) or (layer0_outputs(8611));
    outputs(3225) <= not((layer0_outputs(7609)) xor (layer0_outputs(916)));
    outputs(3226) <= not(layer0_outputs(10194));
    outputs(3227) <= not((layer0_outputs(3539)) xor (layer0_outputs(5224)));
    outputs(3228) <= not(layer0_outputs(9943));
    outputs(3229) <= (layer0_outputs(7449)) xor (layer0_outputs(6365));
    outputs(3230) <= (layer0_outputs(6395)) xor (layer0_outputs(9918));
    outputs(3231) <= (layer0_outputs(5698)) and not (layer0_outputs(6709));
    outputs(3232) <= (layer0_outputs(9300)) xor (layer0_outputs(9140));
    outputs(3233) <= not(layer0_outputs(8093));
    outputs(3234) <= layer0_outputs(1528);
    outputs(3235) <= not(layer0_outputs(2029));
    outputs(3236) <= not((layer0_outputs(5615)) or (layer0_outputs(1702)));
    outputs(3237) <= (layer0_outputs(6820)) xor (layer0_outputs(2921));
    outputs(3238) <= not(layer0_outputs(7667)) or (layer0_outputs(5588));
    outputs(3239) <= layer0_outputs(1969);
    outputs(3240) <= not(layer0_outputs(2862));
    outputs(3241) <= layer0_outputs(105);
    outputs(3242) <= (layer0_outputs(8784)) and not (layer0_outputs(4728));
    outputs(3243) <= (layer0_outputs(7317)) and (layer0_outputs(3257));
    outputs(3244) <= layer0_outputs(6922);
    outputs(3245) <= not((layer0_outputs(9832)) and (layer0_outputs(2025)));
    outputs(3246) <= not(layer0_outputs(5827)) or (layer0_outputs(5812));
    outputs(3247) <= (layer0_outputs(1616)) and not (layer0_outputs(4440));
    outputs(3248) <= not(layer0_outputs(168));
    outputs(3249) <= not((layer0_outputs(5573)) or (layer0_outputs(8402)));
    outputs(3250) <= not((layer0_outputs(6033)) xor (layer0_outputs(9192)));
    outputs(3251) <= layer0_outputs(5918);
    outputs(3252) <= layer0_outputs(8473);
    outputs(3253) <= layer0_outputs(9354);
    outputs(3254) <= (layer0_outputs(2115)) and (layer0_outputs(5169));
    outputs(3255) <= layer0_outputs(4538);
    outputs(3256) <= not((layer0_outputs(1629)) xor (layer0_outputs(5186)));
    outputs(3257) <= (layer0_outputs(341)) xor (layer0_outputs(4578));
    outputs(3258) <= layer0_outputs(9);
    outputs(3259) <= (layer0_outputs(10126)) and (layer0_outputs(2646));
    outputs(3260) <= not(layer0_outputs(5366)) or (layer0_outputs(662));
    outputs(3261) <= not((layer0_outputs(8321)) xor (layer0_outputs(3987)));
    outputs(3262) <= (layer0_outputs(5194)) or (layer0_outputs(7235));
    outputs(3263) <= not(layer0_outputs(1332));
    outputs(3264) <= not(layer0_outputs(4183));
    outputs(3265) <= (layer0_outputs(8949)) or (layer0_outputs(4246));
    outputs(3266) <= layer0_outputs(4172);
    outputs(3267) <= not((layer0_outputs(4444)) or (layer0_outputs(7273)));
    outputs(3268) <= layer0_outputs(3564);
    outputs(3269) <= layer0_outputs(4066);
    outputs(3270) <= (layer0_outputs(1532)) and (layer0_outputs(5102));
    outputs(3271) <= not((layer0_outputs(3558)) xor (layer0_outputs(3316)));
    outputs(3272) <= not(layer0_outputs(3147)) or (layer0_outputs(5910));
    outputs(3273) <= (layer0_outputs(1987)) xor (layer0_outputs(3899));
    outputs(3274) <= layer0_outputs(3922);
    outputs(3275) <= (layer0_outputs(5207)) xor (layer0_outputs(9670));
    outputs(3276) <= layer0_outputs(8073);
    outputs(3277) <= (layer0_outputs(4031)) and not (layer0_outputs(7855));
    outputs(3278) <= (layer0_outputs(8013)) or (layer0_outputs(6321));
    outputs(3279) <= not(layer0_outputs(216));
    outputs(3280) <= layer0_outputs(402);
    outputs(3281) <= not(layer0_outputs(8692)) or (layer0_outputs(10130));
    outputs(3282) <= not(layer0_outputs(9469));
    outputs(3283) <= not(layer0_outputs(3567));
    outputs(3284) <= not(layer0_outputs(4442)) or (layer0_outputs(5383));
    outputs(3285) <= (layer0_outputs(10155)) and not (layer0_outputs(468));
    outputs(3286) <= not(layer0_outputs(41)) or (layer0_outputs(3288));
    outputs(3287) <= not(layer0_outputs(9851));
    outputs(3288) <= layer0_outputs(6524);
    outputs(3289) <= not(layer0_outputs(7178));
    outputs(3290) <= (layer0_outputs(5133)) and (layer0_outputs(10078));
    outputs(3291) <= (layer0_outputs(4608)) xor (layer0_outputs(22));
    outputs(3292) <= (layer0_outputs(4507)) and not (layer0_outputs(8215));
    outputs(3293) <= not((layer0_outputs(4433)) xor (layer0_outputs(4007)));
    outputs(3294) <= (layer0_outputs(7266)) and not (layer0_outputs(90));
    outputs(3295) <= (layer0_outputs(5287)) xor (layer0_outputs(3437));
    outputs(3296) <= not((layer0_outputs(2222)) xor (layer0_outputs(8526)));
    outputs(3297) <= not((layer0_outputs(387)) xor (layer0_outputs(2313)));
    outputs(3298) <= not(layer0_outputs(9955));
    outputs(3299) <= (layer0_outputs(1939)) xor (layer0_outputs(4744));
    outputs(3300) <= (layer0_outputs(2809)) and (layer0_outputs(968));
    outputs(3301) <= layer0_outputs(6679);
    outputs(3302) <= (layer0_outputs(1542)) and not (layer0_outputs(4739));
    outputs(3303) <= (layer0_outputs(3070)) and not (layer0_outputs(9710));
    outputs(3304) <= layer0_outputs(2242);
    outputs(3305) <= not(layer0_outputs(6973)) or (layer0_outputs(3664));
    outputs(3306) <= not((layer0_outputs(1554)) xor (layer0_outputs(4839)));
    outputs(3307) <= (layer0_outputs(2179)) and not (layer0_outputs(777));
    outputs(3308) <= not((layer0_outputs(2171)) xor (layer0_outputs(3285)));
    outputs(3309) <= not(layer0_outputs(3167)) or (layer0_outputs(1617));
    outputs(3310) <= (layer0_outputs(2737)) and not (layer0_outputs(9199));
    outputs(3311) <= (layer0_outputs(2497)) and not (layer0_outputs(9495));
    outputs(3312) <= layer0_outputs(399);
    outputs(3313) <= (layer0_outputs(9183)) or (layer0_outputs(3580));
    outputs(3314) <= layer0_outputs(1238);
    outputs(3315) <= not((layer0_outputs(8403)) xor (layer0_outputs(3115)));
    outputs(3316) <= not(layer0_outputs(6795));
    outputs(3317) <= not((layer0_outputs(2190)) and (layer0_outputs(5455)));
    outputs(3318) <= (layer0_outputs(10035)) or (layer0_outputs(1362));
    outputs(3319) <= not(layer0_outputs(8276));
    outputs(3320) <= not((layer0_outputs(2838)) or (layer0_outputs(8154)));
    outputs(3321) <= not(layer0_outputs(5444));
    outputs(3322) <= (layer0_outputs(3949)) and not (layer0_outputs(7990));
    outputs(3323) <= not((layer0_outputs(1032)) and (layer0_outputs(5170)));
    outputs(3324) <= (layer0_outputs(7738)) and (layer0_outputs(9172));
    outputs(3325) <= not((layer0_outputs(9921)) xor (layer0_outputs(8390)));
    outputs(3326) <= layer0_outputs(4348);
    outputs(3327) <= not(layer0_outputs(9554)) or (layer0_outputs(9387));
    outputs(3328) <= layer0_outputs(885);
    outputs(3329) <= not(layer0_outputs(7612));
    outputs(3330) <= not(layer0_outputs(8560));
    outputs(3331) <= (layer0_outputs(6320)) or (layer0_outputs(2892));
    outputs(3332) <= (layer0_outputs(3845)) xor (layer0_outputs(1056));
    outputs(3333) <= layer0_outputs(4091);
    outputs(3334) <= (layer0_outputs(676)) and not (layer0_outputs(5290));
    outputs(3335) <= not(layer0_outputs(3280));
    outputs(3336) <= not(layer0_outputs(8479));
    outputs(3337) <= not(layer0_outputs(5060));
    outputs(3338) <= (layer0_outputs(7724)) xor (layer0_outputs(4502));
    outputs(3339) <= layer0_outputs(4329);
    outputs(3340) <= (layer0_outputs(378)) or (layer0_outputs(7546));
    outputs(3341) <= (layer0_outputs(1487)) xor (layer0_outputs(3426));
    outputs(3342) <= (layer0_outputs(9905)) xor (layer0_outputs(2751));
    outputs(3343) <= (layer0_outputs(2877)) and not (layer0_outputs(5227));
    outputs(3344) <= not(layer0_outputs(1862));
    outputs(3345) <= not(layer0_outputs(9275));
    outputs(3346) <= layer0_outputs(2114);
    outputs(3347) <= layer0_outputs(176);
    outputs(3348) <= (layer0_outputs(4031)) xor (layer0_outputs(5418));
    outputs(3349) <= (layer0_outputs(4093)) xor (layer0_outputs(545));
    outputs(3350) <= not((layer0_outputs(710)) xor (layer0_outputs(4159)));
    outputs(3351) <= (layer0_outputs(10185)) or (layer0_outputs(9543));
    outputs(3352) <= not(layer0_outputs(4670));
    outputs(3353) <= not((layer0_outputs(7866)) or (layer0_outputs(9047)));
    outputs(3354) <= not(layer0_outputs(586));
    outputs(3355) <= layer0_outputs(3716);
    outputs(3356) <= (layer0_outputs(3706)) or (layer0_outputs(9189));
    outputs(3357) <= not(layer0_outputs(1441));
    outputs(3358) <= not(layer0_outputs(1922));
    outputs(3359) <= not(layer0_outputs(6009)) or (layer0_outputs(9522));
    outputs(3360) <= layer0_outputs(7921);
    outputs(3361) <= not(layer0_outputs(6625));
    outputs(3362) <= not(layer0_outputs(1473));
    outputs(3363) <= layer0_outputs(4104);
    outputs(3364) <= layer0_outputs(7245);
    outputs(3365) <= layer0_outputs(1805);
    outputs(3366) <= (layer0_outputs(5083)) and not (layer0_outputs(5188));
    outputs(3367) <= not(layer0_outputs(596));
    outputs(3368) <= (layer0_outputs(2831)) xor (layer0_outputs(9861));
    outputs(3369) <= (layer0_outputs(7519)) and (layer0_outputs(6425));
    outputs(3370) <= not(layer0_outputs(2048));
    outputs(3371) <= layer0_outputs(5025);
    outputs(3372) <= not(layer0_outputs(10039)) or (layer0_outputs(3397));
    outputs(3373) <= not(layer0_outputs(428)) or (layer0_outputs(7100));
    outputs(3374) <= layer0_outputs(8632);
    outputs(3375) <= (layer0_outputs(6375)) and (layer0_outputs(4293));
    outputs(3376) <= layer0_outputs(8217);
    outputs(3377) <= not(layer0_outputs(4628));
    outputs(3378) <= not((layer0_outputs(7881)) xor (layer0_outputs(4135)));
    outputs(3379) <= not(layer0_outputs(1980));
    outputs(3380) <= not(layer0_outputs(3998));
    outputs(3381) <= not((layer0_outputs(4717)) xor (layer0_outputs(9370)));
    outputs(3382) <= (layer0_outputs(1181)) or (layer0_outputs(5514));
    outputs(3383) <= (layer0_outputs(8060)) xor (layer0_outputs(6418));
    outputs(3384) <= not(layer0_outputs(3534));
    outputs(3385) <= (layer0_outputs(3382)) and (layer0_outputs(5257));
    outputs(3386) <= layer0_outputs(2632);
    outputs(3387) <= not(layer0_outputs(6435)) or (layer0_outputs(2378));
    outputs(3388) <= not((layer0_outputs(1366)) xor (layer0_outputs(765)));
    outputs(3389) <= (layer0_outputs(7781)) xor (layer0_outputs(9094));
    outputs(3390) <= layer0_outputs(8211);
    outputs(3391) <= not(layer0_outputs(4059));
    outputs(3392) <= (layer0_outputs(5008)) xor (layer0_outputs(1339));
    outputs(3393) <= layer0_outputs(2);
    outputs(3394) <= (layer0_outputs(7744)) or (layer0_outputs(964));
    outputs(3395) <= not(layer0_outputs(437));
    outputs(3396) <= (layer0_outputs(4291)) or (layer0_outputs(1243));
    outputs(3397) <= not(layer0_outputs(5052)) or (layer0_outputs(4032));
    outputs(3398) <= (layer0_outputs(1028)) xor (layer0_outputs(7685));
    outputs(3399) <= layer0_outputs(4811);
    outputs(3400) <= (layer0_outputs(1936)) xor (layer0_outputs(4126));
    outputs(3401) <= not(layer0_outputs(1072));
    outputs(3402) <= (layer0_outputs(5941)) and not (layer0_outputs(2608));
    outputs(3403) <= not((layer0_outputs(9283)) or (layer0_outputs(9740)));
    outputs(3404) <= layer0_outputs(5555);
    outputs(3405) <= (layer0_outputs(8462)) and (layer0_outputs(6020));
    outputs(3406) <= not(layer0_outputs(1558));
    outputs(3407) <= (layer0_outputs(7549)) xor (layer0_outputs(7851));
    outputs(3408) <= layer0_outputs(3083);
    outputs(3409) <= layer0_outputs(6005);
    outputs(3410) <= (layer0_outputs(6966)) xor (layer0_outputs(5458));
    outputs(3411) <= not((layer0_outputs(7962)) xor (layer0_outputs(7330)));
    outputs(3412) <= not((layer0_outputs(6208)) xor (layer0_outputs(9946)));
    outputs(3413) <= not((layer0_outputs(6263)) and (layer0_outputs(4767)));
    outputs(3414) <= layer0_outputs(809);
    outputs(3415) <= layer0_outputs(7515);
    outputs(3416) <= not(layer0_outputs(5400));
    outputs(3417) <= not((layer0_outputs(9369)) or (layer0_outputs(477)));
    outputs(3418) <= (layer0_outputs(4048)) xor (layer0_outputs(5618));
    outputs(3419) <= layer0_outputs(4532);
    outputs(3420) <= layer0_outputs(3488);
    outputs(3421) <= layer0_outputs(7690);
    outputs(3422) <= (layer0_outputs(6194)) xor (layer0_outputs(10085));
    outputs(3423) <= not((layer0_outputs(4535)) and (layer0_outputs(5634)));
    outputs(3424) <= not((layer0_outputs(5091)) and (layer0_outputs(730)));
    outputs(3425) <= (layer0_outputs(3773)) xor (layer0_outputs(4492));
    outputs(3426) <= (layer0_outputs(3757)) xor (layer0_outputs(6677));
    outputs(3427) <= not(layer0_outputs(2550));
    outputs(3428) <= not(layer0_outputs(5406)) or (layer0_outputs(7722));
    outputs(3429) <= layer0_outputs(5764);
    outputs(3430) <= (layer0_outputs(5818)) or (layer0_outputs(7522));
    outputs(3431) <= not(layer0_outputs(8330));
    outputs(3432) <= (layer0_outputs(573)) xor (layer0_outputs(4890));
    outputs(3433) <= not((layer0_outputs(9479)) or (layer0_outputs(10082)));
    outputs(3434) <= not((layer0_outputs(6783)) xor (layer0_outputs(2885)));
    outputs(3435) <= not((layer0_outputs(83)) xor (layer0_outputs(9056)));
    outputs(3436) <= (layer0_outputs(278)) and not (layer0_outputs(4368));
    outputs(3437) <= layer0_outputs(8422);
    outputs(3438) <= (layer0_outputs(9099)) and not (layer0_outputs(2463));
    outputs(3439) <= not(layer0_outputs(7360)) or (layer0_outputs(6938));
    outputs(3440) <= layer0_outputs(1167);
    outputs(3441) <= not(layer0_outputs(4787)) or (layer0_outputs(2720));
    outputs(3442) <= (layer0_outputs(4169)) and not (layer0_outputs(9450));
    outputs(3443) <= not(layer0_outputs(6182));
    outputs(3444) <= (layer0_outputs(8386)) and (layer0_outputs(9422));
    outputs(3445) <= not(layer0_outputs(3440));
    outputs(3446) <= not(layer0_outputs(755)) or (layer0_outputs(9644));
    outputs(3447) <= not((layer0_outputs(1530)) or (layer0_outputs(2126)));
    outputs(3448) <= layer0_outputs(5677);
    outputs(3449) <= not((layer0_outputs(9154)) or (layer0_outputs(3981)));
    outputs(3450) <= not(layer0_outputs(3676));
    outputs(3451) <= not(layer0_outputs(7267));
    outputs(3452) <= layer0_outputs(1963);
    outputs(3453) <= (layer0_outputs(483)) and (layer0_outputs(8198));
    outputs(3454) <= not((layer0_outputs(1621)) xor (layer0_outputs(9066)));
    outputs(3455) <= not((layer0_outputs(9418)) xor (layer0_outputs(23)));
    outputs(3456) <= not(layer0_outputs(1410));
    outputs(3457) <= not(layer0_outputs(7985));
    outputs(3458) <= layer0_outputs(4781);
    outputs(3459) <= layer0_outputs(5023);
    outputs(3460) <= (layer0_outputs(7121)) and (layer0_outputs(274));
    outputs(3461) <= (layer0_outputs(7544)) and (layer0_outputs(7752));
    outputs(3462) <= (layer0_outputs(8798)) and not (layer0_outputs(7273));
    outputs(3463) <= not((layer0_outputs(8065)) or (layer0_outputs(5599)));
    outputs(3464) <= (layer0_outputs(4870)) and (layer0_outputs(5904));
    outputs(3465) <= layer0_outputs(644);
    outputs(3466) <= layer0_outputs(746);
    outputs(3467) <= not((layer0_outputs(206)) or (layer0_outputs(6186)));
    outputs(3468) <= not(layer0_outputs(4966));
    outputs(3469) <= (layer0_outputs(6477)) and (layer0_outputs(8438));
    outputs(3470) <= (layer0_outputs(10088)) and not (layer0_outputs(8161));
    outputs(3471) <= not((layer0_outputs(2847)) and (layer0_outputs(1767)));
    outputs(3472) <= not((layer0_outputs(7284)) or (layer0_outputs(3634)));
    outputs(3473) <= not((layer0_outputs(4743)) or (layer0_outputs(5003)));
    outputs(3474) <= not(layer0_outputs(4553));
    outputs(3475) <= not(layer0_outputs(3451));
    outputs(3476) <= layer0_outputs(8994);
    outputs(3477) <= not((layer0_outputs(9500)) xor (layer0_outputs(6683)));
    outputs(3478) <= not(layer0_outputs(3379));
    outputs(3479) <= layer0_outputs(3127);
    outputs(3480) <= (layer0_outputs(4738)) xor (layer0_outputs(4845));
    outputs(3481) <= layer0_outputs(8642);
    outputs(3482) <= layer0_outputs(2902);
    outputs(3483) <= (layer0_outputs(6064)) and not (layer0_outputs(7813));
    outputs(3484) <= not((layer0_outputs(2952)) xor (layer0_outputs(6835)));
    outputs(3485) <= layer0_outputs(4888);
    outputs(3486) <= not(layer0_outputs(10138)) or (layer0_outputs(1929));
    outputs(3487) <= not((layer0_outputs(358)) xor (layer0_outputs(5458)));
    outputs(3488) <= (layer0_outputs(6627)) xor (layer0_outputs(4216));
    outputs(3489) <= not(layer0_outputs(2105));
    outputs(3490) <= not(layer0_outputs(1171));
    outputs(3491) <= not(layer0_outputs(8196));
    outputs(3492) <= not((layer0_outputs(10126)) xor (layer0_outputs(1321)));
    outputs(3493) <= not(layer0_outputs(9301)) or (layer0_outputs(3544));
    outputs(3494) <= not((layer0_outputs(9749)) xor (layer0_outputs(1656)));
    outputs(3495) <= not((layer0_outputs(554)) and (layer0_outputs(7651)));
    outputs(3496) <= layer0_outputs(8863);
    outputs(3497) <= not(layer0_outputs(5814));
    outputs(3498) <= not(layer0_outputs(7602));
    outputs(3499) <= not(layer0_outputs(6924));
    outputs(3500) <= not(layer0_outputs(9173)) or (layer0_outputs(3247));
    outputs(3501) <= (layer0_outputs(9141)) and (layer0_outputs(4016));
    outputs(3502) <= layer0_outputs(8155);
    outputs(3503) <= not(layer0_outputs(6368));
    outputs(3504) <= not(layer0_outputs(392));
    outputs(3505) <= (layer0_outputs(6485)) or (layer0_outputs(250));
    outputs(3506) <= not((layer0_outputs(8019)) or (layer0_outputs(159)));
    outputs(3507) <= not(layer0_outputs(6347));
    outputs(3508) <= layer0_outputs(371);
    outputs(3509) <= not((layer0_outputs(230)) and (layer0_outputs(1506)));
    outputs(3510) <= (layer0_outputs(3283)) and not (layer0_outputs(26));
    outputs(3511) <= not(layer0_outputs(7653)) or (layer0_outputs(566));
    outputs(3512) <= (layer0_outputs(953)) xor (layer0_outputs(5412));
    outputs(3513) <= layer0_outputs(6023);
    outputs(3514) <= not((layer0_outputs(7925)) or (layer0_outputs(2774)));
    outputs(3515) <= layer0_outputs(6382);
    outputs(3516) <= layer0_outputs(781);
    outputs(3517) <= (layer0_outputs(8269)) and not (layer0_outputs(271));
    outputs(3518) <= (layer0_outputs(797)) and (layer0_outputs(4389));
    outputs(3519) <= (layer0_outputs(500)) xor (layer0_outputs(2776));
    outputs(3520) <= (layer0_outputs(46)) xor (layer0_outputs(8848));
    outputs(3521) <= layer0_outputs(4008);
    outputs(3522) <= not(layer0_outputs(6500));
    outputs(3523) <= not(layer0_outputs(1026));
    outputs(3524) <= layer0_outputs(1404);
    outputs(3525) <= (layer0_outputs(8593)) and not (layer0_outputs(6316));
    outputs(3526) <= (layer0_outputs(7546)) or (layer0_outputs(989));
    outputs(3527) <= layer0_outputs(2893);
    outputs(3528) <= layer0_outputs(8654);
    outputs(3529) <= layer0_outputs(3587);
    outputs(3530) <= layer0_outputs(9074);
    outputs(3531) <= (layer0_outputs(982)) and (layer0_outputs(7716));
    outputs(3532) <= (layer0_outputs(1599)) xor (layer0_outputs(8534));
    outputs(3533) <= (layer0_outputs(8517)) and not (layer0_outputs(2124));
    outputs(3534) <= layer0_outputs(5927);
    outputs(3535) <= layer0_outputs(7014);
    outputs(3536) <= layer0_outputs(5256);
    outputs(3537) <= not(layer0_outputs(9886));
    outputs(3538) <= (layer0_outputs(10093)) and not (layer0_outputs(4776));
    outputs(3539) <= (layer0_outputs(8455)) xor (layer0_outputs(5599));
    outputs(3540) <= (layer0_outputs(3614)) or (layer0_outputs(10123));
    outputs(3541) <= not((layer0_outputs(1992)) xor (layer0_outputs(4037)));
    outputs(3542) <= not(layer0_outputs(1102));
    outputs(3543) <= (layer0_outputs(4030)) and not (layer0_outputs(5497));
    outputs(3544) <= not(layer0_outputs(901));
    outputs(3545) <= (layer0_outputs(5163)) and not (layer0_outputs(3439));
    outputs(3546) <= (layer0_outputs(918)) or (layer0_outputs(8868));
    outputs(3547) <= not(layer0_outputs(7175));
    outputs(3548) <= (layer0_outputs(4404)) xor (layer0_outputs(3126));
    outputs(3549) <= (layer0_outputs(7875)) xor (layer0_outputs(9621));
    outputs(3550) <= not(layer0_outputs(1085));
    outputs(3551) <= layer0_outputs(7981);
    outputs(3552) <= (layer0_outputs(142)) and (layer0_outputs(8232));
    outputs(3553) <= layer0_outputs(1212);
    outputs(3554) <= layer0_outputs(9406);
    outputs(3555) <= not(layer0_outputs(7705)) or (layer0_outputs(4209));
    outputs(3556) <= (layer0_outputs(1176)) xor (layer0_outputs(10237));
    outputs(3557) <= not((layer0_outputs(2478)) xor (layer0_outputs(8026)));
    outputs(3558) <= not((layer0_outputs(6532)) or (layer0_outputs(6962)));
    outputs(3559) <= (layer0_outputs(10012)) and not (layer0_outputs(289));
    outputs(3560) <= not((layer0_outputs(4134)) xor (layer0_outputs(6238)));
    outputs(3561) <= not(layer0_outputs(3878));
    outputs(3562) <= layer0_outputs(2392);
    outputs(3563) <= (layer0_outputs(6036)) or (layer0_outputs(5979));
    outputs(3564) <= (layer0_outputs(5091)) xor (layer0_outputs(6377));
    outputs(3565) <= layer0_outputs(8047);
    outputs(3566) <= not(layer0_outputs(796)) or (layer0_outputs(8361));
    outputs(3567) <= not((layer0_outputs(3327)) xor (layer0_outputs(8235)));
    outputs(3568) <= layer0_outputs(8974);
    outputs(3569) <= not(layer0_outputs(5007)) or (layer0_outputs(2663));
    outputs(3570) <= (layer0_outputs(56)) and (layer0_outputs(236));
    outputs(3571) <= not((layer0_outputs(6061)) or (layer0_outputs(7200)));
    outputs(3572) <= not(layer0_outputs(7297)) or (layer0_outputs(9350));
    outputs(3573) <= not((layer0_outputs(2463)) or (layer0_outputs(1135)));
    outputs(3574) <= (layer0_outputs(7298)) and not (layer0_outputs(4972));
    outputs(3575) <= not((layer0_outputs(8398)) xor (layer0_outputs(5099)));
    outputs(3576) <= (layer0_outputs(1412)) and (layer0_outputs(5915));
    outputs(3577) <= not(layer0_outputs(1797)) or (layer0_outputs(5503));
    outputs(3578) <= not((layer0_outputs(8855)) or (layer0_outputs(328)));
    outputs(3579) <= layer0_outputs(6860);
    outputs(3580) <= (layer0_outputs(1792)) and (layer0_outputs(1534));
    outputs(3581) <= layer0_outputs(5217);
    outputs(3582) <= not(layer0_outputs(6169));
    outputs(3583) <= not(layer0_outputs(860));
    outputs(3584) <= layer0_outputs(4080);
    outputs(3585) <= layer0_outputs(5289);
    outputs(3586) <= not(layer0_outputs(9554));
    outputs(3587) <= not(layer0_outputs(7080)) or (layer0_outputs(1588));
    outputs(3588) <= not(layer0_outputs(5757));
    outputs(3589) <= layer0_outputs(503);
    outputs(3590) <= not(layer0_outputs(3320));
    outputs(3591) <= layer0_outputs(8386);
    outputs(3592) <= not(layer0_outputs(2831)) or (layer0_outputs(8913));
    outputs(3593) <= not((layer0_outputs(1820)) or (layer0_outputs(2081)));
    outputs(3594) <= not((layer0_outputs(9563)) xor (layer0_outputs(7457)));
    outputs(3595) <= not(layer0_outputs(2157));
    outputs(3596) <= not(layer0_outputs(104));
    outputs(3597) <= (layer0_outputs(6515)) xor (layer0_outputs(8031));
    outputs(3598) <= (layer0_outputs(8822)) or (layer0_outputs(792));
    outputs(3599) <= not(layer0_outputs(6708));
    outputs(3600) <= (layer0_outputs(4210)) and not (layer0_outputs(4187));
    outputs(3601) <= not((layer0_outputs(2569)) xor (layer0_outputs(8622)));
    outputs(3602) <= (layer0_outputs(5711)) or (layer0_outputs(1565));
    outputs(3603) <= (layer0_outputs(5329)) and (layer0_outputs(3582));
    outputs(3604) <= not(layer0_outputs(7376));
    outputs(3605) <= (layer0_outputs(457)) xor (layer0_outputs(2435));
    outputs(3606) <= not(layer0_outputs(767));
    outputs(3607) <= (layer0_outputs(2248)) and (layer0_outputs(6303));
    outputs(3608) <= not(layer0_outputs(6706));
    outputs(3609) <= not((layer0_outputs(3593)) xor (layer0_outputs(8820)));
    outputs(3610) <= not((layer0_outputs(2444)) xor (layer0_outputs(4120)));
    outputs(3611) <= not((layer0_outputs(10212)) and (layer0_outputs(5402)));
    outputs(3612) <= (layer0_outputs(9675)) xor (layer0_outputs(1080));
    outputs(3613) <= not((layer0_outputs(1924)) or (layer0_outputs(6519)));
    outputs(3614) <= (layer0_outputs(10132)) or (layer0_outputs(7928));
    outputs(3615) <= layer0_outputs(2299);
    outputs(3616) <= layer0_outputs(3552);
    outputs(3617) <= layer0_outputs(7683);
    outputs(3618) <= layer0_outputs(3029);
    outputs(3619) <= not((layer0_outputs(8046)) xor (layer0_outputs(6334)));
    outputs(3620) <= not(layer0_outputs(3527));
    outputs(3621) <= not((layer0_outputs(8575)) xor (layer0_outputs(2689)));
    outputs(3622) <= layer0_outputs(4872);
    outputs(3623) <= not((layer0_outputs(3457)) xor (layer0_outputs(7341)));
    outputs(3624) <= not((layer0_outputs(3433)) xor (layer0_outputs(3695)));
    outputs(3625) <= not(layer0_outputs(9760));
    outputs(3626) <= not((layer0_outputs(6989)) or (layer0_outputs(9630)));
    outputs(3627) <= (layer0_outputs(7421)) xor (layer0_outputs(5404));
    outputs(3628) <= not((layer0_outputs(1409)) xor (layer0_outputs(1823)));
    outputs(3629) <= not(layer0_outputs(3096));
    outputs(3630) <= not(layer0_outputs(243)) or (layer0_outputs(5358));
    outputs(3631) <= not((layer0_outputs(1507)) xor (layer0_outputs(7710)));
    outputs(3632) <= layer0_outputs(611);
    outputs(3633) <= not((layer0_outputs(3089)) xor (layer0_outputs(9879)));
    outputs(3634) <= not(layer0_outputs(1641));
    outputs(3635) <= not(layer0_outputs(1114));
    outputs(3636) <= not(layer0_outputs(8277));
    outputs(3637) <= (layer0_outputs(3073)) xor (layer0_outputs(3919));
    outputs(3638) <= (layer0_outputs(6984)) xor (layer0_outputs(5813));
    outputs(3639) <= not(layer0_outputs(4827));
    outputs(3640) <= not(layer0_outputs(8446));
    outputs(3641) <= not(layer0_outputs(5221));
    outputs(3642) <= not(layer0_outputs(3978));
    outputs(3643) <= not(layer0_outputs(1155));
    outputs(3644) <= (layer0_outputs(704)) and (layer0_outputs(8703));
    outputs(3645) <= not(layer0_outputs(3824)) or (layer0_outputs(7969));
    outputs(3646) <= not((layer0_outputs(8603)) xor (layer0_outputs(7911)));
    outputs(3647) <= (layer0_outputs(9639)) or (layer0_outputs(9249));
    outputs(3648) <= layer0_outputs(8577);
    outputs(3649) <= not((layer0_outputs(248)) or (layer0_outputs(9602)));
    outputs(3650) <= layer0_outputs(7969);
    outputs(3651) <= not(layer0_outputs(1570));
    outputs(3652) <= (layer0_outputs(4386)) and (layer0_outputs(7424));
    outputs(3653) <= layer0_outputs(5392);
    outputs(3654) <= (layer0_outputs(1758)) or (layer0_outputs(7831));
    outputs(3655) <= (layer0_outputs(3590)) xor (layer0_outputs(3216));
    outputs(3656) <= layer0_outputs(1232);
    outputs(3657) <= not((layer0_outputs(9584)) xor (layer0_outputs(182)));
    outputs(3658) <= (layer0_outputs(8201)) and (layer0_outputs(8170));
    outputs(3659) <= layer0_outputs(5115);
    outputs(3660) <= (layer0_outputs(4081)) xor (layer0_outputs(4105));
    outputs(3661) <= not(layer0_outputs(1896));
    outputs(3662) <= layer0_outputs(6291);
    outputs(3663) <= layer0_outputs(9488);
    outputs(3664) <= not(layer0_outputs(4089));
    outputs(3665) <= not(layer0_outputs(1140));
    outputs(3666) <= layer0_outputs(2525);
    outputs(3667) <= layer0_outputs(3425);
    outputs(3668) <= not(layer0_outputs(5320));
    outputs(3669) <= not(layer0_outputs(6011));
    outputs(3670) <= not(layer0_outputs(2984));
    outputs(3671) <= not(layer0_outputs(8794));
    outputs(3672) <= not(layer0_outputs(9290)) or (layer0_outputs(9786));
    outputs(3673) <= not(layer0_outputs(7563));
    outputs(3674) <= not(layer0_outputs(7282));
    outputs(3675) <= not((layer0_outputs(417)) xor (layer0_outputs(1369)));
    outputs(3676) <= not((layer0_outputs(4174)) or (layer0_outputs(5440)));
    outputs(3677) <= not(layer0_outputs(7481));
    outputs(3678) <= (layer0_outputs(1864)) xor (layer0_outputs(4542));
    outputs(3679) <= layer0_outputs(8747);
    outputs(3680) <= not(layer0_outputs(7325));
    outputs(3681) <= not((layer0_outputs(2185)) xor (layer0_outputs(5852)));
    outputs(3682) <= not(layer0_outputs(940)) or (layer0_outputs(9273));
    outputs(3683) <= not(layer0_outputs(9256)) or (layer0_outputs(9069));
    outputs(3684) <= (layer0_outputs(1993)) and not (layer0_outputs(1438));
    outputs(3685) <= not((layer0_outputs(5804)) or (layer0_outputs(2793)));
    outputs(3686) <= (layer0_outputs(2635)) or (layer0_outputs(3422));
    outputs(3687) <= (layer0_outputs(8970)) and not (layer0_outputs(7802));
    outputs(3688) <= not(layer0_outputs(4628));
    outputs(3689) <= not(layer0_outputs(10206)) or (layer0_outputs(4379));
    outputs(3690) <= not((layer0_outputs(3117)) or (layer0_outputs(6265)));
    outputs(3691) <= not(layer0_outputs(6528));
    outputs(3692) <= not(layer0_outputs(6941));
    outputs(3693) <= (layer0_outputs(6353)) and not (layer0_outputs(5000));
    outputs(3694) <= not(layer0_outputs(8024));
    outputs(3695) <= (layer0_outputs(4603)) or (layer0_outputs(7142));
    outputs(3696) <= (layer0_outputs(479)) and not (layer0_outputs(5940));
    outputs(3697) <= (layer0_outputs(7888)) and not (layer0_outputs(1034));
    outputs(3698) <= (layer0_outputs(3602)) and (layer0_outputs(9053));
    outputs(3699) <= (layer0_outputs(6462)) and not (layer0_outputs(594));
    outputs(3700) <= not(layer0_outputs(8558));
    outputs(3701) <= layer0_outputs(3865);
    outputs(3702) <= (layer0_outputs(9512)) and not (layer0_outputs(4838));
    outputs(3703) <= (layer0_outputs(1635)) xor (layer0_outputs(942));
    outputs(3704) <= not(layer0_outputs(8344)) or (layer0_outputs(1469));
    outputs(3705) <= not(layer0_outputs(8068)) or (layer0_outputs(10156));
    outputs(3706) <= (layer0_outputs(853)) and not (layer0_outputs(5816));
    outputs(3707) <= (layer0_outputs(3639)) xor (layer0_outputs(3613));
    outputs(3708) <= not((layer0_outputs(2798)) or (layer0_outputs(5096)));
    outputs(3709) <= not((layer0_outputs(4149)) xor (layer0_outputs(5475)));
    outputs(3710) <= not(layer0_outputs(9362));
    outputs(3711) <= (layer0_outputs(797)) and not (layer0_outputs(9042));
    outputs(3712) <= layer0_outputs(9329);
    outputs(3713) <= not(layer0_outputs(3770));
    outputs(3714) <= (layer0_outputs(928)) xor (layer0_outputs(1363));
    outputs(3715) <= '0';
    outputs(3716) <= not(layer0_outputs(4458));
    outputs(3717) <= layer0_outputs(8972);
    outputs(3718) <= (layer0_outputs(9626)) and not (layer0_outputs(6193));
    outputs(3719) <= not(layer0_outputs(807));
    outputs(3720) <= layer0_outputs(9611);
    outputs(3721) <= not(layer0_outputs(1578));
    outputs(3722) <= not(layer0_outputs(5565));
    outputs(3723) <= (layer0_outputs(3385)) and not (layer0_outputs(198));
    outputs(3724) <= (layer0_outputs(8235)) xor (layer0_outputs(7725));
    outputs(3725) <= not(layer0_outputs(4243)) or (layer0_outputs(5372));
    outputs(3726) <= not(layer0_outputs(3404));
    outputs(3727) <= not((layer0_outputs(7360)) and (layer0_outputs(8833)));
    outputs(3728) <= not((layer0_outputs(7516)) xor (layer0_outputs(9531)));
    outputs(3729) <= (layer0_outputs(2458)) and (layer0_outputs(150));
    outputs(3730) <= not((layer0_outputs(6332)) or (layer0_outputs(3410)));
    outputs(3731) <= not(layer0_outputs(10229)) or (layer0_outputs(5213));
    outputs(3732) <= (layer0_outputs(267)) and not (layer0_outputs(5810));
    outputs(3733) <= layer0_outputs(5760);
    outputs(3734) <= not(layer0_outputs(4662)) or (layer0_outputs(6392));
    outputs(3735) <= layer0_outputs(6136);
    outputs(3736) <= (layer0_outputs(7869)) xor (layer0_outputs(5128));
    outputs(3737) <= not((layer0_outputs(8496)) xor (layer0_outputs(8897)));
    outputs(3738) <= layer0_outputs(3898);
    outputs(3739) <= not((layer0_outputs(6192)) xor (layer0_outputs(9150)));
    outputs(3740) <= (layer0_outputs(6645)) and (layer0_outputs(6952));
    outputs(3741) <= layer0_outputs(7134);
    outputs(3742) <= not(layer0_outputs(3427));
    outputs(3743) <= (layer0_outputs(9320)) xor (layer0_outputs(4010));
    outputs(3744) <= (layer0_outputs(9810)) xor (layer0_outputs(8187));
    outputs(3745) <= not((layer0_outputs(9040)) xor (layer0_outputs(6051)));
    outputs(3746) <= layer0_outputs(370);
    outputs(3747) <= not((layer0_outputs(3237)) xor (layer0_outputs(4250)));
    outputs(3748) <= not(layer0_outputs(7541));
    outputs(3749) <= (layer0_outputs(4350)) and not (layer0_outputs(5290));
    outputs(3750) <= layer0_outputs(5377);
    outputs(3751) <= not((layer0_outputs(2623)) xor (layer0_outputs(2378)));
    outputs(3752) <= not(layer0_outputs(1117));
    outputs(3753) <= not((layer0_outputs(1501)) xor (layer0_outputs(9974)));
    outputs(3754) <= (layer0_outputs(4389)) and (layer0_outputs(2691));
    outputs(3755) <= layer0_outputs(491);
    outputs(3756) <= (layer0_outputs(3772)) and not (layer0_outputs(1696));
    outputs(3757) <= (layer0_outputs(1194)) xor (layer0_outputs(2424));
    outputs(3758) <= layer0_outputs(3385);
    outputs(3759) <= not(layer0_outputs(5721));
    outputs(3760) <= (layer0_outputs(9778)) xor (layer0_outputs(9359));
    outputs(3761) <= not(layer0_outputs(1582));
    outputs(3762) <= layer0_outputs(5979);
    outputs(3763) <= (layer0_outputs(8953)) xor (layer0_outputs(4497));
    outputs(3764) <= not((layer0_outputs(1553)) xor (layer0_outputs(6041)));
    outputs(3765) <= layer0_outputs(5078);
    outputs(3766) <= not(layer0_outputs(1289));
    outputs(3767) <= (layer0_outputs(3243)) and not (layer0_outputs(9987));
    outputs(3768) <= not((layer0_outputs(743)) or (layer0_outputs(6798)));
    outputs(3769) <= not(layer0_outputs(2082)) or (layer0_outputs(1575));
    outputs(3770) <= not(layer0_outputs(5366)) or (layer0_outputs(8737));
    outputs(3771) <= not(layer0_outputs(1580));
    outputs(3772) <= not(layer0_outputs(1450)) or (layer0_outputs(8857));
    outputs(3773) <= (layer0_outputs(7723)) xor (layer0_outputs(4132));
    outputs(3774) <= layer0_outputs(1811);
    outputs(3775) <= not(layer0_outputs(778));
    outputs(3776) <= layer0_outputs(7981);
    outputs(3777) <= not((layer0_outputs(6419)) xor (layer0_outputs(5717)));
    outputs(3778) <= layer0_outputs(5265);
    outputs(3779) <= layer0_outputs(3516);
    outputs(3780) <= not((layer0_outputs(629)) or (layer0_outputs(2323)));
    outputs(3781) <= (layer0_outputs(4009)) and not (layer0_outputs(9191));
    outputs(3782) <= (layer0_outputs(2878)) or (layer0_outputs(836));
    outputs(3783) <= (layer0_outputs(6575)) xor (layer0_outputs(2975));
    outputs(3784) <= not((layer0_outputs(856)) xor (layer0_outputs(6761)));
    outputs(3785) <= not((layer0_outputs(5357)) or (layer0_outputs(3045)));
    outputs(3786) <= not(layer0_outputs(4413));
    outputs(3787) <= layer0_outputs(7880);
    outputs(3788) <= (layer0_outputs(264)) xor (layer0_outputs(7483));
    outputs(3789) <= not(layer0_outputs(5508));
    outputs(3790) <= not(layer0_outputs(9793)) or (layer0_outputs(9453));
    outputs(3791) <= layer0_outputs(8601);
    outputs(3792) <= layer0_outputs(7825);
    outputs(3793) <= (layer0_outputs(2900)) and not (layer0_outputs(8241));
    outputs(3794) <= (layer0_outputs(9681)) or (layer0_outputs(2805));
    outputs(3795) <= layer0_outputs(2533);
    outputs(3796) <= (layer0_outputs(3756)) xor (layer0_outputs(8771));
    outputs(3797) <= layer0_outputs(9084);
    outputs(3798) <= not(layer0_outputs(8071));
    outputs(3799) <= (layer0_outputs(2968)) xor (layer0_outputs(5075));
    outputs(3800) <= (layer0_outputs(8769)) and not (layer0_outputs(2480));
    outputs(3801) <= layer0_outputs(2319);
    outputs(3802) <= (layer0_outputs(8056)) and not (layer0_outputs(8284));
    outputs(3803) <= not((layer0_outputs(5483)) or (layer0_outputs(2065)));
    outputs(3804) <= not(layer0_outputs(7480));
    outputs(3805) <= layer0_outputs(8409);
    outputs(3806) <= layer0_outputs(1598);
    outputs(3807) <= not((layer0_outputs(3103)) xor (layer0_outputs(10228)));
    outputs(3808) <= layer0_outputs(4749);
    outputs(3809) <= not((layer0_outputs(3966)) xor (layer0_outputs(923)));
    outputs(3810) <= layer0_outputs(7872);
    outputs(3811) <= layer0_outputs(2832);
    outputs(3812) <= not(layer0_outputs(8008));
    outputs(3813) <= not(layer0_outputs(374));
    outputs(3814) <= not((layer0_outputs(3720)) xor (layer0_outputs(5324)));
    outputs(3815) <= not(layer0_outputs(3770)) or (layer0_outputs(21));
    outputs(3816) <= not(layer0_outputs(843));
    outputs(3817) <= layer0_outputs(7600);
    outputs(3818) <= not((layer0_outputs(9161)) xor (layer0_outputs(3282)));
    outputs(3819) <= (layer0_outputs(4250)) xor (layer0_outputs(798));
    outputs(3820) <= layer0_outputs(9583);
    outputs(3821) <= not((layer0_outputs(6831)) xor (layer0_outputs(451)));
    outputs(3822) <= (layer0_outputs(2889)) xor (layer0_outputs(2626));
    outputs(3823) <= not((layer0_outputs(1)) xor (layer0_outputs(2878)));
    outputs(3824) <= (layer0_outputs(9097)) and not (layer0_outputs(6708));
    outputs(3825) <= (layer0_outputs(9010)) xor (layer0_outputs(2358));
    outputs(3826) <= layer0_outputs(9953);
    outputs(3827) <= (layer0_outputs(3375)) xor (layer0_outputs(7662));
    outputs(3828) <= (layer0_outputs(4290)) xor (layer0_outputs(3740));
    outputs(3829) <= (layer0_outputs(10010)) xor (layer0_outputs(7070));
    outputs(3830) <= not((layer0_outputs(8334)) xor (layer0_outputs(4582)));
    outputs(3831) <= layer0_outputs(4298);
    outputs(3832) <= not(layer0_outputs(2911));
    outputs(3833) <= not(layer0_outputs(3694)) or (layer0_outputs(1346));
    outputs(3834) <= not(layer0_outputs(3223));
    outputs(3835) <= not((layer0_outputs(5000)) or (layer0_outputs(3526)));
    outputs(3836) <= layer0_outputs(4796);
    outputs(3837) <= layer0_outputs(8853);
    outputs(3838) <= (layer0_outputs(9407)) xor (layer0_outputs(6704));
    outputs(3839) <= not(layer0_outputs(3293));
    outputs(3840) <= (layer0_outputs(3262)) and not (layer0_outputs(9909));
    outputs(3841) <= (layer0_outputs(7822)) and not (layer0_outputs(6702));
    outputs(3842) <= not(layer0_outputs(2851));
    outputs(3843) <= (layer0_outputs(568)) and (layer0_outputs(145));
    outputs(3844) <= (layer0_outputs(4139)) xor (layer0_outputs(3193));
    outputs(3845) <= not(layer0_outputs(6116));
    outputs(3846) <= layer0_outputs(5211);
    outputs(3847) <= (layer0_outputs(3735)) xor (layer0_outputs(8208));
    outputs(3848) <= (layer0_outputs(3991)) xor (layer0_outputs(8502));
    outputs(3849) <= not(layer0_outputs(2851));
    outputs(3850) <= not(layer0_outputs(2659));
    outputs(3851) <= not(layer0_outputs(4438));
    outputs(3852) <= not(layer0_outputs(9230));
    outputs(3853) <= not(layer0_outputs(4933));
    outputs(3854) <= not(layer0_outputs(6695));
    outputs(3855) <= layer0_outputs(5162);
    outputs(3856) <= (layer0_outputs(1215)) xor (layer0_outputs(4123));
    outputs(3857) <= not(layer0_outputs(5500)) or (layer0_outputs(8877));
    outputs(3858) <= not((layer0_outputs(3801)) or (layer0_outputs(2895)));
    outputs(3859) <= layer0_outputs(6412);
    outputs(3860) <= (layer0_outputs(5030)) xor (layer0_outputs(1923));
    outputs(3861) <= (layer0_outputs(7011)) or (layer0_outputs(1986));
    outputs(3862) <= (layer0_outputs(2394)) and (layer0_outputs(4407));
    outputs(3863) <= (layer0_outputs(2982)) and not (layer0_outputs(3973));
    outputs(3864) <= layer0_outputs(253);
    outputs(3865) <= not((layer0_outputs(6928)) or (layer0_outputs(7718)));
    outputs(3866) <= (layer0_outputs(6601)) xor (layer0_outputs(5426));
    outputs(3867) <= (layer0_outputs(9204)) and not (layer0_outputs(9026));
    outputs(3868) <= (layer0_outputs(7269)) or (layer0_outputs(7007));
    outputs(3869) <= (layer0_outputs(3310)) and not (layer0_outputs(3318));
    outputs(3870) <= layer0_outputs(7246);
    outputs(3871) <= not(layer0_outputs(9291)) or (layer0_outputs(6392));
    outputs(3872) <= (layer0_outputs(4017)) and (layer0_outputs(8774));
    outputs(3873) <= not((layer0_outputs(2351)) xor (layer0_outputs(3820)));
    outputs(3874) <= not(layer0_outputs(10183));
    outputs(3875) <= (layer0_outputs(2944)) xor (layer0_outputs(7545));
    outputs(3876) <= not((layer0_outputs(1694)) or (layer0_outputs(8715)));
    outputs(3877) <= layer0_outputs(9542);
    outputs(3878) <= layer0_outputs(8567);
    outputs(3879) <= not(layer0_outputs(5484));
    outputs(3880) <= not(layer0_outputs(3518));
    outputs(3881) <= not(layer0_outputs(4751));
    outputs(3882) <= not(layer0_outputs(4372));
    outputs(3883) <= (layer0_outputs(4522)) and not (layer0_outputs(2509));
    outputs(3884) <= not(layer0_outputs(9924));
    outputs(3885) <= (layer0_outputs(8778)) and not (layer0_outputs(9433));
    outputs(3886) <= (layer0_outputs(9960)) xor (layer0_outputs(2785));
    outputs(3887) <= layer0_outputs(3629);
    outputs(3888) <= not((layer0_outputs(9258)) or (layer0_outputs(7075)));
    outputs(3889) <= layer0_outputs(67);
    outputs(3890) <= not(layer0_outputs(8783));
    outputs(3891) <= not((layer0_outputs(6240)) xor (layer0_outputs(9296)));
    outputs(3892) <= (layer0_outputs(614)) xor (layer0_outputs(3877));
    outputs(3893) <= layer0_outputs(1524);
    outputs(3894) <= (layer0_outputs(3173)) xor (layer0_outputs(3279));
    outputs(3895) <= not((layer0_outputs(669)) xor (layer0_outputs(5582)));
    outputs(3896) <= layer0_outputs(3238);
    outputs(3897) <= not(layer0_outputs(1371));
    outputs(3898) <= not(layer0_outputs(8888));
    outputs(3899) <= (layer0_outputs(1729)) xor (layer0_outputs(7184));
    outputs(3900) <= not((layer0_outputs(4664)) or (layer0_outputs(300)));
    outputs(3901) <= (layer0_outputs(4601)) xor (layer0_outputs(8289));
    outputs(3902) <= not(layer0_outputs(8840));
    outputs(3903) <= not((layer0_outputs(6508)) xor (layer0_outputs(1809)));
    outputs(3904) <= layer0_outputs(6870);
    outputs(3905) <= layer0_outputs(3486);
    outputs(3906) <= (layer0_outputs(6357)) and not (layer0_outputs(5769));
    outputs(3907) <= not((layer0_outputs(8169)) xor (layer0_outputs(2824)));
    outputs(3908) <= layer0_outputs(6520);
    outputs(3909) <= not(layer0_outputs(6931)) or (layer0_outputs(2744));
    outputs(3910) <= (layer0_outputs(2220)) xor (layer0_outputs(8353));
    outputs(3911) <= layer0_outputs(1590);
    outputs(3912) <= not(layer0_outputs(7514)) or (layer0_outputs(8642));
    outputs(3913) <= (layer0_outputs(8877)) and not (layer0_outputs(9730));
    outputs(3914) <= not(layer0_outputs(1360));
    outputs(3915) <= not(layer0_outputs(254)) or (layer0_outputs(8509));
    outputs(3916) <= (layer0_outputs(9894)) and not (layer0_outputs(621));
    outputs(3917) <= not(layer0_outputs(7189));
    outputs(3918) <= not((layer0_outputs(8292)) xor (layer0_outputs(9260)));
    outputs(3919) <= (layer0_outputs(8431)) and not (layer0_outputs(9519));
    outputs(3920) <= not(layer0_outputs(2685));
    outputs(3921) <= layer0_outputs(507);
    outputs(3922) <= (layer0_outputs(4038)) xor (layer0_outputs(296));
    outputs(3923) <= not(layer0_outputs(5708)) or (layer0_outputs(6766));
    outputs(3924) <= not(layer0_outputs(9793)) or (layer0_outputs(9926));
    outputs(3925) <= not(layer0_outputs(7436));
    outputs(3926) <= (layer0_outputs(10061)) xor (layer0_outputs(2268));
    outputs(3927) <= not((layer0_outputs(5676)) xor (layer0_outputs(7333)));
    outputs(3928) <= not(layer0_outputs(1));
    outputs(3929) <= not((layer0_outputs(9947)) xor (layer0_outputs(4980)));
    outputs(3930) <= layer0_outputs(9728);
    outputs(3931) <= not((layer0_outputs(3410)) xor (layer0_outputs(2237)));
    outputs(3932) <= not(layer0_outputs(2071));
    outputs(3933) <= (layer0_outputs(6568)) and (layer0_outputs(1753));
    outputs(3934) <= not(layer0_outputs(9847));
    outputs(3935) <= (layer0_outputs(5722)) and not (layer0_outputs(4956));
    outputs(3936) <= not(layer0_outputs(597)) or (layer0_outputs(5531));
    outputs(3937) <= not(layer0_outputs(7190));
    outputs(3938) <= not((layer0_outputs(5881)) and (layer0_outputs(2150)));
    outputs(3939) <= (layer0_outputs(7977)) and not (layer0_outputs(8237));
    outputs(3940) <= (layer0_outputs(8323)) and not (layer0_outputs(515));
    outputs(3941) <= not(layer0_outputs(681)) or (layer0_outputs(10186));
    outputs(3942) <= (layer0_outputs(1528)) and not (layer0_outputs(5063));
    outputs(3943) <= not((layer0_outputs(1280)) xor (layer0_outputs(6540)));
    outputs(3944) <= (layer0_outputs(2999)) or (layer0_outputs(8303));
    outputs(3945) <= not(layer0_outputs(2935));
    outputs(3946) <= layer0_outputs(1445);
    outputs(3947) <= not(layer0_outputs(4885));
    outputs(3948) <= layer0_outputs(4330);
    outputs(3949) <= not((layer0_outputs(1544)) xor (layer0_outputs(168)));
    outputs(3950) <= not(layer0_outputs(9800));
    outputs(3951) <= not((layer0_outputs(1489)) xor (layer0_outputs(3520)));
    outputs(3952) <= (layer0_outputs(841)) or (layer0_outputs(5107));
    outputs(3953) <= not(layer0_outputs(6511));
    outputs(3954) <= (layer0_outputs(6353)) and (layer0_outputs(506));
    outputs(3955) <= (layer0_outputs(8696)) xor (layer0_outputs(8933));
    outputs(3956) <= not(layer0_outputs(596));
    outputs(3957) <= (layer0_outputs(5682)) and not (layer0_outputs(1762));
    outputs(3958) <= not((layer0_outputs(4311)) xor (layer0_outputs(1652)));
    outputs(3959) <= (layer0_outputs(1006)) and (layer0_outputs(5849));
    outputs(3960) <= not(layer0_outputs(7471));
    outputs(3961) <= layer0_outputs(5955);
    outputs(3962) <= layer0_outputs(8925);
    outputs(3963) <= not((layer0_outputs(7201)) and (layer0_outputs(3515)));
    outputs(3964) <= not(layer0_outputs(1705)) or (layer0_outputs(3179));
    outputs(3965) <= layer0_outputs(8769);
    outputs(3966) <= not(layer0_outputs(1684));
    outputs(3967) <= not((layer0_outputs(10213)) and (layer0_outputs(5430)));
    outputs(3968) <= (layer0_outputs(9005)) xor (layer0_outputs(7553));
    outputs(3969) <= not((layer0_outputs(9519)) and (layer0_outputs(4286)));
    outputs(3970) <= (layer0_outputs(4575)) xor (layer0_outputs(10081));
    outputs(3971) <= layer0_outputs(1912);
    outputs(3972) <= not((layer0_outputs(7104)) or (layer0_outputs(7217)));
    outputs(3973) <= not((layer0_outputs(784)) xor (layer0_outputs(611)));
    outputs(3974) <= not((layer0_outputs(1088)) or (layer0_outputs(8692)));
    outputs(3975) <= layer0_outputs(5913);
    outputs(3976) <= layer0_outputs(754);
    outputs(3977) <= not((layer0_outputs(6917)) and (layer0_outputs(4883)));
    outputs(3978) <= layer0_outputs(4082);
    outputs(3979) <= not(layer0_outputs(5733));
    outputs(3980) <= (layer0_outputs(4316)) and (layer0_outputs(7271));
    outputs(3981) <= (layer0_outputs(9867)) xor (layer0_outputs(2223));
    outputs(3982) <= (layer0_outputs(151)) or (layer0_outputs(7614));
    outputs(3983) <= not(layer0_outputs(5499));
    outputs(3984) <= not((layer0_outputs(6492)) xor (layer0_outputs(8701)));
    outputs(3985) <= (layer0_outputs(3993)) xor (layer0_outputs(7618));
    outputs(3986) <= not((layer0_outputs(5016)) xor (layer0_outputs(4863)));
    outputs(3987) <= (layer0_outputs(2977)) and not (layer0_outputs(2986));
    outputs(3988) <= not(layer0_outputs(3907)) or (layer0_outputs(8229));
    outputs(3989) <= (layer0_outputs(3244)) xor (layer0_outputs(9902));
    outputs(3990) <= not((layer0_outputs(3463)) or (layer0_outputs(1423)));
    outputs(3991) <= not((layer0_outputs(4820)) or (layer0_outputs(5350)));
    outputs(3992) <= not((layer0_outputs(1510)) xor (layer0_outputs(9302)));
    outputs(3993) <= not((layer0_outputs(6495)) or (layer0_outputs(9980)));
    outputs(3994) <= not((layer0_outputs(7944)) xor (layer0_outputs(9629)));
    outputs(3995) <= layer0_outputs(8332);
    outputs(3996) <= not(layer0_outputs(1937));
    outputs(3997) <= not(layer0_outputs(4165)) or (layer0_outputs(5196));
    outputs(3998) <= layer0_outputs(1335);
    outputs(3999) <= not((layer0_outputs(9162)) and (layer0_outputs(8864)));
    outputs(4000) <= not(layer0_outputs(9871));
    outputs(4001) <= layer0_outputs(83);
    outputs(4002) <= layer0_outputs(9636);
    outputs(4003) <= (layer0_outputs(949)) and not (layer0_outputs(926));
    outputs(4004) <= (layer0_outputs(872)) xor (layer0_outputs(5884));
    outputs(4005) <= (layer0_outputs(29)) or (layer0_outputs(8890));
    outputs(4006) <= not(layer0_outputs(5747));
    outputs(4007) <= not((layer0_outputs(5421)) xor (layer0_outputs(2194)));
    outputs(4008) <= not(layer0_outputs(9343));
    outputs(4009) <= not((layer0_outputs(6566)) or (layer0_outputs(6495)));
    outputs(4010) <= not(layer0_outputs(7118)) or (layer0_outputs(5314));
    outputs(4011) <= (layer0_outputs(5756)) and not (layer0_outputs(6073));
    outputs(4012) <= (layer0_outputs(2100)) and not (layer0_outputs(8609));
    outputs(4013) <= not((layer0_outputs(4235)) xor (layer0_outputs(2143)));
    outputs(4014) <= not((layer0_outputs(2302)) xor (layer0_outputs(2381)));
    outputs(4015) <= layer0_outputs(4612);
    outputs(4016) <= (layer0_outputs(6577)) and (layer0_outputs(1966));
    outputs(4017) <= not((layer0_outputs(6789)) xor (layer0_outputs(8483)));
    outputs(4018) <= layer0_outputs(6119);
    outputs(4019) <= (layer0_outputs(455)) xor (layer0_outputs(5125));
    outputs(4020) <= not((layer0_outputs(3553)) or (layer0_outputs(8878)));
    outputs(4021) <= (layer0_outputs(7295)) and not (layer0_outputs(697));
    outputs(4022) <= (layer0_outputs(850)) or (layer0_outputs(1401));
    outputs(4023) <= not(layer0_outputs(6187));
    outputs(4024) <= not(layer0_outputs(3831));
    outputs(4025) <= (layer0_outputs(10182)) and not (layer0_outputs(5476));
    outputs(4026) <= not((layer0_outputs(1325)) xor (layer0_outputs(4838)));
    outputs(4027) <= not(layer0_outputs(871));
    outputs(4028) <= not(layer0_outputs(3983)) or (layer0_outputs(6852));
    outputs(4029) <= not((layer0_outputs(6161)) xor (layer0_outputs(8097)));
    outputs(4030) <= not((layer0_outputs(8582)) xor (layer0_outputs(5454)));
    outputs(4031) <= (layer0_outputs(2017)) xor (layer0_outputs(1035));
    outputs(4032) <= layer0_outputs(9703);
    outputs(4033) <= not(layer0_outputs(8377)) or (layer0_outputs(2217));
    outputs(4034) <= (layer0_outputs(7447)) and not (layer0_outputs(9766));
    outputs(4035) <= not((layer0_outputs(9529)) or (layer0_outputs(8069)));
    outputs(4036) <= not((layer0_outputs(6889)) and (layer0_outputs(4618)));
    outputs(4037) <= layer0_outputs(8298);
    outputs(4038) <= not(layer0_outputs(5388));
    outputs(4039) <= not(layer0_outputs(3591));
    outputs(4040) <= (layer0_outputs(7733)) and (layer0_outputs(3257));
    outputs(4041) <= not(layer0_outputs(8506));
    outputs(4042) <= not((layer0_outputs(5894)) xor (layer0_outputs(186)));
    outputs(4043) <= (layer0_outputs(3241)) and not (layer0_outputs(8545));
    outputs(4044) <= (layer0_outputs(2717)) xor (layer0_outputs(5013));
    outputs(4045) <= (layer0_outputs(7353)) and (layer0_outputs(6583));
    outputs(4046) <= (layer0_outputs(3818)) and not (layer0_outputs(314));
    outputs(4047) <= layer0_outputs(5686);
    outputs(4048) <= not(layer0_outputs(641));
    outputs(4049) <= not((layer0_outputs(7631)) xor (layer0_outputs(355)));
    outputs(4050) <= not(layer0_outputs(3245));
    outputs(4051) <= not(layer0_outputs(8110));
    outputs(4052) <= layer0_outputs(1395);
    outputs(4053) <= not((layer0_outputs(2451)) xor (layer0_outputs(5591)));
    outputs(4054) <= not((layer0_outputs(4646)) xor (layer0_outputs(1249)));
    outputs(4055) <= (layer0_outputs(8389)) or (layer0_outputs(1752));
    outputs(4056) <= (layer0_outputs(3594)) or (layer0_outputs(1940));
    outputs(4057) <= not(layer0_outputs(761));
    outputs(4058) <= not((layer0_outputs(5201)) or (layer0_outputs(7032)));
    outputs(4059) <= layer0_outputs(1467);
    outputs(4060) <= (layer0_outputs(7078)) and not (layer0_outputs(3782));
    outputs(4061) <= layer0_outputs(1859);
    outputs(4062) <= not(layer0_outputs(6782));
    outputs(4063) <= not(layer0_outputs(8682));
    outputs(4064) <= (layer0_outputs(7047)) and not (layer0_outputs(1573));
    outputs(4065) <= not(layer0_outputs(9288));
    outputs(4066) <= not(layer0_outputs(693));
    outputs(4067) <= not(layer0_outputs(5268));
    outputs(4068) <= (layer0_outputs(7735)) and (layer0_outputs(8657));
    outputs(4069) <= not((layer0_outputs(8402)) or (layer0_outputs(8777)));
    outputs(4070) <= not(layer0_outputs(3065));
    outputs(4071) <= layer0_outputs(3765);
    outputs(4072) <= not(layer0_outputs(374));
    outputs(4073) <= (layer0_outputs(4679)) xor (layer0_outputs(3378));
    outputs(4074) <= layer0_outputs(5957);
    outputs(4075) <= layer0_outputs(7133);
    outputs(4076) <= not((layer0_outputs(7040)) xor (layer0_outputs(1981)));
    outputs(4077) <= (layer0_outputs(4884)) and (layer0_outputs(3093));
    outputs(4078) <= (layer0_outputs(629)) xor (layer0_outputs(2493));
    outputs(4079) <= layer0_outputs(4481);
    outputs(4080) <= not(layer0_outputs(4899));
    outputs(4081) <= not(layer0_outputs(325));
    outputs(4082) <= (layer0_outputs(1396)) and (layer0_outputs(8819));
    outputs(4083) <= not(layer0_outputs(8809));
    outputs(4084) <= not(layer0_outputs(2276));
    outputs(4085) <= not(layer0_outputs(7076));
    outputs(4086) <= (layer0_outputs(8157)) xor (layer0_outputs(1874));
    outputs(4087) <= not(layer0_outputs(5461));
    outputs(4088) <= layer0_outputs(7489);
    outputs(4089) <= not(layer0_outputs(2405));
    outputs(4090) <= layer0_outputs(7479);
    outputs(4091) <= not(layer0_outputs(751));
    outputs(4092) <= (layer0_outputs(5298)) and (layer0_outputs(7294));
    outputs(4093) <= not((layer0_outputs(5740)) and (layer0_outputs(8450)));
    outputs(4094) <= (layer0_outputs(9684)) and not (layer0_outputs(4561));
    outputs(4095) <= not(layer0_outputs(7925));
    outputs(4096) <= layer0_outputs(5632);
    outputs(4097) <= layer0_outputs(2727);
    outputs(4098) <= (layer0_outputs(3930)) and (layer0_outputs(2817));
    outputs(4099) <= not((layer0_outputs(6111)) xor (layer0_outputs(2519)));
    outputs(4100) <= not((layer0_outputs(10225)) xor (layer0_outputs(7144)));
    outputs(4101) <= not(layer0_outputs(9289));
    outputs(4102) <= (layer0_outputs(7445)) and not (layer0_outputs(4174));
    outputs(4103) <= not(layer0_outputs(4780)) or (layer0_outputs(91));
    outputs(4104) <= layer0_outputs(1556);
    outputs(4105) <= layer0_outputs(5535);
    outputs(4106) <= (layer0_outputs(791)) and (layer0_outputs(8941));
    outputs(4107) <= layer0_outputs(9585);
    outputs(4108) <= not(layer0_outputs(2800)) or (layer0_outputs(2267));
    outputs(4109) <= (layer0_outputs(2581)) and (layer0_outputs(3747));
    outputs(4110) <= layer0_outputs(7377);
    outputs(4111) <= (layer0_outputs(8138)) and not (layer0_outputs(2968));
    outputs(4112) <= not((layer0_outputs(5644)) or (layer0_outputs(8487)));
    outputs(4113) <= not((layer0_outputs(8317)) xor (layer0_outputs(6534)));
    outputs(4114) <= not((layer0_outputs(5321)) xor (layer0_outputs(8115)));
    outputs(4115) <= not(layer0_outputs(6679));
    outputs(4116) <= (layer0_outputs(1830)) xor (layer0_outputs(1443));
    outputs(4117) <= (layer0_outputs(2219)) and not (layer0_outputs(4207));
    outputs(4118) <= not(layer0_outputs(4287));
    outputs(4119) <= layer0_outputs(7019);
    outputs(4120) <= (layer0_outputs(8805)) and not (layer0_outputs(3794));
    outputs(4121) <= not((layer0_outputs(8931)) xor (layer0_outputs(5042)));
    outputs(4122) <= layer0_outputs(5770);
    outputs(4123) <= not(layer0_outputs(5443)) or (layer0_outputs(6417));
    outputs(4124) <= layer0_outputs(4750);
    outputs(4125) <= not(layer0_outputs(393));
    outputs(4126) <= not(layer0_outputs(9598));
    outputs(4127) <= not(layer0_outputs(5155));
    outputs(4128) <= not((layer0_outputs(3854)) and (layer0_outputs(59)));
    outputs(4129) <= layer0_outputs(1351);
    outputs(4130) <= not(layer0_outputs(1748)) or (layer0_outputs(9772));
    outputs(4131) <= layer0_outputs(7385);
    outputs(4132) <= (layer0_outputs(6748)) or (layer0_outputs(3553));
    outputs(4133) <= (layer0_outputs(10162)) xor (layer0_outputs(9892));
    outputs(4134) <= not(layer0_outputs(9376));
    outputs(4135) <= layer0_outputs(2559);
    outputs(4136) <= not(layer0_outputs(2978));
    outputs(4137) <= not(layer0_outputs(4681));
    outputs(4138) <= (layer0_outputs(7373)) and (layer0_outputs(7139));
    outputs(4139) <= layer0_outputs(3003);
    outputs(4140) <= (layer0_outputs(3280)) and not (layer0_outputs(7331));
    outputs(4141) <= (layer0_outputs(4486)) and not (layer0_outputs(4922));
    outputs(4142) <= not((layer0_outputs(10210)) xor (layer0_outputs(1700)));
    outputs(4143) <= not(layer0_outputs(9704)) or (layer0_outputs(4800));
    outputs(4144) <= not(layer0_outputs(726));
    outputs(4145) <= not((layer0_outputs(814)) and (layer0_outputs(10152)));
    outputs(4146) <= layer0_outputs(51);
    outputs(4147) <= (layer0_outputs(1905)) xor (layer0_outputs(3378));
    outputs(4148) <= not((layer0_outputs(7513)) xor (layer0_outputs(10008)));
    outputs(4149) <= (layer0_outputs(6814)) xor (layer0_outputs(8247));
    outputs(4150) <= (layer0_outputs(10036)) xor (layer0_outputs(7079));
    outputs(4151) <= not(layer0_outputs(2298));
    outputs(4152) <= not((layer0_outputs(4876)) and (layer0_outputs(270)));
    outputs(4153) <= (layer0_outputs(9101)) xor (layer0_outputs(5886));
    outputs(4154) <= not((layer0_outputs(7324)) xor (layer0_outputs(7535)));
    outputs(4155) <= layer0_outputs(3485);
    outputs(4156) <= layer0_outputs(5311);
    outputs(4157) <= not(layer0_outputs(9726));
    outputs(4158) <= (layer0_outputs(7937)) and (layer0_outputs(3374));
    outputs(4159) <= not(layer0_outputs(8728));
    outputs(4160) <= (layer0_outputs(5068)) xor (layer0_outputs(226));
    outputs(4161) <= not(layer0_outputs(1993));
    outputs(4162) <= layer0_outputs(6102);
    outputs(4163) <= layer0_outputs(7268);
    outputs(4164) <= not(layer0_outputs(2046));
    outputs(4165) <= (layer0_outputs(495)) or (layer0_outputs(10063));
    outputs(4166) <= not((layer0_outputs(3320)) xor (layer0_outputs(9608)));
    outputs(4167) <= not(layer0_outputs(6839)) or (layer0_outputs(10080));
    outputs(4168) <= (layer0_outputs(5362)) xor (layer0_outputs(1697));
    outputs(4169) <= (layer0_outputs(8527)) and (layer0_outputs(6699));
    outputs(4170) <= (layer0_outputs(2206)) xor (layer0_outputs(8404));
    outputs(4171) <= not(layer0_outputs(7550));
    outputs(4172) <= (layer0_outputs(2407)) xor (layer0_outputs(1158));
    outputs(4173) <= not(layer0_outputs(680));
    outputs(4174) <= layer0_outputs(4193);
    outputs(4175) <= layer0_outputs(9610);
    outputs(4176) <= not((layer0_outputs(2702)) or (layer0_outputs(8627)));
    outputs(4177) <= layer0_outputs(5880);
    outputs(4178) <= layer0_outputs(9372);
    outputs(4179) <= not(layer0_outputs(4680));
    outputs(4180) <= layer0_outputs(2383);
    outputs(4181) <= not((layer0_outputs(4613)) xor (layer0_outputs(1630)));
    outputs(4182) <= (layer0_outputs(5917)) and not (layer0_outputs(1994));
    outputs(4183) <= not(layer0_outputs(2574));
    outputs(4184) <= (layer0_outputs(7736)) and not (layer0_outputs(7188));
    outputs(4185) <= not(layer0_outputs(2371));
    outputs(4186) <= layer0_outputs(255);
    outputs(4187) <= (layer0_outputs(1053)) and (layer0_outputs(5094));
    outputs(4188) <= (layer0_outputs(5883)) xor (layer0_outputs(4514));
    outputs(4189) <= (layer0_outputs(6252)) xor (layer0_outputs(4752));
    outputs(4190) <= layer0_outputs(2795);
    outputs(4191) <= layer0_outputs(2377);
    outputs(4192) <= not(layer0_outputs(9581)) or (layer0_outputs(1377));
    outputs(4193) <= (layer0_outputs(1104)) and (layer0_outputs(7114));
    outputs(4194) <= (layer0_outputs(212)) and not (layer0_outputs(9739));
    outputs(4195) <= (layer0_outputs(3603)) and not (layer0_outputs(1992));
    outputs(4196) <= (layer0_outputs(5851)) xor (layer0_outputs(6492));
    outputs(4197) <= not(layer0_outputs(2381));
    outputs(4198) <= not((layer0_outputs(4108)) xor (layer0_outputs(8181)));
    outputs(4199) <= (layer0_outputs(8731)) xor (layer0_outputs(6203));
    outputs(4200) <= (layer0_outputs(173)) or (layer0_outputs(172));
    outputs(4201) <= not(layer0_outputs(7476));
    outputs(4202) <= (layer0_outputs(241)) and not (layer0_outputs(9093));
    outputs(4203) <= not(layer0_outputs(3018));
    outputs(4204) <= not(layer0_outputs(6637));
    outputs(4205) <= (layer0_outputs(2411)) and not (layer0_outputs(3517));
    outputs(4206) <= not(layer0_outputs(4454));
    outputs(4207) <= not((layer0_outputs(943)) xor (layer0_outputs(10047)));
    outputs(4208) <= (layer0_outputs(1101)) and not (layer0_outputs(5268));
    outputs(4209) <= not(layer0_outputs(175));
    outputs(4210) <= layer0_outputs(654);
    outputs(4211) <= (layer0_outputs(7958)) and not (layer0_outputs(9548));
    outputs(4212) <= (layer0_outputs(7089)) and (layer0_outputs(5315));
    outputs(4213) <= not((layer0_outputs(5236)) and (layer0_outputs(4411)));
    outputs(4214) <= (layer0_outputs(7370)) xor (layer0_outputs(978));
    outputs(4215) <= layer0_outputs(6138);
    outputs(4216) <= (layer0_outputs(7809)) and (layer0_outputs(7530));
    outputs(4217) <= not((layer0_outputs(1126)) xor (layer0_outputs(6006)));
    outputs(4218) <= not(layer0_outputs(8955));
    outputs(4219) <= not(layer0_outputs(1583));
    outputs(4220) <= (layer0_outputs(164)) and not (layer0_outputs(3018));
    outputs(4221) <= not(layer0_outputs(6275));
    outputs(4222) <= not(layer0_outputs(3602));
    outputs(4223) <= layer0_outputs(4940);
    outputs(4224) <= not(layer0_outputs(8565)) or (layer0_outputs(388));
    outputs(4225) <= not(layer0_outputs(2536));
    outputs(4226) <= not(layer0_outputs(7307));
    outputs(4227) <= (layer0_outputs(7747)) xor (layer0_outputs(1631));
    outputs(4228) <= not(layer0_outputs(8266)) or (layer0_outputs(232));
    outputs(4229) <= not(layer0_outputs(3943));
    outputs(4230) <= (layer0_outputs(4536)) xor (layer0_outputs(8879));
    outputs(4231) <= layer0_outputs(698);
    outputs(4232) <= not(layer0_outputs(6771));
    outputs(4233) <= not((layer0_outputs(1982)) or (layer0_outputs(3583)));
    outputs(4234) <= not(layer0_outputs(4268)) or (layer0_outputs(1227));
    outputs(4235) <= layer0_outputs(4894);
    outputs(4236) <= not(layer0_outputs(2448));
    outputs(4237) <= (layer0_outputs(403)) and not (layer0_outputs(5624));
    outputs(4238) <= (layer0_outputs(9145)) and (layer0_outputs(1641));
    outputs(4239) <= (layer0_outputs(3505)) or (layer0_outputs(6290));
    outputs(4240) <= not((layer0_outputs(3727)) xor (layer0_outputs(1402)));
    outputs(4241) <= not((layer0_outputs(8860)) or (layer0_outputs(4945)));
    outputs(4242) <= (layer0_outputs(3905)) xor (layer0_outputs(2866));
    outputs(4243) <= (layer0_outputs(1504)) and not (layer0_outputs(5121));
    outputs(4244) <= not(layer0_outputs(4100));
    outputs(4245) <= not((layer0_outputs(4813)) or (layer0_outputs(801)));
    outputs(4246) <= layer0_outputs(3503);
    outputs(4247) <= not((layer0_outputs(4641)) and (layer0_outputs(8859)));
    outputs(4248) <= not((layer0_outputs(139)) xor (layer0_outputs(6421)));
    outputs(4249) <= layer0_outputs(1316);
    outputs(4250) <= not((layer0_outputs(9110)) and (layer0_outputs(2881)));
    outputs(4251) <= (layer0_outputs(6985)) and not (layer0_outputs(2648));
    outputs(4252) <= (layer0_outputs(2530)) xor (layer0_outputs(6432));
    outputs(4253) <= not((layer0_outputs(7427)) xor (layer0_outputs(8100)));
    outputs(4254) <= not(layer0_outputs(4110));
    outputs(4255) <= layer0_outputs(8445);
    outputs(4256) <= not(layer0_outputs(905));
    outputs(4257) <= not(layer0_outputs(6473)) or (layer0_outputs(4571));
    outputs(4258) <= not(layer0_outputs(8978));
    outputs(4259) <= layer0_outputs(1721);
    outputs(4260) <= (layer0_outputs(3299)) and (layer0_outputs(10109));
    outputs(4261) <= layer0_outputs(2974);
    outputs(4262) <= (layer0_outputs(4082)) or (layer0_outputs(8459));
    outputs(4263) <= layer0_outputs(8391);
    outputs(4264) <= layer0_outputs(7300);
    outputs(4265) <= not(layer0_outputs(6160));
    outputs(4266) <= not((layer0_outputs(2166)) or (layer0_outputs(7092)));
    outputs(4267) <= (layer0_outputs(4760)) and not (layer0_outputs(9970));
    outputs(4268) <= not((layer0_outputs(157)) or (layer0_outputs(9067)));
    outputs(4269) <= not(layer0_outputs(8210));
    outputs(4270) <= not(layer0_outputs(4380)) or (layer0_outputs(8602));
    outputs(4271) <= not((layer0_outputs(1943)) and (layer0_outputs(995)));
    outputs(4272) <= (layer0_outputs(304)) or (layer0_outputs(4859));
    outputs(4273) <= not((layer0_outputs(7587)) xor (layer0_outputs(7719)));
    outputs(4274) <= not((layer0_outputs(8501)) and (layer0_outputs(4963)));
    outputs(4275) <= not(layer0_outputs(2738)) or (layer0_outputs(653));
    outputs(4276) <= (layer0_outputs(6807)) xor (layer0_outputs(2660));
    outputs(4277) <= layer0_outputs(2998);
    outputs(4278) <= not((layer0_outputs(7998)) and (layer0_outputs(7586)));
    outputs(4279) <= layer0_outputs(2146);
    outputs(4280) <= (layer0_outputs(1374)) xor (layer0_outputs(1323));
    outputs(4281) <= not(layer0_outputs(7680));
    outputs(4282) <= not((layer0_outputs(5704)) xor (layer0_outputs(2053)));
    outputs(4283) <= not(layer0_outputs(723));
    outputs(4284) <= not(layer0_outputs(8256));
    outputs(4285) <= not((layer0_outputs(9017)) xor (layer0_outputs(1541)));
    outputs(4286) <= layer0_outputs(5661);
    outputs(4287) <= not(layer0_outputs(1398)) or (layer0_outputs(768));
    outputs(4288) <= not(layer0_outputs(6658));
    outputs(4289) <= layer0_outputs(3988);
    outputs(4290) <= (layer0_outputs(1815)) xor (layer0_outputs(3205));
    outputs(4291) <= layer0_outputs(1519);
    outputs(4292) <= not((layer0_outputs(4644)) xor (layer0_outputs(2984)));
    outputs(4293) <= not(layer0_outputs(5876));
    outputs(4294) <= layer0_outputs(8760);
    outputs(4295) <= (layer0_outputs(5499)) or (layer0_outputs(2806));
    outputs(4296) <= (layer0_outputs(8439)) and (layer0_outputs(3960));
    outputs(4297) <= not(layer0_outputs(1845)) or (layer0_outputs(9337));
    outputs(4298) <= not((layer0_outputs(9562)) xor (layer0_outputs(8250)));
    outputs(4299) <= not(layer0_outputs(9966));
    outputs(4300) <= not(layer0_outputs(6580));
    outputs(4301) <= not(layer0_outputs(6030));
    outputs(4302) <= (layer0_outputs(7170)) and (layer0_outputs(5137));
    outputs(4303) <= layer0_outputs(1222);
    outputs(4304) <= (layer0_outputs(8463)) and (layer0_outputs(9362));
    outputs(4305) <= (layer0_outputs(9575)) or (layer0_outputs(5909));
    outputs(4306) <= not(layer0_outputs(8274));
    outputs(4307) <= not((layer0_outputs(5312)) or (layer0_outputs(8136)));
    outputs(4308) <= not((layer0_outputs(6199)) xor (layer0_outputs(8862)));
    outputs(4309) <= (layer0_outputs(1517)) xor (layer0_outputs(7601));
    outputs(4310) <= (layer0_outputs(3645)) and (layer0_outputs(7067));
    outputs(4311) <= layer0_outputs(1566);
    outputs(4312) <= (layer0_outputs(1386)) xor (layer0_outputs(9130));
    outputs(4313) <= not(layer0_outputs(3693)) or (layer0_outputs(9486));
    outputs(4314) <= not((layer0_outputs(6758)) and (layer0_outputs(4510)));
    outputs(4315) <= not((layer0_outputs(1518)) xor (layer0_outputs(2132)));
    outputs(4316) <= not(layer0_outputs(2008));
    outputs(4317) <= not(layer0_outputs(828));
    outputs(4318) <= (layer0_outputs(4014)) and (layer0_outputs(6267));
    outputs(4319) <= (layer0_outputs(5894)) or (layer0_outputs(192));
    outputs(4320) <= layer0_outputs(7810);
    outputs(4321) <= layer0_outputs(6013);
    outputs(4322) <= (layer0_outputs(1802)) and not (layer0_outputs(5435));
    outputs(4323) <= not(layer0_outputs(6943));
    outputs(4324) <= (layer0_outputs(4572)) or (layer0_outputs(4754));
    outputs(4325) <= layer0_outputs(1142);
    outputs(4326) <= layer0_outputs(2942);
    outputs(4327) <= not((layer0_outputs(1334)) and (layer0_outputs(9991)));
    outputs(4328) <= (layer0_outputs(5336)) and not (layer0_outputs(1765));
    outputs(4329) <= not((layer0_outputs(6301)) xor (layer0_outputs(2848)));
    outputs(4330) <= not(layer0_outputs(9688));
    outputs(4331) <= (layer0_outputs(3694)) and (layer0_outputs(7254));
    outputs(4332) <= (layer0_outputs(7393)) xor (layer0_outputs(4957));
    outputs(4333) <= layer0_outputs(2971);
    outputs(4334) <= (layer0_outputs(5392)) or (layer0_outputs(419));
    outputs(4335) <= (layer0_outputs(4467)) or (layer0_outputs(6159));
    outputs(4336) <= not((layer0_outputs(1615)) xor (layer0_outputs(769)));
    outputs(4337) <= not(layer0_outputs(5845)) or (layer0_outputs(3855));
    outputs(4338) <= (layer0_outputs(9046)) and (layer0_outputs(2825));
    outputs(4339) <= not(layer0_outputs(6710));
    outputs(4340) <= (layer0_outputs(7213)) and (layer0_outputs(1356));
    outputs(4341) <= (layer0_outputs(9637)) and not (layer0_outputs(9590));
    outputs(4342) <= not((layer0_outputs(9166)) or (layer0_outputs(3813)));
    outputs(4343) <= (layer0_outputs(2965)) xor (layer0_outputs(8548));
    outputs(4344) <= not((layer0_outputs(5993)) xor (layer0_outputs(4388)));
    outputs(4345) <= (layer0_outputs(4645)) and (layer0_outputs(4716));
    outputs(4346) <= (layer0_outputs(271)) xor (layer0_outputs(9403));
    outputs(4347) <= layer0_outputs(3125);
    outputs(4348) <= not(layer0_outputs(5842));
    outputs(4349) <= not(layer0_outputs(9025));
    outputs(4350) <= (layer0_outputs(5052)) xor (layer0_outputs(8406));
    outputs(4351) <= (layer0_outputs(3186)) and not (layer0_outputs(3215));
    outputs(4352) <= not(layer0_outputs(4962));
    outputs(4353) <= (layer0_outputs(6048)) xor (layer0_outputs(4602));
    outputs(4354) <= layer0_outputs(1853);
    outputs(4355) <= not((layer0_outputs(303)) and (layer0_outputs(23)));
    outputs(4356) <= (layer0_outputs(8401)) and not (layer0_outputs(1306));
    outputs(4357) <= not((layer0_outputs(4489)) xor (layer0_outputs(9688)));
    outputs(4358) <= not(layer0_outputs(4778)) or (layer0_outputs(206));
    outputs(4359) <= layer0_outputs(1608);
    outputs(4360) <= not(layer0_outputs(6091)) or (layer0_outputs(4859));
    outputs(4361) <= not((layer0_outputs(1737)) xor (layer0_outputs(8281)));
    outputs(4362) <= not(layer0_outputs(5081));
    outputs(4363) <= (layer0_outputs(260)) and not (layer0_outputs(5799));
    outputs(4364) <= layer0_outputs(68);
    outputs(4365) <= (layer0_outputs(8517)) or (layer0_outputs(3318));
    outputs(4366) <= not(layer0_outputs(5465));
    outputs(4367) <= not(layer0_outputs(6294));
    outputs(4368) <= (layer0_outputs(1436)) and (layer0_outputs(3744));
    outputs(4369) <= not(layer0_outputs(719));
    outputs(4370) <= layer0_outputs(4636);
    outputs(4371) <= layer0_outputs(906);
    outputs(4372) <= not(layer0_outputs(183)) or (layer0_outputs(7845));
    outputs(4373) <= not(layer0_outputs(7012));
    outputs(4374) <= not(layer0_outputs(6335));
    outputs(4375) <= (layer0_outputs(2261)) xor (layer0_outputs(2844));
    outputs(4376) <= layer0_outputs(3139);
    outputs(4377) <= not(layer0_outputs(5195)) or (layer0_outputs(4764));
    outputs(4378) <= layer0_outputs(5183);
    outputs(4379) <= (layer0_outputs(7845)) xor (layer0_outputs(2454));
    outputs(4380) <= layer0_outputs(7397);
    outputs(4381) <= layer0_outputs(4331);
    outputs(4382) <= layer0_outputs(6128);
    outputs(4383) <= (layer0_outputs(5901)) and not (layer0_outputs(9576));
    outputs(4384) <= not((layer0_outputs(579)) and (layer0_outputs(5996)));
    outputs(4385) <= layer0_outputs(3293);
    outputs(4386) <= not(layer0_outputs(3708));
    outputs(4387) <= (layer0_outputs(7080)) and not (layer0_outputs(47));
    outputs(4388) <= (layer0_outputs(3114)) and (layer0_outputs(6873));
    outputs(4389) <= not((layer0_outputs(421)) xor (layer0_outputs(830)));
    outputs(4390) <= not((layer0_outputs(6233)) or (layer0_outputs(4661)));
    outputs(4391) <= not((layer0_outputs(9754)) xor (layer0_outputs(4796)));
    outputs(4392) <= not((layer0_outputs(6333)) xor (layer0_outputs(9201)));
    outputs(4393) <= not((layer0_outputs(8418)) xor (layer0_outputs(773)));
    outputs(4394) <= layer0_outputs(4559);
    outputs(4395) <= not((layer0_outputs(580)) xor (layer0_outputs(1521)));
    outputs(4396) <= (layer0_outputs(1667)) and (layer0_outputs(4941));
    outputs(4397) <= (layer0_outputs(8171)) xor (layer0_outputs(2637));
    outputs(4398) <= (layer0_outputs(4095)) and (layer0_outputs(9347));
    outputs(4399) <= not(layer0_outputs(7679));
    outputs(4400) <= (layer0_outputs(6686)) and (layer0_outputs(8631));
    outputs(4401) <= not(layer0_outputs(6196)) or (layer0_outputs(3055));
    outputs(4402) <= not(layer0_outputs(558));
    outputs(4403) <= (layer0_outputs(9349)) xor (layer0_outputs(684));
    outputs(4404) <= not((layer0_outputs(2698)) or (layer0_outputs(152)));
    outputs(4405) <= not(layer0_outputs(7440));
    outputs(4406) <= (layer0_outputs(5005)) and (layer0_outputs(1736));
    outputs(4407) <= not((layer0_outputs(511)) xor (layer0_outputs(5678)));
    outputs(4408) <= (layer0_outputs(5384)) and not (layer0_outputs(6617));
    outputs(4409) <= (layer0_outputs(4257)) and not (layer0_outputs(6251));
    outputs(4410) <= layer0_outputs(4119);
    outputs(4411) <= not(layer0_outputs(5309)) or (layer0_outputs(454));
    outputs(4412) <= (layer0_outputs(2922)) xor (layer0_outputs(4446));
    outputs(4413) <= not(layer0_outputs(5723)) or (layer0_outputs(4157));
    outputs(4414) <= not(layer0_outputs(9041));
    outputs(4415) <= layer0_outputs(3118);
    outputs(4416) <= layer0_outputs(2078);
    outputs(4417) <= layer0_outputs(7837);
    outputs(4418) <= (layer0_outputs(7574)) xor (layer0_outputs(7354));
    outputs(4419) <= (layer0_outputs(10104)) xor (layer0_outputs(4747));
    outputs(4420) <= not(layer0_outputs(8139)) or (layer0_outputs(6792));
    outputs(4421) <= not(layer0_outputs(4366));
    outputs(4422) <= not((layer0_outputs(5716)) and (layer0_outputs(8158)));
    outputs(4423) <= (layer0_outputs(1705)) and not (layer0_outputs(4922));
    outputs(4424) <= not(layer0_outputs(2347));
    outputs(4425) <= '0';
    outputs(4426) <= (layer0_outputs(2936)) and not (layer0_outputs(6436));
    outputs(4427) <= not(layer0_outputs(3689)) or (layer0_outputs(4726));
    outputs(4428) <= not(layer0_outputs(8505)) or (layer0_outputs(7063));
    outputs(4429) <= not(layer0_outputs(3181));
    outputs(4430) <= layer0_outputs(140);
    outputs(4431) <= (layer0_outputs(10125)) xor (layer0_outputs(8579));
    outputs(4432) <= (layer0_outputs(7703)) and not (layer0_outputs(1925));
    outputs(4433) <= layer0_outputs(7124);
    outputs(4434) <= not((layer0_outputs(2700)) or (layer0_outputs(4310)));
    outputs(4435) <= layer0_outputs(2030);
    outputs(4436) <= layer0_outputs(7517);
    outputs(4437) <= not(layer0_outputs(9945));
    outputs(4438) <= not((layer0_outputs(832)) or (layer0_outputs(6976)));
    outputs(4439) <= layer0_outputs(9331);
    outputs(4440) <= not(layer0_outputs(293));
    outputs(4441) <= (layer0_outputs(8777)) xor (layer0_outputs(7185));
    outputs(4442) <= (layer0_outputs(4808)) and (layer0_outputs(4997));
    outputs(4443) <= not((layer0_outputs(5869)) xor (layer0_outputs(2542)));
    outputs(4444) <= (layer0_outputs(391)) xor (layer0_outputs(4117));
    outputs(4445) <= not(layer0_outputs(8006));
    outputs(4446) <= (layer0_outputs(4115)) xor (layer0_outputs(4412));
    outputs(4447) <= not(layer0_outputs(6664));
    outputs(4448) <= (layer0_outputs(8655)) xor (layer0_outputs(2129));
    outputs(4449) <= not((layer0_outputs(8987)) xor (layer0_outputs(4528)));
    outputs(4450) <= not((layer0_outputs(8568)) xor (layer0_outputs(7650)));
    outputs(4451) <= not(layer0_outputs(5273));
    outputs(4452) <= (layer0_outputs(4671)) xor (layer0_outputs(1983));
    outputs(4453) <= not(layer0_outputs(1387));
    outputs(4454) <= not((layer0_outputs(4803)) or (layer0_outputs(32)));
    outputs(4455) <= not(layer0_outputs(6963));
    outputs(4456) <= not((layer0_outputs(605)) xor (layer0_outputs(1138)));
    outputs(4457) <= not(layer0_outputs(3336));
    outputs(4458) <= not((layer0_outputs(4984)) or (layer0_outputs(492)));
    outputs(4459) <= (layer0_outputs(1378)) and not (layer0_outputs(3078));
    outputs(4460) <= layer0_outputs(4910);
    outputs(4461) <= not(layer0_outputs(8198));
    outputs(4462) <= layer0_outputs(802);
    outputs(4463) <= not((layer0_outputs(3304)) xor (layer0_outputs(3377)));
    outputs(4464) <= layer0_outputs(4108);
    outputs(4465) <= layer0_outputs(7194);
    outputs(4466) <= not((layer0_outputs(1406)) xor (layer0_outputs(5844)));
    outputs(4467) <= (layer0_outputs(2862)) xor (layer0_outputs(1258));
    outputs(4468) <= not(layer0_outputs(3821));
    outputs(4469) <= not((layer0_outputs(2017)) and (layer0_outputs(5768)));
    outputs(4470) <= layer0_outputs(6846);
    outputs(4471) <= not((layer0_outputs(2575)) xor (layer0_outputs(4737)));
    outputs(4472) <= layer0_outputs(3389);
    outputs(4473) <= layer0_outputs(3761);
    outputs(4474) <= not((layer0_outputs(9277)) xor (layer0_outputs(8223)));
    outputs(4475) <= not(layer0_outputs(9212));
    outputs(4476) <= (layer0_outputs(710)) and not (layer0_outputs(8605));
    outputs(4477) <= (layer0_outputs(4821)) and (layer0_outputs(8035));
    outputs(4478) <= (layer0_outputs(4724)) and not (layer0_outputs(10008));
    outputs(4479) <= (layer0_outputs(7463)) and (layer0_outputs(4332));
    outputs(4480) <= not((layer0_outputs(6605)) xor (layer0_outputs(7744)));
    outputs(4481) <= layer0_outputs(2475);
    outputs(4482) <= (layer0_outputs(4911)) and (layer0_outputs(285));
    outputs(4483) <= not(layer0_outputs(7818));
    outputs(4484) <= layer0_outputs(1837);
    outputs(4485) <= not(layer0_outputs(6311));
    outputs(4486) <= not((layer0_outputs(3804)) or (layer0_outputs(8195)));
    outputs(4487) <= (layer0_outputs(7111)) and not (layer0_outputs(7258));
    outputs(4488) <= not(layer0_outputs(9763)) or (layer0_outputs(3551));
    outputs(4489) <= not(layer0_outputs(9968));
    outputs(4490) <= (layer0_outputs(627)) or (layer0_outputs(4164));
    outputs(4491) <= not(layer0_outputs(9135));
    outputs(4492) <= (layer0_outputs(7125)) xor (layer0_outputs(6552));
    outputs(4493) <= not(layer0_outputs(799));
    outputs(4494) <= (layer0_outputs(6394)) and not (layer0_outputs(4321));
    outputs(4495) <= (layer0_outputs(5997)) and not (layer0_outputs(941));
    outputs(4496) <= not(layer0_outputs(9660));
    outputs(4497) <= not((layer0_outputs(3522)) xor (layer0_outputs(5961)));
    outputs(4498) <= layer0_outputs(129);
    outputs(4499) <= layer0_outputs(3464);
    outputs(4500) <= (layer0_outputs(6167)) and not (layer0_outputs(7948));
    outputs(4501) <= not(layer0_outputs(3471));
    outputs(4502) <= not((layer0_outputs(8078)) xor (layer0_outputs(7685)));
    outputs(4503) <= (layer0_outputs(4850)) and not (layer0_outputs(5055));
    outputs(4504) <= layer0_outputs(357);
    outputs(4505) <= not(layer0_outputs(6521));
    outputs(4506) <= not((layer0_outputs(536)) xor (layer0_outputs(818)));
    outputs(4507) <= not((layer0_outputs(8470)) or (layer0_outputs(3807)));
    outputs(4508) <= layer0_outputs(5866);
    outputs(4509) <= layer0_outputs(7132);
    outputs(4510) <= layer0_outputs(7580);
    outputs(4511) <= not((layer0_outputs(9341)) or (layer0_outputs(6371)));
    outputs(4512) <= not(layer0_outputs(7382));
    outputs(4513) <= layer0_outputs(2762);
    outputs(4514) <= not(layer0_outputs(3638));
    outputs(4515) <= (layer0_outputs(2760)) and not (layer0_outputs(3218));
    outputs(4516) <= not((layer0_outputs(4360)) xor (layer0_outputs(8089)));
    outputs(4517) <= not(layer0_outputs(6697)) or (layer0_outputs(344));
    outputs(4518) <= not((layer0_outputs(8072)) or (layer0_outputs(2010)));
    outputs(4519) <= not((layer0_outputs(8572)) xor (layer0_outputs(4008)));
    outputs(4520) <= not((layer0_outputs(2527)) xor (layer0_outputs(2348)));
    outputs(4521) <= not((layer0_outputs(3609)) or (layer0_outputs(8983)));
    outputs(4522) <= (layer0_outputs(6296)) and not (layer0_outputs(3706));
    outputs(4523) <= not(layer0_outputs(8859)) or (layer0_outputs(773));
    outputs(4524) <= layer0_outputs(5301);
    outputs(4525) <= (layer0_outputs(1505)) and not (layer0_outputs(1919));
    outputs(4526) <= not(layer0_outputs(5441));
    outputs(4527) <= (layer0_outputs(3954)) xor (layer0_outputs(6370));
    outputs(4528) <= layer0_outputs(300);
    outputs(4529) <= (layer0_outputs(7069)) xor (layer0_outputs(6050));
    outputs(4530) <= not(layer0_outputs(10192));
    outputs(4531) <= (layer0_outputs(6684)) xor (layer0_outputs(1734));
    outputs(4532) <= not((layer0_outputs(10102)) xor (layer0_outputs(7676)));
    outputs(4533) <= layer0_outputs(6072);
    outputs(4534) <= not(layer0_outputs(4178));
    outputs(4535) <= not(layer0_outputs(9686));
    outputs(4536) <= not(layer0_outputs(721)) or (layer0_outputs(8647));
    outputs(4537) <= (layer0_outputs(7961)) and not (layer0_outputs(6466));
    outputs(4538) <= layer0_outputs(9709);
    outputs(4539) <= (layer0_outputs(6010)) and (layer0_outputs(6328));
    outputs(4540) <= not(layer0_outputs(1991));
    outputs(4541) <= not(layer0_outputs(871));
    outputs(4542) <= layer0_outputs(2311);
    outputs(4543) <= not(layer0_outputs(9660));
    outputs(4544) <= not(layer0_outputs(4914));
    outputs(4545) <= (layer0_outputs(3220)) and (layer0_outputs(1753));
    outputs(4546) <= (layer0_outputs(9791)) and (layer0_outputs(3262));
    outputs(4547) <= (layer0_outputs(3364)) xor (layer0_outputs(5874));
    outputs(4548) <= not((layer0_outputs(2152)) and (layer0_outputs(475)));
    outputs(4549) <= (layer0_outputs(6377)) and not (layer0_outputs(9771));
    outputs(4550) <= layer0_outputs(1236);
    outputs(4551) <= (layer0_outputs(9211)) and (layer0_outputs(989));
    outputs(4552) <= not(layer0_outputs(10021));
    outputs(4553) <= (layer0_outputs(4701)) and not (layer0_outputs(155));
    outputs(4554) <= layer0_outputs(5344);
    outputs(4555) <= layer0_outputs(5560);
    outputs(4556) <= (layer0_outputs(1384)) and not (layer0_outputs(10085));
    outputs(4557) <= not((layer0_outputs(4284)) xor (layer0_outputs(1403)));
    outputs(4558) <= not((layer0_outputs(9506)) xor (layer0_outputs(4063)));
    outputs(4559) <= layer0_outputs(4844);
    outputs(4560) <= not(layer0_outputs(4139));
    outputs(4561) <= layer0_outputs(6200);
    outputs(4562) <= not((layer0_outputs(4481)) and (layer0_outputs(3411)));
    outputs(4563) <= not(layer0_outputs(2639));
    outputs(4564) <= not(layer0_outputs(4731));
    outputs(4565) <= layer0_outputs(733);
    outputs(4566) <= (layer0_outputs(7950)) and (layer0_outputs(2308));
    outputs(4567) <= not((layer0_outputs(2228)) xor (layer0_outputs(9018)));
    outputs(4568) <= (layer0_outputs(4354)) xor (layer0_outputs(2168));
    outputs(4569) <= (layer0_outputs(2175)) and (layer0_outputs(4211));
    outputs(4570) <= not(layer0_outputs(4512)) or (layer0_outputs(2539));
    outputs(4571) <= layer0_outputs(701);
    outputs(4572) <= layer0_outputs(4324);
    outputs(4573) <= (layer0_outputs(8947)) and not (layer0_outputs(1404));
    outputs(4574) <= not(layer0_outputs(2934)) or (layer0_outputs(3251));
    outputs(4575) <= not(layer0_outputs(4905));
    outputs(4576) <= (layer0_outputs(4315)) and (layer0_outputs(2770));
    outputs(4577) <= not(layer0_outputs(10));
    outputs(4578) <= not(layer0_outputs(3992));
    outputs(4579) <= layer0_outputs(2798);
    outputs(4580) <= not((layer0_outputs(9614)) and (layer0_outputs(3735)));
    outputs(4581) <= not(layer0_outputs(504)) or (layer0_outputs(3771));
    outputs(4582) <= (layer0_outputs(7434)) or (layer0_outputs(5662));
    outputs(4583) <= not((layer0_outputs(3559)) xor (layer0_outputs(4537)));
    outputs(4584) <= (layer0_outputs(4844)) and not (layer0_outputs(8349));
    outputs(4585) <= (layer0_outputs(405)) xor (layer0_outputs(963));
    outputs(4586) <= not((layer0_outputs(3468)) xor (layer0_outputs(5027)));
    outputs(4587) <= (layer0_outputs(9733)) and not (layer0_outputs(583));
    outputs(4588) <= not(layer0_outputs(632));
    outputs(4589) <= layer0_outputs(3315);
    outputs(4590) <= layer0_outputs(5066);
    outputs(4591) <= (layer0_outputs(9185)) xor (layer0_outputs(3973));
    outputs(4592) <= not(layer0_outputs(4727)) or (layer0_outputs(9711));
    outputs(4593) <= layer0_outputs(6088);
    outputs(4594) <= layer0_outputs(6661);
    outputs(4595) <= not((layer0_outputs(7305)) xor (layer0_outputs(2369)));
    outputs(4596) <= (layer0_outputs(1750)) xor (layer0_outputs(9672));
    outputs(4597) <= not(layer0_outputs(8978));
    outputs(4598) <= (layer0_outputs(6011)) xor (layer0_outputs(1121));
    outputs(4599) <= (layer0_outputs(8688)) and (layer0_outputs(5666));
    outputs(4600) <= not(layer0_outputs(8670)) or (layer0_outputs(3231));
    outputs(4601) <= not(layer0_outputs(6983));
    outputs(4602) <= not(layer0_outputs(2734));
    outputs(4603) <= (layer0_outputs(2003)) xor (layer0_outputs(2251));
    outputs(4604) <= not((layer0_outputs(2386)) xor (layer0_outputs(5074)));
    outputs(4605) <= (layer0_outputs(3026)) xor (layer0_outputs(991));
    outputs(4606) <= (layer0_outputs(220)) xor (layer0_outputs(5532));
    outputs(4607) <= not(layer0_outputs(2767));
    outputs(4608) <= layer0_outputs(6669);
    outputs(4609) <= (layer0_outputs(8550)) and (layer0_outputs(2796));
    outputs(4610) <= (layer0_outputs(193)) and not (layer0_outputs(7570));
    outputs(4611) <= not(layer0_outputs(8662));
    outputs(4612) <= not((layer0_outputs(272)) xor (layer0_outputs(3132)));
    outputs(4613) <= not(layer0_outputs(6831));
    outputs(4614) <= (layer0_outputs(7073)) xor (layer0_outputs(1955));
    outputs(4615) <= layer0_outputs(9048);
    outputs(4616) <= (layer0_outputs(5805)) and not (layer0_outputs(3861));
    outputs(4617) <= layer0_outputs(5857);
    outputs(4618) <= layer0_outputs(3951);
    outputs(4619) <= not((layer0_outputs(5725)) xor (layer0_outputs(8851)));
    outputs(4620) <= (layer0_outputs(9329)) xor (layer0_outputs(5225));
    outputs(4621) <= (layer0_outputs(3824)) xor (layer0_outputs(1835));
    outputs(4622) <= layer0_outputs(2192);
    outputs(4623) <= not((layer0_outputs(5070)) or (layer0_outputs(2193)));
    outputs(4624) <= not((layer0_outputs(397)) xor (layer0_outputs(3306)));
    outputs(4625) <= not(layer0_outputs(5630));
    outputs(4626) <= layer0_outputs(1673);
    outputs(4627) <= not(layer0_outputs(6066)) or (layer0_outputs(6586));
    outputs(4628) <= not((layer0_outputs(3054)) xor (layer0_outputs(2693)));
    outputs(4629) <= (layer0_outputs(5177)) xor (layer0_outputs(6435));
    outputs(4630) <= (layer0_outputs(1587)) and not (layer0_outputs(7499));
    outputs(4631) <= not((layer0_outputs(2253)) xor (layer0_outputs(438)));
    outputs(4632) <= not((layer0_outputs(2930)) or (layer0_outputs(4129)));
    outputs(4633) <= not(layer0_outputs(9936));
    outputs(4634) <= (layer0_outputs(2553)) xor (layer0_outputs(750));
    outputs(4635) <= layer0_outputs(9508);
    outputs(4636) <= layer0_outputs(5335);
    outputs(4637) <= not(layer0_outputs(3803));
    outputs(4638) <= layer0_outputs(1480);
    outputs(4639) <= layer0_outputs(4281);
    outputs(4640) <= layer0_outputs(9647);
    outputs(4641) <= not((layer0_outputs(7351)) or (layer0_outputs(6524)));
    outputs(4642) <= not(layer0_outputs(7426)) or (layer0_outputs(9276));
    outputs(4643) <= (layer0_outputs(9785)) xor (layer0_outputs(3573));
    outputs(4644) <= (layer0_outputs(6766)) xor (layer0_outputs(1429));
    outputs(4645) <= (layer0_outputs(382)) and not (layer0_outputs(8754));
    outputs(4646) <= not(layer0_outputs(8480));
    outputs(4647) <= not((layer0_outputs(6086)) xor (layer0_outputs(9352)));
    outputs(4648) <= not(layer0_outputs(496));
    outputs(4649) <= (layer0_outputs(7713)) xor (layer0_outputs(9497));
    outputs(4650) <= (layer0_outputs(5378)) and (layer0_outputs(1663));
    outputs(4651) <= layer0_outputs(6942);
    outputs(4652) <= (layer0_outputs(2160)) and not (layer0_outputs(5796));
    outputs(4653) <= not((layer0_outputs(4993)) or (layer0_outputs(10222)));
    outputs(4654) <= not((layer0_outputs(895)) xor (layer0_outputs(7224)));
    outputs(4655) <= layer0_outputs(2749);
    outputs(4656) <= not(layer0_outputs(3836)) or (layer0_outputs(7795));
    outputs(4657) <= not(layer0_outputs(4426));
    outputs(4658) <= (layer0_outputs(2310)) xor (layer0_outputs(1977));
    outputs(4659) <= layer0_outputs(5263);
    outputs(4660) <= (layer0_outputs(7434)) and not (layer0_outputs(9483));
    outputs(4661) <= (layer0_outputs(7534)) or (layer0_outputs(6049));
    outputs(4662) <= layer0_outputs(9027);
    outputs(4663) <= (layer0_outputs(6706)) or (layer0_outputs(1778));
    outputs(4664) <= (layer0_outputs(6806)) and not (layer0_outputs(888));
    outputs(4665) <= (layer0_outputs(1817)) and not (layer0_outputs(7460));
    outputs(4666) <= (layer0_outputs(9533)) xor (layer0_outputs(7770));
    outputs(4667) <= layer0_outputs(6034);
    outputs(4668) <= not(layer0_outputs(5029));
    outputs(4669) <= not((layer0_outputs(4593)) or (layer0_outputs(5675)));
    outputs(4670) <= not(layer0_outputs(1368));
    outputs(4671) <= not(layer0_outputs(5032));
    outputs(4672) <= (layer0_outputs(2446)) and not (layer0_outputs(1192));
    outputs(4673) <= not((layer0_outputs(1511)) xor (layer0_outputs(2705)));
    outputs(4674) <= (layer0_outputs(2954)) xor (layer0_outputs(1058));
    outputs(4675) <= not(layer0_outputs(9527));
    outputs(4676) <= layer0_outputs(2180);
    outputs(4677) <= layer0_outputs(8656);
    outputs(4678) <= not(layer0_outputs(8333));
    outputs(4679) <= (layer0_outputs(6828)) and not (layer0_outputs(10158));
    outputs(4680) <= (layer0_outputs(6893)) xor (layer0_outputs(7378));
    outputs(4681) <= layer0_outputs(1873);
    outputs(4682) <= layer0_outputs(735);
    outputs(4683) <= layer0_outputs(6010);
    outputs(4684) <= not(layer0_outputs(9351));
    outputs(4685) <= layer0_outputs(7795);
    outputs(4686) <= layer0_outputs(1134);
    outputs(4687) <= not(layer0_outputs(4959)) or (layer0_outputs(4674));
    outputs(4688) <= not(layer0_outputs(7840));
    outputs(4689) <= layer0_outputs(5365);
    outputs(4690) <= not((layer0_outputs(5303)) xor (layer0_outputs(5779)));
    outputs(4691) <= layer0_outputs(3074);
    outputs(4692) <= not(layer0_outputs(1148));
    outputs(4693) <= (layer0_outputs(5417)) or (layer0_outputs(8042));
    outputs(4694) <= not(layer0_outputs(4672));
    outputs(4695) <= not(layer0_outputs(8359));
    outputs(4696) <= not((layer0_outputs(5254)) xor (layer0_outputs(9635)));
    outputs(4697) <= not(layer0_outputs(6224));
    outputs(4698) <= (layer0_outputs(5060)) and not (layer0_outputs(5279));
    outputs(4699) <= not((layer0_outputs(4383)) xor (layer0_outputs(1015)));
    outputs(4700) <= layer0_outputs(7066);
    outputs(4701) <= (layer0_outputs(29)) xor (layer0_outputs(10206));
    outputs(4702) <= (layer0_outputs(963)) or (layer0_outputs(9839));
    outputs(4703) <= not((layer0_outputs(8024)) xor (layer0_outputs(7683)));
    outputs(4704) <= not(layer0_outputs(10059));
    outputs(4705) <= (layer0_outputs(6791)) xor (layer0_outputs(4852));
    outputs(4706) <= (layer0_outputs(5506)) xor (layer0_outputs(951));
    outputs(4707) <= not((layer0_outputs(8719)) xor (layer0_outputs(1947)));
    outputs(4708) <= not(layer0_outputs(2839));
    outputs(4709) <= not((layer0_outputs(3834)) xor (layer0_outputs(753)));
    outputs(4710) <= (layer0_outputs(3722)) and not (layer0_outputs(10013));
    outputs(4711) <= (layer0_outputs(3588)) xor (layer0_outputs(6354));
    outputs(4712) <= not((layer0_outputs(8910)) xor (layer0_outputs(7715)));
    outputs(4713) <= not(layer0_outputs(3230));
    outputs(4714) <= (layer0_outputs(7508)) and not (layer0_outputs(8582));
    outputs(4715) <= not((layer0_outputs(6502)) xor (layer0_outputs(951)));
    outputs(4716) <= (layer0_outputs(6539)) xor (layer0_outputs(2016));
    outputs(4717) <= not(layer0_outputs(9706));
    outputs(4718) <= layer0_outputs(2493);
    outputs(4719) <= not((layer0_outputs(6480)) or (layer0_outputs(812)));
    outputs(4720) <= not((layer0_outputs(9466)) xor (layer0_outputs(7243)));
    outputs(4721) <= not((layer0_outputs(4072)) or (layer0_outputs(2028)));
    outputs(4722) <= not((layer0_outputs(683)) or (layer0_outputs(4100)));
    outputs(4723) <= not((layer0_outputs(3008)) xor (layer0_outputs(10093)));
    outputs(4724) <= layer0_outputs(4048);
    outputs(4725) <= not(layer0_outputs(3956));
    outputs(4726) <= (layer0_outputs(4375)) or (layer0_outputs(4447));
    outputs(4727) <= not(layer0_outputs(3935));
    outputs(4728) <= layer0_outputs(9241);
    outputs(4729) <= layer0_outputs(5105);
    outputs(4730) <= (layer0_outputs(7751)) and not (layer0_outputs(1612));
    outputs(4731) <= (layer0_outputs(8773)) xor (layer0_outputs(9013));
    outputs(4732) <= (layer0_outputs(7578)) and (layer0_outputs(3870));
    outputs(4733) <= (layer0_outputs(4569)) xor (layer0_outputs(4047));
    outputs(4734) <= (layer0_outputs(3946)) and not (layer0_outputs(5799));
    outputs(4735) <= not(layer0_outputs(2523));
    outputs(4736) <= not(layer0_outputs(7843));
    outputs(4737) <= (layer0_outputs(5009)) xor (layer0_outputs(5443));
    outputs(4738) <= layer0_outputs(9782);
    outputs(4739) <= layer0_outputs(5490);
    outputs(4740) <= (layer0_outputs(9492)) or (layer0_outputs(6586));
    outputs(4741) <= (layer0_outputs(6328)) and (layer0_outputs(6378));
    outputs(4742) <= (layer0_outputs(7905)) xor (layer0_outputs(7640));
    outputs(4743) <= not((layer0_outputs(8419)) or (layer0_outputs(2980)));
    outputs(4744) <= not(layer0_outputs(1111));
    outputs(4745) <= not(layer0_outputs(10151));
    outputs(4746) <= not(layer0_outputs(4127));
    outputs(4747) <= not(layer0_outputs(8775)) or (layer0_outputs(2955));
    outputs(4748) <= not(layer0_outputs(2517));
    outputs(4749) <= not((layer0_outputs(3022)) or (layer0_outputs(6809)));
    outputs(4750) <= (layer0_outputs(9268)) xor (layer0_outputs(1330));
    outputs(4751) <= (layer0_outputs(10205)) xor (layer0_outputs(1579));
    outputs(4752) <= (layer0_outputs(5167)) and not (layer0_outputs(6273));
    outputs(4753) <= not((layer0_outputs(780)) xor (layer0_outputs(8618)));
    outputs(4754) <= layer0_outputs(5820);
    outputs(4755) <= (layer0_outputs(260)) and (layer0_outputs(505));
    outputs(4756) <= (layer0_outputs(4985)) and not (layer0_outputs(1023));
    outputs(4757) <= not((layer0_outputs(6379)) and (layer0_outputs(4395)));
    outputs(4758) <= (layer0_outputs(8341)) xor (layer0_outputs(1850));
    outputs(4759) <= not((layer0_outputs(4339)) xor (layer0_outputs(1254)));
    outputs(4760) <= not((layer0_outputs(7758)) or (layer0_outputs(3827)));
    outputs(4761) <= (layer0_outputs(6909)) and not (layer0_outputs(8325));
    outputs(4762) <= (layer0_outputs(634)) xor (layer0_outputs(2598));
    outputs(4763) <= layer0_outputs(3647);
    outputs(4764) <= layer0_outputs(8313);
    outputs(4765) <= layer0_outputs(40);
    outputs(4766) <= not(layer0_outputs(2506));
    outputs(4767) <= (layer0_outputs(3842)) and not (layer0_outputs(8765));
    outputs(4768) <= not(layer0_outputs(7929));
    outputs(4769) <= not(layer0_outputs(911));
    outputs(4770) <= layer0_outputs(1936);
    outputs(4771) <= not(layer0_outputs(3355));
    outputs(4772) <= layer0_outputs(8282);
    outputs(4773) <= layer0_outputs(8012);
    outputs(4774) <= not(layer0_outputs(8002)) or (layer0_outputs(5673));
    outputs(4775) <= not(layer0_outputs(4125));
    outputs(4776) <= not(layer0_outputs(1967)) or (layer0_outputs(2066));
    outputs(4777) <= (layer0_outputs(3635)) xor (layer0_outputs(6754));
    outputs(4778) <= not(layer0_outputs(5905));
    outputs(4779) <= layer0_outputs(6643);
    outputs(4780) <= not(layer0_outputs(4143));
    outputs(4781) <= not(layer0_outputs(8083));
    outputs(4782) <= not(layer0_outputs(2576));
    outputs(4783) <= not(layer0_outputs(37)) or (layer0_outputs(1449));
    outputs(4784) <= layer0_outputs(1585);
    outputs(4785) <= layer0_outputs(63);
    outputs(4786) <= (layer0_outputs(2088)) and not (layer0_outputs(5640));
    outputs(4787) <= layer0_outputs(2951);
    outputs(4788) <= not(layer0_outputs(9795));
    outputs(4789) <= not(layer0_outputs(9391)) or (layer0_outputs(8468));
    outputs(4790) <= (layer0_outputs(6176)) or (layer0_outputs(6908));
    outputs(4791) <= layer0_outputs(2887);
    outputs(4792) <= not(layer0_outputs(5065));
    outputs(4793) <= layer0_outputs(3681);
    outputs(4794) <= layer0_outputs(5774);
    outputs(4795) <= not(layer0_outputs(2572));
    outputs(4796) <= not(layer0_outputs(8624)) or (layer0_outputs(8898));
    outputs(4797) <= not(layer0_outputs(1376));
    outputs(4798) <= not(layer0_outputs(2279));
    outputs(4799) <= (layer0_outputs(6166)) and not (layer0_outputs(3807));
    outputs(4800) <= not(layer0_outputs(6946));
    outputs(4801) <= (layer0_outputs(9947)) and not (layer0_outputs(9917));
    outputs(4802) <= not((layer0_outputs(7486)) or (layer0_outputs(5117)));
    outputs(4803) <= layer0_outputs(1209);
    outputs(4804) <= (layer0_outputs(2417)) xor (layer0_outputs(6120));
    outputs(4805) <= not((layer0_outputs(840)) xor (layer0_outputs(3972)));
    outputs(4806) <= not(layer0_outputs(5330));
    outputs(4807) <= (layer0_outputs(2260)) xor (layer0_outputs(8014));
    outputs(4808) <= layer0_outputs(1952);
    outputs(4809) <= not((layer0_outputs(1863)) xor (layer0_outputs(2163)));
    outputs(4810) <= (layer0_outputs(5062)) and (layer0_outputs(8793));
    outputs(4811) <= (layer0_outputs(7288)) xor (layer0_outputs(9197));
    outputs(4812) <= not(layer0_outputs(9478)) or (layer0_outputs(4994));
    outputs(4813) <= not(layer0_outputs(3811));
    outputs(4814) <= not((layer0_outputs(7228)) or (layer0_outputs(2310)));
    outputs(4815) <= layer0_outputs(5841);
    outputs(4816) <= not((layer0_outputs(9145)) xor (layer0_outputs(874)));
    outputs(4817) <= not((layer0_outputs(5930)) xor (layer0_outputs(1950)));
    outputs(4818) <= not(layer0_outputs(3623));
    outputs(4819) <= layer0_outputs(1744);
    outputs(4820) <= (layer0_outputs(6046)) or (layer0_outputs(3586));
    outputs(4821) <= not((layer0_outputs(220)) xor (layer0_outputs(2252)));
    outputs(4822) <= not(layer0_outputs(2999));
    outputs(4823) <= not((layer0_outputs(7078)) xor (layer0_outputs(8079)));
    outputs(4824) <= (layer0_outputs(7624)) and (layer0_outputs(8827));
    outputs(4825) <= (layer0_outputs(5229)) and (layer0_outputs(9915));
    outputs(4826) <= not(layer0_outputs(6056));
    outputs(4827) <= not(layer0_outputs(6444));
    outputs(4828) <= not(layer0_outputs(2826));
    outputs(4829) <= (layer0_outputs(8109)) xor (layer0_outputs(5311));
    outputs(4830) <= not((layer0_outputs(2361)) xor (layer0_outputs(8723)));
    outputs(4831) <= not(layer0_outputs(1794));
    outputs(4832) <= not(layer0_outputs(8457));
    outputs(4833) <= layer0_outputs(10018);
    outputs(4834) <= not((layer0_outputs(9990)) xor (layer0_outputs(6840)));
    outputs(4835) <= not((layer0_outputs(335)) xor (layer0_outputs(5246)));
    outputs(4836) <= layer0_outputs(10179);
    outputs(4837) <= not(layer0_outputs(3473));
    outputs(4838) <= (layer0_outputs(9158)) xor (layer0_outputs(3170));
    outputs(4839) <= layer0_outputs(3574);
    outputs(4840) <= not((layer0_outputs(8708)) or (layer0_outputs(7652)));
    outputs(4841) <= layer0_outputs(2719);
    outputs(4842) <= (layer0_outputs(3303)) and not (layer0_outputs(9417));
    outputs(4843) <= layer0_outputs(705);
    outputs(4844) <= (layer0_outputs(89)) xor (layer0_outputs(6779));
    outputs(4845) <= not(layer0_outputs(6953));
    outputs(4846) <= (layer0_outputs(5777)) and not (layer0_outputs(4402));
    outputs(4847) <= (layer0_outputs(9577)) xor (layer0_outputs(2380));
    outputs(4848) <= not(layer0_outputs(8318));
    outputs(4849) <= not(layer0_outputs(4712));
    outputs(4850) <= layer0_outputs(7942);
    outputs(4851) <= (layer0_outputs(5574)) xor (layer0_outputs(1829));
    outputs(4852) <= (layer0_outputs(7291)) xor (layer0_outputs(71));
    outputs(4853) <= (layer0_outputs(4817)) and (layer0_outputs(993));
    outputs(4854) <= (layer0_outputs(221)) xor (layer0_outputs(2002));
    outputs(4855) <= (layer0_outputs(1546)) or (layer0_outputs(10118));
    outputs(4856) <= (layer0_outputs(1259)) and not (layer0_outputs(7741));
    outputs(4857) <= (layer0_outputs(6796)) xor (layer0_outputs(5652));
    outputs(4858) <= not(layer0_outputs(2319));
    outputs(4859) <= not((layer0_outputs(2055)) or (layer0_outputs(7758)));
    outputs(4860) <= not(layer0_outputs(1344));
    outputs(4861) <= (layer0_outputs(3149)) and (layer0_outputs(6936));
    outputs(4862) <= not(layer0_outputs(8714));
    outputs(4863) <= (layer0_outputs(3504)) xor (layer0_outputs(6032));
    outputs(4864) <= layer0_outputs(5508);
    outputs(4865) <= not((layer0_outputs(3489)) and (layer0_outputs(7368)));
    outputs(4866) <= not(layer0_outputs(2963)) or (layer0_outputs(5994));
    outputs(4867) <= layer0_outputs(9384);
    outputs(4868) <= not((layer0_outputs(8360)) xor (layer0_outputs(2897)));
    outputs(4869) <= not((layer0_outputs(9891)) xor (layer0_outputs(616)));
    outputs(4870) <= not((layer0_outputs(3324)) xor (layer0_outputs(2068)));
    outputs(4871) <= layer0_outputs(1043);
    outputs(4872) <= (layer0_outputs(1690)) or (layer0_outputs(5491));
    outputs(4873) <= (layer0_outputs(9419)) xor (layer0_outputs(5432));
    outputs(4874) <= not(layer0_outputs(4177));
    outputs(4875) <= (layer0_outputs(386)) and not (layer0_outputs(1208));
    outputs(4876) <= (layer0_outputs(4807)) and (layer0_outputs(1938));
    outputs(4877) <= not(layer0_outputs(1072)) or (layer0_outputs(4573));
    outputs(4878) <= layer0_outputs(411);
    outputs(4879) <= (layer0_outputs(9382)) and (layer0_outputs(8885));
    outputs(4880) <= not((layer0_outputs(8340)) and (layer0_outputs(6201)));
    outputs(4881) <= not(layer0_outputs(6888)) or (layer0_outputs(7238));
    outputs(4882) <= not((layer0_outputs(1555)) xor (layer0_outputs(6268)));
    outputs(4883) <= not(layer0_outputs(3095));
    outputs(4884) <= layer0_outputs(6548);
    outputs(4885) <= (layer0_outputs(6550)) xor (layer0_outputs(3894));
    outputs(4886) <= (layer0_outputs(5495)) and not (layer0_outputs(9951));
    outputs(4887) <= (layer0_outputs(5258)) xor (layer0_outputs(6296));
    outputs(4888) <= layer0_outputs(2941);
    outputs(4889) <= layer0_outputs(3980);
    outputs(4890) <= not((layer0_outputs(8917)) and (layer0_outputs(8243)));
    outputs(4891) <= (layer0_outputs(2477)) and not (layer0_outputs(5837));
    outputs(4892) <= not((layer0_outputs(5141)) xor (layer0_outputs(5066)));
    outputs(4893) <= (layer0_outputs(1191)) and (layer0_outputs(5462));
    outputs(4894) <= (layer0_outputs(3261)) and (layer0_outputs(5022));
    outputs(4895) <= layer0_outputs(5389);
    outputs(4896) <= (layer0_outputs(6344)) and (layer0_outputs(9493));
    outputs(4897) <= (layer0_outputs(3159)) and (layer0_outputs(6108));
    outputs(4898) <= layer0_outputs(1066);
    outputs(4899) <= not((layer0_outputs(9416)) xor (layer0_outputs(3829)));
    outputs(4900) <= not(layer0_outputs(7193)) or (layer0_outputs(8908));
    outputs(4901) <= not((layer0_outputs(9648)) and (layer0_outputs(6799)));
    outputs(4902) <= layer0_outputs(6083);
    outputs(4903) <= layer0_outputs(9809);
    outputs(4904) <= (layer0_outputs(3882)) and not (layer0_outputs(5524));
    outputs(4905) <= layer0_outputs(1489);
    outputs(4906) <= layer0_outputs(3847);
    outputs(4907) <= not((layer0_outputs(6149)) or (layer0_outputs(5426)));
    outputs(4908) <= not((layer0_outputs(9691)) xor (layer0_outputs(6149)));
    outputs(4909) <= not((layer0_outputs(8604)) xor (layer0_outputs(4387)));
    outputs(4910) <= layer0_outputs(2022);
    outputs(4911) <= not(layer0_outputs(4505));
    outputs(4912) <= not(layer0_outputs(5764));
    outputs(4913) <= not(layer0_outputs(2200));
    outputs(4914) <= not(layer0_outputs(3110));
    outputs(4915) <= (layer0_outputs(9463)) xor (layer0_outputs(4625));
    outputs(4916) <= (layer0_outputs(5006)) xor (layer0_outputs(2211));
    outputs(4917) <= not(layer0_outputs(3965));
    outputs(4918) <= (layer0_outputs(1998)) and not (layer0_outputs(7611));
    outputs(4919) <= not(layer0_outputs(5731));
    outputs(4920) <= not(layer0_outputs(2654));
    outputs(4921) <= not(layer0_outputs(8929));
    outputs(4922) <= (layer0_outputs(7436)) and not (layer0_outputs(3638));
    outputs(4923) <= layer0_outputs(10177);
    outputs(4924) <= layer0_outputs(7734);
    outputs(4925) <= layer0_outputs(10005);
    outputs(4926) <= (layer0_outputs(6911)) and not (layer0_outputs(5822));
    outputs(4927) <= not((layer0_outputs(8257)) or (layer0_outputs(2004)));
    outputs(4928) <= not(layer0_outputs(835));
    outputs(4929) <= (layer0_outputs(8464)) and not (layer0_outputs(229));
    outputs(4930) <= not(layer0_outputs(8610));
    outputs(4931) <= (layer0_outputs(1095)) xor (layer0_outputs(1645));
    outputs(4932) <= layer0_outputs(2174);
    outputs(4933) <= (layer0_outputs(3488)) xor (layer0_outputs(7871));
    outputs(4934) <= not(layer0_outputs(10047)) or (layer0_outputs(9405));
    outputs(4935) <= not((layer0_outputs(6727)) and (layer0_outputs(1931)));
    outputs(4936) <= layer0_outputs(9377);
    outputs(4937) <= not(layer0_outputs(2558)) or (layer0_outputs(6756));
    outputs(4938) <= not(layer0_outputs(6351));
    outputs(4939) <= not((layer0_outputs(6522)) or (layer0_outputs(2698)));
    outputs(4940) <= not(layer0_outputs(1947));
    outputs(4941) <= not((layer0_outputs(3830)) xor (layer0_outputs(1165)));
    outputs(4942) <= (layer0_outputs(2214)) xor (layer0_outputs(5629));
    outputs(4943) <= (layer0_outputs(5385)) and not (layer0_outputs(8954));
    outputs(4944) <= layer0_outputs(7279);
    outputs(4945) <= (layer0_outputs(3665)) and (layer0_outputs(8227));
    outputs(4946) <= (layer0_outputs(2861)) xor (layer0_outputs(4006));
    outputs(4947) <= not(layer0_outputs(314));
    outputs(4948) <= not(layer0_outputs(2594));
    outputs(4949) <= not(layer0_outputs(1407));
    outputs(4950) <= not(layer0_outputs(161));
    outputs(4951) <= not(layer0_outputs(4456));
    outputs(4952) <= not((layer0_outputs(4466)) xor (layer0_outputs(7498)));
    outputs(4953) <= not(layer0_outputs(9342));
    outputs(4954) <= (layer0_outputs(3634)) or (layer0_outputs(4328));
    outputs(4955) <= (layer0_outputs(2431)) and not (layer0_outputs(1521));
    outputs(4956) <= not(layer0_outputs(1825)) or (layer0_outputs(607));
    outputs(4957) <= layer0_outputs(2117);
    outputs(4958) <= (layer0_outputs(3102)) xor (layer0_outputs(9088));
    outputs(4959) <= (layer0_outputs(4675)) and not (layer0_outputs(6702));
    outputs(4960) <= (layer0_outputs(2554)) and (layer0_outputs(8437));
    outputs(4961) <= not(layer0_outputs(141));
    outputs(4962) <= not((layer0_outputs(9666)) xor (layer0_outputs(3740)));
    outputs(4963) <= (layer0_outputs(7673)) and (layer0_outputs(4788));
    outputs(4964) <= layer0_outputs(4978);
    outputs(4965) <= not((layer0_outputs(2757)) xor (layer0_outputs(1855)));
    outputs(4966) <= not((layer0_outputs(751)) or (layer0_outputs(308)));
    outputs(4967) <= not((layer0_outputs(3502)) xor (layer0_outputs(7667)));
    outputs(4968) <= layer0_outputs(4925);
    outputs(4969) <= (layer0_outputs(6472)) xor (layer0_outputs(7616));
    outputs(4970) <= layer0_outputs(10103);
    outputs(4971) <= not(layer0_outputs(274));
    outputs(4972) <= not((layer0_outputs(6781)) xor (layer0_outputs(6217)));
    outputs(4973) <= not(layer0_outputs(1542));
    outputs(4974) <= not((layer0_outputs(6796)) or (layer0_outputs(9008)));
    outputs(4975) <= not((layer0_outputs(3963)) xor (layer0_outputs(2612)));
    outputs(4976) <= (layer0_outputs(5474)) and (layer0_outputs(3752));
    outputs(4977) <= (layer0_outputs(4853)) xor (layer0_outputs(1544));
    outputs(4978) <= (layer0_outputs(460)) and not (layer0_outputs(6292));
    outputs(4979) <= (layer0_outputs(4168)) xor (layer0_outputs(922));
    outputs(4980) <= not((layer0_outputs(253)) xor (layer0_outputs(5031)));
    outputs(4981) <= (layer0_outputs(4684)) xor (layer0_outputs(858));
    outputs(4982) <= (layer0_outputs(5338)) and not (layer0_outputs(8180));
    outputs(4983) <= (layer0_outputs(6636)) and not (layer0_outputs(9689));
    outputs(4984) <= not(layer0_outputs(8300));
    outputs(4985) <= (layer0_outputs(10207)) and (layer0_outputs(14));
    outputs(4986) <= (layer0_outputs(3686)) and not (layer0_outputs(4123));
    outputs(4987) <= (layer0_outputs(7375)) xor (layer0_outputs(251));
    outputs(4988) <= not((layer0_outputs(9286)) or (layer0_outputs(27)));
    outputs(4989) <= not((layer0_outputs(1015)) xor (layer0_outputs(6838)));
    outputs(4990) <= layer0_outputs(9205);
    outputs(4991) <= not(layer0_outputs(4658));
    outputs(4992) <= (layer0_outputs(2290)) and not (layer0_outputs(7627));
    outputs(4993) <= layer0_outputs(5007);
    outputs(4994) <= not((layer0_outputs(8645)) xor (layer0_outputs(7438)));
    outputs(4995) <= layer0_outputs(10096);
    outputs(4996) <= not(layer0_outputs(5639));
    outputs(4997) <= not(layer0_outputs(9680));
    outputs(4998) <= (layer0_outputs(5993)) xor (layer0_outputs(740));
    outputs(4999) <= not((layer0_outputs(1701)) xor (layer0_outputs(1196)));
    outputs(5000) <= layer0_outputs(9132);
    outputs(5001) <= (layer0_outputs(0)) xor (layer0_outputs(4161));
    outputs(5002) <= (layer0_outputs(8821)) and not (layer0_outputs(8719));
    outputs(5003) <= not((layer0_outputs(9390)) xor (layer0_outputs(7648)));
    outputs(5004) <= (layer0_outputs(6151)) xor (layer0_outputs(9679));
    outputs(5005) <= not((layer0_outputs(3497)) xor (layer0_outputs(1898)));
    outputs(5006) <= layer0_outputs(6438);
    outputs(5007) <= not((layer0_outputs(4791)) xor (layer0_outputs(947)));
    outputs(5008) <= layer0_outputs(9674);
    outputs(5009) <= (layer0_outputs(4868)) and not (layer0_outputs(7097));
    outputs(5010) <= layer0_outputs(9654);
    outputs(5011) <= (layer0_outputs(7979)) and (layer0_outputs(3810));
    outputs(5012) <= not(layer0_outputs(9448));
    outputs(5013) <= (layer0_outputs(9544)) xor (layer0_outputs(8466));
    outputs(5014) <= (layer0_outputs(6598)) and (layer0_outputs(7442));
    outputs(5015) <= (layer0_outputs(6824)) and not (layer0_outputs(8592));
    outputs(5016) <= not((layer0_outputs(3496)) xor (layer0_outputs(2022)));
    outputs(5017) <= (layer0_outputs(9282)) and not (layer0_outputs(10003));
    outputs(5018) <= layer0_outputs(8441);
    outputs(5019) <= not((layer0_outputs(7314)) xor (layer0_outputs(8537)));
    outputs(5020) <= layer0_outputs(1893);
    outputs(5021) <= not((layer0_outputs(9034)) or (layer0_outputs(1093)));
    outputs(5022) <= not(layer0_outputs(3832));
    outputs(5023) <= not(layer0_outputs(2562));
    outputs(5024) <= (layer0_outputs(4214)) and (layer0_outputs(2541));
    outputs(5025) <= (layer0_outputs(2326)) and not (layer0_outputs(6619));
    outputs(5026) <= (layer0_outputs(2051)) xor (layer0_outputs(6191));
    outputs(5027) <= not(layer0_outputs(5509));
    outputs(5028) <= not(layer0_outputs(2231));
    outputs(5029) <= layer0_outputs(5724);
    outputs(5030) <= layer0_outputs(6277);
    outputs(5031) <= not((layer0_outputs(584)) or (layer0_outputs(3798)));
    outputs(5032) <= not((layer0_outputs(3960)) xor (layer0_outputs(10036)));
    outputs(5033) <= (layer0_outputs(7016)) and not (layer0_outputs(7288));
    outputs(5034) <= not(layer0_outputs(8876)) or (layer0_outputs(1727));
    outputs(5035) <= not(layer0_outputs(7094)) or (layer0_outputs(725));
    outputs(5036) <= not(layer0_outputs(2067));
    outputs(5037) <= (layer0_outputs(9537)) or (layer0_outputs(10188));
    outputs(5038) <= layer0_outputs(8319);
    outputs(5039) <= not(layer0_outputs(9510));
    outputs(5040) <= not((layer0_outputs(7739)) xor (layer0_outputs(4566)));
    outputs(5041) <= not(layer0_outputs(1518));
    outputs(5042) <= layer0_outputs(598);
    outputs(5043) <= layer0_outputs(4610);
    outputs(5044) <= layer0_outputs(1732);
    outputs(5045) <= layer0_outputs(5567);
    outputs(5046) <= (layer0_outputs(9651)) and not (layer0_outputs(6186));
    outputs(5047) <= not(layer0_outputs(1163));
    outputs(5048) <= not((layer0_outputs(5154)) xor (layer0_outputs(9392)));
    outputs(5049) <= not((layer0_outputs(6570)) or (layer0_outputs(686)));
    outputs(5050) <= not((layer0_outputs(8229)) xor (layer0_outputs(124)));
    outputs(5051) <= (layer0_outputs(6804)) and (layer0_outputs(4580));
    outputs(5052) <= not((layer0_outputs(8396)) xor (layer0_outputs(771)));
    outputs(5053) <= (layer0_outputs(6955)) and (layer0_outputs(5920));
    outputs(5054) <= not(layer0_outputs(3016)) or (layer0_outputs(7821));
    outputs(5055) <= not(layer0_outputs(3863)) or (layer0_outputs(2397));
    outputs(5056) <= not((layer0_outputs(8897)) and (layer0_outputs(8278)));
    outputs(5057) <= not(layer0_outputs(9025));
    outputs(5058) <= not((layer0_outputs(736)) and (layer0_outputs(6676)));
    outputs(5059) <= not((layer0_outputs(1515)) xor (layer0_outputs(9909)));
    outputs(5060) <= layer0_outputs(1274);
    outputs(5061) <= (layer0_outputs(2396)) and (layer0_outputs(5528));
    outputs(5062) <= (layer0_outputs(2775)) and not (layer0_outputs(6499));
    outputs(5063) <= not(layer0_outputs(3123));
    outputs(5064) <= not(layer0_outputs(8554));
    outputs(5065) <= layer0_outputs(899);
    outputs(5066) <= layer0_outputs(8711);
    outputs(5067) <= not(layer0_outputs(89));
    outputs(5068) <= not(layer0_outputs(87)) or (layer0_outputs(8391));
    outputs(5069) <= not(layer0_outputs(6269));
    outputs(5070) <= layer0_outputs(7388);
    outputs(5071) <= layer0_outputs(7029);
    outputs(5072) <= not(layer0_outputs(3521));
    outputs(5073) <= (layer0_outputs(5530)) or (layer0_outputs(7425));
    outputs(5074) <= not(layer0_outputs(5425)) or (layer0_outputs(1324));
    outputs(5075) <= (layer0_outputs(8819)) and not (layer0_outputs(1749));
    outputs(5076) <= layer0_outputs(10038);
    outputs(5077) <= layer0_outputs(6977);
    outputs(5078) <= not((layer0_outputs(8050)) xor (layer0_outputs(533)));
    outputs(5079) <= (layer0_outputs(3002)) and not (layer0_outputs(8574));
    outputs(5080) <= layer0_outputs(2502);
    outputs(5081) <= not(layer0_outputs(6649));
    outputs(5082) <= layer0_outputs(2325);
    outputs(5083) <= not(layer0_outputs(3197));
    outputs(5084) <= not((layer0_outputs(5318)) xor (layer0_outputs(5136)));
    outputs(5085) <= not(layer0_outputs(1428));
    outputs(5086) <= not(layer0_outputs(356));
    outputs(5087) <= (layer0_outputs(4907)) xor (layer0_outputs(3680));
    outputs(5088) <= (layer0_outputs(6189)) xor (layer0_outputs(7764));
    outputs(5089) <= not(layer0_outputs(7263));
    outputs(5090) <= not((layer0_outputs(10104)) or (layer0_outputs(2826)));
    outputs(5091) <= layer0_outputs(1678);
    outputs(5092) <= not(layer0_outputs(5275));
    outputs(5093) <= (layer0_outputs(6326)) and (layer0_outputs(8331));
    outputs(5094) <= layer0_outputs(9816);
    outputs(5095) <= not((layer0_outputs(4752)) or (layer0_outputs(4280)));
    outputs(5096) <= not(layer0_outputs(728));
    outputs(5097) <= not(layer0_outputs(7422));
    outputs(5098) <= not(layer0_outputs(3381));
    outputs(5099) <= not((layer0_outputs(3168)) xor (layer0_outputs(3085)));
    outputs(5100) <= not(layer0_outputs(9867));
    outputs(5101) <= not(layer0_outputs(2244));
    outputs(5102) <= not(layer0_outputs(5215));
    outputs(5103) <= (layer0_outputs(6541)) xor (layer0_outputs(4794));
    outputs(5104) <= layer0_outputs(106);
    outputs(5105) <= layer0_outputs(7371);
    outputs(5106) <= (layer0_outputs(7665)) xor (layer0_outputs(240));
    outputs(5107) <= not(layer0_outputs(5699)) or (layer0_outputs(7152));
    outputs(5108) <= (layer0_outputs(108)) and not (layer0_outputs(5077));
    outputs(5109) <= (layer0_outputs(4221)) and not (layer0_outputs(5640));
    outputs(5110) <= not(layer0_outputs(6207));
    outputs(5111) <= not(layer0_outputs(5524));
    outputs(5112) <= not(layer0_outputs(6743)) or (layer0_outputs(6930));
    outputs(5113) <= not(layer0_outputs(646)) or (layer0_outputs(8718));
    outputs(5114) <= not(layer0_outputs(3798));
    outputs(5115) <= not(layer0_outputs(4466));
    outputs(5116) <= not(layer0_outputs(8454));
    outputs(5117) <= not(layer0_outputs(7526)) or (layer0_outputs(2376));
    outputs(5118) <= (layer0_outputs(9133)) and not (layer0_outputs(9423));
    outputs(5119) <= layer0_outputs(7576);
    outputs(5120) <= layer0_outputs(4021);
    outputs(5121) <= not((layer0_outputs(578)) xor (layer0_outputs(8746)));
    outputs(5122) <= layer0_outputs(4809);
    outputs(5123) <= not(layer0_outputs(6827));
    outputs(5124) <= not((layer0_outputs(10111)) xor (layer0_outputs(2047)));
    outputs(5125) <= (layer0_outputs(9928)) and not (layer0_outputs(4877));
    outputs(5126) <= (layer0_outputs(5558)) and (layer0_outputs(9146));
    outputs(5127) <= not((layer0_outputs(1162)) or (layer0_outputs(8191)));
    outputs(5128) <= layer0_outputs(5629);
    outputs(5129) <= (layer0_outputs(7715)) xor (layer0_outputs(4023));
    outputs(5130) <= (layer0_outputs(9795)) xor (layer0_outputs(8045));
    outputs(5131) <= (layer0_outputs(7736)) xor (layer0_outputs(3684));
    outputs(5132) <= (layer0_outputs(1247)) and (layer0_outputs(2823));
    outputs(5133) <= (layer0_outputs(8081)) xor (layer0_outputs(10217));
    outputs(5134) <= not((layer0_outputs(171)) xor (layer0_outputs(2020)));
    outputs(5135) <= not(layer0_outputs(4864));
    outputs(5136) <= not(layer0_outputs(5436));
    outputs(5137) <= layer0_outputs(494);
    outputs(5138) <= (layer0_outputs(4242)) xor (layer0_outputs(3985));
    outputs(5139) <= layer0_outputs(3455);
    outputs(5140) <= not(layer0_outputs(422));
    outputs(5141) <= layer0_outputs(687);
    outputs(5142) <= not(layer0_outputs(3674));
    outputs(5143) <= not((layer0_outputs(52)) or (layer0_outputs(6750)));
    outputs(5144) <= layer0_outputs(4812);
    outputs(5145) <= not(layer0_outputs(1150)) or (layer0_outputs(3751));
    outputs(5146) <= layer0_outputs(7699);
    outputs(5147) <= not(layer0_outputs(8031)) or (layer0_outputs(7849));
    outputs(5148) <= not((layer0_outputs(7302)) or (layer0_outputs(7162)));
    outputs(5149) <= not((layer0_outputs(969)) xor (layer0_outputs(2292)));
    outputs(5150) <= (layer0_outputs(6470)) and not (layer0_outputs(4400));
    outputs(5151) <= (layer0_outputs(118)) xor (layer0_outputs(7340));
    outputs(5152) <= layer0_outputs(3483);
    outputs(5153) <= not(layer0_outputs(1372)) or (layer0_outputs(5978));
    outputs(5154) <= not((layer0_outputs(9820)) and (layer0_outputs(7592)));
    outputs(5155) <= layer0_outputs(3169);
    outputs(5156) <= not(layer0_outputs(9324));
    outputs(5157) <= not(layer0_outputs(6927));
    outputs(5158) <= not(layer0_outputs(9015));
    outputs(5159) <= not((layer0_outputs(930)) xor (layer0_outputs(9409)));
    outputs(5160) <= layer0_outputs(7472);
    outputs(5161) <= layer0_outputs(5265);
    outputs(5162) <= not(layer0_outputs(4792));
    outputs(5163) <= not((layer0_outputs(9267)) xor (layer0_outputs(2243)));
    outputs(5164) <= layer0_outputs(8939);
    outputs(5165) <= layer0_outputs(131);
    outputs(5166) <= layer0_outputs(6527);
    outputs(5167) <= (layer0_outputs(2938)) xor (layer0_outputs(6670));
    outputs(5168) <= not(layer0_outputs(5317)) or (layer0_outputs(7573));
    outputs(5169) <= not((layer0_outputs(1786)) xor (layer0_outputs(8519)));
    outputs(5170) <= layer0_outputs(360);
    outputs(5171) <= (layer0_outputs(8994)) xor (layer0_outputs(4335));
    outputs(5172) <= not(layer0_outputs(10172));
    outputs(5173) <= not((layer0_outputs(2808)) xor (layer0_outputs(1189)));
    outputs(5174) <= not(layer0_outputs(1869));
    outputs(5175) <= (layer0_outputs(2429)) xor (layer0_outputs(8383));
    outputs(5176) <= not(layer0_outputs(9471));
    outputs(5177) <= (layer0_outputs(485)) xor (layer0_outputs(1883));
    outputs(5178) <= not(layer0_outputs(3180));
    outputs(5179) <= layer0_outputs(6275);
    outputs(5180) <= not(layer0_outputs(8263));
    outputs(5181) <= (layer0_outputs(7594)) xor (layer0_outputs(6062));
    outputs(5182) <= not((layer0_outputs(8959)) or (layer0_outputs(8314)));
    outputs(5183) <= (layer0_outputs(3133)) and not (layer0_outputs(4309));
    outputs(5184) <= not((layer0_outputs(3268)) xor (layer0_outputs(3462)));
    outputs(5185) <= not((layer0_outputs(1455)) xor (layer0_outputs(4882)));
    outputs(5186) <= not((layer0_outputs(5141)) xor (layer0_outputs(10016)));
    outputs(5187) <= not(layer0_outputs(9306));
    outputs(5188) <= (layer0_outputs(6968)) and (layer0_outputs(5694));
    outputs(5189) <= not(layer0_outputs(7394)) or (layer0_outputs(523));
    outputs(5190) <= not(layer0_outputs(882));
    outputs(5191) <= (layer0_outputs(8884)) and not (layer0_outputs(2101));
    outputs(5192) <= not(layer0_outputs(1657));
    outputs(5193) <= not(layer0_outputs(8544));
    outputs(5194) <= layer0_outputs(2571);
    outputs(5195) <= (layer0_outputs(5695)) xor (layer0_outputs(2850));
    outputs(5196) <= not(layer0_outputs(6188));
    outputs(5197) <= (layer0_outputs(5950)) xor (layer0_outputs(5605));
    outputs(5198) <= not(layer0_outputs(8908));
    outputs(5199) <= layer0_outputs(346);
    outputs(5200) <= not(layer0_outputs(4009));
    outputs(5201) <= not(layer0_outputs(970)) or (layer0_outputs(10086));
    outputs(5202) <= layer0_outputs(4274);
    outputs(5203) <= not((layer0_outputs(6137)) xor (layer0_outputs(9885)));
    outputs(5204) <= not(layer0_outputs(685)) or (layer0_outputs(8208));
    outputs(5205) <= layer0_outputs(9920);
    outputs(5206) <= layer0_outputs(3598);
    outputs(5207) <= not((layer0_outputs(2272)) xor (layer0_outputs(6308)));
    outputs(5208) <= not((layer0_outputs(8997)) xor (layer0_outputs(8907)));
    outputs(5209) <= (layer0_outputs(5706)) and not (layer0_outputs(7219));
    outputs(5210) <= not(layer0_outputs(3536)) or (layer0_outputs(8755));
    outputs(5211) <= not((layer0_outputs(7367)) xor (layer0_outputs(9530)));
    outputs(5212) <= not(layer0_outputs(4598));
    outputs(5213) <= not(layer0_outputs(6846));
    outputs(5214) <= (layer0_outputs(2972)) and not (layer0_outputs(1788));
    outputs(5215) <= (layer0_outputs(9120)) or (layer0_outputs(10041));
    outputs(5216) <= not((layer0_outputs(9912)) xor (layer0_outputs(8946)));
    outputs(5217) <= not(layer0_outputs(4668));
    outputs(5218) <= not(layer0_outputs(8499));
    outputs(5219) <= (layer0_outputs(1329)) xor (layer0_outputs(1297));
    outputs(5220) <= layer0_outputs(8276);
    outputs(5221) <= not((layer0_outputs(4099)) xor (layer0_outputs(6703)));
    outputs(5222) <= not((layer0_outputs(556)) or (layer0_outputs(7819)));
    outputs(5223) <= layer0_outputs(2023);
    outputs(5224) <= (layer0_outputs(5274)) xor (layer0_outputs(2481));
    outputs(5225) <= (layer0_outputs(7216)) xor (layer0_outputs(1679));
    outputs(5226) <= (layer0_outputs(9561)) or (layer0_outputs(5228));
    outputs(5227) <= not(layer0_outputs(5436));
    outputs(5228) <= not(layer0_outputs(85));
    outputs(5229) <= not((layer0_outputs(7516)) or (layer0_outputs(3546)));
    outputs(5230) <= not(layer0_outputs(8680)) or (layer0_outputs(9695));
    outputs(5231) <= not(layer0_outputs(4312));
    outputs(5232) <= (layer0_outputs(2084)) xor (layer0_outputs(8519));
    outputs(5233) <= not((layer0_outputs(6912)) xor (layer0_outputs(3405)));
    outputs(5234) <= not((layer0_outputs(9564)) or (layer0_outputs(6046)));
    outputs(5235) <= (layer0_outputs(229)) xor (layer0_outputs(4359));
    outputs(5236) <= not((layer0_outputs(899)) and (layer0_outputs(656)));
    outputs(5237) <= layer0_outputs(8430);
    outputs(5238) <= not(layer0_outputs(5981)) or (layer0_outputs(7839));
    outputs(5239) <= not(layer0_outputs(2131));
    outputs(5240) <= (layer0_outputs(7259)) xor (layer0_outputs(4657));
    outputs(5241) <= not((layer0_outputs(6698)) or (layer0_outputs(6510)));
    outputs(5242) <= (layer0_outputs(4337)) and (layer0_outputs(6198));
    outputs(5243) <= not((layer0_outputs(4633)) or (layer0_outputs(5202)));
    outputs(5244) <= not((layer0_outputs(7946)) or (layer0_outputs(422)));
    outputs(5245) <= not(layer0_outputs(5602));
    outputs(5246) <= not(layer0_outputs(110));
    outputs(5247) <= (layer0_outputs(270)) and (layer0_outputs(9776));
    outputs(5248) <= layer0_outputs(7482);
    outputs(5249) <= not(layer0_outputs(9790));
    outputs(5250) <= (layer0_outputs(7499)) and not (layer0_outputs(8647));
    outputs(5251) <= (layer0_outputs(7944)) xor (layer0_outputs(7366));
    outputs(5252) <= layer0_outputs(8297);
    outputs(5253) <= layer0_outputs(6063);
    outputs(5254) <= not((layer0_outputs(528)) and (layer0_outputs(1181)));
    outputs(5255) <= (layer0_outputs(8629)) xor (layer0_outputs(5455));
    outputs(5256) <= (layer0_outputs(4711)) xor (layer0_outputs(6869));
    outputs(5257) <= not(layer0_outputs(3642)) or (layer0_outputs(8418));
    outputs(5258) <= not(layer0_outputs(6029));
    outputs(5259) <= not(layer0_outputs(7357)) or (layer0_outputs(3112));
    outputs(5260) <= not(layer0_outputs(6833)) or (layer0_outputs(1062));
    outputs(5261) <= layer0_outputs(7147);
    outputs(5262) <= not(layer0_outputs(2496));
    outputs(5263) <= (layer0_outputs(9614)) and (layer0_outputs(850));
    outputs(5264) <= not(layer0_outputs(5415));
    outputs(5265) <= layer0_outputs(8000);
    outputs(5266) <= layer0_outputs(2678);
    outputs(5267) <= (layer0_outputs(4612)) xor (layer0_outputs(1080));
    outputs(5268) <= (layer0_outputs(6687)) and not (layer0_outputs(8732));
    outputs(5269) <= not(layer0_outputs(5282));
    outputs(5270) <= (layer0_outputs(3557)) xor (layer0_outputs(4476));
    outputs(5271) <= (layer0_outputs(8401)) xor (layer0_outputs(685));
    outputs(5272) <= not((layer0_outputs(7383)) and (layer0_outputs(320)));
    outputs(5273) <= not(layer0_outputs(7812));
    outputs(5274) <= not(layer0_outputs(6885)) or (layer0_outputs(7699));
    outputs(5275) <= layer0_outputs(613);
    outputs(5276) <= (layer0_outputs(8797)) xor (layer0_outputs(6337));
    outputs(5277) <= not(layer0_outputs(3014));
    outputs(5278) <= not(layer0_outputs(5226));
    outputs(5279) <= not(layer0_outputs(6818));
    outputs(5280) <= not(layer0_outputs(3895));
    outputs(5281) <= not(layer0_outputs(2755));
    outputs(5282) <= (layer0_outputs(3975)) xor (layer0_outputs(2972));
    outputs(5283) <= not(layer0_outputs(214));
    outputs(5284) <= layer0_outputs(4950);
    outputs(5285) <= (layer0_outputs(5333)) xor (layer0_outputs(9516));
    outputs(5286) <= layer0_outputs(6141);
    outputs(5287) <= not(layer0_outputs(2699));
    outputs(5288) <= not(layer0_outputs(4525));
    outputs(5289) <= (layer0_outputs(3715)) xor (layer0_outputs(5574));
    outputs(5290) <= layer0_outputs(7794);
    outputs(5291) <= (layer0_outputs(5754)) and (layer0_outputs(446));
    outputs(5292) <= not(layer0_outputs(5973)) or (layer0_outputs(6929));
    outputs(5293) <= (layer0_outputs(9071)) and not (layer0_outputs(1175));
    outputs(5294) <= layer0_outputs(9062);
    outputs(5295) <= not((layer0_outputs(7010)) xor (layer0_outputs(5151)));
    outputs(5296) <= layer0_outputs(1611);
    outputs(5297) <= not((layer0_outputs(2860)) or (layer0_outputs(6572)));
    outputs(5298) <= not(layer0_outputs(5343));
    outputs(5299) <= (layer0_outputs(4857)) and not (layer0_outputs(1068));
    outputs(5300) <= (layer0_outputs(3589)) or (layer0_outputs(572));
    outputs(5301) <= layer0_outputs(636);
    outputs(5302) <= (layer0_outputs(3969)) xor (layer0_outputs(5110));
    outputs(5303) <= (layer0_outputs(3169)) and not (layer0_outputs(6270));
    outputs(5304) <= not(layer0_outputs(8412));
    outputs(5305) <= not(layer0_outputs(4517));
    outputs(5306) <= not((layer0_outputs(1363)) xor (layer0_outputs(9462)));
    outputs(5307) <= not(layer0_outputs(5208));
    outputs(5308) <= (layer0_outputs(1429)) xor (layer0_outputs(9520));
    outputs(5309) <= (layer0_outputs(5083)) and not (layer0_outputs(5427));
    outputs(5310) <= not((layer0_outputs(7971)) and (layer0_outputs(2449)));
    outputs(5311) <= not(layer0_outputs(3234)) or (layer0_outputs(4990));
    outputs(5312) <= not(layer0_outputs(3252));
    outputs(5313) <= (layer0_outputs(1102)) xor (layer0_outputs(5092));
    outputs(5314) <= layer0_outputs(4461);
    outputs(5315) <= (layer0_outputs(6493)) xor (layer0_outputs(4202));
    outputs(5316) <= not(layer0_outputs(852));
    outputs(5317) <= layer0_outputs(415);
    outputs(5318) <= layer0_outputs(4351);
    outputs(5319) <= not(layer0_outputs(9676));
    outputs(5320) <= (layer0_outputs(588)) and not (layer0_outputs(4252));
    outputs(5321) <= not(layer0_outputs(2003));
    outputs(5322) <= not((layer0_outputs(207)) and (layer0_outputs(531)));
    outputs(5323) <= not(layer0_outputs(6573));
    outputs(5324) <= (layer0_outputs(3321)) xor (layer0_outputs(3688));
    outputs(5325) <= not((layer0_outputs(1016)) xor (layer0_outputs(7773)));
    outputs(5326) <= layer0_outputs(9012);
    outputs(5327) <= layer0_outputs(4161);
    outputs(5328) <= (layer0_outputs(758)) and not (layer0_outputs(5912));
    outputs(5329) <= (layer0_outputs(9750)) xor (layer0_outputs(4516));
    outputs(5330) <= layer0_outputs(2186);
    outputs(5331) <= layer0_outputs(601);
    outputs(5332) <= (layer0_outputs(7671)) or (layer0_outputs(3048));
    outputs(5333) <= (layer0_outputs(3232)) xor (layer0_outputs(4315));
    outputs(5334) <= not(layer0_outputs(2649));
    outputs(5335) <= (layer0_outputs(2433)) xor (layer0_outputs(10122));
    outputs(5336) <= layer0_outputs(7081);
    outputs(5337) <= not(layer0_outputs(9767));
    outputs(5338) <= (layer0_outputs(889)) xor (layer0_outputs(2280));
    outputs(5339) <= layer0_outputs(6990);
    outputs(5340) <= (layer0_outputs(2929)) and not (layer0_outputs(1034));
    outputs(5341) <= layer0_outputs(610);
    outputs(5342) <= (layer0_outputs(2081)) xor (layer0_outputs(5001));
    outputs(5343) <= layer0_outputs(6498);
    outputs(5344) <= (layer0_outputs(9973)) or (layer0_outputs(10153));
    outputs(5345) <= not(layer0_outputs(6547)) or (layer0_outputs(8815));
    outputs(5346) <= not(layer0_outputs(6388));
    outputs(5347) <= layer0_outputs(7985);
    outputs(5348) <= not(layer0_outputs(8894));
    outputs(5349) <= not((layer0_outputs(3803)) or (layer0_outputs(2136)));
    outputs(5350) <= layer0_outputs(7684);
    outputs(5351) <= not((layer0_outputs(9949)) and (layer0_outputs(1689)));
    outputs(5352) <= (layer0_outputs(10228)) and not (layer0_outputs(3300));
    outputs(5353) <= not((layer0_outputs(6825)) or (layer0_outputs(5728)));
    outputs(5354) <= layer0_outputs(4418);
    outputs(5355) <= not((layer0_outputs(933)) and (layer0_outputs(1665)));
    outputs(5356) <= (layer0_outputs(7737)) xor (layer0_outputs(7887));
    outputs(5357) <= not(layer0_outputs(39));
    outputs(5358) <= (layer0_outputs(4364)) or (layer0_outputs(9126));
    outputs(5359) <= not(layer0_outputs(4902));
    outputs(5360) <= not(layer0_outputs(805));
    outputs(5361) <= not(layer0_outputs(9880));
    outputs(5362) <= (layer0_outputs(5836)) xor (layer0_outputs(1775));
    outputs(5363) <= not(layer0_outputs(4409)) or (layer0_outputs(8076));
    outputs(5364) <= (layer0_outputs(3916)) xor (layer0_outputs(5796));
    outputs(5365) <= layer0_outputs(7386);
    outputs(5366) <= (layer0_outputs(2863)) xor (layer0_outputs(8335));
    outputs(5367) <= layer0_outputs(8027);
    outputs(5368) <= (layer0_outputs(7938)) xor (layer0_outputs(7853));
    outputs(5369) <= (layer0_outputs(992)) xor (layer0_outputs(1493));
    outputs(5370) <= (layer0_outputs(750)) and not (layer0_outputs(2253));
    outputs(5371) <= (layer0_outputs(4606)) xor (layer0_outputs(3900));
    outputs(5372) <= (layer0_outputs(4578)) xor (layer0_outputs(742));
    outputs(5373) <= (layer0_outputs(1643)) and not (layer0_outputs(7193));
    outputs(5374) <= (layer0_outputs(5398)) or (layer0_outputs(5024));
    outputs(5375) <= (layer0_outputs(9071)) and not (layer0_outputs(5053));
    outputs(5376) <= (layer0_outputs(7659)) and (layer0_outputs(5127));
    outputs(5377) <= not((layer0_outputs(5205)) and (layer0_outputs(3445)));
    outputs(5378) <= (layer0_outputs(5160)) and (layer0_outputs(9228));
    outputs(5379) <= not(layer0_outputs(6382));
    outputs(5380) <= not(layer0_outputs(10181));
    outputs(5381) <= not((layer0_outputs(9276)) xor (layer0_outputs(8353)));
    outputs(5382) <= (layer0_outputs(1620)) xor (layer0_outputs(4148));
    outputs(5383) <= (layer0_outputs(1205)) xor (layer0_outputs(3336));
    outputs(5384) <= not((layer0_outputs(9339)) xor (layer0_outputs(8496)));
    outputs(5385) <= layer0_outputs(4052);
    outputs(5386) <= (layer0_outputs(9054)) and not (layer0_outputs(306));
    outputs(5387) <= not(layer0_outputs(7721));
    outputs(5388) <= layer0_outputs(1997);
    outputs(5389) <= layer0_outputs(3382);
    outputs(5390) <= not((layer0_outputs(9842)) xor (layer0_outputs(2092)));
    outputs(5391) <= (layer0_outputs(4741)) xor (layer0_outputs(6722));
    outputs(5392) <= layer0_outputs(3121);
    outputs(5393) <= not(layer0_outputs(4015)) or (layer0_outputs(8839));
    outputs(5394) <= not(layer0_outputs(2229));
    outputs(5395) <= (layer0_outputs(6262)) xor (layer0_outputs(8566));
    outputs(5396) <= not(layer0_outputs(4079));
    outputs(5397) <= not(layer0_outputs(776));
    outputs(5398) <= not(layer0_outputs(700)) or (layer0_outputs(4770));
    outputs(5399) <= not(layer0_outputs(8370));
    outputs(5400) <= not((layer0_outputs(8358)) xor (layer0_outputs(9469)));
    outputs(5401) <= (layer0_outputs(7941)) xor (layer0_outputs(9996));
    outputs(5402) <= layer0_outputs(7552);
    outputs(5403) <= (layer0_outputs(7700)) and not (layer0_outputs(9352));
    outputs(5404) <= not((layer0_outputs(6309)) xor (layer0_outputs(8452)));
    outputs(5405) <= not(layer0_outputs(6341));
    outputs(5406) <= layer0_outputs(4872);
    outputs(5407) <= layer0_outputs(4026);
    outputs(5408) <= not((layer0_outputs(7577)) xor (layer0_outputs(7384)));
    outputs(5409) <= (layer0_outputs(6636)) xor (layer0_outputs(7444));
    outputs(5410) <= not((layer0_outputs(3443)) xor (layer0_outputs(8871)));
    outputs(5411) <= not(layer0_outputs(5759)) or (layer0_outputs(652));
    outputs(5412) <= layer0_outputs(6568);
    outputs(5413) <= not(layer0_outputs(6245));
    outputs(5414) <= layer0_outputs(1471);
    outputs(5415) <= not(layer0_outputs(326)) or (layer0_outputs(8932));
    outputs(5416) <= (layer0_outputs(212)) xor (layer0_outputs(6977));
    outputs(5417) <= not(layer0_outputs(317));
    outputs(5418) <= not(layer0_outputs(10098));
    outputs(5419) <= not((layer0_outputs(6950)) and (layer0_outputs(2318)));
    outputs(5420) <= (layer0_outputs(6604)) xor (layer0_outputs(1486));
    outputs(5421) <= layer0_outputs(427);
    outputs(5422) <= (layer0_outputs(3864)) and not (layer0_outputs(697));
    outputs(5423) <= not((layer0_outputs(5675)) xor (layer0_outputs(1483)));
    outputs(5424) <= (layer0_outputs(5761)) xor (layer0_outputs(7084));
    outputs(5425) <= layer0_outputs(6674);
    outputs(5426) <= not((layer0_outputs(10077)) xor (layer0_outputs(3426)));
    outputs(5427) <= (layer0_outputs(1741)) xor (layer0_outputs(7169));
    outputs(5428) <= not(layer0_outputs(2210));
    outputs(5429) <= not((layer0_outputs(3846)) and (layer0_outputs(815)));
    outputs(5430) <= not(layer0_outputs(9674));
    outputs(5431) <= not(layer0_outputs(4996));
    outputs(5432) <= (layer0_outputs(8757)) xor (layer0_outputs(811));
    outputs(5433) <= (layer0_outputs(561)) xor (layer0_outputs(8480));
    outputs(5434) <= not(layer0_outputs(7757));
    outputs(5435) <= not(layer0_outputs(5094)) or (layer0_outputs(5383));
    outputs(5436) <= layer0_outputs(4057);
    outputs(5437) <= not(layer0_outputs(5995));
    outputs(5438) <= (layer0_outputs(7311)) or (layer0_outputs(9859));
    outputs(5439) <= not((layer0_outputs(3604)) xor (layer0_outputs(2537)));
    outputs(5440) <= (layer0_outputs(4144)) xor (layer0_outputs(2524));
    outputs(5441) <= not(layer0_outputs(4746));
    outputs(5442) <= not(layer0_outputs(6792));
    outputs(5443) <= layer0_outputs(8207);
    outputs(5444) <= (layer0_outputs(569)) and not (layer0_outputs(7395));
    outputs(5445) <= not(layer0_outputs(7227));
    outputs(5446) <= not((layer0_outputs(9224)) and (layer0_outputs(2482)));
    outputs(5447) <= layer0_outputs(6122);
    outputs(5448) <= layer0_outputs(1298);
    outputs(5449) <= layer0_outputs(8533);
    outputs(5450) <= not(layer0_outputs(2617));
    outputs(5451) <= not(layer0_outputs(2633));
    outputs(5452) <= (layer0_outputs(7780)) xor (layer0_outputs(235));
    outputs(5453) <= layer0_outputs(5577);
    outputs(5454) <= layer0_outputs(2847);
    outputs(5455) <= (layer0_outputs(6976)) or (layer0_outputs(5541));
    outputs(5456) <= not((layer0_outputs(3976)) xor (layer0_outputs(9429)));
    outputs(5457) <= layer0_outputs(1169);
    outputs(5458) <= layer0_outputs(3087);
    outputs(5459) <= not(layer0_outputs(5889));
    outputs(5460) <= not(layer0_outputs(9629));
    outputs(5461) <= not(layer0_outputs(1424)) or (layer0_outputs(7978));
    outputs(5462) <= not(layer0_outputs(9000));
    outputs(5463) <= (layer0_outputs(9568)) and not (layer0_outputs(1625));
    outputs(5464) <= (layer0_outputs(8763)) xor (layer0_outputs(3190));
    outputs(5465) <= not((layer0_outputs(1549)) xor (layer0_outputs(3366)));
    outputs(5466) <= not(layer0_outputs(5755)) or (layer0_outputs(619));
    outputs(5467) <= not((layer0_outputs(8052)) xor (layer0_outputs(8641)));
    outputs(5468) <= (layer0_outputs(2614)) xor (layer0_outputs(8228));
    outputs(5469) <= layer0_outputs(6222);
    outputs(5470) <= (layer0_outputs(970)) xor (layer0_outputs(1357));
    outputs(5471) <= not(layer0_outputs(8221));
    outputs(5472) <= not(layer0_outputs(9339));
    outputs(5473) <= (layer0_outputs(1204)) xor (layer0_outputs(9755));
    outputs(5474) <= not((layer0_outputs(983)) xor (layer0_outputs(6398)));
    outputs(5475) <= (layer0_outputs(1259)) xor (layer0_outputs(4946));
    outputs(5476) <= (layer0_outputs(7745)) xor (layer0_outputs(7456));
    outputs(5477) <= (layer0_outputs(5165)) xor (layer0_outputs(5879));
    outputs(5478) <= not((layer0_outputs(10214)) xor (layer0_outputs(8489)));
    outputs(5479) <= layer0_outputs(5605);
    outputs(5480) <= not((layer0_outputs(4501)) xor (layer0_outputs(3842)));
    outputs(5481) <= not(layer0_outputs(3534));
    outputs(5482) <= layer0_outputs(1366);
    outputs(5483) <= (layer0_outputs(5274)) xor (layer0_outputs(4297));
    outputs(5484) <= not(layer0_outputs(8972)) or (layer0_outputs(8073));
    outputs(5485) <= not((layer0_outputs(7865)) xor (layer0_outputs(8491)));
    outputs(5486) <= (layer0_outputs(2718)) xor (layer0_outputs(221));
    outputs(5487) <= not(layer0_outputs(6583));
    outputs(5488) <= layer0_outputs(10048);
    outputs(5489) <= not((layer0_outputs(9541)) or (layer0_outputs(8668)));
    outputs(5490) <= (layer0_outputs(5332)) xor (layer0_outputs(4832));
    outputs(5491) <= layer0_outputs(616);
    outputs(5492) <= layer0_outputs(1458);
    outputs(5493) <= not(layer0_outputs(608));
    outputs(5494) <= layer0_outputs(3707);
    outputs(5495) <= (layer0_outputs(5306)) or (layer0_outputs(2427));
    outputs(5496) <= not((layer0_outputs(195)) xor (layer0_outputs(2540)));
    outputs(5497) <= (layer0_outputs(7740)) and not (layer0_outputs(3671));
    outputs(5498) <= not((layer0_outputs(2801)) xor (layer0_outputs(3507)));
    outputs(5499) <= layer0_outputs(5856);
    outputs(5500) <= layer0_outputs(5960);
    outputs(5501) <= layer0_outputs(1548);
    outputs(5502) <= (layer0_outputs(4979)) xor (layer0_outputs(7926));
    outputs(5503) <= not(layer0_outputs(2695));
    outputs(5504) <= (layer0_outputs(525)) xor (layer0_outputs(6535));
    outputs(5505) <= (layer0_outputs(3512)) or (layer0_outputs(3998));
    outputs(5506) <= (layer0_outputs(2307)) and not (layer0_outputs(6588));
    outputs(5507) <= (layer0_outputs(2207)) xor (layer0_outputs(9618));
    outputs(5508) <= layer0_outputs(5163);
    outputs(5509) <= not(layer0_outputs(1061));
    outputs(5510) <= (layer0_outputs(5288)) xor (layer0_outputs(6988));
    outputs(5511) <= (layer0_outputs(1874)) and not (layer0_outputs(6352));
    outputs(5512) <= layer0_outputs(5898);
    outputs(5513) <= (layer0_outputs(4705)) and (layer0_outputs(2729));
    outputs(5514) <= (layer0_outputs(7492)) xor (layer0_outputs(3502));
    outputs(5515) <= (layer0_outputs(3670)) xor (layer0_outputs(514));
    outputs(5516) <= not((layer0_outputs(8752)) xor (layer0_outputs(2197)));
    outputs(5517) <= not(layer0_outputs(3576));
    outputs(5518) <= (layer0_outputs(8484)) and not (layer0_outputs(2552));
    outputs(5519) <= (layer0_outputs(807)) and (layer0_outputs(1806));
    outputs(5520) <= not(layer0_outputs(5922));
    outputs(5521) <= layer0_outputs(5861);
    outputs(5522) <= (layer0_outputs(4192)) or (layer0_outputs(4952));
    outputs(5523) <= not(layer0_outputs(5389));
    outputs(5524) <= layer0_outputs(3864);
    outputs(5525) <= (layer0_outputs(2766)) xor (layer0_outputs(4344));
    outputs(5526) <= not(layer0_outputs(5868));
    outputs(5527) <= not((layer0_outputs(9003)) xor (layer0_outputs(5337)));
    outputs(5528) <= not((layer0_outputs(9890)) or (layer0_outputs(2835)));
    outputs(5529) <= (layer0_outputs(4680)) and (layer0_outputs(7472));
    outputs(5530) <= not((layer0_outputs(8245)) or (layer0_outputs(7435)));
    outputs(5531) <= not((layer0_outputs(2573)) xor (layer0_outputs(5811)));
    outputs(5532) <= (layer0_outputs(2848)) xor (layer0_outputs(1856));
    outputs(5533) <= not((layer0_outputs(7060)) xor (layer0_outputs(4114)));
    outputs(5534) <= (layer0_outputs(7310)) xor (layer0_outputs(891));
    outputs(5535) <= not((layer0_outputs(1785)) xor (layer0_outputs(4668)));
    outputs(5536) <= not((layer0_outputs(8372)) and (layer0_outputs(10099)));
    outputs(5537) <= (layer0_outputs(1863)) xor (layer0_outputs(5264));
    outputs(5538) <= not((layer0_outputs(9190)) or (layer0_outputs(9779)));
    outputs(5539) <= layer0_outputs(7829);
    outputs(5540) <= not((layer0_outputs(2989)) xor (layer0_outputs(7586)));
    outputs(5541) <= not(layer0_outputs(9567)) or (layer0_outputs(6143));
    outputs(5542) <= layer0_outputs(6770);
    outputs(5543) <= not((layer0_outputs(8022)) xor (layer0_outputs(8168)));
    outputs(5544) <= layer0_outputs(2965);
    outputs(5545) <= not((layer0_outputs(665)) xor (layer0_outputs(3463)));
    outputs(5546) <= layer0_outputs(7560);
    outputs(5547) <= (layer0_outputs(9729)) xor (layer0_outputs(561));
    outputs(5548) <= layer0_outputs(3528);
    outputs(5549) <= not((layer0_outputs(8621)) xor (layer0_outputs(6155)));
    outputs(5550) <= (layer0_outputs(6851)) and (layer0_outputs(7615));
    outputs(5551) <= not((layer0_outputs(4151)) xor (layer0_outputs(4958)));
    outputs(5552) <= (layer0_outputs(4469)) and (layer0_outputs(1401));
    outputs(5553) <= (layer0_outputs(6657)) and not (layer0_outputs(4034));
    outputs(5554) <= layer0_outputs(223);
    outputs(5555) <= layer0_outputs(1801);
    outputs(5556) <= layer0_outputs(1975);
    outputs(5557) <= not(layer0_outputs(6417)) or (layer0_outputs(2547));
    outputs(5558) <= not((layer0_outputs(5305)) xor (layer0_outputs(6031)));
    outputs(5559) <= layer0_outputs(4319);
    outputs(5560) <= not((layer0_outputs(7165)) and (layer0_outputs(324)));
    outputs(5561) <= (layer0_outputs(8892)) xor (layer0_outputs(3482));
    outputs(5562) <= (layer0_outputs(2810)) xor (layer0_outputs(6797));
    outputs(5563) <= not(layer0_outputs(7067));
    outputs(5564) <= not((layer0_outputs(425)) xor (layer0_outputs(2591)));
    outputs(5565) <= layer0_outputs(5518);
    outputs(5566) <= not((layer0_outputs(420)) xor (layer0_outputs(3061)));
    outputs(5567) <= not((layer0_outputs(3400)) xor (layer0_outputs(3515)));
    outputs(5568) <= not((layer0_outputs(5646)) xor (layer0_outputs(3367)));
    outputs(5569) <= layer0_outputs(8061);
    outputs(5570) <= layer0_outputs(1904);
    outputs(5571) <= not(layer0_outputs(5347));
    outputs(5572) <= not(layer0_outputs(9395)) or (layer0_outputs(2134));
    outputs(5573) <= (layer0_outputs(7285)) xor (layer0_outputs(7884));
    outputs(5574) <= layer0_outputs(2086);
    outputs(5575) <= not(layer0_outputs(5718));
    outputs(5576) <= not(layer0_outputs(6096));
    outputs(5577) <= (layer0_outputs(2018)) and not (layer0_outputs(3850));
    outputs(5578) <= (layer0_outputs(609)) or (layer0_outputs(8754));
    outputs(5579) <= not((layer0_outputs(7168)) or (layer0_outputs(4924)));
    outputs(5580) <= not(layer0_outputs(854)) or (layer0_outputs(3743));
    outputs(5581) <= not((layer0_outputs(6211)) or (layer0_outputs(1736)));
    outputs(5582) <= (layer0_outputs(4543)) and not (layer0_outputs(5686));
    outputs(5583) <= (layer0_outputs(6510)) xor (layer0_outputs(8442));
    outputs(5584) <= not((layer0_outputs(5089)) xor (layer0_outputs(800)));
    outputs(5585) <= not(layer0_outputs(6425)) or (layer0_outputs(4135));
    outputs(5586) <= not(layer0_outputs(9802));
    outputs(5587) <= layer0_outputs(9438);
    outputs(5588) <= (layer0_outputs(2178)) and not (layer0_outputs(3667));
    outputs(5589) <= (layer0_outputs(3090)) xor (layer0_outputs(8119));
    outputs(5590) <= not(layer0_outputs(9401));
    outputs(5591) <= not(layer0_outputs(5017));
    outputs(5592) <= (layer0_outputs(5434)) and (layer0_outputs(4774));
    outputs(5593) <= not((layer0_outputs(7705)) xor (layer0_outputs(5737)));
    outputs(5594) <= not(layer0_outputs(5604));
    outputs(5595) <= (layer0_outputs(3977)) xor (layer0_outputs(6379));
    outputs(5596) <= (layer0_outputs(2719)) xor (layer0_outputs(3938));
    outputs(5597) <= not(layer0_outputs(2315));
    outputs(5598) <= not((layer0_outputs(10)) xor (layer0_outputs(9512)));
    outputs(5599) <= not((layer0_outputs(9471)) xor (layer0_outputs(5123)));
    outputs(5600) <= not(layer0_outputs(1143));
    outputs(5601) <= layer0_outputs(2661);
    outputs(5602) <= (layer0_outputs(3017)) xor (layer0_outputs(6937));
    outputs(5603) <= not(layer0_outputs(2137));
    outputs(5604) <= not((layer0_outputs(1756)) xor (layer0_outputs(7133)));
    outputs(5605) <= not(layer0_outputs(9940));
    outputs(5606) <= not(layer0_outputs(5855));
    outputs(5607) <= not((layer0_outputs(595)) xor (layer0_outputs(8748)));
    outputs(5608) <= layer0_outputs(5496);
    outputs(5609) <= layer0_outputs(7157);
    outputs(5610) <= not(layer0_outputs(4030));
    outputs(5611) <= not((layer0_outputs(1287)) xor (layer0_outputs(6748)));
    outputs(5612) <= not((layer0_outputs(8247)) xor (layer0_outputs(5672)));
    outputs(5613) <= not(layer0_outputs(4205)) or (layer0_outputs(3951));
    outputs(5614) <= not((layer0_outputs(7122)) xor (layer0_outputs(6823)));
    outputs(5615) <= (layer0_outputs(7148)) or (layer0_outputs(9106));
    outputs(5616) <= not((layer0_outputs(8080)) or (layer0_outputs(11)));
    outputs(5617) <= (layer0_outputs(5543)) xor (layer0_outputs(8671));
    outputs(5618) <= not(layer0_outputs(8366));
    outputs(5619) <= not(layer0_outputs(9967));
    outputs(5620) <= not((layer0_outputs(6623)) and (layer0_outputs(10213)));
    outputs(5621) <= not(layer0_outputs(6023));
    outputs(5622) <= not(layer0_outputs(1453));
    outputs(5623) <= not(layer0_outputs(5463)) or (layer0_outputs(6855));
    outputs(5624) <= (layer0_outputs(2513)) xor (layer0_outputs(3365));
    outputs(5625) <= layer0_outputs(353);
    outputs(5626) <= layer0_outputs(7230);
    outputs(5627) <= (layer0_outputs(6872)) xor (layer0_outputs(4325));
    outputs(5628) <= not(layer0_outputs(6306));
    outputs(5629) <= not((layer0_outputs(9033)) xor (layer0_outputs(128)));
    outputs(5630) <= (layer0_outputs(2830)) and not (layer0_outputs(934));
    outputs(5631) <= layer0_outputs(10208);
    outputs(5632) <= not((layer0_outputs(4984)) and (layer0_outputs(8325)));
    outputs(5633) <= not(layer0_outputs(3232));
    outputs(5634) <= layer0_outputs(9583);
    outputs(5635) <= (layer0_outputs(4579)) xor (layer0_outputs(3004));
    outputs(5636) <= not((layer0_outputs(3844)) or (layer0_outputs(3338)));
    outputs(5637) <= not((layer0_outputs(6104)) xor (layer0_outputs(10004)));
    outputs(5638) <= not(layer0_outputs(521));
    outputs(5639) <= layer0_outputs(8988);
    outputs(5640) <= (layer0_outputs(1403)) or (layer0_outputs(7416));
    outputs(5641) <= not(layer0_outputs(8044));
    outputs(5642) <= not(layer0_outputs(8355)) or (layer0_outputs(2014));
    outputs(5643) <= layer0_outputs(7031);
    outputs(5644) <= not(layer0_outputs(4467));
    outputs(5645) <= (layer0_outputs(19)) xor (layer0_outputs(5153));
    outputs(5646) <= layer0_outputs(8410);
    outputs(5647) <= (layer0_outputs(7776)) or (layer0_outputs(8679));
    outputs(5648) <= not((layer0_outputs(9351)) xor (layer0_outputs(9781)));
    outputs(5649) <= not((layer0_outputs(6659)) xor (layer0_outputs(1968)));
    outputs(5650) <= layer0_outputs(4577);
    outputs(5651) <= not((layer0_outputs(4562)) or (layer0_outputs(2281)));
    outputs(5652) <= not(layer0_outputs(1052)) or (layer0_outputs(4130));
    outputs(5653) <= not((layer0_outputs(1704)) xor (layer0_outputs(7562)));
    outputs(5654) <= (layer0_outputs(3163)) xor (layer0_outputs(7906));
    outputs(5655) <= not((layer0_outputs(5598)) xor (layer0_outputs(1481)));
    outputs(5656) <= not((layer0_outputs(843)) xor (layer0_outputs(3468)));
    outputs(5657) <= layer0_outputs(8958);
    outputs(5658) <= (layer0_outputs(8726)) xor (layer0_outputs(9701));
    outputs(5659) <= (layer0_outputs(4713)) and (layer0_outputs(4272));
    outputs(5660) <= not((layer0_outputs(2531)) xor (layer0_outputs(2568)));
    outputs(5661) <= not((layer0_outputs(4074)) xor (layer0_outputs(8923)));
    outputs(5662) <= not(layer0_outputs(9594)) or (layer0_outputs(9433));
    outputs(5663) <= (layer0_outputs(4431)) xor (layer0_outputs(8841));
    outputs(5664) <= not(layer0_outputs(5298));
    outputs(5665) <= not((layer0_outputs(1850)) xor (layer0_outputs(3579)));
    outputs(5666) <= not(layer0_outputs(4907));
    outputs(5667) <= not((layer0_outputs(8290)) xor (layer0_outputs(9502)));
    outputs(5668) <= (layer0_outputs(921)) xor (layer0_outputs(4822));
    outputs(5669) <= (layer0_outputs(7891)) xor (layer0_outputs(8346));
    outputs(5670) <= (layer0_outputs(258)) or (layer0_outputs(6595));
    outputs(5671) <= layer0_outputs(6060);
    outputs(5672) <= not((layer0_outputs(2174)) xor (layer0_outputs(4292)));
    outputs(5673) <= not(layer0_outputs(5251)) or (layer0_outputs(3736));
    outputs(5674) <= not((layer0_outputs(7276)) xor (layer0_outputs(7292)));
    outputs(5675) <= not((layer0_outputs(8740)) xor (layer0_outputs(7470)));
    outputs(5676) <= not((layer0_outputs(7865)) xor (layer0_outputs(8625)));
    outputs(5677) <= not(layer0_outputs(7917));
    outputs(5678) <= layer0_outputs(6055);
    outputs(5679) <= layer0_outputs(2686);
    outputs(5680) <= (layer0_outputs(4327)) and not (layer0_outputs(4340));
    outputs(5681) <= layer0_outputs(311);
    outputs(5682) <= layer0_outputs(3001);
    outputs(5683) <= layer0_outputs(9104);
    outputs(5684) <= (layer0_outputs(8683)) xor (layer0_outputs(7250));
    outputs(5685) <= (layer0_outputs(5280)) xor (layer0_outputs(164));
    outputs(5686) <= layer0_outputs(5479);
    outputs(5687) <= not(layer0_outputs(9375));
    outputs(5688) <= (layer0_outputs(6214)) xor (layer0_outputs(9166));
    outputs(5689) <= not((layer0_outputs(7110)) xor (layer0_outputs(5736)));
    outputs(5690) <= not(layer0_outputs(7204));
    outputs(5691) <= (layer0_outputs(774)) or (layer0_outputs(8881));
    outputs(5692) <= not((layer0_outputs(3076)) xor (layer0_outputs(6472)));
    outputs(5693) <= not((layer0_outputs(3388)) xor (layer0_outputs(2546)));
    outputs(5694) <= layer0_outputs(7521);
    outputs(5695) <= not((layer0_outputs(6349)) or (layer0_outputs(8810)));
    outputs(5696) <= not((layer0_outputs(6808)) xor (layer0_outputs(1470)));
    outputs(5697) <= not((layer0_outputs(9317)) or (layer0_outputs(6894)));
    outputs(5698) <= (layer0_outputs(3795)) xor (layer0_outputs(108));
    outputs(5699) <= not((layer0_outputs(1361)) or (layer0_outputs(8927)));
    outputs(5700) <= layer0_outputs(5082);
    outputs(5701) <= (layer0_outputs(6876)) or (layer0_outputs(3236));
    outputs(5702) <= not((layer0_outputs(3990)) xor (layer0_outputs(4002)));
    outputs(5703) <= (layer0_outputs(1142)) xor (layer0_outputs(4732));
    outputs(5704) <= layer0_outputs(6264);
    outputs(5705) <= not((layer0_outputs(692)) and (layer0_outputs(9973)));
    outputs(5706) <= not(layer0_outputs(9065));
    outputs(5707) <= (layer0_outputs(671)) xor (layer0_outputs(3300));
    outputs(5708) <= (layer0_outputs(7802)) xor (layer0_outputs(1286));
    outputs(5709) <= not(layer0_outputs(4120));
    outputs(5710) <= layer0_outputs(7694);
    outputs(5711) <= not(layer0_outputs(881)) or (layer0_outputs(3651));
    outputs(5712) <= not(layer0_outputs(3979)) or (layer0_outputs(8745));
    outputs(5713) <= not((layer0_outputs(1097)) xor (layer0_outputs(3892)));
    outputs(5714) <= not(layer0_outputs(639));
    outputs(5715) <= layer0_outputs(1148);
    outputs(5716) <= layer0_outputs(9756);
    outputs(5717) <= layer0_outputs(6995);
    outputs(5718) <= not((layer0_outputs(4429)) or (layer0_outputs(6581)));
    outputs(5719) <= not(layer0_outputs(833));
    outputs(5720) <= layer0_outputs(4261);
    outputs(5721) <= (layer0_outputs(6272)) and (layer0_outputs(3342));
    outputs(5722) <= layer0_outputs(1854);
    outputs(5723) <= not((layer0_outputs(1331)) xor (layer0_outputs(8282)));
    outputs(5724) <= not((layer0_outputs(816)) xor (layer0_outputs(3042)));
    outputs(5725) <= (layer0_outputs(2922)) xor (layer0_outputs(6156));
    outputs(5726) <= (layer0_outputs(9703)) and not (layer0_outputs(4296));
    outputs(5727) <= layer0_outputs(2332);
    outputs(5728) <= not(layer0_outputs(2482)) or (layer0_outputs(1399));
    outputs(5729) <= (layer0_outputs(661)) or (layer0_outputs(8337));
    outputs(5730) <= not(layer0_outputs(3535));
    outputs(5731) <= (layer0_outputs(7988)) xor (layer0_outputs(5413));
    outputs(5732) <= not(layer0_outputs(9646)) or (layer0_outputs(7040));
    outputs(5733) <= not(layer0_outputs(5250));
    outputs(5734) <= not(layer0_outputs(2857)) or (layer0_outputs(1367));
    outputs(5735) <= layer0_outputs(8179);
    outputs(5736) <= not(layer0_outputs(8597));
    outputs(5737) <= layer0_outputs(5539);
    outputs(5738) <= (layer0_outputs(9878)) and (layer0_outputs(6236));
    outputs(5739) <= (layer0_outputs(2627)) and not (layer0_outputs(1280));
    outputs(5740) <= not(layer0_outputs(5437));
    outputs(5741) <= not((layer0_outputs(4152)) xor (layer0_outputs(5684)));
    outputs(5742) <= layer0_outputs(9080);
    outputs(5743) <= not((layer0_outputs(7018)) xor (layer0_outputs(5431)));
    outputs(5744) <= not(layer0_outputs(9461));
    outputs(5745) <= not((layer0_outputs(2943)) xor (layer0_outputs(2996)));
    outputs(5746) <= not((layer0_outputs(6350)) and (layer0_outputs(10142)));
    outputs(5747) <= (layer0_outputs(1248)) xor (layer0_outputs(1110));
    outputs(5748) <= (layer0_outputs(6742)) xor (layer0_outputs(1952));
    outputs(5749) <= (layer0_outputs(6375)) xor (layer0_outputs(4398));
    outputs(5750) <= (layer0_outputs(1646)) and not (layer0_outputs(9252));
    outputs(5751) <= (layer0_outputs(5380)) xor (layer0_outputs(8010));
    outputs(5752) <= not(layer0_outputs(165));
    outputs(5753) <= (layer0_outputs(746)) xor (layer0_outputs(3390));
    outputs(5754) <= (layer0_outputs(535)) xor (layer0_outputs(8845));
    outputs(5755) <= (layer0_outputs(1056)) xor (layer0_outputs(5808));
    outputs(5756) <= layer0_outputs(4688);
    outputs(5757) <= (layer0_outputs(1760)) and not (layer0_outputs(9905));
    outputs(5758) <= not((layer0_outputs(8319)) or (layer0_outputs(5100)));
    outputs(5759) <= not((layer0_outputs(3667)) xor (layer0_outputs(6801)));
    outputs(5760) <= (layer0_outputs(4322)) xor (layer0_outputs(7317));
    outputs(5761) <= (layer0_outputs(10112)) and not (layer0_outputs(8316));
    outputs(5762) <= not(layer0_outputs(3253)) or (layer0_outputs(6438));
    outputs(5763) <= not(layer0_outputs(2680));
    outputs(5764) <= not((layer0_outputs(130)) xor (layer0_outputs(1320)));
    outputs(5765) <= (layer0_outputs(2695)) xor (layer0_outputs(2356));
    outputs(5766) <= (layer0_outputs(9877)) xor (layer0_outputs(5301));
    outputs(5767) <= (layer0_outputs(8242)) xor (layer0_outputs(230));
    outputs(5768) <= not(layer0_outputs(5604));
    outputs(5769) <= layer0_outputs(6072);
    outputs(5770) <= not(layer0_outputs(2160));
    outputs(5771) <= (layer0_outputs(8200)) xor (layer0_outputs(4394));
    outputs(5772) <= not((layer0_outputs(4981)) xor (layer0_outputs(3993)));
    outputs(5773) <= not(layer0_outputs(9184));
    outputs(5774) <= not(layer0_outputs(3550));
    outputs(5775) <= not(layer0_outputs(78)) or (layer0_outputs(1364));
    outputs(5776) <= not(layer0_outputs(3397));
    outputs(5777) <= layer0_outputs(6343);
    outputs(5778) <= not((layer0_outputs(2841)) and (layer0_outputs(2781)));
    outputs(5779) <= not((layer0_outputs(2184)) and (layer0_outputs(6624)));
    outputs(5780) <= (layer0_outputs(7832)) xor (layer0_outputs(2929));
    outputs(5781) <= (layer0_outputs(4873)) xor (layer0_outputs(7457));
    outputs(5782) <= (layer0_outputs(8827)) xor (layer0_outputs(9913));
    outputs(5783) <= (layer0_outputs(4494)) or (layer0_outputs(9043));
    outputs(5784) <= not((layer0_outputs(2775)) xor (layer0_outputs(5826)));
    outputs(5785) <= layer0_outputs(9245);
    outputs(5786) <= not(layer0_outputs(2758));
    outputs(5787) <= (layer0_outputs(7559)) xor (layer0_outputs(976));
    outputs(5788) <= layer0_outputs(6486);
    outputs(5789) <= not((layer0_outputs(6106)) xor (layer0_outputs(9805)));
    outputs(5790) <= layer0_outputs(8939);
    outputs(5791) <= not(layer0_outputs(5442));
    outputs(5792) <= not(layer0_outputs(3595)) or (layer0_outputs(7742));
    outputs(5793) <= (layer0_outputs(4151)) xor (layer0_outputs(9640));
    outputs(5794) <= not((layer0_outputs(9373)) and (layer0_outputs(52)));
    outputs(5795) <= not((layer0_outputs(5316)) xor (layer0_outputs(6000)));
    outputs(5796) <= not((layer0_outputs(4326)) xor (layer0_outputs(1816)));
    outputs(5797) <= (layer0_outputs(7336)) xor (layer0_outputs(4683));
    outputs(5798) <= layer0_outputs(1514);
    outputs(5799) <= not((layer0_outputs(7)) or (layer0_outputs(7903)));
    outputs(5800) <= not(layer0_outputs(211));
    outputs(5801) <= (layer0_outputs(2416)) or (layer0_outputs(1087));
    outputs(5802) <= (layer0_outputs(255)) or (layer0_outputs(4364));
    outputs(5803) <= not(layer0_outputs(5616));
    outputs(5804) <= not((layer0_outputs(1822)) or (layer0_outputs(659)));
    outputs(5805) <= not(layer0_outputs(1601));
    outputs(5806) <= (layer0_outputs(4381)) xor (layer0_outputs(2080));
    outputs(5807) <= not(layer0_outputs(4050));
    outputs(5808) <= layer0_outputs(7232);
    outputs(5809) <= not(layer0_outputs(8385));
    outputs(5810) <= not(layer0_outputs(440));
    outputs(5811) <= (layer0_outputs(8570)) xor (layer0_outputs(6461));
    outputs(5812) <= not(layer0_outputs(6008));
    outputs(5813) <= not(layer0_outputs(4742));
    outputs(5814) <= layer0_outputs(5325);
    outputs(5815) <= layer0_outputs(2158);
    outputs(5816) <= (layer0_outputs(5564)) xor (layer0_outputs(1030));
    outputs(5817) <= not(layer0_outputs(5873)) or (layer0_outputs(6565));
    outputs(5818) <= not(layer0_outputs(7868)) or (layer0_outputs(51));
    outputs(5819) <= (layer0_outputs(8101)) xor (layer0_outputs(3809));
    outputs(5820) <= (layer0_outputs(9620)) or (layer0_outputs(4790));
    outputs(5821) <= (layer0_outputs(5384)) and (layer0_outputs(2924));
    outputs(5822) <= (layer0_outputs(6698)) xor (layer0_outputs(4427));
    outputs(5823) <= (layer0_outputs(8474)) and not (layer0_outputs(2189));
    outputs(5824) <= layer0_outputs(6184);
    outputs(5825) <= layer0_outputs(1955);
    outputs(5826) <= (layer0_outputs(8133)) xor (layer0_outputs(3177));
    outputs(5827) <= (layer0_outputs(6550)) xor (layer0_outputs(7584));
    outputs(5828) <= layer0_outputs(5556);
    outputs(5829) <= (layer0_outputs(1552)) or (layer0_outputs(5522));
    outputs(5830) <= layer0_outputs(9245);
    outputs(5831) <= not(layer0_outputs(5180));
    outputs(5832) <= (layer0_outputs(1131)) and not (layer0_outputs(190));
    outputs(5833) <= layer0_outputs(4463);
    outputs(5834) <= (layer0_outputs(7126)) or (layer0_outputs(1773));
    outputs(5835) <= not((layer0_outputs(5278)) or (layer0_outputs(2279)));
    outputs(5836) <= (layer0_outputs(7445)) xor (layer0_outputs(322));
    outputs(5837) <= layer0_outputs(3940);
    outputs(5838) <= (layer0_outputs(9064)) xor (layer0_outputs(2270));
    outputs(5839) <= (layer0_outputs(8125)) and (layer0_outputs(6122));
    outputs(5840) <= (layer0_outputs(3890)) or (layer0_outputs(5069));
    outputs(5841) <= not((layer0_outputs(10239)) xor (layer0_outputs(4620)));
    outputs(5842) <= not(layer0_outputs(4023));
    outputs(5843) <= (layer0_outputs(5147)) xor (layer0_outputs(6642));
    outputs(5844) <= (layer0_outputs(9210)) and not (layer0_outputs(3425));
    outputs(5845) <= not(layer0_outputs(1677));
    outputs(5846) <= not(layer0_outputs(4581));
    outputs(5847) <= not((layer0_outputs(4288)) xor (layer0_outputs(7554)));
    outputs(5848) <= not((layer0_outputs(1904)) xor (layer0_outputs(9242)));
    outputs(5849) <= not(layer0_outputs(7923));
    outputs(5850) <= not(layer0_outputs(8524));
    outputs(5851) <= not((layer0_outputs(9214)) and (layer0_outputs(1762)));
    outputs(5852) <= (layer0_outputs(3183)) and not (layer0_outputs(4034));
    outputs(5853) <= (layer0_outputs(3363)) xor (layer0_outputs(2021));
    outputs(5854) <= not(layer0_outputs(2162)) or (layer0_outputs(5517));
    outputs(5855) <= layer0_outputs(1342);
    outputs(5856) <= (layer0_outputs(8329)) or (layer0_outputs(1439));
    outputs(5857) <= layer0_outputs(4367);
    outputs(5858) <= not(layer0_outputs(5365));
    outputs(5859) <= layer0_outputs(3439);
    outputs(5860) <= not(layer0_outputs(791));
    outputs(5861) <= not(layer0_outputs(13));
    outputs(5862) <= not((layer0_outputs(2588)) xor (layer0_outputs(1352)));
    outputs(5863) <= (layer0_outputs(2235)) xor (layer0_outputs(1310));
    outputs(5864) <= (layer0_outputs(9939)) xor (layer0_outputs(2256));
    outputs(5865) <= not(layer0_outputs(7115)) or (layer0_outputs(3423));
    outputs(5866) <= not((layer0_outputs(3616)) xor (layer0_outputs(9099)));
    outputs(5867) <= not(layer0_outputs(1541));
    outputs(5868) <= not(layer0_outputs(2490)) or (layer0_outputs(695));
    outputs(5869) <= (layer0_outputs(8305)) and not (layer0_outputs(9037));
    outputs(5870) <= not(layer0_outputs(4718));
    outputs(5871) <= not(layer0_outputs(8195));
    outputs(5872) <= not((layer0_outputs(2905)) and (layer0_outputs(9714)));
    outputs(5873) <= (layer0_outputs(9193)) xor (layer0_outputs(6785));
    outputs(5874) <= layer0_outputs(2116);
    outputs(5875) <= not((layer0_outputs(974)) xor (layer0_outputs(5794)));
    outputs(5876) <= not((layer0_outputs(505)) xor (layer0_outputs(5667)));
    outputs(5877) <= layer0_outputs(9044);
    outputs(5878) <= not(layer0_outputs(2064));
    outputs(5879) <= not(layer0_outputs(9006));
    outputs(5880) <= (layer0_outputs(1202)) or (layer0_outputs(10217));
    outputs(5881) <= not(layer0_outputs(2584));
    outputs(5882) <= (layer0_outputs(8962)) and not (layer0_outputs(1937));
    outputs(5883) <= not((layer0_outputs(7682)) xor (layer0_outputs(3517)));
    outputs(5884) <= (layer0_outputs(243)) xor (layer0_outputs(1088));
    outputs(5885) <= not((layer0_outputs(1211)) xor (layer0_outputs(1508)));
    outputs(5886) <= (layer0_outputs(2487)) or (layer0_outputs(2085));
    outputs(5887) <= not(layer0_outputs(2037));
    outputs(5888) <= layer0_outputs(4234);
    outputs(5889) <= not((layer0_outputs(2043)) xor (layer0_outputs(4603)));
    outputs(5890) <= not((layer0_outputs(10198)) xor (layer0_outputs(4349)));
    outputs(5891) <= layer0_outputs(5306);
    outputs(5892) <= (layer0_outputs(2411)) or (layer0_outputs(5821));
    outputs(5893) <= not(layer0_outputs(5705));
    outputs(5894) <= (layer0_outputs(8612)) xor (layer0_outputs(3046));
    outputs(5895) <= not(layer0_outputs(2039));
    outputs(5896) <= (layer0_outputs(9332)) xor (layer0_outputs(1711));
    outputs(5897) <= not(layer0_outputs(2488)) or (layer0_outputs(8832));
    outputs(5898) <= not(layer0_outputs(5735));
    outputs(5899) <= not(layer0_outputs(7846)) or (layer0_outputs(2224));
    outputs(5900) <= not(layer0_outputs(8163)) or (layer0_outputs(1499));
    outputs(5901) <= layer0_outputs(10227);
    outputs(5902) <= not(layer0_outputs(7023));
    outputs(5903) <= not(layer0_outputs(8912));
    outputs(5904) <= (layer0_outputs(4408)) and (layer0_outputs(8141));
    outputs(5905) <= (layer0_outputs(2563)) and not (layer0_outputs(6944));
    outputs(5906) <= not((layer0_outputs(10133)) and (layer0_outputs(5243)));
    outputs(5907) <= layer0_outputs(4696);
    outputs(5908) <= not((layer0_outputs(7920)) xor (layer0_outputs(9496)));
    outputs(5909) <= not(layer0_outputs(9770));
    outputs(5910) <= not((layer0_outputs(1359)) and (layer0_outputs(7915)));
    outputs(5911) <= not((layer0_outputs(7146)) xor (layer0_outputs(10030)));
    outputs(5912) <= not(layer0_outputs(1141));
    outputs(5913) <= not(layer0_outputs(9051)) or (layer0_outputs(2714));
    outputs(5914) <= not((layer0_outputs(6228)) xor (layer0_outputs(762)));
    outputs(5915) <= (layer0_outputs(3447)) xor (layer0_outputs(6054));
    outputs(5916) <= not((layer0_outputs(8065)) and (layer0_outputs(10121)));
    outputs(5917) <= (layer0_outputs(10009)) xor (layer0_outputs(5800));
    outputs(5918) <= (layer0_outputs(8950)) xor (layer0_outputs(2787));
    outputs(5919) <= layer0_outputs(7835);
    outputs(5920) <= not((layer0_outputs(4929)) xor (layer0_outputs(7670)));
    outputs(5921) <= (layer0_outputs(2900)) and (layer0_outputs(3789));
    outputs(5922) <= not((layer0_outputs(3755)) xor (layer0_outputs(9447)));
    outputs(5923) <= not((layer0_outputs(6258)) xor (layer0_outputs(9811)));
    outputs(5924) <= not((layer0_outputs(7113)) xor (layer0_outputs(6829)));
    outputs(5925) <= layer0_outputs(5420);
    outputs(5926) <= (layer0_outputs(7039)) xor (layer0_outputs(3009));
    outputs(5927) <= not((layer0_outputs(242)) or (layer0_outputs(2107)));
    outputs(5928) <= not(layer0_outputs(2495));
    outputs(5929) <= not((layer0_outputs(2067)) xor (layer0_outputs(2199)));
    outputs(5930) <= (layer0_outputs(1984)) and (layer0_outputs(8087));
    outputs(5931) <= layer0_outputs(4987);
    outputs(5932) <= layer0_outputs(7615);
    outputs(5933) <= not(layer0_outputs(4666));
    outputs(5934) <= (layer0_outputs(5448)) xor (layer0_outputs(351));
    outputs(5935) <= not(layer0_outputs(10033));
    outputs(5936) <= not((layer0_outputs(2484)) xor (layer0_outputs(1945)));
    outputs(5937) <= (layer0_outputs(6461)) or (layer0_outputs(1051));
    outputs(5938) <= (layer0_outputs(2182)) xor (layer0_outputs(3978));
    outputs(5939) <= (layer0_outputs(7788)) xor (layer0_outputs(8589));
    outputs(5940) <= layer0_outputs(9478);
    outputs(5941) <= (layer0_outputs(6564)) xor (layer0_outputs(185));
    outputs(5942) <= layer0_outputs(9414);
    outputs(5943) <= layer0_outputs(4495);
    outputs(5944) <= layer0_outputs(3419);
    outputs(5945) <= (layer0_outputs(7847)) and not (layer0_outputs(2579));
    outputs(5946) <= not((layer0_outputs(7218)) xor (layer0_outputs(6725)));
    outputs(5947) <= not((layer0_outputs(5619)) xor (layer0_outputs(9050)));
    outputs(5948) <= not(layer0_outputs(8214));
    outputs(5949) <= layer0_outputs(237);
    outputs(5950) <= not((layer0_outputs(7728)) xor (layer0_outputs(7824)));
    outputs(5951) <= not((layer0_outputs(9159)) xor (layer0_outputs(3184)));
    outputs(5952) <= (layer0_outputs(30)) xor (layer0_outputs(4851));
    outputs(5953) <= not(layer0_outputs(10052));
    outputs(5954) <= not(layer0_outputs(9217));
    outputs(5955) <= not(layer0_outputs(2010));
    outputs(5956) <= not(layer0_outputs(1129)) or (layer0_outputs(6715));
    outputs(5957) <= not(layer0_outputs(1853));
    outputs(5958) <= (layer0_outputs(4064)) xor (layer0_outputs(8844));
    outputs(5959) <= not(layer0_outputs(9585));
    outputs(5960) <= not((layer0_outputs(5276)) xor (layer0_outputs(3990)));
    outputs(5961) <= (layer0_outputs(9584)) xor (layer0_outputs(5042));
    outputs(5962) <= layer0_outputs(6112);
    outputs(5963) <= not(layer0_outputs(5580));
    outputs(5964) <= not(layer0_outputs(6080)) or (layer0_outputs(2639));
    outputs(5965) <= layer0_outputs(6804);
    outputs(5966) <= (layer0_outputs(7637)) and not (layer0_outputs(9775));
    outputs(5967) <= layer0_outputs(2444);
    outputs(5968) <= not(layer0_outputs(3799)) or (layer0_outputs(3970));
    outputs(5969) <= not((layer0_outputs(5692)) xor (layer0_outputs(4998)));
    outputs(5970) <= (layer0_outputs(9150)) and (layer0_outputs(6307));
    outputs(5971) <= not((layer0_outputs(7185)) xor (layer0_outputs(6213)));
    outputs(5972) <= (layer0_outputs(8640)) xor (layer0_outputs(6322));
    outputs(5973) <= (layer0_outputs(962)) xor (layer0_outputs(4959));
    outputs(5974) <= not(layer0_outputs(1790)) or (layer0_outputs(961));
    outputs(5975) <= not((layer0_outputs(8639)) xor (layer0_outputs(511)));
    outputs(5976) <= (layer0_outputs(3974)) and not (layer0_outputs(4095));
    outputs(5977) <= layer0_outputs(3500);
    outputs(5978) <= (layer0_outputs(350)) and not (layer0_outputs(701));
    outputs(5979) <= layer0_outputs(880);
    outputs(5980) <= (layer0_outputs(4725)) xor (layer0_outputs(5325));
    outputs(5981) <= not((layer0_outputs(6095)) xor (layer0_outputs(5972)));
    outputs(5982) <= layer0_outputs(631);
    outputs(5983) <= not((layer0_outputs(2419)) xor (layer0_outputs(1836)));
    outputs(5984) <= not(layer0_outputs(3407)) or (layer0_outputs(10202));
    outputs(5985) <= not((layer0_outputs(6673)) xor (layer0_outputs(4482)));
    outputs(5986) <= layer0_outputs(7887);
    outputs(5987) <= not((layer0_outputs(9018)) xor (layer0_outputs(430)));
    outputs(5988) <= not((layer0_outputs(3504)) and (layer0_outputs(6671)));
    outputs(5989) <= (layer0_outputs(5643)) xor (layer0_outputs(396));
    outputs(5990) <= (layer0_outputs(2009)) xor (layer0_outputs(331));
    outputs(5991) <= (layer0_outputs(5768)) xor (layer0_outputs(1255));
    outputs(5992) <= layer0_outputs(2971);
    outputs(5993) <= not((layer0_outputs(3535)) or (layer0_outputs(2340)));
    outputs(5994) <= not(layer0_outputs(4251));
    outputs(5995) <= (layer0_outputs(9459)) xor (layer0_outputs(8293));
    outputs(5996) <= not((layer0_outputs(8967)) xor (layer0_outputs(8234)));
    outputs(5997) <= not(layer0_outputs(8148));
    outputs(5998) <= layer0_outputs(654);
    outputs(5999) <= (layer0_outputs(8484)) or (layer0_outputs(5374));
    outputs(6000) <= layer0_outputs(2034);
    outputs(6001) <= not(layer0_outputs(3292));
    outputs(6002) <= (layer0_outputs(9999)) and not (layer0_outputs(1924));
    outputs(6003) <= not((layer0_outputs(4476)) xor (layer0_outputs(3117)));
    outputs(6004) <= (layer0_outputs(10113)) and (layer0_outputs(9213));
    outputs(6005) <= not(layer0_outputs(6440));
    outputs(6006) <= not((layer0_outputs(9843)) xor (layer0_outputs(1953)));
    outputs(6007) <= not((layer0_outputs(3858)) xor (layer0_outputs(8013)));
    outputs(6008) <= not(layer0_outputs(8324)) or (layer0_outputs(6136));
    outputs(6009) <= not((layer0_outputs(1919)) xor (layer0_outputs(5510)));
    outputs(6010) <= not(layer0_outputs(8528)) or (layer0_outputs(3008));
    outputs(6011) <= not(layer0_outputs(293));
    outputs(6012) <= (layer0_outputs(3510)) xor (layer0_outputs(4738));
    outputs(6013) <= not((layer0_outputs(6093)) xor (layer0_outputs(1571)));
    outputs(6014) <= not(layer0_outputs(6634));
    outputs(6015) <= not(layer0_outputs(3548));
    outputs(6016) <= layer0_outputs(9399);
    outputs(6017) <= (layer0_outputs(3806)) xor (layer0_outputs(6641));
    outputs(6018) <= layer0_outputs(10018);
    outputs(6019) <= (layer0_outputs(772)) xor (layer0_outputs(3588));
    outputs(6020) <= layer0_outputs(6190);
    outputs(6021) <= layer0_outputs(8488);
    outputs(6022) <= layer0_outputs(6897);
    outputs(6023) <= not((layer0_outputs(1043)) xor (layer0_outputs(5540)));
    outputs(6024) <= not(layer0_outputs(8112));
    outputs(6025) <= (layer0_outputs(4505)) and not (layer0_outputs(1289));
    outputs(6026) <= not(layer0_outputs(3422)) or (layer0_outputs(6618));
    outputs(6027) <= not((layer0_outputs(3033)) xor (layer0_outputs(4690)));
    outputs(6028) <= (layer0_outputs(3566)) xor (layer0_outputs(9794));
    outputs(6029) <= layer0_outputs(1419);
    outputs(6030) <= not((layer0_outputs(3747)) and (layer0_outputs(397)));
    outputs(6031) <= not(layer0_outputs(8802)) or (layer0_outputs(95));
    outputs(6032) <= (layer0_outputs(4689)) and not (layer0_outputs(1626));
    outputs(6033) <= (layer0_outputs(7948)) and not (layer0_outputs(6462));
    outputs(6034) <= layer0_outputs(2207);
    outputs(6035) <= (layer0_outputs(9783)) or (layer0_outputs(2041));
    outputs(6036) <= (layer0_outputs(2165)) xor (layer0_outputs(8201));
    outputs(6037) <= not(layer0_outputs(8572)) or (layer0_outputs(6101));
    outputs(6038) <= (layer0_outputs(3233)) xor (layer0_outputs(10216));
    outputs(6039) <= layer0_outputs(5964);
    outputs(6040) <= (layer0_outputs(3822)) xor (layer0_outputs(180));
    outputs(6041) <= (layer0_outputs(9963)) and not (layer0_outputs(9164));
    outputs(6042) <= layer0_outputs(7842);
    outputs(6043) <= (layer0_outputs(10064)) xor (layer0_outputs(8966));
    outputs(6044) <= layer0_outputs(7928);
    outputs(6045) <= not((layer0_outputs(4800)) or (layer0_outputs(1586)));
    outputs(6046) <= not(layer0_outputs(7893));
    outputs(6047) <= (layer0_outputs(6360)) and (layer0_outputs(1816));
    outputs(6048) <= not(layer0_outputs(2586));
    outputs(6049) <= not((layer0_outputs(7897)) xor (layer0_outputs(513)));
    outputs(6050) <= (layer0_outputs(9288)) and not (layer0_outputs(3111));
    outputs(6051) <= layer0_outputs(10061);
    outputs(6052) <= not(layer0_outputs(4536));
    outputs(6053) <= not(layer0_outputs(79)) or (layer0_outputs(1910));
    outputs(6054) <= not((layer0_outputs(8750)) xor (layer0_outputs(6836)));
    outputs(6055) <= not((layer0_outputs(2990)) xor (layer0_outputs(1931)));
    outputs(6056) <= not(layer0_outputs(5600));
    outputs(6057) <= not(layer0_outputs(6549));
    outputs(6058) <= not((layer0_outputs(8907)) xor (layer0_outputs(2263)));
    outputs(6059) <= layer0_outputs(2819);
    outputs(6060) <= layer0_outputs(3472);
    outputs(6061) <= layer0_outputs(3831);
    outputs(6062) <= not(layer0_outputs(5054));
    outputs(6063) <= layer0_outputs(7521);
    outputs(6064) <= (layer0_outputs(3266)) and not (layer0_outputs(3822));
    outputs(6065) <= not(layer0_outputs(2226));
    outputs(6066) <= not((layer0_outputs(510)) xor (layer0_outputs(20)));
    outputs(6067) <= layer0_outputs(7515);
    outputs(6068) <= not((layer0_outputs(3512)) xor (layer0_outputs(4951)));
    outputs(6069) <= (layer0_outputs(4153)) and (layer0_outputs(3630));
    outputs(6070) <= not(layer0_outputs(8525));
    outputs(6071) <= layer0_outputs(4626);
    outputs(6072) <= not(layer0_outputs(3958));
    outputs(6073) <= not(layer0_outputs(8965));
    outputs(6074) <= layer0_outputs(4697);
    outputs(6075) <= (layer0_outputs(9287)) xor (layer0_outputs(2520));
    outputs(6076) <= not((layer0_outputs(268)) xor (layer0_outputs(7327)));
    outputs(6077) <= (layer0_outputs(93)) and (layer0_outputs(1051));
    outputs(6078) <= not((layer0_outputs(1242)) xor (layer0_outputs(4521)));
    outputs(6079) <= not(layer0_outputs(6043)) or (layer0_outputs(5313));
    outputs(6080) <= not(layer0_outputs(1875));
    outputs(6081) <= not(layer0_outputs(3681));
    outputs(6082) <= (layer0_outputs(2684)) and not (layer0_outputs(6115));
    outputs(6083) <= layer0_outputs(4348);
    outputs(6084) <= not((layer0_outputs(3321)) xor (layer0_outputs(4410)));
    outputs(6085) <= layer0_outputs(4374);
    outputs(6086) <= layer0_outputs(7678);
    outputs(6087) <= (layer0_outputs(5197)) and (layer0_outputs(5090));
    outputs(6088) <= (layer0_outputs(3176)) xor (layer0_outputs(5304));
    outputs(6089) <= not((layer0_outputs(745)) xor (layer0_outputs(4896)));
    outputs(6090) <= not((layer0_outputs(5562)) xor (layer0_outputs(1543)));
    outputs(6091) <= not(layer0_outputs(6812));
    outputs(6092) <= (layer0_outputs(9741)) xor (layer0_outputs(6262));
    outputs(6093) <= not((layer0_outputs(1703)) xor (layer0_outputs(3961)));
    outputs(6094) <= layer0_outputs(5145);
    outputs(6095) <= (layer0_outputs(1132)) xor (layer0_outputs(1899));
    outputs(6096) <= not((layer0_outputs(6085)) xor (layer0_outputs(2516)));
    outputs(6097) <= not((layer0_outputs(1923)) xor (layer0_outputs(9479)));
    outputs(6098) <= not(layer0_outputs(177)) or (layer0_outputs(2615));
    outputs(6099) <= not((layer0_outputs(3035)) xor (layer0_outputs(10230)));
    outputs(6100) <= (layer0_outputs(6286)) and not (layer0_outputs(2348));
    outputs(6101) <= (layer0_outputs(9177)) and not (layer0_outputs(5968));
    outputs(6102) <= not((layer0_outputs(2092)) xor (layer0_outputs(10114)));
    outputs(6103) <= not(layer0_outputs(2281));
    outputs(6104) <= not(layer0_outputs(1353));
    outputs(6105) <= (layer0_outputs(5089)) and not (layer0_outputs(2354));
    outputs(6106) <= (layer0_outputs(2809)) xor (layer0_outputs(2339));
    outputs(6107) <= not(layer0_outputs(5490)) or (layer0_outputs(8992));
    outputs(6108) <= not(layer0_outputs(5293));
    outputs(6109) <= (layer0_outputs(2079)) xor (layer0_outputs(9751));
    outputs(6110) <= layer0_outputs(9481);
    outputs(6111) <= (layer0_outputs(5657)) xor (layer0_outputs(2425));
    outputs(6112) <= (layer0_outputs(693)) or (layer0_outputs(7561));
    outputs(6113) <= not(layer0_outputs(1407));
    outputs(6114) <= (layer0_outputs(4648)) xor (layer0_outputs(7939));
    outputs(6115) <= (layer0_outputs(8602)) xor (layer0_outputs(2153));
    outputs(6116) <= not((layer0_outputs(8686)) and (layer0_outputs(2933)));
    outputs(6117) <= not(layer0_outputs(3088));
    outputs(6118) <= not(layer0_outputs(1361));
    outputs(6119) <= layer0_outputs(3554);
    outputs(6120) <= layer0_outputs(9737);
    outputs(6121) <= layer0_outputs(8563);
    outputs(6122) <= not(layer0_outputs(8203));
    outputs(6123) <= layer0_outputs(6719);
    outputs(6124) <= not(layer0_outputs(3333)) or (layer0_outputs(5327));
    outputs(6125) <= (layer0_outputs(9762)) xor (layer0_outputs(6834));
    outputs(6126) <= (layer0_outputs(2578)) or (layer0_outputs(45));
    outputs(6127) <= not((layer0_outputs(6604)) or (layer0_outputs(3792)));
    outputs(6128) <= not(layer0_outputs(2837));
    outputs(6129) <= not((layer0_outputs(1467)) xor (layer0_outputs(4888)));
    outputs(6130) <= not((layer0_outputs(544)) xor (layer0_outputs(2448)));
    outputs(6131) <= not((layer0_outputs(6560)) and (layer0_outputs(9525)));
    outputs(6132) <= not((layer0_outputs(8888)) xor (layer0_outputs(8048)));
    outputs(6133) <= not(layer0_outputs(9641));
    outputs(6134) <= (layer0_outputs(9837)) xor (layer0_outputs(10197));
    outputs(6135) <= layer0_outputs(5917);
    outputs(6136) <= (layer0_outputs(3626)) or (layer0_outputs(3208));
    outputs(6137) <= layer0_outputs(4183);
    outputs(6138) <= not(layer0_outputs(5820));
    outputs(6139) <= not((layer0_outputs(5732)) or (layer0_outputs(9827)));
    outputs(6140) <= not(layer0_outputs(3235));
    outputs(6141) <= (layer0_outputs(2280)) xor (layer0_outputs(4114));
    outputs(6142) <= (layer0_outputs(8)) xor (layer0_outputs(9911));
    outputs(6143) <= (layer0_outputs(9738)) xor (layer0_outputs(5310));
    outputs(6144) <= layer0_outputs(7858);
    outputs(6145) <= (layer0_outputs(9425)) xor (layer0_outputs(4529));
    outputs(6146) <= not(layer0_outputs(9019));
    outputs(6147) <= (layer0_outputs(2133)) and not (layer0_outputs(8969));
    outputs(6148) <= (layer0_outputs(8557)) or (layer0_outputs(1918));
    outputs(6149) <= (layer0_outputs(4511)) and (layer0_outputs(8150));
    outputs(6150) <= not(layer0_outputs(184)) or (layer0_outputs(5323));
    outputs(6151) <= (layer0_outputs(3077)) and not (layer0_outputs(8906));
    outputs(6152) <= not(layer0_outputs(6934));
    outputs(6153) <= layer0_outputs(669);
    outputs(6154) <= not((layer0_outputs(9696)) and (layer0_outputs(9705)));
    outputs(6155) <= not(layer0_outputs(6506));
    outputs(6156) <= layer0_outputs(1308);
    outputs(6157) <= layer0_outputs(1496);
    outputs(6158) <= not(layer0_outputs(3641));
    outputs(6159) <= not(layer0_outputs(6966));
    outputs(6160) <= layer0_outputs(9416);
    outputs(6161) <= not(layer0_outputs(4676));
    outputs(6162) <= (layer0_outputs(7610)) and not (layer0_outputs(3296));
    outputs(6163) <= not(layer0_outputs(8442));
    outputs(6164) <= not((layer0_outputs(9534)) or (layer0_outputs(4041)));
    outputs(6165) <= (layer0_outputs(579)) xor (layer0_outputs(9113));
    outputs(6166) <= (layer0_outputs(3194)) and (layer0_outputs(3950));
    outputs(6167) <= layer0_outputs(4140);
    outputs(6168) <= not(layer0_outputs(8394));
    outputs(6169) <= layer0_outputs(3832);
    outputs(6170) <= layer0_outputs(4182);
    outputs(6171) <= not(layer0_outputs(793));
    outputs(6172) <= layer0_outputs(7398);
    outputs(6173) <= not((layer0_outputs(9200)) xor (layer0_outputs(2910)));
    outputs(6174) <= not(layer0_outputs(2326));
    outputs(6175) <= not(layer0_outputs(1687));
    outputs(6176) <= layer0_outputs(1480);
    outputs(6177) <= (layer0_outputs(8469)) and (layer0_outputs(2556));
    outputs(6178) <= not(layer0_outputs(3478));
    outputs(6179) <= not(layer0_outputs(3185));
    outputs(6180) <= (layer0_outputs(7386)) and (layer0_outputs(3481));
    outputs(6181) <= (layer0_outputs(167)) and not (layer0_outputs(7164));
    outputs(6182) <= not(layer0_outputs(3234));
    outputs(6183) <= not(layer0_outputs(1389)) or (layer0_outputs(9286));
    outputs(6184) <= layer0_outputs(8259);
    outputs(6185) <= not(layer0_outputs(4945));
    outputs(6186) <= not((layer0_outputs(1568)) xor (layer0_outputs(9400)));
    outputs(6187) <= (layer0_outputs(8528)) xor (layer0_outputs(2283));
    outputs(6188) <= layer0_outputs(1584);
    outputs(6189) <= not(layer0_outputs(4184));
    outputs(6190) <= (layer0_outputs(2640)) and not (layer0_outputs(3759));
    outputs(6191) <= layer0_outputs(2780);
    outputs(6192) <= layer0_outputs(8395);
    outputs(6193) <= layer0_outputs(1083);
    outputs(6194) <= (layer0_outputs(430)) xor (layer0_outputs(6319));
    outputs(6195) <= layer0_outputs(4846);
    outputs(6196) <= (layer0_outputs(1095)) and not (layer0_outputs(7192));
    outputs(6197) <= not((layer0_outputs(947)) and (layer0_outputs(2366)));
    outputs(6198) <= not((layer0_outputs(6534)) or (layer0_outputs(4470)));
    outputs(6199) <= not(layer0_outputs(562));
    outputs(6200) <= layer0_outputs(6884);
    outputs(6201) <= not((layer0_outputs(3555)) or (layer0_outputs(5616)));
    outputs(6202) <= layer0_outputs(32);
    outputs(6203) <= (layer0_outputs(4438)) or (layer0_outputs(59));
    outputs(6204) <= (layer0_outputs(8432)) and not (layer0_outputs(7924));
    outputs(6205) <= layer0_outputs(40);
    outputs(6206) <= (layer0_outputs(6393)) and (layer0_outputs(2821));
    outputs(6207) <= not(layer0_outputs(2786)) or (layer0_outputs(10073));
    outputs(6208) <= (layer0_outputs(3181)) and not (layer0_outputs(7742));
    outputs(6209) <= (layer0_outputs(7041)) and not (layer0_outputs(9075));
    outputs(6210) <= (layer0_outputs(3794)) and not (layer0_outputs(8838));
    outputs(6211) <= (layer0_outputs(2269)) or (layer0_outputs(1942));
    outputs(6212) <= (layer0_outputs(5767)) xor (layer0_outputs(658));
    outputs(6213) <= layer0_outputs(9813);
    outputs(6214) <= (layer0_outputs(1530)) and not (layer0_outputs(8101));
    outputs(6215) <= not(layer0_outputs(5633));
    outputs(6216) <= not(layer0_outputs(8087));
    outputs(6217) <= (layer0_outputs(6621)) and (layer0_outputs(9962));
    outputs(6218) <= layer0_outputs(4283);
    outputs(6219) <= not(layer0_outputs(5157));
    outputs(6220) <= not(layer0_outputs(6082));
    outputs(6221) <= layer0_outputs(6879);
    outputs(6222) <= layer0_outputs(7577);
    outputs(6223) <= layer0_outputs(6050);
    outputs(6224) <= layer0_outputs(289);
    outputs(6225) <= (layer0_outputs(9668)) and not (layer0_outputs(6276));
    outputs(6226) <= (layer0_outputs(1614)) and not (layer0_outputs(6147));
    outputs(6227) <= not((layer0_outputs(7785)) or (layer0_outputs(4955)));
    outputs(6228) <= not((layer0_outputs(6930)) or (layer0_outputs(4827)));
    outputs(6229) <= (layer0_outputs(7878)) and (layer0_outputs(1049));
    outputs(6230) <= not(layer0_outputs(4146));
    outputs(6231) <= (layer0_outputs(7830)) xor (layer0_outputs(2774));
    outputs(6232) <= not(layer0_outputs(3514));
    outputs(6233) <= layer0_outputs(7181);
    outputs(6234) <= layer0_outputs(671);
    outputs(6235) <= (layer0_outputs(5670)) and (layer0_outputs(1121));
    outputs(6236) <= not((layer0_outputs(6711)) and (layer0_outputs(1233)));
    outputs(6237) <= not(layer0_outputs(9993)) or (layer0_outputs(256));
    outputs(6238) <= (layer0_outputs(7435)) and not (layer0_outputs(2843));
    outputs(6239) <= not((layer0_outputs(589)) or (layer0_outputs(3399)));
    outputs(6240) <= not(layer0_outputs(2450)) or (layer0_outputs(7204));
    outputs(6241) <= layer0_outputs(7122);
    outputs(6242) <= layer0_outputs(9327);
    outputs(6243) <= (layer0_outputs(5360)) xor (layer0_outputs(1269));
    outputs(6244) <= not(layer0_outputs(2027)) or (layer0_outputs(4631));
    outputs(6245) <= layer0_outputs(459);
    outputs(6246) <= not(layer0_outputs(1179));
    outputs(6247) <= (layer0_outputs(127)) and (layer0_outputs(4624));
    outputs(6248) <= not(layer0_outputs(2284));
    outputs(6249) <= (layer0_outputs(1473)) and not (layer0_outputs(7642));
    outputs(6250) <= (layer0_outputs(3150)) and (layer0_outputs(2252));
    outputs(6251) <= not(layer0_outputs(4024));
    outputs(6252) <= (layer0_outputs(708)) and not (layer0_outputs(9415));
    outputs(6253) <= layer0_outputs(5056);
    outputs(6254) <= not((layer0_outputs(5815)) xor (layer0_outputs(6662)));
    outputs(6255) <= not((layer0_outputs(6267)) xor (layer0_outputs(4538)));
    outputs(6256) <= not(layer0_outputs(664));
    outputs(6257) <= not((layer0_outputs(7400)) xor (layer0_outputs(7486)));
    outputs(6258) <= not(layer0_outputs(2331));
    outputs(6259) <= (layer0_outputs(3079)) and (layer0_outputs(6369));
    outputs(6260) <= not(layer0_outputs(9635));
    outputs(6261) <= layer0_outputs(6312);
    outputs(6262) <= not(layer0_outputs(2671));
    outputs(6263) <= not(layer0_outputs(3604));
    outputs(6264) <= layer0_outputs(4362);
    outputs(6265) <= layer0_outputs(8151);
    outputs(6266) <= (layer0_outputs(2705)) or (layer0_outputs(9085));
    outputs(6267) <= not(layer0_outputs(6500));
    outputs(6268) <= not(layer0_outputs(811)) or (layer0_outputs(50));
    outputs(6269) <= (layer0_outputs(3545)) and not (layer0_outputs(9207));
    outputs(6270) <= (layer0_outputs(5395)) and not (layer0_outputs(3058));
    outputs(6271) <= not(layer0_outputs(8532));
    outputs(6272) <= (layer0_outputs(9553)) and not (layer0_outputs(5947));
    outputs(6273) <= (layer0_outputs(2839)) and not (layer0_outputs(5005));
    outputs(6274) <= not(layer0_outputs(4618));
    outputs(6275) <= not((layer0_outputs(10148)) and (layer0_outputs(3910)));
    outputs(6276) <= not(layer0_outputs(4856));
    outputs(6277) <= not(layer0_outputs(1759));
    outputs(6278) <= layer0_outputs(5099);
    outputs(6279) <= not(layer0_outputs(7638));
    outputs(6280) <= not(layer0_outputs(3655));
    outputs(6281) <= not((layer0_outputs(3755)) xor (layer0_outputs(1040)));
    outputs(6282) <= (layer0_outputs(3868)) or (layer0_outputs(4440));
    outputs(6283) <= not(layer0_outputs(7712)) or (layer0_outputs(9719));
    outputs(6284) <= (layer0_outputs(1451)) and (layer0_outputs(9991));
    outputs(6285) <= layer0_outputs(1300);
    outputs(6286) <= not((layer0_outputs(8423)) xor (layer0_outputs(1883)));
    outputs(6287) <= (layer0_outputs(7343)) xor (layer0_outputs(9248));
    outputs(6288) <= not(layer0_outputs(3370)) or (layer0_outputs(3816));
    outputs(6289) <= not(layer0_outputs(461));
    outputs(6290) <= layer0_outputs(9198);
    outputs(6291) <= not((layer0_outputs(7351)) or (layer0_outputs(4215)));
    outputs(6292) <= not(layer0_outputs(6794));
    outputs(6293) <= layer0_outputs(3750);
    outputs(6294) <= (layer0_outputs(134)) and (layer0_outputs(9242));
    outputs(6295) <= (layer0_outputs(1348)) xor (layer0_outputs(2897));
    outputs(6296) <= (layer0_outputs(519)) and not (layer0_outputs(8344));
    outputs(6297) <= not(layer0_outputs(7421));
    outputs(6298) <= not(layer0_outputs(8460)) or (layer0_outputs(133));
    outputs(6299) <= not(layer0_outputs(8816));
    outputs(6300) <= not(layer0_outputs(2928)) or (layer0_outputs(6114));
    outputs(6301) <= not(layer0_outputs(2255));
    outputs(6302) <= layer0_outputs(4537);
    outputs(6303) <= not(layer0_outputs(6997));
    outputs(6304) <= (layer0_outputs(7664)) xor (layer0_outputs(5014));
    outputs(6305) <= (layer0_outputs(1615)) and (layer0_outputs(2932));
    outputs(6306) <= layer0_outputs(5899);
    outputs(6307) <= (layer0_outputs(5939)) xor (layer0_outputs(7775));
    outputs(6308) <= not((layer0_outputs(8916)) or (layer0_outputs(7030)));
    outputs(6309) <= not(layer0_outputs(1006));
    outputs(6310) <= not((layer0_outputs(6416)) xor (layer0_outputs(1341)));
    outputs(6311) <= layer0_outputs(3028);
    outputs(6312) <= (layer0_outputs(5310)) and not (layer0_outputs(2779));
    outputs(6313) <= (layer0_outputs(2338)) or (layer0_outputs(6978));
    outputs(6314) <= layer0_outputs(5048);
    outputs(6315) <= not(layer0_outputs(6243));
    outputs(6316) <= (layer0_outputs(1828)) xor (layer0_outputs(7021));
    outputs(6317) <= not((layer0_outputs(3182)) and (layer0_outputs(6529)));
    outputs(6318) <= layer0_outputs(7601);
    outputs(6319) <= layer0_outputs(8835);
    outputs(6320) <= not(layer0_outputs(2083));
    outputs(6321) <= (layer0_outputs(3307)) and (layer0_outputs(9032));
    outputs(6322) <= not(layer0_outputs(4027)) or (layer0_outputs(484));
    outputs(6323) <= layer0_outputs(3452);
    outputs(6324) <= (layer0_outputs(4733)) and not (layer0_outputs(1743));
    outputs(6325) <= not(layer0_outputs(1728)) or (layer0_outputs(572));
    outputs(6326) <= not(layer0_outputs(6566));
    outputs(6327) <= not(layer0_outputs(2520));
    outputs(6328) <= not(layer0_outputs(4482));
    outputs(6329) <= not(layer0_outputs(10056));
    outputs(6330) <= (layer0_outputs(6300)) and not (layer0_outputs(7274));
    outputs(6331) <= not(layer0_outputs(7977));
    outputs(6332) <= layer0_outputs(1312);
    outputs(6333) <= not(layer0_outputs(5403));
    outputs(6334) <= (layer0_outputs(1987)) and not (layer0_outputs(3465));
    outputs(6335) <= layer0_outputs(4459);
    outputs(6336) <= not((layer0_outputs(6142)) or (layer0_outputs(7389)));
    outputs(6337) <= (layer0_outputs(8332)) and not (layer0_outputs(3799));
    outputs(6338) <= not(layer0_outputs(9375)) or (layer0_outputs(9377));
    outputs(6339) <= layer0_outputs(4116);
    outputs(6340) <= (layer0_outputs(5709)) and not (layer0_outputs(458));
    outputs(6341) <= not(layer0_outputs(3849));
    outputs(6342) <= not((layer0_outputs(6699)) xor (layer0_outputs(3288)));
    outputs(6343) <= (layer0_outputs(9661)) or (layer0_outputs(7415));
    outputs(6344) <= layer0_outputs(6060);
    outputs(6345) <= not(layer0_outputs(5424));
    outputs(6346) <= not(layer0_outputs(1206)) or (layer0_outputs(715));
    outputs(6347) <= layer0_outputs(500);
    outputs(6348) <= (layer0_outputs(6589)) and (layer0_outputs(958));
    outputs(6349) <= not(layer0_outputs(8051)) or (layer0_outputs(5244));
    outputs(6350) <= layer0_outputs(7177);
    outputs(6351) <= not((layer0_outputs(909)) xor (layer0_outputs(6409)));
    outputs(6352) <= not(layer0_outputs(5409));
    outputs(6353) <= not((layer0_outputs(2532)) xor (layer0_outputs(5784)));
    outputs(6354) <= not((layer0_outputs(2118)) or (layer0_outputs(4576)));
    outputs(6355) <= (layer0_outputs(5844)) and not (layer0_outputs(1338));
    outputs(6356) <= layer0_outputs(6692);
    outputs(6357) <= not(layer0_outputs(2097));
    outputs(6358) <= not((layer0_outputs(7264)) and (layer0_outputs(5948)));
    outputs(6359) <= layer0_outputs(7431);
    outputs(6360) <= (layer0_outputs(48)) and not (layer0_outputs(5177));
    outputs(6361) <= (layer0_outputs(1497)) xor (layer0_outputs(8240));
    outputs(6362) <= not((layer0_outputs(2794)) xor (layer0_outputs(1019)));
    outputs(6363) <= (layer0_outputs(6910)) and not (layer0_outputs(879));
    outputs(6364) <= not(layer0_outputs(10102));
    outputs(6365) <= layer0_outputs(702);
    outputs(6366) <= not(layer0_outputs(8145));
    outputs(6367) <= not((layer0_outputs(5828)) xor (layer0_outputs(6)));
    outputs(6368) <= not((layer0_outputs(7446)) or (layer0_outputs(1468)));
    outputs(6369) <= (layer0_outputs(8399)) xor (layer0_outputs(1665));
    outputs(6370) <= layer0_outputs(9400);
    outputs(6371) <= (layer0_outputs(9528)) and not (layer0_outputs(3677));
    outputs(6372) <= not((layer0_outputs(8089)) and (layer0_outputs(6570)));
    outputs(6373) <= not(layer0_outputs(2400)) or (layer0_outputs(5420));
    outputs(6374) <= not((layer0_outputs(1374)) xor (layer0_outputs(10125)));
    outputs(6375) <= not(layer0_outputs(1622));
    outputs(6376) <= layer0_outputs(2159);
    outputs(6377) <= (layer0_outputs(6994)) xor (layer0_outputs(2464));
    outputs(6378) <= (layer0_outputs(312)) xor (layer0_outputs(3143));
    outputs(6379) <= not(layer0_outputs(9456));
    outputs(6380) <= (layer0_outputs(2472)) and not (layer0_outputs(504));
    outputs(6381) <= (layer0_outputs(5051)) and not (layer0_outputs(5860));
    outputs(6382) <= not(layer0_outputs(6126));
    outputs(6383) <= not((layer0_outputs(9829)) and (layer0_outputs(4212)));
    outputs(6384) <= (layer0_outputs(6428)) and (layer0_outputs(6357));
    outputs(6385) <= layer0_outputs(7101);
    outputs(6386) <= layer0_outputs(2166);
    outputs(6387) <= not((layer0_outputs(4699)) and (layer0_outputs(7579)));
    outputs(6388) <= not(layer0_outputs(2443));
    outputs(6389) <= layer0_outputs(4233);
    outputs(6390) <= not(layer0_outputs(9089));
    outputs(6391) <= not(layer0_outputs(1440));
    outputs(6392) <= not((layer0_outputs(446)) and (layer0_outputs(890)));
    outputs(6393) <= layer0_outputs(6489);
    outputs(6394) <= (layer0_outputs(8891)) and not (layer0_outputs(1756));
    outputs(6395) <= layer0_outputs(9235);
    outputs(6396) <= not(layer0_outputs(6666));
    outputs(6397) <= not(layer0_outputs(9724));
    outputs(6398) <= layer0_outputs(2883);
    outputs(6399) <= not(layer0_outputs(7557));
    outputs(6400) <= layer0_outputs(3714);
    outputs(6401) <= not(layer0_outputs(9785));
    outputs(6402) <= not(layer0_outputs(8904));
    outputs(6403) <= not(layer0_outputs(6257));
    outputs(6404) <= (layer0_outputs(9454)) xor (layer0_outputs(5181));
    outputs(6405) <= not((layer0_outputs(8918)) or (layer0_outputs(9093)));
    outputs(6406) <= not(layer0_outputs(3082));
    outputs(6407) <= (layer0_outputs(2628)) or (layer0_outputs(179));
    outputs(6408) <= not(layer0_outputs(4483));
    outputs(6409) <= layer0_outputs(9219);
    outputs(6410) <= not(layer0_outputs(3699));
    outputs(6411) <= not((layer0_outputs(3317)) or (layer0_outputs(7344)));
    outputs(6412) <= not((layer0_outputs(10094)) or (layer0_outputs(7838)));
    outputs(6413) <= not((layer0_outputs(2097)) or (layer0_outputs(3531)));
    outputs(6414) <= layer0_outputs(9151);
    outputs(6415) <= not(layer0_outputs(8904));
    outputs(6416) <= (layer0_outputs(8613)) xor (layer0_outputs(732));
    outputs(6417) <= not(layer0_outputs(6028));
    outputs(6418) <= (layer0_outputs(1315)) or (layer0_outputs(2438));
    outputs(6419) <= layer0_outputs(3806);
    outputs(6420) <= layer0_outputs(4342);
    outputs(6421) <= not(layer0_outputs(5517));
    outputs(6422) <= (layer0_outputs(1105)) and (layer0_outputs(3658));
    outputs(6423) <= layer0_outputs(6501);
    outputs(6424) <= (layer0_outputs(1370)) and not (layer0_outputs(6518));
    outputs(6425) <= (layer0_outputs(1086)) or (layer0_outputs(7131));
    outputs(6426) <= not((layer0_outputs(8049)) or (layer0_outputs(4076)));
    outputs(6427) <= (layer0_outputs(9461)) and not (layer0_outputs(1991));
    outputs(6428) <= not((layer0_outputs(2655)) xor (layer0_outputs(9889)));
    outputs(6429) <= layer0_outputs(9298);
    outputs(6430) <= not(layer0_outputs(10184));
    outputs(6431) <= (layer0_outputs(2116)) and not (layer0_outputs(3048));
    outputs(6432) <= not((layer0_outputs(1681)) or (layer0_outputs(10068)));
    outputs(6433) <= layer0_outputs(9270);
    outputs(6434) <= (layer0_outputs(5120)) and (layer0_outputs(1152));
    outputs(6435) <= layer0_outputs(4101);
    outputs(6436) <= layer0_outputs(1694);
    outputs(6437) <= (layer0_outputs(1415)) or (layer0_outputs(9862));
    outputs(6438) <= layer0_outputs(4577);
    outputs(6439) <= (layer0_outputs(5246)) and not (layer0_outputs(5372));
    outputs(6440) <= (layer0_outputs(4919)) and not (layer0_outputs(7613));
    outputs(6441) <= not(layer0_outputs(3458));
    outputs(6442) <= not((layer0_outputs(7654)) and (layer0_outputs(7950)));
    outputs(6443) <= not((layer0_outputs(4333)) or (layer0_outputs(9662)));
    outputs(6444) <= layer0_outputs(529);
    outputs(6445) <= not(layer0_outputs(3292));
    outputs(6446) <= layer0_outputs(6454);
    outputs(6447) <= not(layer0_outputs(8659));
    outputs(6448) <= not((layer0_outputs(7313)) xor (layer0_outputs(4921)));
    outputs(6449) <= not((layer0_outputs(6676)) or (layer0_outputs(5785)));
    outputs(6450) <= not(layer0_outputs(6458)) or (layer0_outputs(3722));
    outputs(6451) <= not(layer0_outputs(5219));
    outputs(6452) <= not(layer0_outputs(8858));
    outputs(6453) <= not((layer0_outputs(1664)) xor (layer0_outputs(3843)));
    outputs(6454) <= not(layer0_outputs(1581));
    outputs(6455) <= (layer0_outputs(3483)) and not (layer0_outputs(8216));
    outputs(6456) <= (layer0_outputs(1739)) xor (layer0_outputs(6163));
    outputs(6457) <= layer0_outputs(1954);
    outputs(6458) <= (layer0_outputs(5973)) and not (layer0_outputs(4063));
    outputs(6459) <= not(layer0_outputs(6012));
    outputs(6460) <= not((layer0_outputs(1465)) or (layer0_outputs(9634)));
    outputs(6461) <= not(layer0_outputs(1482));
    outputs(6462) <= not(layer0_outputs(6739));
    outputs(6463) <= (layer0_outputs(605)) and not (layer0_outputs(1179));
    outputs(6464) <= layer0_outputs(2073);
    outputs(6465) <= not(layer0_outputs(2243));
    outputs(6466) <= not(layer0_outputs(2470)) or (layer0_outputs(6585));
    outputs(6467) <= layer0_outputs(8320);
    outputs(6468) <= not((layer0_outputs(2600)) or (layer0_outputs(867)));
    outputs(6469) <= not(layer0_outputs(5126));
    outputs(6470) <= not((layer0_outputs(6227)) or (layer0_outputs(7664)));
    outputs(6471) <= not(layer0_outputs(4520));
    outputs(6472) <= (layer0_outputs(8886)) and (layer0_outputs(8935));
    outputs(6473) <= not((layer0_outputs(5303)) or (layer0_outputs(4355)));
    outputs(6474) <= (layer0_outputs(3470)) xor (layer0_outputs(9322));
    outputs(6475) <= (layer0_outputs(1081)) xor (layer0_outputs(4526));
    outputs(6476) <= not(layer0_outputs(7729));
    outputs(6477) <= layer0_outputs(8663);
    outputs(6478) <= not(layer0_outputs(4997));
    outputs(6479) <= (layer0_outputs(1557)) and (layer0_outputs(9881));
    outputs(6480) <= not(layer0_outputs(598));
    outputs(6481) <= layer0_outputs(2357);
    outputs(6482) <= (layer0_outputs(5974)) or (layer0_outputs(3075));
    outputs(6483) <= not(layer0_outputs(2392));
    outputs(6484) <= layer0_outputs(7633);
    outputs(6485) <= not(layer0_outputs(10117));
    outputs(6486) <= (layer0_outputs(7658)) and not (layer0_outputs(6986));
    outputs(6487) <= layer0_outputs(1921);
    outputs(6488) <= (layer0_outputs(3200)) and not (layer0_outputs(2681));
    outputs(6489) <= not((layer0_outputs(8858)) or (layer0_outputs(4667)));
    outputs(6490) <= (layer0_outputs(1538)) and (layer0_outputs(5421));
    outputs(6491) <= (layer0_outputs(200)) and (layer0_outputs(8388));
    outputs(6492) <= (layer0_outputs(9730)) and not (layer0_outputs(2584));
    outputs(6493) <= not(layer0_outputs(3583));
    outputs(6494) <= not((layer0_outputs(6027)) or (layer0_outputs(6741)));
    outputs(6495) <= not(layer0_outputs(9945));
    outputs(6496) <= not((layer0_outputs(6996)) or (layer0_outputs(2219)));
    outputs(6497) <= not((layer0_outputs(6225)) and (layer0_outputs(1766)));
    outputs(6498) <= layer0_outputs(9933);
    outputs(6499) <= not(layer0_outputs(4113));
    outputs(6500) <= not(layer0_outputs(7429)) or (layer0_outputs(9483));
    outputs(6501) <= layer0_outputs(6892);
    outputs(6502) <= layer0_outputs(2398);
    outputs(6503) <= not((layer0_outputs(7935)) or (layer0_outputs(10189)));
    outputs(6504) <= (layer0_outputs(976)) or (layer0_outputs(1927));
    outputs(6505) <= not(layer0_outputs(6157));
    outputs(6506) <= not(layer0_outputs(5010));
    outputs(6507) <= layer0_outputs(4944);
    outputs(6508) <= not(layer0_outputs(6345));
    outputs(6509) <= layer0_outputs(772);
    outputs(6510) <= layer0_outputs(4745);
    outputs(6511) <= (layer0_outputs(7208)) xor (layer0_outputs(5425));
    outputs(6512) <= layer0_outputs(357);
    outputs(6513) <= not((layer0_outputs(8425)) xor (layer0_outputs(5283)));
    outputs(6514) <= not(layer0_outputs(1577));
    outputs(6515) <= layer0_outputs(3203);
    outputs(6516) <= not(layer0_outputs(7991));
    outputs(6517) <= (layer0_outputs(3975)) and not (layer0_outputs(4691));
    outputs(6518) <= not((layer0_outputs(2947)) xor (layer0_outputs(7197)));
    outputs(6519) <= not(layer0_outputs(9659));
    outputs(6520) <= not((layer0_outputs(4895)) xor (layer0_outputs(7029)));
    outputs(6521) <= layer0_outputs(8514);
    outputs(6522) <= not(layer0_outputs(633)) or (layer0_outputs(3933));
    outputs(6523) <= (layer0_outputs(5608)) and not (layer0_outputs(1799));
    outputs(6524) <= (layer0_outputs(3213)) and not (layer0_outputs(2000));
    outputs(6525) <= not((layer0_outputs(7550)) xor (layer0_outputs(4791)));
    outputs(6526) <= layer0_outputs(9774);
    outputs(6527) <= (layer0_outputs(223)) and not (layer0_outputs(6587));
    outputs(6528) <= layer0_outputs(2597);
    outputs(6529) <= not((layer0_outputs(3548)) xor (layer0_outputs(9294)));
    outputs(6530) <= not((layer0_outputs(4378)) and (layer0_outputs(9964)));
    outputs(6531) <= not((layer0_outputs(6441)) or (layer0_outputs(6876)));
    outputs(6532) <= not(layer0_outputs(5185));
    outputs(6533) <= (layer0_outputs(8963)) and not (layer0_outputs(2000));
    outputs(6534) <= layer0_outputs(5688);
    outputs(6535) <= not((layer0_outputs(262)) xor (layer0_outputs(3161)));
    outputs(6536) <= (layer0_outputs(7325)) and (layer0_outputs(3392));
    outputs(6537) <= layer0_outputs(4940);
    outputs(6538) <= not((layer0_outputs(7927)) or (layer0_outputs(9333)));
    outputs(6539) <= not(layer0_outputs(5986)) or (layer0_outputs(7019));
    outputs(6540) <= (layer0_outputs(3893)) or (layer0_outputs(4806));
    outputs(6541) <= (layer0_outputs(2388)) and not (layer0_outputs(1421));
    outputs(6542) <= layer0_outputs(3710);
    outputs(6543) <= not(layer0_outputs(4024));
    outputs(6544) <= (layer0_outputs(5087)) xor (layer0_outputs(5471));
    outputs(6545) <= layer0_outputs(3312);
    outputs(6546) <= (layer0_outputs(4695)) and (layer0_outputs(9578));
    outputs(6547) <= (layer0_outputs(5943)) and not (layer0_outputs(5391));
    outputs(6548) <= not((layer0_outputs(3519)) or (layer0_outputs(4720)));
    outputs(6549) <= not(layer0_outputs(1309)) or (layer0_outputs(645));
    outputs(6550) <= (layer0_outputs(709)) and not (layer0_outputs(8309));
    outputs(6551) <= layer0_outputs(4669);
    outputs(6552) <= layer0_outputs(3863);
    outputs(6553) <= not(layer0_outputs(732));
    outputs(6554) <= (layer0_outputs(3599)) and not (layer0_outputs(6759));
    outputs(6555) <= (layer0_outputs(3763)) and not (layer0_outputs(3362));
    outputs(6556) <= layer0_outputs(8721);
    outputs(6557) <= not((layer0_outputs(6979)) or (layer0_outputs(1215)));
    outputs(6558) <= (layer0_outputs(2389)) xor (layer0_outputs(2637));
    outputs(6559) <= (layer0_outputs(4652)) and (layer0_outputs(9386));
    outputs(6560) <= layer0_outputs(9695);
    outputs(6561) <= layer0_outputs(6651);
    outputs(6562) <= not((layer0_outputs(7048)) xor (layer0_outputs(9422)));
    outputs(6563) <= (layer0_outputs(4035)) xor (layer0_outputs(2314));
    outputs(6564) <= layer0_outputs(5688);
    outputs(6565) <= layer0_outputs(6079);
    outputs(6566) <= not((layer0_outputs(1670)) or (layer0_outputs(8717)));
    outputs(6567) <= not(layer0_outputs(3615)) or (layer0_outputs(5441));
    outputs(6568) <= not((layer0_outputs(7506)) and (layer0_outputs(9852)));
    outputs(6569) <= (layer0_outputs(6965)) and not (layer0_outputs(2394));
    outputs(6570) <= layer0_outputs(5494);
    outputs(6571) <= (layer0_outputs(3416)) and not (layer0_outputs(7827));
    outputs(6572) <= layer0_outputs(5650);
    outputs(6573) <= not(layer0_outputs(1699));
    outputs(6574) <= (layer0_outputs(6202)) and not (layer0_outputs(5401));
    outputs(6575) <= not(layer0_outputs(4215));
    outputs(6576) <= not((layer0_outputs(7163)) or (layer0_outputs(4957)));
    outputs(6577) <= not(layer0_outputs(5630));
    outputs(6578) <= (layer0_outputs(2566)) xor (layer0_outputs(6075));
    outputs(6579) <= (layer0_outputs(6224)) and (layer0_outputs(7839));
    outputs(6580) <= not(layer0_outputs(8975));
    outputs(6581) <= (layer0_outputs(1360)) and not (layer0_outputs(7400));
    outputs(6582) <= not(layer0_outputs(183)) or (layer0_outputs(9753));
    outputs(6583) <= not(layer0_outputs(3240)) or (layer0_outputs(4655));
    outputs(6584) <= not((layer0_outputs(1391)) or (layer0_outputs(2238)));
    outputs(6585) <= layer0_outputs(10155);
    outputs(6586) <= (layer0_outputs(3690)) and not (layer0_outputs(9996));
    outputs(6587) <= (layer0_outputs(6505)) or (layer0_outputs(9330));
    outputs(6588) <= not(layer0_outputs(7135));
    outputs(6589) <= not(layer0_outputs(7784));
    outputs(6590) <= layer0_outputs(6007);
    outputs(6591) <= not(layer0_outputs(5980));
    outputs(6592) <= layer0_outputs(2154);
    outputs(6593) <= layer0_outputs(4594);
    outputs(6594) <= (layer0_outputs(2973)) xor (layer0_outputs(6067));
    outputs(6595) <= layer0_outputs(449);
    outputs(6596) <= not((layer0_outputs(3922)) or (layer0_outputs(7134)));
    outputs(6597) <= (layer0_outputs(3829)) and not (layer0_outputs(9175));
    outputs(6598) <= (layer0_outputs(3852)) and not (layer0_outputs(6026));
    outputs(6599) <= not(layer0_outputs(5097));
    outputs(6600) <= not((layer0_outputs(2863)) xor (layer0_outputs(7798)));
    outputs(6601) <= (layer0_outputs(8995)) or (layer0_outputs(7983));
    outputs(6602) <= layer0_outputs(700);
    outputs(6603) <= not(layer0_outputs(7868));
    outputs(6604) <= (layer0_outputs(9116)) xor (layer0_outputs(3717));
    outputs(6605) <= not(layer0_outputs(9234));
    outputs(6606) <= not(layer0_outputs(8295)) or (layer0_outputs(1500));
    outputs(6607) <= (layer0_outputs(9382)) xor (layer0_outputs(8830));
    outputs(6608) <= layer0_outputs(6358);
    outputs(6609) <= layer0_outputs(8238);
    outputs(6610) <= layer0_outputs(5547);
    outputs(6611) <= not(layer0_outputs(4159));
    outputs(6612) <= (layer0_outputs(7870)) xor (layer0_outputs(5581));
    outputs(6613) <= not(layer0_outputs(2726));
    outputs(6614) <= not(layer0_outputs(10178));
    outputs(6615) <= layer0_outputs(1520);
    outputs(6616) <= not(layer0_outputs(4252));
    outputs(6617) <= not((layer0_outputs(147)) or (layer0_outputs(3465)));
    outputs(6618) <= layer0_outputs(586);
    outputs(6619) <= (layer0_outputs(9156)) or (layer0_outputs(2832));
    outputs(6620) <= not(layer0_outputs(5875));
    outputs(6621) <= not((layer0_outputs(6838)) xor (layer0_outputs(6649)));
    outputs(6622) <= not(layer0_outputs(9699));
    outputs(6623) <= layer0_outputs(2856);
    outputs(6624) <= not(layer0_outputs(3877));
    outputs(6625) <= (layer0_outputs(6746)) and not (layer0_outputs(10187));
    outputs(6626) <= not(layer0_outputs(6956));
    outputs(6627) <= (layer0_outputs(997)) and (layer0_outputs(3409));
    outputs(6628) <= layer0_outputs(8114);
    outputs(6629) <= layer0_outputs(3508);
    outputs(6630) <= not(layer0_outputs(3133));
    outputs(6631) <= not(layer0_outputs(485));
    outputs(6632) <= layer0_outputs(1377);
    outputs(6633) <= not(layer0_outputs(3041));
    outputs(6634) <= (layer0_outputs(3909)) xor (layer0_outputs(427));
    outputs(6635) <= not((layer0_outputs(9185)) or (layer0_outputs(2167)));
    outputs(6636) <= not(layer0_outputs(4003));
    outputs(6637) <= (layer0_outputs(2924)) and (layer0_outputs(4977));
    outputs(6638) <= not((layer0_outputs(6611)) or (layer0_outputs(2502)));
    outputs(6639) <= (layer0_outputs(6471)) and (layer0_outputs(1100));
    outputs(6640) <= not((layer0_outputs(9084)) or (layer0_outputs(908)));
    outputs(6641) <= layer0_outputs(1559);
    outputs(6642) <= not(layer0_outputs(4616));
    outputs(6643) <= (layer0_outputs(9938)) or (layer0_outputs(8813));
    outputs(6644) <= (layer0_outputs(1446)) and not (layer0_outputs(2354));
    outputs(6645) <= (layer0_outputs(8883)) xor (layer0_outputs(149));
    outputs(6646) <= not(layer0_outputs(3193));
    outputs(6647) <= (layer0_outputs(7413)) and (layer0_outputs(7121));
    outputs(6648) <= not(layer0_outputs(3939));
    outputs(6649) <= (layer0_outputs(6851)) and not (layer0_outputs(9744));
    outputs(6650) <= not(layer0_outputs(6756));
    outputs(6651) <= not(layer0_outputs(8805));
    outputs(6652) <= layer0_outputs(225);
    outputs(6653) <= not(layer0_outputs(5209));
    outputs(6654) <= layer0_outputs(1353);
    outputs(6655) <= layer0_outputs(6879);
    outputs(6656) <= not(layer0_outputs(8925));
    outputs(6657) <= (layer0_outputs(295)) and (layer0_outputs(4619));
    outputs(6658) <= (layer0_outputs(8735)) and not (layer0_outputs(6542));
    outputs(6659) <= not(layer0_outputs(7280));
    outputs(6660) <= layer0_outputs(6972);
    outputs(6661) <= layer0_outputs(1478);
    outputs(6662) <= layer0_outputs(4942);
    outputs(6663) <= layer0_outputs(4807);
    outputs(6664) <= layer0_outputs(4870);
    outputs(6665) <= layer0_outputs(6411);
    outputs(6666) <= not(layer0_outputs(5826));
    outputs(6667) <= not(layer0_outputs(2869));
    outputs(6668) <= not(layer0_outputs(1777)) or (layer0_outputs(7677));
    outputs(6669) <= (layer0_outputs(8488)) and not (layer0_outputs(10025));
    outputs(6670) <= not((layer0_outputs(6590)) or (layer0_outputs(1183)));
    outputs(6671) <= not(layer0_outputs(2611));
    outputs(6672) <= (layer0_outputs(10226)) or (layer0_outputs(527));
    outputs(6673) <= not(layer0_outputs(6198));
    outputs(6674) <= not(layer0_outputs(3937));
    outputs(6675) <= (layer0_outputs(6701)) xor (layer0_outputs(249));
    outputs(6676) <= not(layer0_outputs(1648));
    outputs(6677) <= (layer0_outputs(6063)) and not (layer0_outputs(3524));
    outputs(6678) <= (layer0_outputs(1945)) or (layer0_outputs(1809));
    outputs(6679) <= (layer0_outputs(1197)) xor (layer0_outputs(5198));
    outputs(6680) <= not((layer0_outputs(4493)) and (layer0_outputs(4295)));
    outputs(6681) <= not(layer0_outputs(334));
    outputs(6682) <= not(layer0_outputs(2938)) or (layer0_outputs(4866));
    outputs(6683) <= not((layer0_outputs(8486)) and (layer0_outputs(9845)));
    outputs(6684) <= not(layer0_outputs(7836));
    outputs(6685) <= (layer0_outputs(7763)) and not (layer0_outputs(8047));
    outputs(6686) <= not(layer0_outputs(7035));
    outputs(6687) <= (layer0_outputs(4227)) and not (layer0_outputs(1029));
    outputs(6688) <= layer0_outputs(920);
    outputs(6689) <= (layer0_outputs(7694)) and not (layer0_outputs(4587));
    outputs(6690) <= (layer0_outputs(7819)) xor (layer0_outputs(9318));
    outputs(6691) <= layer0_outputs(9539);
    outputs(6692) <= (layer0_outputs(9162)) xor (layer0_outputs(1230));
    outputs(6693) <= not(layer0_outputs(8456));
    outputs(6694) <= (layer0_outputs(1103)) and (layer0_outputs(8259));
    outputs(6695) <= (layer0_outputs(7234)) xor (layer0_outputs(4196));
    outputs(6696) <= layer0_outputs(1225);
    outputs(6697) <= (layer0_outputs(4133)) and not (layer0_outputs(4994));
    outputs(6698) <= not((layer0_outputs(666)) xor (layer0_outputs(2910)));
    outputs(6699) <= not(layer0_outputs(4450)) or (layer0_outputs(3196));
    outputs(6700) <= (layer0_outputs(7544)) and not (layer0_outputs(3869));
    outputs(6701) <= layer0_outputs(9906);
    outputs(6702) <= not(layer0_outputs(4558));
    outputs(6703) <= not((layer0_outputs(7935)) xor (layer0_outputs(10051)));
    outputs(6704) <= (layer0_outputs(7329)) and (layer0_outputs(4666));
    outputs(6705) <= not(layer0_outputs(7092));
    outputs(6706) <= layer0_outputs(7011);
    outputs(6707) <= layer0_outputs(4288);
    outputs(6708) <= (layer0_outputs(1470)) and not (layer0_outputs(7826));
    outputs(6709) <= not((layer0_outputs(7675)) xor (layer0_outputs(480)));
    outputs(6710) <= (layer0_outputs(6476)) xor (layer0_outputs(9934));
    outputs(6711) <= (layer0_outputs(9613)) and (layer0_outputs(9345));
    outputs(6712) <= not(layer0_outputs(1444)) or (layer0_outputs(9766));
    outputs(6713) <= (layer0_outputs(3139)) and not (layer0_outputs(5440));
    outputs(6714) <= not(layer0_outputs(2360));
    outputs(6715) <= layer0_outputs(8042);
    outputs(6716) <= layer0_outputs(3920);
    outputs(6717) <= not(layer0_outputs(6226));
    outputs(6718) <= (layer0_outputs(758)) and not (layer0_outputs(5519));
    outputs(6719) <= not(layer0_outputs(93)) or (layer0_outputs(7109));
    outputs(6720) <= (layer0_outputs(8213)) xor (layer0_outputs(1441));
    outputs(6721) <= layer0_outputs(9844);
    outputs(6722) <= not(layer0_outputs(338)) or (layer0_outputs(9136));
    outputs(6723) <= not(layer0_outputs(2988));
    outputs(6724) <= not(layer0_outputs(5783));
    outputs(6725) <= not(layer0_outputs(8768));
    outputs(6726) <= layer0_outputs(1894);
    outputs(6727) <= not(layer0_outputs(5234));
    outputs(6728) <= (layer0_outputs(5887)) and not (layer0_outputs(6744));
    outputs(6729) <= not(layer0_outputs(4909)) or (layer0_outputs(1672));
    outputs(6730) <= not(layer0_outputs(8236));
    outputs(6731) <= not((layer0_outputs(6497)) or (layer0_outputs(124)));
    outputs(6732) <= layer0_outputs(581);
    outputs(6733) <= not((layer0_outputs(6874)) xor (layer0_outputs(1060)));
    outputs(6734) <= not(layer0_outputs(8985));
    outputs(6735) <= layer0_outputs(167);
    outputs(6736) <= (layer0_outputs(2814)) and not (layer0_outputs(3309));
    outputs(6737) <= (layer0_outputs(8576)) xor (layer0_outputs(9619));
    outputs(6738) <= not((layer0_outputs(2957)) xor (layer0_outputs(9547)));
    outputs(6739) <= not((layer0_outputs(7255)) xor (layer0_outputs(5778)));
    outputs(6740) <= (layer0_outputs(9213)) and (layer0_outputs(1089));
    outputs(6741) <= not(layer0_outputs(3192));
    outputs(6742) <= not(layer0_outputs(8581)) or (layer0_outputs(7897));
    outputs(6743) <= (layer0_outputs(1301)) and (layer0_outputs(6069));
    outputs(6744) <= layer0_outputs(4912);
    outputs(6745) <= not(layer0_outputs(3210));
    outputs(6746) <= (layer0_outputs(5165)) and not (layer0_outputs(7022));
    outputs(6747) <= layer0_outputs(7312);
    outputs(6748) <= not(layer0_outputs(10078)) or (layer0_outputs(10058));
    outputs(6749) <= not(layer0_outputs(7014));
    outputs(6750) <= (layer0_outputs(601)) xor (layer0_outputs(8264));
    outputs(6751) <= layer0_outputs(3788);
    outputs(6752) <= (layer0_outputs(3084)) and not (layer0_outputs(2589));
    outputs(6753) <= (layer0_outputs(7538)) xor (layer0_outputs(747));
    outputs(6754) <= not(layer0_outputs(9622));
    outputs(6755) <= not((layer0_outputs(3027)) or (layer0_outputs(570)));
    outputs(6756) <= not(layer0_outputs(9744));
    outputs(6757) <= not(layer0_outputs(909));
    outputs(6758) <= not((layer0_outputs(8677)) xor (layer0_outputs(5475)));
    outputs(6759) <= not(layer0_outputs(4203));
    outputs(6760) <= layer0_outputs(9271);
    outputs(6761) <= (layer0_outputs(8917)) and (layer0_outputs(7438));
    outputs(6762) <= (layer0_outputs(8212)) and not (layer0_outputs(8784));
    outputs(6763) <= layer0_outputs(7052);
    outputs(6764) <= layer0_outputs(6975);
    outputs(6765) <= not(layer0_outputs(9617)) or (layer0_outputs(4464));
    outputs(6766) <= not(layer0_outputs(6739));
    outputs(6767) <= (layer0_outputs(6177)) or (layer0_outputs(6317));
    outputs(6768) <= not(layer0_outputs(120)) or (layer0_outputs(5952));
    outputs(6769) <= not(layer0_outputs(896));
    outputs(6770) <= (layer0_outputs(9824)) and not (layer0_outputs(4172));
    outputs(6771) <= (layer0_outputs(4733)) and not (layer0_outputs(2738));
    outputs(6772) <= not((layer0_outputs(2206)) or (layer0_outputs(6219)));
    outputs(6773) <= not((layer0_outputs(2162)) and (layer0_outputs(1628)));
    outputs(6774) <= not(layer0_outputs(3835));
    outputs(6775) <= not(layer0_outputs(2080));
    outputs(6776) <= (layer0_outputs(4590)) and (layer0_outputs(10048));
    outputs(6777) <= layer0_outputs(8140);
    outputs(6778) <= not(layer0_outputs(8129));
    outputs(6779) <= not(layer0_outputs(55)) or (layer0_outputs(8018));
    outputs(6780) <= (layer0_outputs(3885)) and not (layer0_outputs(8850));
    outputs(6781) <= not((layer0_outputs(827)) or (layer0_outputs(4143)));
    outputs(6782) <= (layer0_outputs(4191)) and (layer0_outputs(2861));
    outputs(6783) <= not(layer0_outputs(8393));
    outputs(6784) <= not((layer0_outputs(9679)) or (layer0_outputs(1107)));
    outputs(6785) <= (layer0_outputs(343)) and not (layer0_outputs(3650));
    outputs(6786) <= layer0_outputs(8114);
    outputs(6787) <= layer0_outputs(5575);
    outputs(6788) <= not(layer0_outputs(8741));
    outputs(6789) <= (layer0_outputs(3212)) and not (layer0_outputs(6787));
    outputs(6790) <= (layer0_outputs(1545)) and not (layer0_outputs(3695));
    outputs(6791) <= layer0_outputs(3821);
    outputs(6792) <= (layer0_outputs(5916)) and not (layer0_outputs(9409));
    outputs(6793) <= (layer0_outputs(9963)) and not (layer0_outputs(476));
    outputs(6794) <= not((layer0_outputs(6355)) or (layer0_outputs(72)));
    outputs(6795) <= (layer0_outputs(2335)) xor (layer0_outputs(3964));
    outputs(6796) <= (layer0_outputs(9627)) or (layer0_outputs(9757));
    outputs(6797) <= (layer0_outputs(4564)) or (layer0_outputs(6066));
    outputs(6798) <= layer0_outputs(340);
    outputs(6799) <= (layer0_outputs(8046)) and not (layer0_outputs(7));
    outputs(6800) <= not((layer0_outputs(7016)) or (layer0_outputs(8720)));
    outputs(6801) <= not(layer0_outputs(1033));
    outputs(6802) <= (layer0_outputs(7021)) xor (layer0_outputs(1344));
    outputs(6803) <= layer0_outputs(4499);
    outputs(6804) <= layer0_outputs(5709);
    outputs(6805) <= not((layer0_outputs(5642)) or (layer0_outputs(4005)));
    outputs(6806) <= not(layer0_outputs(3809));
    outputs(6807) <= (layer0_outputs(201)) and (layer0_outputs(1970));
    outputs(6808) <= (layer0_outputs(7015)) xor (layer0_outputs(6414));
    outputs(6809) <= (layer0_outputs(5591)) or (layer0_outputs(498));
    outputs(6810) <= (layer0_outputs(4468)) xor (layer0_outputs(3201));
    outputs(6811) <= not((layer0_outputs(6768)) xor (layer0_outputs(9907)));
    outputs(6812) <= layer0_outputs(1261);
    outputs(6813) <= not(layer0_outputs(2182));
    outputs(6814) <= layer0_outputs(3357);
    outputs(6815) <= not(layer0_outputs(9723));
    outputs(6816) <= not(layer0_outputs(6215));
    outputs(6817) <= (layer0_outputs(3830)) and not (layer0_outputs(4106));
    outputs(6818) <= (layer0_outputs(5352)) and not (layer0_outputs(6355));
    outputs(6819) <= not(layer0_outputs(1710));
    outputs(6820) <= (layer0_outputs(6501)) and not (layer0_outputs(3880));
    outputs(6821) <= (layer0_outputs(8552)) and (layer0_outputs(493));
    outputs(6822) <= not(layer0_outputs(7411));
    outputs(6823) <= not((layer0_outputs(8016)) and (layer0_outputs(205)));
    outputs(6824) <= layer0_outputs(864);
    outputs(6825) <= (layer0_outputs(1770)) xor (layer0_outputs(7388));
    outputs(6826) <= layer0_outputs(3673);
    outputs(6827) <= (layer0_outputs(4599)) and (layer0_outputs(8555));
    outputs(6828) <= not(layer0_outputs(4439)) or (layer0_outputs(2593));
    outputs(6829) <= (layer0_outputs(7462)) and not (layer0_outputs(787));
    outputs(6830) <= not(layer0_outputs(2749)) or (layer0_outputs(1959));
    outputs(6831) <= (layer0_outputs(822)) and not (layer0_outputs(9822));
    outputs(6832) <= not(layer0_outputs(2457)) or (layer0_outputs(4886));
    outputs(6833) <= (layer0_outputs(1535)) and (layer0_outputs(8092));
    outputs(6834) <= (layer0_outputs(7509)) xor (layer0_outputs(7426));
    outputs(6835) <= not((layer0_outputs(5011)) or (layer0_outputs(7821)));
    outputs(6836) <= not(layer0_outputs(4510));
    outputs(6837) <= (layer0_outputs(3157)) and not (layer0_outputs(6955));
    outputs(6838) <= not(layer0_outputs(699));
    outputs(6839) <= (layer0_outputs(9732)) and (layer0_outputs(8762));
    outputs(6840) <= layer0_outputs(10053);
    outputs(6841) <= (layer0_outputs(5906)) and (layer0_outputs(4570));
    outputs(6842) <= (layer0_outputs(9685)) and (layer0_outputs(4163));
    outputs(6843) <= not((layer0_outputs(19)) or (layer0_outputs(7532)));
    outputs(6844) <= (layer0_outputs(9492)) or (layer0_outputs(8275));
    outputs(6845) <= not((layer0_outputs(5302)) xor (layer0_outputs(234)));
    outputs(6846) <= not(layer0_outputs(2672));
    outputs(6847) <= not(layer0_outputs(2907));
    outputs(6848) <= not((layer0_outputs(8174)) xor (layer0_outputs(6682)));
    outputs(6849) <= not(layer0_outputs(1044));
    outputs(6850) <= not(layer0_outputs(4766));
    outputs(6851) <= not(layer0_outputs(1531));
    outputs(6852) <= (layer0_outputs(8199)) and not (layer0_outputs(1696));
    outputs(6853) <= (layer0_outputs(2297)) xor (layer0_outputs(3702));
    outputs(6854) <= not(layer0_outputs(1540));
    outputs(6855) <= not(layer0_outputs(1531));
    outputs(6856) <= not(layer0_outputs(2331));
    outputs(6857) <= not(layer0_outputs(1781));
    outputs(6858) <= (layer0_outputs(1409)) and not (layer0_outputs(5045));
    outputs(6859) <= not((layer0_outputs(7310)) or (layer0_outputs(8553)));
    outputs(6860) <= not((layer0_outputs(1184)) xor (layer0_outputs(3044)));
    outputs(6861) <= layer0_outputs(2218);
    outputs(6862) <= not(layer0_outputs(1901));
    outputs(6863) <= layer0_outputs(3091);
    outputs(6864) <= not(layer0_outputs(5674)) or (layer0_outputs(1949));
    outputs(6865) <= (layer0_outputs(7713)) xor (layer0_outputs(9031));
    outputs(6866) <= (layer0_outputs(119)) and not (layer0_outputs(557));
    outputs(6867) <= (layer0_outputs(6980)) and not (layer0_outputs(8590));
    outputs(6868) <= layer0_outputs(25);
    outputs(6869) <= (layer0_outputs(3660)) and (layer0_outputs(2593));
    outputs(6870) <= not(layer0_outputs(6410));
    outputs(6871) <= not((layer0_outputs(9430)) and (layer0_outputs(3637)));
    outputs(6872) <= (layer0_outputs(2171)) and not (layer0_outputs(4719));
    outputs(6873) <= layer0_outputs(914);
    outputs(6874) <= layer0_outputs(3825);
    outputs(6875) <= (layer0_outputs(8823)) and not (layer0_outputs(10026));
    outputs(6876) <= (layer0_outputs(9852)) xor (layer0_outputs(245));
    outputs(6877) <= (layer0_outputs(6074)) and not (layer0_outputs(694));
    outputs(6878) <= (layer0_outputs(8072)) xor (layer0_outputs(2146));
    outputs(6879) <= (layer0_outputs(4091)) and not (layer0_outputs(9835));
    outputs(6880) <= (layer0_outputs(6053)) or (layer0_outputs(9434));
    outputs(6881) <= not(layer0_outputs(410));
    outputs(6882) <= (layer0_outputs(1645)) or (layer0_outputs(3530));
    outputs(6883) <= (layer0_outputs(2472)) and not (layer0_outputs(3968));
    outputs(6884) <= not((layer0_outputs(4113)) xor (layer0_outputs(7258)));
    outputs(6885) <= not(layer0_outputs(7094));
    outputs(6886) <= layer0_outputs(2168);
    outputs(6887) <= not(layer0_outputs(7666)) or (layer0_outputs(2480));
    outputs(6888) <= not(layer0_outputs(6056));
    outputs(6889) <= not((layer0_outputs(4333)) or (layer0_outputs(8136)));
    outputs(6890) <= not(layer0_outputs(5516));
    outputs(6891) <= not(layer0_outputs(7180)) or (layer0_outputs(1672));
    outputs(6892) <= (layer0_outputs(7346)) and not (layer0_outputs(9942));
    outputs(6893) <= (layer0_outputs(8187)) and (layer0_outputs(2145));
    outputs(6894) <= not(layer0_outputs(106));
    outputs(6895) <= not(layer0_outputs(2402));
    outputs(6896) <= (layer0_outputs(2115)) and (layer0_outputs(4560));
    outputs(6897) <= not(layer0_outputs(8414));
    outputs(6898) <= not(layer0_outputs(8547));
    outputs(6899) <= not(layer0_outputs(3276));
    outputs(6900) <= not(layer0_outputs(1618)) or (layer0_outputs(1552));
    outputs(6901) <= (layer0_outputs(2736)) or (layer0_outputs(9319));
    outputs(6902) <= not(layer0_outputs(9643));
    outputs(6903) <= layer0_outputs(9957);
    outputs(6904) <= not(layer0_outputs(3876));
    outputs(6905) <= not(layer0_outputs(2926)) or (layer0_outputs(9460));
    outputs(6906) <= not(layer0_outputs(5978));
    outputs(6907) <= (layer0_outputs(3267)) xor (layer0_outputs(7348));
    outputs(6908) <= not(layer0_outputs(9727));
    outputs(6909) <= layer0_outputs(4892);
    outputs(6910) <= not(layer0_outputs(5144));
    outputs(6911) <= layer0_outputs(2797);
    outputs(6912) <= layer0_outputs(5598);
    outputs(6913) <= layer0_outputs(3779);
    outputs(6914) <= not(layer0_outputs(1096));
    outputs(6915) <= not(layer0_outputs(3861));
    outputs(6916) <= layer0_outputs(1589);
    outputs(6917) <= (layer0_outputs(404)) or (layer0_outputs(1928));
    outputs(6918) <= not(layer0_outputs(8375));
    outputs(6919) <= not((layer0_outputs(3613)) xor (layer0_outputs(8937)));
    outputs(6920) <= layer0_outputs(6762);
    outputs(6921) <= not((layer0_outputs(2069)) xor (layer0_outputs(1456)));
    outputs(6922) <= layer0_outputs(3751);
    outputs(6923) <= not(layer0_outputs(9593));
    outputs(6924) <= not(layer0_outputs(3227));
    outputs(6925) <= (layer0_outputs(1564)) xor (layer0_outputs(1011));
    outputs(6926) <= not(layer0_outputs(4316)) or (layer0_outputs(7156));
    outputs(6927) <= not((layer0_outputs(10071)) xor (layer0_outputs(5264)));
    outputs(6928) <= not((layer0_outputs(6906)) and (layer0_outputs(6467)));
    outputs(6929) <= (layer0_outputs(3340)) and (layer0_outputs(4424));
    outputs(6930) <= layer0_outputs(4248);
    outputs(6931) <= (layer0_outputs(9118)) and not (layer0_outputs(5010));
    outputs(6932) <= layer0_outputs(1274);
    outputs(6933) <= layer0_outputs(4836);
    outputs(6934) <= not(layer0_outputs(1106));
    outputs(6935) <= layer0_outputs(3452);
    outputs(6936) <= layer0_outputs(6881);
    outputs(6937) <= (layer0_outputs(2666)) or (layer0_outputs(4375));
    outputs(6938) <= (layer0_outputs(4584)) and (layer0_outputs(3066));
    outputs(6939) <= (layer0_outputs(9983)) and not (layer0_outputs(9105));
    outputs(6940) <= (layer0_outputs(4758)) and not (layer0_outputs(8938));
    outputs(6941) <= not(layer0_outputs(9285)) or (layer0_outputs(2836));
    outputs(6942) <= layer0_outputs(4230);
    outputs(6943) <= not(layer0_outputs(9563)) or (layer0_outputs(6978));
    outputs(6944) <= layer0_outputs(3101);
    outputs(6945) <= not((layer0_outputs(713)) or (layer0_outputs(7738)));
    outputs(6946) <= layer0_outputs(1070);
    outputs(6947) <= not(layer0_outputs(7114)) or (layer0_outputs(424));
    outputs(6948) <= not((layer0_outputs(10037)) xor (layer0_outputs(10175)));
    outputs(6949) <= (layer0_outputs(8220)) and not (layer0_outputs(9221));
    outputs(6950) <= not(layer0_outputs(8540));
    outputs(6951) <= (layer0_outputs(143)) and not (layer0_outputs(5869));
    outputs(6952) <= (layer0_outputs(1870)) and not (layer0_outputs(4378));
    outputs(6953) <= layer0_outputs(979);
    outputs(6954) <= not((layer0_outputs(6677)) and (layer0_outputs(2203)));
    outputs(6955) <= (layer0_outputs(5156)) xor (layer0_outputs(674));
    outputs(6956) <= not(layer0_outputs(10025));
    outputs(6957) <= (layer0_outputs(762)) and not (layer0_outputs(218));
    outputs(6958) <= not(layer0_outputs(9056)) or (layer0_outputs(5156));
    outputs(6959) <= (layer0_outputs(7968)) and not (layer0_outputs(6286));
    outputs(6960) <= layer0_outputs(8886);
    outputs(6961) <= not(layer0_outputs(563)) or (layer0_outputs(4790));
    outputs(6962) <= not(layer0_outputs(2009));
    outputs(6963) <= not((layer0_outputs(1839)) and (layer0_outputs(6479)));
    outputs(6964) <= (layer0_outputs(2455)) and not (layer0_outputs(5115));
    outputs(6965) <= layer0_outputs(9147);
    outputs(6966) <= (layer0_outputs(7692)) xor (layer0_outputs(8686));
    outputs(6967) <= not(layer0_outputs(8166));
    outputs(6968) <= not((layer0_outputs(607)) or (layer0_outputs(2164)));
    outputs(6969) <= (layer0_outputs(2303)) and not (layer0_outputs(9931));
    outputs(6970) <= layer0_outputs(2811);
    outputs(6971) <= layer0_outputs(5919);
    outputs(6972) <= layer0_outputs(913);
    outputs(6973) <= not(layer0_outputs(192));
    outputs(6974) <= layer0_outputs(7220);
    outputs(6975) <= layer0_outputs(2674);
    outputs(6976) <= (layer0_outputs(9568)) and not (layer0_outputs(3531));
    outputs(6977) <= not(layer0_outputs(5846));
    outputs(6978) <= (layer0_outputs(9893)) and not (layer0_outputs(6227));
    outputs(6979) <= not((layer0_outputs(5179)) or (layer0_outputs(7669)));
    outputs(6980) <= not((layer0_outputs(8414)) or (layer0_outputs(5435)));
    outputs(6981) <= layer0_outputs(2330);
    outputs(6982) <= not(layer0_outputs(6044));
    outputs(6983) <= (layer0_outputs(7009)) and not (layer0_outputs(9812));
    outputs(6984) <= not((layer0_outputs(730)) and (layer0_outputs(3491)));
    outputs(6985) <= (layer0_outputs(8697)) and (layer0_outputs(4663));
    outputs(6986) <= not(layer0_outputs(8509));
    outputs(6987) <= layer0_outputs(6185);
    outputs(6988) <= layer0_outputs(6384);
    outputs(6989) <= not(layer0_outputs(7817));
    outputs(6990) <= not(layer0_outputs(8223));
    outputs(6991) <= layer0_outputs(6138);
    outputs(6992) <= not(layer0_outputs(10127)) or (layer0_outputs(3712));
    outputs(6993) <= layer0_outputs(5250);
    outputs(6994) <= not(layer0_outputs(1692));
    outputs(6995) <= not((layer0_outputs(8525)) or (layer0_outputs(5614)));
    outputs(6996) <= not(layer0_outputs(867));
    outputs(6997) <= (layer0_outputs(7289)) xor (layer0_outputs(5742));
    outputs(6998) <= layer0_outputs(1073);
    outputs(6999) <= not(layer0_outputs(3793));
    outputs(7000) <= (layer0_outputs(456)) and (layer0_outputs(4799));
    outputs(7001) <= not(layer0_outputs(9845)) or (layer0_outputs(950));
    outputs(7002) <= not((layer0_outputs(8095)) xor (layer0_outputs(2585)));
    outputs(7003) <= (layer0_outputs(6588)) xor (layer0_outputs(7176));
    outputs(7004) <= not(layer0_outputs(5695));
    outputs(7005) <= not((layer0_outputs(3476)) or (layer0_outputs(4677)));
    outputs(7006) <= layer0_outputs(3352);
    outputs(7007) <= (layer0_outputs(2953)) and not (layer0_outputs(363));
    outputs(7008) <= layer0_outputs(9863);
    outputs(7009) <= not((layer0_outputs(1283)) and (layer0_outputs(4399)));
    outputs(7010) <= layer0_outputs(7501);
    outputs(7011) <= not(layer0_outputs(5642));
    outputs(7012) <= layer0_outputs(2209);
    outputs(7013) <= (layer0_outputs(2667)) and (layer0_outputs(2126));
    outputs(7014) <= not((layer0_outputs(5854)) xor (layer0_outputs(1790)));
    outputs(7015) <= (layer0_outputs(6947)) and not (layer0_outputs(10067));
    outputs(7016) <= (layer0_outputs(6970)) and not (layer0_outputs(4819));
    outputs(7017) <= layer0_outputs(6491);
    outputs(7018) <= (layer0_outputs(1970)) and not (layer0_outputs(309));
    outputs(7019) <= not((layer0_outputs(6622)) xor (layer0_outputs(9613)));
    outputs(7020) <= (layer0_outputs(7407)) xor (layer0_outputs(5921));
    outputs(7021) <= not(layer0_outputs(1276));
    outputs(7022) <= (layer0_outputs(7668)) xor (layer0_outputs(8524));
    outputs(7023) <= not((layer0_outputs(4156)) xor (layer0_outputs(3909)));
    outputs(7024) <= (layer0_outputs(6424)) xor (layer0_outputs(7330));
    outputs(7025) <= not(layer0_outputs(3709));
    outputs(7026) <= not(layer0_outputs(8311));
    outputs(7027) <= not(layer0_outputs(994)) or (layer0_outputs(308));
    outputs(7028) <= not((layer0_outputs(4518)) or (layer0_outputs(2665)));
    outputs(7029) <= (layer0_outputs(9919)) xor (layer0_outputs(1054));
    outputs(7030) <= (layer0_outputs(4928)) xor (layer0_outputs(4475));
    outputs(7031) <= layer0_outputs(5428);
    outputs(7032) <= (layer0_outputs(7329)) and not (layer0_outputs(8558));
    outputs(7033) <= not((layer0_outputs(8064)) and (layer0_outputs(1071)));
    outputs(7034) <= not(layer0_outputs(2491));
    outputs(7035) <= not(layer0_outputs(9658));
    outputs(7036) <= not(layer0_outputs(2843));
    outputs(7037) <= not((layer0_outputs(7688)) or (layer0_outputs(6205)));
    outputs(7038) <= not((layer0_outputs(3632)) and (layer0_outputs(7058)));
    outputs(7039) <= layer0_outputs(6762);
    outputs(7040) <= (layer0_outputs(9761)) and (layer0_outputs(2974));
    outputs(7041) <= not(layer0_outputs(679));
    outputs(7042) <= layer0_outputs(9073);
    outputs(7043) <= layer0_outputs(7101);
    outputs(7044) <= layer0_outputs(4461);
    outputs(7045) <= (layer0_outputs(6780)) or (layer0_outputs(9875));
    outputs(7046) <= (layer0_outputs(7860)) and (layer0_outputs(429));
    outputs(7047) <= not((layer0_outputs(489)) or (layer0_outputs(8967)));
    outputs(7048) <= layer0_outputs(2273);
    outputs(7049) <= not(layer0_outputs(3625));
    outputs(7050) <= not((layer0_outputs(2876)) or (layer0_outputs(7792)));
    outputs(7051) <= (layer0_outputs(2461)) and (layer0_outputs(1504));
    outputs(7052) <= not(layer0_outputs(2817));
    outputs(7053) <= not((layer0_outputs(1459)) or (layer0_outputs(10013)));
    outputs(7054) <= layer0_outputs(721);
    outputs(7055) <= (layer0_outputs(4610)) and not (layer0_outputs(10136));
    outputs(7056) <= layer0_outputs(1219);
    outputs(7057) <= not((layer0_outputs(670)) and (layer0_outputs(1129)));
    outputs(7058) <= not(layer0_outputs(9178));
    outputs(7059) <= (layer0_outputs(9720)) and not (layer0_outputs(5292));
    outputs(7060) <= (layer0_outputs(10041)) xor (layer0_outputs(672));
    outputs(7061) <= layer0_outputs(541);
    outputs(7062) <= (layer0_outputs(7510)) and not (layer0_outputs(6329));
    outputs(7063) <= (layer0_outputs(9799)) and (layer0_outputs(1768));
    outputs(7064) <= layer0_outputs(642);
    outputs(7065) <= not((layer0_outputs(8196)) and (layer0_outputs(8478)));
    outputs(7066) <= not(layer0_outputs(5706));
    outputs(7067) <= layer0_outputs(9032);
    outputs(7068) <= (layer0_outputs(9129)) and (layer0_outputs(292));
    outputs(7069) <= not(layer0_outputs(1778));
    outputs(7070) <= layer0_outputs(6912);
    outputs(7071) <= not((layer0_outputs(4784)) and (layer0_outputs(9536)));
    outputs(7072) <= layer0_outputs(3782);
    outputs(7073) <= not(layer0_outputs(7638));
    outputs(7074) <= layer0_outputs(7361);
    outputs(7075) <= not((layer0_outputs(6926)) and (layer0_outputs(1810)));
    outputs(7076) <= (layer0_outputs(5974)) or (layer0_outputs(2059));
    outputs(7077) <= (layer0_outputs(5273)) xor (layer0_outputs(4182));
    outputs(7078) <= not(layer0_outputs(8130));
    outputs(7079) <= not(layer0_outputs(1621));
    outputs(7080) <= not(layer0_outputs(2423));
    outputs(7081) <= not((layer0_outputs(2485)) xor (layer0_outputs(3401)));
    outputs(7082) <= not(layer0_outputs(1943));
    outputs(7083) <= (layer0_outputs(4831)) and not (layer0_outputs(4412));
    outputs(7084) <= (layer0_outputs(9799)) and not (layer0_outputs(6359));
    outputs(7085) <= layer0_outputs(8736);
    outputs(7086) <= not(layer0_outputs(3313));
    outputs(7087) <= (layer0_outputs(10168)) and not (layer0_outputs(1962));
    outputs(7088) <= not(layer0_outputs(313));
    outputs(7089) <= not(layer0_outputs(3148));
    outputs(7090) <= (layer0_outputs(3776)) and not (layer0_outputs(3326));
    outputs(7091) <= (layer0_outputs(793)) xor (layer0_outputs(8304));
    outputs(7092) <= layer0_outputs(8074);
    outputs(7093) <= not((layer0_outputs(4804)) and (layer0_outputs(7072)));
    outputs(7094) <= not((layer0_outputs(3971)) or (layer0_outputs(9043)));
    outputs(7095) <= not(layer0_outputs(4426));
    outputs(7096) <= not(layer0_outputs(1128)) or (layer0_outputs(3122));
    outputs(7097) <= (layer0_outputs(5004)) and not (layer0_outputs(3441));
    outputs(7098) <= not((layer0_outputs(7790)) and (layer0_outputs(2188)));
    outputs(7099) <= (layer0_outputs(10154)) or (layer0_outputs(9203));
    outputs(7100) <= not(layer0_outputs(296)) or (layer0_outputs(3089));
    outputs(7101) <= not(layer0_outputs(7759));
    outputs(7102) <= not((layer0_outputs(7393)) or (layer0_outputs(347)));
    outputs(7103) <= not((layer0_outputs(9833)) or (layer0_outputs(8284)));
    outputs(7104) <= not(layer0_outputs(9122)) or (layer0_outputs(3893));
    outputs(7105) <= layer0_outputs(5585);
    outputs(7106) <= (layer0_outputs(6175)) and not (layer0_outputs(2106));
    outputs(7107) <= not(layer0_outputs(135));
    outputs(7108) <= (layer0_outputs(8318)) and not (layer0_outputs(1440));
    outputs(7109) <= layer0_outputs(3390);
    outputs(7110) <= not(layer0_outputs(786));
    outputs(7111) <= layer0_outputs(2105);
    outputs(7112) <= (layer0_outputs(2648)) and not (layer0_outputs(6901));
    outputs(7113) <= not(layer0_outputs(8295)) or (layer0_outputs(8373));
    outputs(7114) <= layer0_outputs(6716);
    outputs(7115) <= not((layer0_outputs(1981)) and (layer0_outputs(7856)));
    outputs(7116) <= (layer0_outputs(3119)) and not (layer0_outputs(646));
    outputs(7117) <= not((layer0_outputs(3028)) xor (layer0_outputs(3660)));
    outputs(7118) <= (layer0_outputs(2421)) xor (layer0_outputs(8999));
    outputs(7119) <= (layer0_outputs(1706)) xor (layer0_outputs(4871));
    outputs(7120) <= not(layer0_outputs(8905));
    outputs(7121) <= not(layer0_outputs(3055));
    outputs(7122) <= layer0_outputs(7678);
    outputs(7123) <= (layer0_outputs(6689)) and not (layer0_outputs(4960));
    outputs(7124) <= layer0_outputs(9378);
    outputs(7125) <= not(layer0_outputs(3780));
    outputs(7126) <= not(layer0_outputs(7509));
    outputs(7127) <= (layer0_outputs(2530)) or (layer0_outputs(2154));
    outputs(7128) <= (layer0_outputs(2679)) or (layer0_outputs(8390));
    outputs(7129) <= not(layer0_outputs(3063));
    outputs(7130) <= (layer0_outputs(3237)) and (layer0_outputs(320));
    outputs(7131) <= layer0_outputs(7171);
    outputs(7132) <= not(layer0_outputs(3585));
    outputs(7133) <= not(layer0_outputs(8412));
    outputs(7134) <= (layer0_outputs(3595)) and not (layer0_outputs(8649));
    outputs(7135) <= not((layer0_outputs(10094)) and (layer0_outputs(215)));
    outputs(7136) <= not(layer0_outputs(5255));
    outputs(7137) <= (layer0_outputs(5892)) and (layer0_outputs(1454));
    outputs(7138) <= (layer0_outputs(5690)) and not (layer0_outputs(3415));
    outputs(7139) <= layer0_outputs(137);
    outputs(7140) <= not((layer0_outputs(2440)) or (layer0_outputs(5326)));
    outputs(7141) <= layer0_outputs(5760);
    outputs(7142) <= not((layer0_outputs(1338)) or (layer0_outputs(2993)));
    outputs(7143) <= (layer0_outputs(9059)) and not (layer0_outputs(7124));
    outputs(7144) <= not(layer0_outputs(6562));
    outputs(7145) <= (layer0_outputs(4387)) and not (layer0_outputs(6468));
    outputs(7146) <= not(layer0_outputs(1178));
    outputs(7147) <= layer0_outputs(7593);
    outputs(7148) <= not(layer0_outputs(4282));
    outputs(7149) <= (layer0_outputs(4763)) and not (layer0_outputs(7127));
    outputs(7150) <= (layer0_outputs(7008)) and not (layer0_outputs(10108));
    outputs(7151) <= not(layer0_outputs(1221));
    outputs(7152) <= layer0_outputs(4494);
    outputs(7153) <= (layer0_outputs(8738)) and not (layer0_outputs(10136));
    outputs(7154) <= (layer0_outputs(5342)) xor (layer0_outputs(7209));
    outputs(7155) <= layer0_outputs(2373);
    outputs(7156) <= not((layer0_outputs(4960)) or (layer0_outputs(448)));
    outputs(7157) <= (layer0_outputs(7659)) and not (layer0_outputs(4711));
    outputs(7158) <= layer0_outputs(7507);
    outputs(7159) <= not(layer0_outputs(8654)) or (layer0_outputs(377));
    outputs(7160) <= layer0_outputs(7316);
    outputs(7161) <= (layer0_outputs(1824)) and not (layer0_outputs(8217));
    outputs(7162) <= not((layer0_outputs(3376)) xor (layer0_outputs(4609)));
    outputs(7163) <= not(layer0_outputs(3224));
    outputs(7164) <= not(layer0_outputs(2285));
    outputs(7165) <= not((layer0_outputs(1234)) or (layer0_outputs(9558)));
    outputs(7166) <= (layer0_outputs(9773)) and (layer0_outputs(4584));
    outputs(7167) <= not((layer0_outputs(4248)) xor (layer0_outputs(7239)));
    outputs(7168) <= (layer0_outputs(1716)) and not (layer0_outputs(8184));
    outputs(7169) <= (layer0_outputs(9633)) and not (layer0_outputs(4062));
    outputs(7170) <= layer0_outputs(2543);
    outputs(7171) <= not(layer0_outputs(3072)) or (layer0_outputs(2920));
    outputs(7172) <= (layer0_outputs(6047)) and not (layer0_outputs(5552));
    outputs(7173) <= not((layer0_outputs(9612)) and (layer0_outputs(8034)));
    outputs(7174) <= layer0_outputs(8716);
    outputs(7175) <= not(layer0_outputs(8143));
    outputs(7176) <= not(layer0_outputs(494));
    outputs(7177) <= not((layer0_outputs(1717)) xor (layer0_outputs(5697)));
    outputs(7178) <= layer0_outputs(4547);
    outputs(7179) <= not(layer0_outputs(1627));
    outputs(7180) <= not(layer0_outputs(3705));
    outputs(7181) <= layer0_outputs(8495);
    outputs(7182) <= not((layer0_outputs(9124)) xor (layer0_outputs(6204)));
    outputs(7183) <= (layer0_outputs(5281)) and not (layer0_outputs(10080));
    outputs(7184) <= layer0_outputs(4488);
    outputs(7185) <= (layer0_outputs(7882)) and not (layer0_outputs(3456));
    outputs(7186) <= not(layer0_outputs(1049));
    outputs(7187) <= not(layer0_outputs(1596));
    outputs(7188) <= layer0_outputs(4700);
    outputs(7189) <= not(layer0_outputs(4020));
    outputs(7190) <= layer0_outputs(7644);
    outputs(7191) <= not((layer0_outputs(3575)) or (layer0_outputs(1199)));
    outputs(7192) <= (layer0_outputs(9948)) and not (layer0_outputs(8471));
    outputs(7193) <= (layer0_outputs(3661)) and (layer0_outputs(9737));
    outputs(7194) <= layer0_outputs(9923);
    outputs(7195) <= not(layer0_outputs(5623));
    outputs(7196) <= not(layer0_outputs(9655));
    outputs(7197) <= not(layer0_outputs(463));
    outputs(7198) <= (layer0_outputs(8581)) and (layer0_outputs(5062));
    outputs(7199) <= not(layer0_outputs(6682));
    outputs(7200) <= (layer0_outputs(4559)) or (layer0_outputs(6087));
    outputs(7201) <= not((layer0_outputs(2669)) or (layer0_outputs(39)));
    outputs(7202) <= layer0_outputs(476);
    outputs(7203) <= (layer0_outputs(5997)) and not (layer0_outputs(5231));
    outputs(7204) <= (layer0_outputs(5885)) and (layer0_outputs(283));
    outputs(7205) <= layer0_outputs(4814);
    outputs(7206) <= layer0_outputs(5418);
    outputs(7207) <= layer0_outputs(8834);
    outputs(7208) <= layer0_outputs(6729);
    outputs(7209) <= (layer0_outputs(261)) and not (layer0_outputs(802));
    outputs(7210) <= (layer0_outputs(9559)) xor (layer0_outputs(5659));
    outputs(7211) <= not((layer0_outputs(298)) or (layer0_outputs(9470)));
    outputs(7212) <= not(layer0_outputs(328));
    outputs(7213) <= layer0_outputs(8683);
    outputs(7214) <= not((layer0_outputs(8242)) and (layer0_outputs(6935)));
    outputs(7215) <= (layer0_outputs(670)) and not (layer0_outputs(8557));
    outputs(7216) <= not((layer0_outputs(9831)) or (layer0_outputs(5080)));
    outputs(7217) <= layer0_outputs(6397);
    outputs(7218) <= (layer0_outputs(6161)) and not (layer0_outputs(2249));
    outputs(7219) <= not((layer0_outputs(9648)) xor (layer0_outputs(5043)));
    outputs(7220) <= layer0_outputs(2363);
    outputs(7221) <= (layer0_outputs(5116)) and not (layer0_outputs(6271));
    outputs(7222) <= not((layer0_outputs(3508)) and (layer0_outputs(8448)));
    outputs(7223) <= layer0_outputs(4995);
    outputs(7224) <= not(layer0_outputs(3174));
    outputs(7225) <= (layer0_outputs(3649)) xor (layer0_outputs(2289));
    outputs(7226) <= layer0_outputs(6482);
    outputs(7227) <= not((layer0_outputs(8388)) and (layer0_outputs(6183)));
    outputs(7228) <= (layer0_outputs(8990)) and (layer0_outputs(5019));
    outputs(7229) <= (layer0_outputs(1726)) or (layer0_outputs(6945));
    outputs(7230) <= not((layer0_outputs(2810)) xor (layer0_outputs(3628)));
    outputs(7231) <= not((layer0_outputs(6951)) or (layer0_outputs(2723)));
    outputs(7232) <= not((layer0_outputs(634)) and (layer0_outputs(4604)));
    outputs(7233) <= not((layer0_outputs(2213)) or (layer0_outputs(1147)));
    outputs(7234) <= layer0_outputs(7781);
    outputs(7235) <= not((layer0_outputs(10083)) or (layer0_outputs(3350)));
    outputs(7236) <= not((layer0_outputs(9001)) or (layer0_outputs(6565)));
    outputs(7237) <= layer0_outputs(2930);
    outputs(7238) <= layer0_outputs(2866);
    outputs(7239) <= not(layer0_outputs(7772));
    outputs(7240) <= layer0_outputs(7254);
    outputs(7241) <= (layer0_outputs(6730)) xor (layer0_outputs(3757));
    outputs(7242) <= not(layer0_outputs(5542)) or (layer0_outputs(625));
    outputs(7243) <= layer0_outputs(1245);
    outputs(7244) <= not(layer0_outputs(1765));
    outputs(7245) <= (layer0_outputs(4530)) xor (layer0_outputs(4647));
    outputs(7246) <= layer0_outputs(8812);
    outputs(7247) <= (layer0_outputs(6839)) xor (layer0_outputs(3582));
    outputs(7248) <= layer0_outputs(3498);
    outputs(7249) <= (layer0_outputs(5557)) and not (layer0_outputs(877));
    outputs(7250) <= not((layer0_outputs(2495)) xor (layer0_outputs(5931)));
    outputs(7251) <= (layer0_outputs(6513)) and (layer0_outputs(9215));
    outputs(7252) <= (layer0_outputs(973)) and not (layer0_outputs(5405));
    outputs(7253) <= not(layer0_outputs(456));
    outputs(7254) <= layer0_outputs(349);
    outputs(7255) <= (layer0_outputs(4469)) and (layer0_outputs(6188));
    outputs(7256) <= not((layer0_outputs(10167)) xor (layer0_outputs(330)));
    outputs(7257) <= layer0_outputs(4723);
    outputs(7258) <= (layer0_outputs(8234)) and (layer0_outputs(8041));
    outputs(7259) <= (layer0_outputs(9882)) and (layer0_outputs(4278));
    outputs(7260) <= layer0_outputs(2223);
    outputs(7261) <= (layer0_outputs(8547)) or (layer0_outputs(384));
    outputs(7262) <= (layer0_outputs(6514)) and not (layer0_outputs(4068));
    outputs(7263) <= not((layer0_outputs(2135)) xor (layer0_outputs(590)));
    outputs(7264) <= not(layer0_outputs(10168)) or (layer0_outputs(8973));
    outputs(7265) <= not(layer0_outputs(7581));
    outputs(7266) <= not((layer0_outputs(3927)) xor (layer0_outputs(986)));
    outputs(7267) <= not(layer0_outputs(7905));
    outputs(7268) <= layer0_outputs(1013);
    outputs(7269) <= (layer0_outputs(9872)) xor (layer0_outputs(2824));
    outputs(7270) <= not((layer0_outputs(4529)) xor (layer0_outputs(5730)));
    outputs(7271) <= (layer0_outputs(3131)) and not (layer0_outputs(5879));
    outputs(7272) <= not((layer0_outputs(2217)) xor (layer0_outputs(7240)));
    outputs(7273) <= layer0_outputs(4039);
    outputs(7274) <= (layer0_outputs(1349)) xor (layer0_outputs(9030));
    outputs(7275) <= layer0_outputs(8934);
    outputs(7276) <= (layer0_outputs(9176)) xor (layer0_outputs(4948));
    outputs(7277) <= (layer0_outputs(2473)) or (layer0_outputs(5476));
    outputs(7278) <= layer0_outputs(4294);
    outputs(7279) <= not(layer0_outputs(2461)) or (layer0_outputs(6100));
    outputs(7280) <= (layer0_outputs(643)) and not (layer0_outputs(9462));
    outputs(7281) <= not(layer0_outputs(7771));
    outputs(7282) <= layer0_outputs(7082);
    outputs(7283) <= (layer0_outputs(5356)) and not (layer0_outputs(2209));
    outputs(7284) <= layer0_outputs(6529);
    outputs(7285) <= not((layer0_outputs(1635)) or (layer0_outputs(484)));
    outputs(7286) <= (layer0_outputs(2722)) or (layer0_outputs(10106));
    outputs(7287) <= (layer0_outputs(1881)) xor (layer0_outputs(5457));
    outputs(7288) <= not(layer0_outputs(6223));
    outputs(7289) <= (layer0_outputs(7135)) and (layer0_outputs(285));
    outputs(7290) <= layer0_outputs(6158);
    outputs(7291) <= layer0_outputs(6348);
    outputs(7292) <= layer0_outputs(7769);
    outputs(7293) <= not((layer0_outputs(9538)) xor (layer0_outputs(5784)));
    outputs(7294) <= (layer0_outputs(7293)) or (layer0_outputs(8091));
    outputs(7295) <= layer0_outputs(7859);
    outputs(7296) <= not(layer0_outputs(6717));
    outputs(7297) <= (layer0_outputs(2786)) and not (layer0_outputs(9063));
    outputs(7298) <= layer0_outputs(5877);
    outputs(7299) <= not(layer0_outputs(1946));
    outputs(7300) <= (layer0_outputs(9279)) xor (layer0_outputs(10034));
    outputs(7301) <= (layer0_outputs(6131)) xor (layer0_outputs(6176));
    outputs(7302) <= not(layer0_outputs(5408));
    outputs(7303) <= not((layer0_outputs(1351)) or (layer0_outputs(5407)));
    outputs(7304) <= (layer0_outputs(4425)) xor (layer0_outputs(7055));
    outputs(7305) <= not(layer0_outputs(10107));
    outputs(7306) <= (layer0_outputs(9137)) and not (layer0_outputs(4860));
    outputs(7307) <= (layer0_outputs(5040)) and not (layer0_outputs(9263));
    outputs(7308) <= layer0_outputs(5970);
    outputs(7309) <= not(layer0_outputs(9255));
    outputs(7310) <= layer0_outputs(5790);
    outputs(7311) <= (layer0_outputs(5913)) and not (layer0_outputs(4090));
    outputs(7312) <= layer0_outputs(1750);
    outputs(7313) <= not(layer0_outputs(170));
    outputs(7314) <= not((layer0_outputs(8202)) xor (layer0_outputs(4974)));
    outputs(7315) <= (layer0_outputs(1944)) xor (layer0_outputs(3138));
    outputs(7316) <= not(layer0_outputs(1661)) or (layer0_outputs(5603));
    outputs(7317) <= (layer0_outputs(5773)) xor (layer0_outputs(7525));
    outputs(7318) <= layer0_outputs(9404);
    outputs(7319) <= layer0_outputs(8083);
    outputs(7320) <= (layer0_outputs(5376)) xor (layer0_outputs(4614));
    outputs(7321) <= not((layer0_outputs(8870)) and (layer0_outputs(9214)));
    outputs(7322) <= (layer0_outputs(8596)) and not (layer0_outputs(7932));
    outputs(7323) <= (layer0_outputs(4894)) xor (layer0_outputs(7047));
    outputs(7324) <= (layer0_outputs(9174)) and (layer0_outputs(5701));
    outputs(7325) <= not((layer0_outputs(8986)) xor (layer0_outputs(3263)));
    outputs(7326) <= (layer0_outputs(9195)) and not (layer0_outputs(7494));
    outputs(7327) <= not(layer0_outputs(8648));
    outputs(7328) <= layer0_outputs(8882);
    outputs(7329) <= not(layer0_outputs(2908));
    outputs(7330) <= layer0_outputs(6669);
    outputs(7331) <= not((layer0_outputs(4906)) xor (layer0_outputs(2425)));
    outputs(7332) <= not(layer0_outputs(4756));
    outputs(7333) <= not(layer0_outputs(5038));
    outputs(7334) <= layer0_outputs(10020);
    outputs(7335) <= (layer0_outputs(8263)) and not (layer0_outputs(9136));
    outputs(7336) <= layer0_outputs(290);
    outputs(7337) <= layer0_outputs(1016);
    outputs(7338) <= not(layer0_outputs(1205));
    outputs(7339) <= layer0_outputs(3442);
    outputs(7340) <= not((layer0_outputs(6039)) xor (layer0_outputs(2201)));
    outputs(7341) <= not(layer0_outputs(9752));
    outputs(7342) <= (layer0_outputs(2563)) and (layer0_outputs(72));
    outputs(7343) <= (layer0_outputs(1113)) xor (layer0_outputs(3997));
    outputs(7344) <= layer0_outputs(9815);
    outputs(7345) <= layer0_outputs(696);
    outputs(7346) <= layer0_outputs(5248);
    outputs(7347) <= (layer0_outputs(2384)) xor (layer0_outputs(7350));
    outputs(7348) <= not(layer0_outputs(6004));
    outputs(7349) <= not(layer0_outputs(5898));
    outputs(7350) <= not(layer0_outputs(8664));
    outputs(7351) <= not((layer0_outputs(8181)) xor (layer0_outputs(7607)));
    outputs(7352) <= not(layer0_outputs(3189));
    outputs(7353) <= layer0_outputs(3688);
    outputs(7354) <= not(layer0_outputs(3238));
    outputs(7355) <= not(layer0_outputs(5825));
    outputs(7356) <= layer0_outputs(9964);
    outputs(7357) <= not(layer0_outputs(10170));
    outputs(7358) <= (layer0_outputs(176)) and (layer0_outputs(4554));
    outputs(7359) <= not(layer0_outputs(9916));
    outputs(7360) <= (layer0_outputs(9808)) and (layer0_outputs(667));
    outputs(7361) <= layer0_outputs(1941);
    outputs(7362) <= not((layer0_outputs(4693)) and (layer0_outputs(5831)));
    outputs(7363) <= (layer0_outputs(349)) and not (layer0_outputs(2697));
    outputs(7364) <= layer0_outputs(6603);
    outputs(7365) <= (layer0_outputs(252)) and not (layer0_outputs(5559));
    outputs(7366) <= (layer0_outputs(1230)) xor (layer0_outputs(9097));
    outputs(7367) <= not(layer0_outputs(8770));
    outputs(7368) <= layer0_outputs(9070);
    outputs(7369) <= not((layer0_outputs(7396)) xor (layer0_outputs(645)));
    outputs(7370) <= (layer0_outputs(3522)) and not (layer0_outputs(3020));
    outputs(7371) <= not((layer0_outputs(6526)) xor (layer0_outputs(45)));
    outputs(7372) <= not((layer0_outputs(1197)) xor (layer0_outputs(197)));
    outputs(7373) <= layer0_outputs(1012);
    outputs(7374) <= layer0_outputs(3436);
    outputs(7375) <= layer0_outputs(7432);
    outputs(7376) <= layer0_outputs(1172);
    outputs(7377) <= not(layer0_outputs(6863));
    outputs(7378) <= layer0_outputs(3584);
    outputs(7379) <= (layer0_outputs(887)) and (layer0_outputs(996));
    outputs(7380) <= (layer0_outputs(2136)) and not (layer0_outputs(5583));
    outputs(7381) <= (layer0_outputs(3823)) and not (layer0_outputs(4801));
    outputs(7382) <= not(layer0_outputs(1897));
    outputs(7383) <= layer0_outputs(87);
    outputs(7384) <= not(layer0_outputs(6222));
    outputs(7385) <= layer0_outputs(3996);
    outputs(7386) <= not(layer0_outputs(6094));
    outputs(7387) <= (layer0_outputs(3936)) and (layer0_outputs(5954));
    outputs(7388) <= not(layer0_outputs(5461));
    outputs(7389) <= (layer0_outputs(5139)) or (layer0_outputs(8098));
    outputs(7390) <= not(layer0_outputs(5923));
    outputs(7391) <= not(layer0_outputs(4861));
    outputs(7392) <= not((layer0_outputs(5722)) xor (layer0_outputs(6003)));
    outputs(7393) <= not(layer0_outputs(1968));
    outputs(7394) <= not(layer0_outputs(8989));
    outputs(7395) <= (layer0_outputs(7216)) and not (layer0_outputs(2690));
    outputs(7396) <= (layer0_outputs(10039)) and (layer0_outputs(9455));
    outputs(7397) <= not(layer0_outputs(1711));
    outputs(7398) <= (layer0_outputs(1413)) and not (layer0_outputs(4567));
    outputs(7399) <= not(layer0_outputs(6515)) or (layer0_outputs(8658));
    outputs(7400) <= layer0_outputs(1310);
    outputs(7401) <= not((layer0_outputs(7610)) xor (layer0_outputs(9114)));
    outputs(7402) <= not(layer0_outputs(3430));
    outputs(7403) <= not(layer0_outputs(9982));
    outputs(7404) <= not(layer0_outputs(6716));
    outputs(7405) <= not((layer0_outputs(2580)) xor (layer0_outputs(777)));
    outputs(7406) <= not(layer0_outputs(5908));
    outputs(7407) <= (layer0_outputs(4908)) or (layer0_outputs(6211));
    outputs(7408) <= not(layer0_outputs(501));
    outputs(7409) <= not(layer0_outputs(9211));
    outputs(7410) <= not(layer0_outputs(7954));
    outputs(7411) <= not((layer0_outputs(24)) xor (layer0_outputs(4948)));
    outputs(7412) <= not(layer0_outputs(3373)) or (layer0_outputs(4470));
    outputs(7413) <= layer0_outputs(885);
    outputs(7414) <= (layer0_outputs(2129)) and (layer0_outputs(8559));
    outputs(7415) <= not((layer0_outputs(8624)) and (layer0_outputs(4748)));
    outputs(7416) <= layer0_outputs(4779);
    outputs(7417) <= (layer0_outputs(5945)) xor (layer0_outputs(1717));
    outputs(7418) <= not(layer0_outputs(8513)) or (layer0_outputs(8890));
    outputs(7419) <= not((layer0_outputs(845)) or (layer0_outputs(6938)));
    outputs(7420) <= not(layer0_outputs(2422));
    outputs(7421) <= layer0_outputs(6137);
    outputs(7422) <= not((layer0_outputs(4377)) xor (layer0_outputs(6750)));
    outputs(7423) <= not((layer0_outputs(7606)) or (layer0_outputs(10004)));
    outputs(7424) <= not(layer0_outputs(2244));
    outputs(7425) <= (layer0_outputs(6852)) xor (layer0_outputs(8521));
    outputs(7426) <= layer0_outputs(3026);
    outputs(7427) <= (layer0_outputs(9197)) xor (layer0_outputs(2442));
    outputs(7428) <= layer0_outputs(3641);
    outputs(7429) <= layer0_outputs(6040);
    outputs(7430) <= not((layer0_outputs(3796)) or (layer0_outputs(757)));
    outputs(7431) <= (layer0_outputs(2869)) and not (layer0_outputs(3308));
    outputs(7432) <= (layer0_outputs(9531)) and (layer0_outputs(332));
    outputs(7433) <= layer0_outputs(4376);
    outputs(7434) <= layer0_outputs(5895);
    outputs(7435) <= (layer0_outputs(6856)) and not (layer0_outputs(10097));
    outputs(7436) <= (layer0_outputs(9318)) and not (layer0_outputs(1369));
    outputs(7437) <= (layer0_outputs(8003)) and not (layer0_outputs(3350));
    outputs(7438) <= (layer0_outputs(8451)) or (layer0_outputs(2543));
    outputs(7439) <= not((layer0_outputs(1125)) xor (layer0_outputs(6902)));
    outputs(7440) <= not((layer0_outputs(7804)) xor (layer0_outputs(9857)));
    outputs(7441) <= not(layer0_outputs(2177));
    outputs(7442) <= layer0_outputs(8772);
    outputs(7443) <= not((layer0_outputs(3469)) or (layer0_outputs(10161)));
    outputs(7444) <= not((layer0_outputs(3703)) xor (layer0_outputs(7138)));
    outputs(7445) <= not(layer0_outputs(6775));
    outputs(7446) <= (layer0_outputs(2977)) and not (layer0_outputs(92));
    outputs(7447) <= not(layer0_outputs(8982));
    outputs(7448) <= layer0_outputs(7219);
    outputs(7449) <= (layer0_outputs(3106)) and (layer0_outputs(7223));
    outputs(7450) <= layer0_outputs(8321);
    outputs(7451) <= (layer0_outputs(1453)) and not (layer0_outputs(512));
    outputs(7452) <= layer0_outputs(4854);
    outputs(7453) <= not((layer0_outputs(4175)) or (layer0_outputs(2408)));
    outputs(7454) <= layer0_outputs(8564);
    outputs(7455) <= not((layer0_outputs(8032)) or (layer0_outputs(3905)));
    outputs(7456) <= not(layer0_outputs(957));
    outputs(7457) <= layer0_outputs(9206);
    outputs(7458) <= not((layer0_outputs(7487)) xor (layer0_outputs(4673)));
    outputs(7459) <= (layer0_outputs(6158)) and (layer0_outputs(844));
    outputs(7460) <= (layer0_outputs(7459)) and (layer0_outputs(1302));
    outputs(7461) <= (layer0_outputs(5872)) xor (layer0_outputs(651));
    outputs(7462) <= (layer0_outputs(9020)) xor (layer0_outputs(6141));
    outputs(7463) <= not((layer0_outputs(5747)) xor (layer0_outputs(7399)));
    outputs(7464) <= layer0_outputs(6160);
    outputs(7465) <= layer0_outputs(2741);
    outputs(7466) <= layer0_outputs(9437);
    outputs(7467) <= (layer0_outputs(1698)) and not (layer0_outputs(9394));
    outputs(7468) <= layer0_outputs(2324);
    outputs(7469) <= not(layer0_outputs(6880));
    outputs(7470) <= layer0_outputs(4569);
    outputs(7471) <= not(layer0_outputs(3497));
    outputs(7472) <= not(layer0_outputs(7797)) or (layer0_outputs(5617));
    outputs(7473) <= layer0_outputs(7450);
    outputs(7474) <= (layer0_outputs(1823)) and not (layer0_outputs(6463));
    outputs(7475) <= not(layer0_outputs(7064));
    outputs(7476) <= not(layer0_outputs(3788)) or (layer0_outputs(4654));
    outputs(7477) <= layer0_outputs(5493);
    outputs(7478) <= (layer0_outputs(8128)) or (layer0_outputs(1577));
    outputs(7479) <= not((layer0_outputs(5477)) xor (layer0_outputs(4337)));
    outputs(7480) <= (layer0_outputs(6256)) and not (layer0_outputs(2264));
    outputs(7481) <= not((layer0_outputs(2261)) xor (layer0_outputs(2156)));
    outputs(7482) <= (layer0_outputs(7010)) or (layer0_outputs(9440));
    outputs(7483) <= (layer0_outputs(4293)) and (layer0_outputs(6187));
    outputs(7484) <= (layer0_outputs(1958)) or (layer0_outputs(2981));
    outputs(7485) <= not((layer0_outputs(5080)) and (layer0_outputs(9481)));
    outputs(7486) <= layer0_outputs(1963);
    outputs(7487) <= layer0_outputs(1488);
    outputs(7488) <= layer0_outputs(1836);
    outputs(7489) <= (layer0_outputs(8443)) xor (layer0_outputs(8423));
    outputs(7490) <= (layer0_outputs(4471)) and not (layer0_outputs(6947));
    outputs(7491) <= layer0_outputs(6998);
    outputs(7492) <= (layer0_outputs(9505)) or (layer0_outputs(1708));
    outputs(7493) <= not((layer0_outputs(114)) or (layer0_outputs(5431)));
    outputs(7494) <= (layer0_outputs(1164)) xor (layer0_outputs(9217));
    outputs(7495) <= not(layer0_outputs(1335));
    outputs(7496) <= (layer0_outputs(6422)) xor (layer0_outputs(9016));
    outputs(7497) <= not((layer0_outputs(7461)) xor (layer0_outputs(7608)));
    outputs(7498) <= layer0_outputs(9924);
    outputs(7499) <= (layer0_outputs(2966)) and not (layer0_outputs(9320));
    outputs(7500) <= not(layer0_outputs(5748));
    outputs(7501) <= layer0_outputs(306);
    outputs(7502) <= layer0_outputs(3108);
    outputs(7503) <= not(layer0_outputs(2454));
    outputs(7504) <= layer0_outputs(2692);
    outputs(7505) <= (layer0_outputs(3843)) and (layer0_outputs(1463));
    outputs(7506) <= (layer0_outputs(2526)) xor (layer0_outputs(3507));
    outputs(7507) <= layer0_outputs(2510);
    outputs(7508) <= (layer0_outputs(2447)) xor (layer0_outputs(5870));
    outputs(7509) <= (layer0_outputs(4269)) and (layer0_outputs(2917));
    outputs(7510) <= (layer0_outputs(9115)) xor (layer0_outputs(4245));
    outputs(7511) <= not((layer0_outputs(1690)) xor (layer0_outputs(9698)));
    outputs(7512) <= (layer0_outputs(3790)) xor (layer0_outputs(9754));
    outputs(7513) <= not((layer0_outputs(4060)) or (layer0_outputs(3771)));
    outputs(7514) <= layer0_outputs(5888);
    outputs(7515) <= (layer0_outputs(5459)) and not (layer0_outputs(1466));
    outputs(7516) <= layer0_outputs(3418);
    outputs(7517) <= not(layer0_outputs(4136));
    outputs(7518) <= not(layer0_outputs(5048));
    outputs(7519) <= (layer0_outputs(1634)) xor (layer0_outputs(2906));
    outputs(7520) <= not(layer0_outputs(8113));
    outputs(7521) <= not(layer0_outputs(3532));
    outputs(7522) <= not((layer0_outputs(9615)) xor (layer0_outputs(10203)));
    outputs(7523) <= not((layer0_outputs(1025)) or (layer0_outputs(9606)));
    outputs(7524) <= not((layer0_outputs(5484)) or (layer0_outputs(9716)));
    outputs(7525) <= layer0_outputs(1314);
    outputs(7526) <= (layer0_outputs(6728)) and (layer0_outputs(8078));
    outputs(7527) <= not((layer0_outputs(10027)) and (layer0_outputs(2750)));
    outputs(7528) <= (layer0_outputs(5349)) and not (layer0_outputs(4861));
    outputs(7529) <= not(layer0_outputs(6139));
    outputs(7530) <= (layer0_outputs(486)) and (layer0_outputs(5323));
    outputs(7531) <= (layer0_outputs(7901)) and (layer0_outputs(3615));
    outputs(7532) <= (layer0_outputs(7099)) and not (layer0_outputs(2923));
    outputs(7533) <= not(layer0_outputs(7052));
    outputs(7534) <= (layer0_outputs(8606)) or (layer0_outputs(10101));
    outputs(7535) <= (layer0_outputs(599)) and not (layer0_outputs(8585));
    outputs(7536) <= (layer0_outputs(6473)) and (layer0_outputs(6129));
    outputs(7537) <= not(layer0_outputs(4546));
    outputs(7538) <= not(layer0_outputs(8932));
    outputs(7539) <= not((layer0_outputs(4062)) or (layer0_outputs(4902)));
    outputs(7540) <= not(layer0_outputs(9336)) or (layer0_outputs(8790));
    outputs(7541) <= (layer0_outputs(4178)) xor (layer0_outputs(4484));
    outputs(7542) <= layer0_outputs(5534);
    outputs(7543) <= (layer0_outputs(147)) and (layer0_outputs(4992));
    outputs(7544) <= (layer0_outputs(10200)) and not (layer0_outputs(362));
    outputs(7545) <= (layer0_outputs(10089)) xor (layer0_outputs(892));
    outputs(7546) <= not(layer0_outputs(7442));
    outputs(7547) <= layer0_outputs(4785);
    outputs(7548) <= (layer0_outputs(2077)) xor (layer0_outputs(417));
    outputs(7549) <= not(layer0_outputs(8873)) or (layer0_outputs(8029));
    outputs(7550) <= not(layer0_outputs(2250));
    outputs(7551) <= layer0_outputs(1087);
    outputs(7552) <= not(layer0_outputs(668));
    outputs(7553) <= (layer0_outputs(3691)) xor (layer0_outputs(9509));
    outputs(7554) <= not((layer0_outputs(4991)) xor (layer0_outputs(8646)));
    outputs(7555) <= layer0_outputs(9119);
    outputs(7556) <= (layer0_outputs(1962)) xor (layer0_outputs(2113));
    outputs(7557) <= layer0_outputs(8787);
    outputs(7558) <= not(layer0_outputs(4619)) or (layer0_outputs(495));
    outputs(7559) <= not(layer0_outputs(7627));
    outputs(7560) <= (layer0_outputs(766)) and not (layer0_outputs(4649));
    outputs(7561) <= not((layer0_outputs(630)) xor (layer0_outputs(1347)));
    outputs(7562) <= not(layer0_outputs(3954));
    outputs(7563) <= not((layer0_outputs(2990)) xor (layer0_outputs(5612)));
    outputs(7564) <= not(layer0_outputs(156));
    outputs(7565) <= layer0_outputs(8781);
    outputs(7566) <= layer0_outputs(9331);
    outputs(7567) <= (layer0_outputs(9995)) xor (layer0_outputs(10193));
    outputs(7568) <= layer0_outputs(904);
    outputs(7569) <= not((layer0_outputs(3802)) or (layer0_outputs(3920)));
    outputs(7570) <= not(layer0_outputs(3023));
    outputs(7571) <= layer0_outputs(128);
    outputs(7572) <= (layer0_outputs(4190)) and not (layer0_outputs(3255));
    outputs(7573) <= not(layer0_outputs(6116)) or (layer0_outputs(2246));
    outputs(7574) <= not((layer0_outputs(5155)) or (layer0_outputs(2151)));
    outputs(7575) <= not((layer0_outputs(7593)) or (layer0_outputs(3225)));
    outputs(7576) <= layer0_outputs(1116);
    outputs(7577) <= layer0_outputs(6340);
    outputs(7578) <= not(layer0_outputs(7374));
    outputs(7579) <= not(layer0_outputs(3915)) or (layer0_outputs(4231));
    outputs(7580) <= not(layer0_outputs(9669));
    outputs(7581) <= not((layer0_outputs(4001)) or (layer0_outputs(8630)));
    outputs(7582) <= (layer0_outputs(2093)) xor (layer0_outputs(5982));
    outputs(7583) <= not(layer0_outputs(907));
    outputs(7584) <= not((layer0_outputs(5976)) xor (layer0_outputs(5584)));
    outputs(7585) <= (layer0_outputs(5281)) and not (layer0_outputs(482));
    outputs(7586) <= layer0_outputs(5132);
    outputs(7587) <= not(layer0_outputs(10203));
    outputs(7588) <= not((layer0_outputs(1291)) and (layer0_outputs(5446)));
    outputs(7589) <= not(layer0_outputs(5118));
    outputs(7590) <= not(layer0_outputs(4934));
    outputs(7591) <= not((layer0_outputs(7470)) and (layer0_outputs(411)));
    outputs(7592) <= (layer0_outputs(2677)) and not (layer0_outputs(6763));
    outputs(7593) <= not(layer0_outputs(5638));
    outputs(7594) <= layer0_outputs(2052);
    outputs(7595) <= layer0_outputs(8950);
    outputs(7596) <= (layer0_outputs(7697)) and not (layer0_outputs(10186));
    outputs(7597) <= not((layer0_outputs(7049)) or (layer0_outputs(1436)));
    outputs(7598) <= layer0_outputs(5947);
    outputs(7599) <= layer0_outputs(9368);
    outputs(7600) <= layer0_outputs(4778);
    outputs(7601) <= not(layer0_outputs(1350));
    outputs(7602) <= not(layer0_outputs(9472));
    outputs(7603) <= layer0_outputs(4490);
    outputs(7604) <= not((layer0_outputs(7918)) or (layer0_outputs(8117)));
    outputs(7605) <= (layer0_outputs(7265)) xor (layer0_outputs(7674));
    outputs(7606) <= not((layer0_outputs(513)) xor (layer0_outputs(9886)));
    outputs(7607) <= layer0_outputs(8626);
    outputs(7608) <= not(layer0_outputs(8621)) or (layer0_outputs(9253));
    outputs(7609) <= (layer0_outputs(1638)) and not (layer0_outputs(3171));
    outputs(7610) <= (layer0_outputs(9273)) and not (layer0_outputs(10040));
    outputs(7611) <= not(layer0_outputs(2058));
    outputs(7612) <= not((layer0_outputs(6104)) xor (layer0_outputs(4403)));
    outputs(7613) <= not((layer0_outputs(6873)) xor (layer0_outputs(6290)));
    outputs(7614) <= not((layer0_outputs(203)) or (layer0_outputs(10163)));
    outputs(7615) <= not((layer0_outputs(6822)) or (layer0_outputs(8956)));
    outputs(7616) <= (layer0_outputs(3633)) and not (layer0_outputs(2002));
    outputs(7617) <= (layer0_outputs(6496)) or (layer0_outputs(834));
    outputs(7618) <= (layer0_outputs(8649)) and not (layer0_outputs(789));
    outputs(7619) <= not((layer0_outputs(1365)) or (layer0_outputs(7720)));
    outputs(7620) <= not(layer0_outputs(5905));
    outputs(7621) <= not(layer0_outputs(2748));
    outputs(7622) <= not(layer0_outputs(8664));
    outputs(7623) <= not((layer0_outputs(6420)) xor (layer0_outputs(3228)));
    outputs(7624) <= not(layer0_outputs(3509));
    outputs(7625) <= not(layer0_outputs(3494));
    outputs(7626) <= layer0_outputs(8440);
    outputs(7627) <= not(layer0_outputs(3433));
    outputs(7628) <= not(layer0_outputs(6230));
    outputs(7629) <= not((layer0_outputs(5302)) xor (layer0_outputs(2760)));
    outputs(7630) <= not(layer0_outputs(9665));
    outputs(7631) <= (layer0_outputs(3105)) xor (layer0_outputs(1039));
    outputs(7632) <= not(layer0_outputs(6504));
    outputs(7633) <= layer0_outputs(9829);
    outputs(7634) <= layer0_outputs(5622);
    outputs(7635) <= (layer0_outputs(5150)) and (layer0_outputs(5012));
    outputs(7636) <= (layer0_outputs(3953)) xor (layer0_outputs(4874));
    outputs(7637) <= (layer0_outputs(6780)) and not (layer0_outputs(4765));
    outputs(7638) <= layer0_outputs(5811);
    outputs(7639) <= (layer0_outputs(936)) and not (layer0_outputs(1847));
    outputs(7640) <= layer0_outputs(4436);
    outputs(7641) <= (layer0_outputs(8363)) or (layer0_outputs(1609));
    outputs(7642) <= (layer0_outputs(2035)) and not (layer0_outputs(6605));
    outputs(7643) <= layer0_outputs(5794);
    outputs(7644) <= not((layer0_outputs(6420)) xor (layer0_outputs(4839)));
    outputs(7645) <= layer0_outputs(543);
    outputs(7646) <= (layer0_outputs(7531)) and not (layer0_outputs(1512));
    outputs(7647) <= not(layer0_outputs(8836));
    outputs(7648) <= not((layer0_outputs(8960)) or (layer0_outputs(9736)));
    outputs(7649) <= (layer0_outputs(2167)) xor (layer0_outputs(3568));
    outputs(7650) <= not(layer0_outputs(9399));
    outputs(7651) <= (layer0_outputs(9676)) and (layer0_outputs(6957));
    outputs(7652) <= not((layer0_outputs(2257)) xor (layer0_outputs(1592)));
    outputs(7653) <= layer0_outputs(2525);
    outputs(7654) <= layer0_outputs(7387);
    outputs(7655) <= layer0_outputs(8945);
    outputs(7656) <= (layer0_outputs(6578)) and (layer0_outputs(9222));
    outputs(7657) <= layer0_outputs(400);
    outputs(7658) <= (layer0_outputs(9550)) and (layer0_outputs(2368));
    outputs(7659) <= (layer0_outputs(4035)) and not (layer0_outputs(8628));
    outputs(7660) <= not(layer0_outputs(3003));
    outputs(7661) <= layer0_outputs(9098);
    outputs(7662) <= (layer0_outputs(2169)) and (layer0_outputs(3644));
    outputs(7663) <= not((layer0_outputs(1972)) and (layer0_outputs(4197)));
    outputs(7664) <= not((layer0_outputs(5521)) or (layer0_outputs(9182)));
    outputs(7665) <= not((layer0_outputs(1198)) and (layer0_outputs(7448)));
    outputs(7666) <= not(layer0_outputs(8476));
    outputs(7667) <= not(layer0_outputs(5623));
    outputs(7668) <= not((layer0_outputs(6691)) xor (layer0_outputs(540)));
    outputs(7669) <= (layer0_outputs(8749)) xor (layer0_outputs(7334));
    outputs(7670) <= layer0_outputs(583);
    outputs(7671) <= (layer0_outputs(1058)) xor (layer0_outputs(8492));
    outputs(7672) <= not(layer0_outputs(4532)) or (layer0_outputs(2232));
    outputs(7673) <= layer0_outputs(3337);
    outputs(7674) <= (layer0_outputs(5571)) and not (layer0_outputs(2815));
    outputs(7675) <= not((layer0_outputs(9147)) or (layer0_outputs(6216)));
    outputs(7676) <= (layer0_outputs(9374)) xor (layer0_outputs(3346));
    outputs(7677) <= (layer0_outputs(2293)) and (layer0_outputs(2535));
    outputs(7678) <= not(layer0_outputs(8556)) or (layer0_outputs(1201));
    outputs(7679) <= not(layer0_outputs(7440));
    outputs(7680) <= (layer0_outputs(8717)) xor (layer0_outputs(5865));
    outputs(7681) <= not((layer0_outputs(6671)) xor (layer0_outputs(9647)));
    outputs(7682) <= (layer0_outputs(3752)) and (layer0_outputs(163));
    outputs(7683) <= (layer0_outputs(694)) and not (layer0_outputs(9243));
    outputs(7684) <= not(layer0_outputs(4433));
    outputs(7685) <= layer0_outputs(4025);
    outputs(7686) <= layer0_outputs(78);
    outputs(7687) <= not((layer0_outputs(9820)) xor (layer0_outputs(9196)));
    outputs(7688) <= layer0_outputs(8193);
    outputs(7689) <= (layer0_outputs(1935)) and (layer0_outputs(2340));
    outputs(7690) <= layer0_outputs(5140);
    outputs(7691) <= layer0_outputs(1789);
    outputs(7692) <= layer0_outputs(2033);
    outputs(7693) <= (layer0_outputs(9480)) and (layer0_outputs(3731));
    outputs(7694) <= layer0_outputs(9051);
    outputs(7695) <= (layer0_outputs(4443)) and not (layer0_outputs(8993));
    outputs(7696) <= layer0_outputs(400);
    outputs(7697) <= (layer0_outputs(3737)) xor (layer0_outputs(1776));
    outputs(7698) <= not((layer0_outputs(3569)) xor (layer0_outputs(4640)));
    outputs(7699) <= (layer0_outputs(8285)) and not (layer0_outputs(5355));
    outputs(7700) <= (layer0_outputs(7423)) xor (layer0_outputs(8115));
    outputs(7701) <= (layer0_outputs(1682)) and not (layer0_outputs(9529));
    outputs(7702) <= (layer0_outputs(7936)) xor (layer0_outputs(9240));
    outputs(7703) <= not((layer0_outputs(8936)) xor (layer0_outputs(9993)));
    outputs(7704) <= not(layer0_outputs(3932));
    outputs(7705) <= (layer0_outputs(2942)) and not (layer0_outputs(6883));
    outputs(7706) <= not((layer0_outputs(8404)) or (layer0_outputs(6877)));
    outputs(7707) <= not((layer0_outputs(8129)) or (layer0_outputs(1868)));
    outputs(7708) <= not(layer0_outputs(9735));
    outputs(7709) <= layer0_outputs(6207);
    outputs(7710) <= not(layer0_outputs(7620)) or (layer0_outputs(8533));
    outputs(7711) <= (layer0_outputs(1709)) or (layer0_outputs(1037));
    outputs(7712) <= (layer0_outputs(1507)) xor (layer0_outputs(9437));
    outputs(7713) <= not(layer0_outputs(7585));
    outputs(7714) <= (layer0_outputs(9898)) xor (layer0_outputs(6968));
    outputs(7715) <= (layer0_outputs(1864)) or (layer0_outputs(8746));
    outputs(7716) <= not((layer0_outputs(8815)) or (layer0_outputs(1795)));
    outputs(7717) <= (layer0_outputs(7245)) xor (layer0_outputs(5498));
    outputs(7718) <= (layer0_outputs(2103)) and not (layer0_outputs(6724));
    outputs(7719) <= (layer0_outputs(3224)) xor (layer0_outputs(3994));
    outputs(7720) <= (layer0_outputs(1655)) and not (layer0_outputs(5367));
    outputs(7721) <= (layer0_outputs(2928)) and not (layer0_outputs(3012));
    outputs(7722) <= (layer0_outputs(1606)) and (layer0_outputs(6626));
    outputs(7723) <= not(layer0_outputs(9220));
    outputs(7724) <= not((layer0_outputs(4638)) or (layer0_outputs(5022)));
    outputs(7725) <= not(layer0_outputs(623));
    outputs(7726) <= (layer0_outputs(2395)) xor (layer0_outputs(6100));
    outputs(7727) <= not(layer0_outputs(8993));
    outputs(7728) <= (layer0_outputs(334)) and not (layer0_outputs(10190));
    outputs(7729) <= (layer0_outputs(1428)) and not (layer0_outputs(8156));
    outputs(7730) <= not(layer0_outputs(2464)) or (layer0_outputs(1692));
    outputs(7731) <= not(layer0_outputs(7502));
    outputs(7732) <= layer0_outputs(6061);
    outputs(7733) <= not((layer0_outputs(1371)) and (layer0_outputs(3076)));
    outputs(7734) <= (layer0_outputs(3576)) and not (layer0_outputs(8681));
    outputs(7735) <= (layer0_outputs(7198)) and (layer0_outputs(6697));
    outputs(7736) <= (layer0_outputs(6513)) and (layer0_outputs(9152));
    outputs(7737) <= not(layer0_outputs(2479));
    outputs(7738) <= not(layer0_outputs(2364));
    outputs(7739) <= not((layer0_outputs(1738)) or (layer0_outputs(1900)));
    outputs(7740) <= layer0_outputs(6823);
    outputs(7741) <= (layer0_outputs(7895)) xor (layer0_outputs(2269));
    outputs(7742) <= (layer0_outputs(4689)) and not (layer0_outputs(1686));
    outputs(7743) <= (layer0_outputs(7342)) and not (layer0_outputs(10083));
    outputs(7744) <= (layer0_outputs(3371)) xor (layer0_outputs(5660));
    outputs(7745) <= not(layer0_outputs(4249)) or (layer0_outputs(5659));
    outputs(7746) <= not(layer0_outputs(8889));
    outputs(7747) <= not(layer0_outputs(6167)) or (layer0_outputs(644));
    outputs(7748) <= (layer0_outputs(650)) and (layer0_outputs(10069));
    outputs(7749) <= not((layer0_outputs(7583)) xor (layer0_outputs(955)));
    outputs(7750) <= (layer0_outputs(3910)) and (layer0_outputs(6688));
    outputs(7751) <= (layer0_outputs(5793)) and (layer0_outputs(9172));
    outputs(7752) <= (layer0_outputs(9545)) and (layer0_outputs(8806));
    outputs(7753) <= (layer0_outputs(1117)) or (layer0_outputs(3231));
    outputs(7754) <= (layer0_outputs(4373)) xor (layer0_outputs(7179));
    outputs(7755) <= not(layer0_outputs(5550)) or (layer0_outputs(810));
    outputs(7756) <= layer0_outputs(7038);
    outputs(7757) <= not(layer0_outputs(534));
    outputs(7758) <= (layer0_outputs(6729)) and not (layer0_outputs(180));
    outputs(7759) <= layer0_outputs(9027);
    outputs(7760) <= not(layer0_outputs(9248));
    outputs(7761) <= (layer0_outputs(7180)) and not (layer0_outputs(4416));
    outputs(7762) <= (layer0_outputs(3223)) and (layer0_outputs(2901));
    outputs(7763) <= not(layer0_outputs(5370));
    outputs(7764) <= layer0_outputs(5802);
    outputs(7765) <= not((layer0_outputs(10144)) or (layer0_outputs(5710)));
    outputs(7766) <= layer0_outputs(2350);
    outputs(7767) <= not((layer0_outputs(6455)) or (layer0_outputs(9972)));
    outputs(7768) <= not((layer0_outputs(924)) or (layer0_outputs(8264)));
    outputs(7769) <= not(layer0_outputs(7630));
    outputs(7770) <= (layer0_outputs(3254)) and (layer0_outputs(557));
    outputs(7771) <= layer0_outputs(4818);
    outputs(7772) <= not(layer0_outputs(2558));
    outputs(7773) <= layer0_outputs(5472);
    outputs(7774) <= not(layer0_outputs(9238));
    outputs(7775) <= layer0_outputs(7741);
    outputs(7776) <= not(layer0_outputs(1135));
    outputs(7777) <= (layer0_outputs(9170)) and not (layer0_outputs(4890));
    outputs(7778) <= not((layer0_outputs(778)) xor (layer0_outputs(8108)));
    outputs(7779) <= (layer0_outputs(9821)) and not (layer0_outputs(6443));
    outputs(7780) <= (layer0_outputs(2204)) xor (layer0_outputs(4726));
    outputs(7781) <= (layer0_outputs(8707)) and not (layer0_outputs(6074));
    outputs(7782) <= not(layer0_outputs(1343));
    outputs(7783) <= (layer0_outputs(5547)) xor (layer0_outputs(353));
    outputs(7784) <= not(layer0_outputs(2496));
    outputs(7785) <= (layer0_outputs(6253)) and (layer0_outputs(4396));
    outputs(7786) <= not(layer0_outputs(9235));
    outputs(7787) <= not(layer0_outputs(9623));
    outputs(7788) <= not(layer0_outputs(8422));
    outputs(7789) <= (layer0_outputs(2123)) or (layer0_outputs(2683));
    outputs(7790) <= not(layer0_outputs(272));
    outputs(7791) <= layer0_outputs(7945);
    outputs(7792) <= layer0_outputs(517);
    outputs(7793) <= (layer0_outputs(9296)) and not (layer0_outputs(5037));
    outputs(7794) <= layer0_outputs(4111);
    outputs(7795) <= not((layer0_outputs(1060)) xor (layer0_outputs(6225)));
    outputs(7796) <= layer0_outputs(4434);
    outputs(7797) <= not(layer0_outputs(7205));
    outputs(7798) <= layer0_outputs(4);
    outputs(7799) <= not((layer0_outputs(1195)) or (layer0_outputs(5498)));
    outputs(7800) <= not((layer0_outputs(9765)) xor (layer0_outputs(6542)));
    outputs(7801) <= (layer0_outputs(8059)) and (layer0_outputs(1540));
    outputs(7802) <= (layer0_outputs(512)) xor (layer0_outputs(2321));
    outputs(7803) <= layer0_outputs(5992);
    outputs(7804) <= (layer0_outputs(4126)) and (layer0_outputs(5932));
    outputs(7805) <= not((layer0_outputs(3996)) xor (layer0_outputs(5195)));
    outputs(7806) <= not((layer0_outputs(10239)) xor (layer0_outputs(4816)));
    outputs(7807) <= layer0_outputs(6205);
    outputs(7808) <= layer0_outputs(8057);
    outputs(7809) <= (layer0_outputs(8790)) xor (layer0_outputs(2294));
    outputs(7810) <= not(layer0_outputs(8791));
    outputs(7811) <= layer0_outputs(8872);
    outputs(7812) <= (layer0_outputs(3903)) and not (layer0_outputs(9620));
    outputs(7813) <= not(layer0_outputs(971)) or (layer0_outputs(3161));
    outputs(7814) <= (layer0_outputs(496)) xor (layer0_outputs(3766));
    outputs(7815) <= not(layer0_outputs(9450));
    outputs(7816) <= (layer0_outputs(684)) and not (layer0_outputs(9655));
    outputs(7817) <= not(layer0_outputs(9988));
    outputs(7818) <= (layer0_outputs(7158)) and not (layer0_outputs(4635));
    outputs(7819) <= (layer0_outputs(1333)) and not (layer0_outputs(4052));
    outputs(7820) <= not(layer0_outputs(4005));
    outputs(7821) <= not(layer0_outputs(8943));
    outputs(7822) <= (layer0_outputs(2061)) and not (layer0_outputs(4413));
    outputs(7823) <= layer0_outputs(3685);
    outputs(7824) <= not(layer0_outputs(8222));
    outputs(7825) <= (layer0_outputs(5397)) and (layer0_outputs(8279));
    outputs(7826) <= not((layer0_outputs(98)) or (layer0_outputs(133)));
    outputs(7827) <= layer0_outputs(1108);
    outputs(7828) <= (layer0_outputs(6150)) or (layer0_outputs(1381));
    outputs(7829) <= (layer0_outputs(2906)) xor (layer0_outputs(8690));
    outputs(7830) <= not(layer0_outputs(6465));
    outputs(7831) <= layer0_outputs(4996);
    outputs(7832) <= not((layer0_outputs(2036)) xor (layer0_outputs(5878)));
    outputs(7833) <= layer0_outputs(829);
    outputs(7834) <= layer0_outputs(2688);
    outputs(7835) <= layer0_outputs(4736);
    outputs(7836) <= layer0_outputs(4920);
    outputs(7837) <= not((layer0_outputs(5277)) xor (layer0_outputs(1380)));
    outputs(7838) <= (layer0_outputs(2624)) and not (layer0_outputs(8171));
    outputs(7839) <= (layer0_outputs(7069)) and not (layer0_outputs(6819));
    outputs(7840) <= (layer0_outputs(6247)) and not (layer0_outputs(7921));
    outputs(7841) <= not(layer0_outputs(8244));
    outputs(7842) <= layer0_outputs(3252);
    outputs(7843) <= (layer0_outputs(1334)) and not (layer0_outputs(2499));
    outputs(7844) <= not(layer0_outputs(9014));
    outputs(7845) <= not(layer0_outputs(10072));
    outputs(7846) <= (layer0_outputs(2517)) and (layer0_outputs(4388));
    outputs(7847) <= not((layer0_outputs(6490)) and (layer0_outputs(5694)));
    outputs(7848) <= not(layer0_outputs(6312));
    outputs(7849) <= layer0_outputs(4847);
    outputs(7850) <= not(layer0_outputs(5926));
    outputs(7851) <= not((layer0_outputs(7876)) or (layer0_outputs(3585)));
    outputs(7852) <= layer0_outputs(8394);
    outputs(7853) <= (layer0_outputs(8911)) xor (layer0_outputs(193));
    outputs(7854) <= not((layer0_outputs(10118)) xor (layer0_outputs(4259)));
    outputs(7855) <= not(layer0_outputs(5184));
    outputs(7856) <= layer0_outputs(5962);
    outputs(7857) <= layer0_outputs(2344);
    outputs(7858) <= not(layer0_outputs(10095));
    outputs(7859) <= (layer0_outputs(5780)) and (layer0_outputs(8501));
    outputs(7860) <= not(layer0_outputs(7933));
    outputs(7861) <= not(layer0_outputs(7879)) or (layer0_outputs(8084));
    outputs(7862) <= not(layer0_outputs(5043));
    outputs(7863) <= not(layer0_outputs(5862)) or (layer0_outputs(9517));
    outputs(7864) <= not(layer0_outputs(5410));
    outputs(7865) <= layer0_outputs(9290);
    outputs(7866) <= (layer0_outputs(9335)) xor (layer0_outputs(3929));
    outputs(7867) <= not(layer0_outputs(6932));
    outputs(7868) <= layer0_outputs(4975);
    outputs(7869) <= (layer0_outputs(6606)) and not (layer0_outputs(186));
    outputs(7870) <= layer0_outputs(2620);
    outputs(7871) <= layer0_outputs(931);
    outputs(7872) <= layer0_outputs(5519);
    outputs(7873) <= (layer0_outputs(5374)) xor (layer0_outputs(3098));
    outputs(7874) <= (layer0_outputs(8906)) and not (layer0_outputs(9748));
    outputs(7875) <= (layer0_outputs(407)) and not (layer0_outputs(3413));
    outputs(7876) <= layer0_outputs(1784);
    outputs(7877) <= (layer0_outputs(2325)) and not (layer0_outputs(1354));
    outputs(7878) <= (layer0_outputs(4971)) xor (layer0_outputs(3852));
    outputs(7879) <= (layer0_outputs(4725)) and not (layer0_outputs(7093));
    outputs(7880) <= (layer0_outputs(4939)) and not (layer0_outputs(7720));
    outputs(7881) <= not(layer0_outputs(2352));
    outputs(7882) <= not(layer0_outputs(9371));
    outputs(7883) <= not(layer0_outputs(6170));
    outputs(7884) <= not(layer0_outputs(3683));
    outputs(7885) <= (layer0_outputs(10030)) xor (layer0_outputs(673));
    outputs(7886) <= not(layer0_outputs(924));
    outputs(7887) <= not((layer0_outputs(3354)) xor (layer0_outputs(1633)));
    outputs(7888) <= (layer0_outputs(3654)) and not (layer0_outputs(4196));
    outputs(7889) <= (layer0_outputs(10137)) and not (layer0_outputs(7973));
    outputs(7890) <= not((layer0_outputs(9607)) xor (layer0_outputs(506)));
    outputs(7891) <= not(layer0_outputs(9657));
    outputs(7892) <= layer0_outputs(560);
    outputs(7893) <= (layer0_outputs(5464)) and not (layer0_outputs(3841));
    outputs(7894) <= not((layer0_outputs(6732)) and (layer0_outputs(8796)));
    outputs(7895) <= not(layer0_outputs(916)) or (layer0_outputs(5788));
    outputs(7896) <= (layer0_outputs(9763)) and not (layer0_outputs(4171));
    outputs(7897) <= not(layer0_outputs(8331)) or (layer0_outputs(7975));
    outputs(7898) <= layer0_outputs(5963);
    outputs(7899) <= not((layer0_outputs(9117)) xor (layer0_outputs(8053)));
    outputs(7900) <= layer0_outputs(117);
    outputs(7901) <= (layer0_outputs(1206)) and (layer0_outputs(3052));
    outputs(7902) <= not(layer0_outputs(4119));
    outputs(7903) <= (layer0_outputs(5674)) and not (layer0_outputs(10145));
    outputs(7904) <= not(layer0_outputs(3073));
    outputs(7905) <= layer0_outputs(9573);
    outputs(7906) <= not(layer0_outputs(4211));
    outputs(7907) <= (layer0_outputs(9369)) and not (layer0_outputs(6164));
    outputs(7908) <= not(layer0_outputs(9326));
    outputs(7909) <= not(layer0_outputs(8365));
    outputs(7910) <= not(layer0_outputs(5853));
    outputs(7911) <= not((layer0_outputs(6981)) or (layer0_outputs(9021)));
    outputs(7912) <= not((layer0_outputs(3848)) and (layer0_outputs(2939)));
    outputs(7913) <= not((layer0_outputs(7730)) or (layer0_outputs(6969)));
    outputs(7914) <= layer0_outputs(1457);
    outputs(7915) <= not(layer0_outputs(9582));
    outputs(7916) <= layer0_outputs(7568);
    outputs(7917) <= not((layer0_outputs(5269)) or (layer0_outputs(2544)));
    outputs(7918) <= (layer0_outputs(1304)) and not (layer0_outputs(4773));
    outputs(7919) <= (layer0_outputs(991)) and not (layer0_outputs(2531));
    outputs(7920) <= layer0_outputs(8205);
    outputs(7921) <= (layer0_outputs(10148)) and (layer0_outputs(4634));
    outputs(7922) <= not((layer0_outputs(3400)) and (layer0_outputs(5795)));
    outputs(7923) <= not(layer0_outputs(9254));
    outputs(7924) <= not(layer0_outputs(3081));
    outputs(7925) <= layer0_outputs(2570);
    outputs(7926) <= not((layer0_outputs(9801)) xor (layer0_outputs(1562)));
    outputs(7927) <= not(layer0_outputs(3718));
    outputs(7928) <= not((layer0_outputs(8186)) or (layer0_outputs(9858)));
    outputs(7929) <= layer0_outputs(2709);
    outputs(7930) <= (layer0_outputs(8473)) and not (layer0_outputs(7318));
    outputs(7931) <= layer0_outputs(4153);
    outputs(7932) <= (layer0_outputs(9671)) and not (layer0_outputs(404));
    outputs(7933) <= layer0_outputs(1685);
    outputs(7934) <= (layer0_outputs(2913)) and not (layer0_outputs(659));
    outputs(7935) <= layer0_outputs(6813);
    outputs(7936) <= (layer0_outputs(5890)) xor (layer0_outputs(8659));
    outputs(7937) <= (layer0_outputs(1172)) and (layer0_outputs(5191));
    outputs(7938) <= (layer0_outputs(2992)) and not (layer0_outputs(6939));
    outputs(7939) <= layer0_outputs(10218);
    outputs(7940) <= not((layer0_outputs(5271)) and (layer0_outputs(2996)));
    outputs(7941) <= layer0_outputs(10122);
    outputs(7942) <= not(layer0_outputs(8648));
    outputs(7943) <= not(layer0_outputs(7525));
    outputs(7944) <= not(layer0_outputs(2431)) or (layer0_outputs(1182));
    outputs(7945) <= not(layer0_outputs(8305)) or (layer0_outputs(8239));
    outputs(7946) <= not((layer0_outputs(7511)) xor (layer0_outputs(6768)));
    outputs(7947) <= not((layer0_outputs(2650)) and (layer0_outputs(4300)));
    outputs(7948) <= (layer0_outputs(3021)) or (layer0_outputs(3869));
    outputs(7949) <= layer0_outputs(85);
    outputs(7950) <= not(layer0_outputs(2645));
    outputs(7951) <= layer0_outputs(898);
    outputs(7952) <= not((layer0_outputs(939)) xor (layer0_outputs(960)));
    outputs(7953) <= layer0_outputs(8779);
    outputs(7954) <= not(layer0_outputs(7375)) or (layer0_outputs(5801));
    outputs(7955) <= not((layer0_outputs(43)) and (layer0_outputs(1731)));
    outputs(7956) <= (layer0_outputs(9842)) xor (layer0_outputs(3080));
    outputs(7957) <= not(layer0_outputs(9919));
    outputs(7958) <= not((layer0_outputs(3267)) and (layer0_outputs(9219)));
    outputs(7959) <= not(layer0_outputs(7519));
    outputs(7960) <= layer0_outputs(7130);
    outputs(7961) <= not(layer0_outputs(7306));
    outputs(7962) <= not((layer0_outputs(2541)) xor (layer0_outputs(3970)));
    outputs(7963) <= not((layer0_outputs(4602)) xor (layer0_outputs(604)));
    outputs(7964) <= (layer0_outputs(2605)) xor (layer0_outputs(7294));
    outputs(7965) <= not((layer0_outputs(8215)) xor (layer0_outputs(5411)));
    outputs(7966) <= layer0_outputs(8676);
    outputs(7967) <= not(layer0_outputs(3673));
    outputs(7968) <= layer0_outputs(4730);
    outputs(7969) <= layer0_outputs(2316);
    outputs(7970) <= layer0_outputs(5503);
    outputs(7971) <= not(layer0_outputs(9487));
    outputs(7972) <= layer0_outputs(10224);
    outputs(7973) <= layer0_outputs(803);
    outputs(7974) <= not(layer0_outputs(9514));
    outputs(7975) <= not(layer0_outputs(3586));
    outputs(7976) <= not(layer0_outputs(3980));
    outputs(7977) <= (layer0_outputs(2492)) and (layer0_outputs(7490));
    outputs(7978) <= (layer0_outputs(7463)) xor (layer0_outputs(6594));
    outputs(7979) <= not(layer0_outputs(8660));
    outputs(7980) <= (layer0_outputs(3453)) and not (layer0_outputs(7148));
    outputs(7981) <= not((layer0_outputs(7201)) xor (layer0_outputs(9227)));
    outputs(7982) <= not(layer0_outputs(4253));
    outputs(7983) <= (layer0_outputs(584)) xor (layer0_outputs(3123));
    outputs(7984) <= layer0_outputs(2570);
    outputs(7985) <= (layer0_outputs(8044)) and not (layer0_outputs(7536));
    outputs(7986) <= (layer0_outputs(8426)) and not (layer0_outputs(2765));
    outputs(7987) <= not(layer0_outputs(3701));
    outputs(7988) <= (layer0_outputs(897)) xor (layer0_outputs(959));
    outputs(7989) <= (layer0_outputs(3654)) and not (layer0_outputs(4697));
    outputs(7990) <= not(layer0_outputs(4523));
    outputs(7991) <= (layer0_outputs(9977)) and (layer0_outputs(3056));
    outputs(7992) <= not(layer0_outputs(4441));
    outputs(7993) <= layer0_outputs(7345);
    outputs(7994) <= (layer0_outputs(2458)) xor (layer0_outputs(7710));
    outputs(7995) <= not(layer0_outputs(336)) or (layer0_outputs(4653));
    outputs(7996) <= (layer0_outputs(96)) xor (layer0_outputs(7982));
    outputs(7997) <= not(layer0_outputs(4836));
    outputs(7998) <= layer0_outputs(8364);
    outputs(7999) <= not((layer0_outputs(9572)) or (layer0_outputs(6973)));
    outputs(8000) <= (layer0_outputs(5493)) and (layer0_outputs(2561));
    outputs(8001) <= (layer0_outputs(4054)) and (layer0_outputs(2662));
    outputs(8002) <= layer0_outputs(5085);
    outputs(8003) <= not(layer0_outputs(6512));
    outputs(8004) <= layer0_outputs(5975);
    outputs(8005) <= layer0_outputs(3260);
    outputs(8006) <= layer0_outputs(2469);
    outputs(8007) <= (layer0_outputs(5481)) and (layer0_outputs(3254));
    outputs(8008) <= (layer0_outputs(8102)) and not (layer0_outputs(2950));
    outputs(8009) <= (layer0_outputs(5025)) xor (layer0_outputs(8571));
    outputs(8010) <= not(layer0_outputs(6279));
    outputs(8011) <= layer0_outputs(1464);
    outputs(8012) <= not(layer0_outputs(5253));
    outputs(8013) <= (layer0_outputs(3097)) and (layer0_outputs(1971));
    outputs(8014) <= (layer0_outputs(559)) and not (layer0_outputs(7757));
    outputs(8015) <= not(layer0_outputs(4046));
    outputs(8016) <= (layer0_outputs(7496)) or (layer0_outputs(4106));
    outputs(8017) <= (layer0_outputs(1570)) xor (layer0_outputs(2891));
    outputs(8018) <= not(layer0_outputs(1961));
    outputs(8019) <= (layer0_outputs(7214)) and not (layer0_outputs(8837));
    outputs(8020) <= (layer0_outputs(7505)) and not (layer0_outputs(2148));
    outputs(8021) <= not((layer0_outputs(6233)) xor (layer0_outputs(4755)));
    outputs(8022) <= layer0_outputs(8283);
    outputs(8023) <= layer0_outputs(1375);
    outputs(8024) <= layer0_outputs(5149);
    outputs(8025) <= (layer0_outputs(8054)) or (layer0_outputs(242));
    outputs(8026) <= (layer0_outputs(10010)) and not (layer0_outputs(1888));
    outputs(8027) <= not(layer0_outputs(4227));
    outputs(8028) <= not(layer0_outputs(7753)) or (layer0_outputs(831));
    outputs(8029) <= (layer0_outputs(3069)) and not (layer0_outputs(4853));
    outputs(8030) <= not((layer0_outputs(8971)) or (layer0_outputs(8425)));
    outputs(8031) <= not(layer0_outputs(2948));
    outputs(8032) <= (layer0_outputs(4361)) and not (layer0_outputs(362));
    outputs(8033) <= (layer0_outputs(2462)) and not (layer0_outputs(1078));
    outputs(8034) <= not(layer0_outputs(9460));
    outputs(8035) <= not((layer0_outputs(3469)) or (layer0_outputs(8896)));
    outputs(8036) <= not(layer0_outputs(3800)) or (layer0_outputs(6815));
    outputs(8037) <= layer0_outputs(8262);
    outputs(8038) <= (layer0_outputs(9125)) and (layer0_outputs(6084));
    outputs(8039) <= (layer0_outputs(8934)) and not (layer0_outputs(2056));
    outputs(8040) <= not(layer0_outputs(8974));
    outputs(8041) <= (layer0_outputs(1721)) xor (layer0_outputs(6304));
    outputs(8042) <= not(layer0_outputs(2751));
    outputs(8043) <= (layer0_outputs(581)) xor (layer0_outputs(8976));
    outputs(8044) <= layer0_outputs(3474);
    outputs(8045) <= layer0_outputs(8670);
    outputs(8046) <= not((layer0_outputs(5134)) xor (layer0_outputs(3175)));
    outputs(8047) <= (layer0_outputs(3839)) xor (layer0_outputs(993));
    outputs(8048) <= not(layer0_outputs(3912));
    outputs(8049) <= (layer0_outputs(9004)) and not (layer0_outputs(6543));
    outputs(8050) <= (layer0_outputs(2713)) xor (layer0_outputs(9859));
    outputs(8051) <= (layer0_outputs(4011)) and not (layer0_outputs(9028));
    outputs(8052) <= (layer0_outputs(603)) and not (layer0_outputs(166));
    outputs(8053) <= not(layer0_outputs(4029));
    outputs(8054) <= (layer0_outputs(9265)) and (layer0_outputs(9715));
    outputs(8055) <= (layer0_outputs(1128)) and not (layer0_outputs(6025));
    outputs(8056) <= not(layer0_outputs(9350));
    outputs(8057) <= (layer0_outputs(4382)) and (layer0_outputs(6019));
    outputs(8058) <= not((layer0_outputs(10208)) xor (layer0_outputs(1629)));
    outputs(8059) <= layer0_outputs(2663);
    outputs(8060) <= (layer0_outputs(3817)) xor (layer0_outputs(8628));
    outputs(8061) <= not((layer0_outputs(4237)) or (layer0_outputs(5024)));
    outputs(8062) <= not(layer0_outputs(8455)) or (layer0_outputs(5333));
    outputs(8063) <= not(layer0_outputs(9379));
    outputs(8064) <= not(layer0_outputs(5200));
    outputs(8065) <= (layer0_outputs(682)) and not (layer0_outputs(8225));
    outputs(8066) <= not((layer0_outputs(9580)) or (layer0_outputs(9499)));
    outputs(8067) <= layer0_outputs(6850);
    outputs(8068) <= (layer0_outputs(7831)) xor (layer0_outputs(8782));
    outputs(8069) <= layer0_outputs(6544);
    outputs(8070) <= (layer0_outputs(307)) xor (layer0_outputs(8949));
    outputs(8071) <= not((layer0_outputs(9472)) or (layer0_outputs(3560)));
    outputs(8072) <= layer0_outputs(4198);
    outputs(8073) <= (layer0_outputs(8806)) and (layer0_outputs(1194));
    outputs(8074) <= (layer0_outputs(3605)) and (layer0_outputs(6346));
    outputs(8075) <= (layer0_outputs(5772)) and not (layer0_outputs(8387));
    outputs(8076) <= (layer0_outputs(9814)) and not (layer0_outputs(6021));
    outputs(8077) <= (layer0_outputs(3865)) and not (layer0_outputs(8839));
    outputs(8078) <= not((layer0_outputs(3330)) or (layer0_outputs(3429)));
    outputs(8079) <= (layer0_outputs(8595)) xor (layer0_outputs(9075));
    outputs(8080) <= layer0_outputs(5076);
    outputs(8081) <= layer0_outputs(2523);
    outputs(8082) <= not((layer0_outputs(1331)) xor (layer0_outputs(8077)));
    outputs(8083) <= (layer0_outputs(4067)) xor (layer0_outputs(2613));
    outputs(8084) <= (layer0_outputs(6755)) and not (layer0_outputs(3963));
    outputs(8085) <= not((layer0_outputs(5991)) and (layer0_outputs(9109)));
    outputs(8086) <= not((layer0_outputs(6287)) or (layer0_outputs(6144)));
    outputs(8087) <= (layer0_outputs(10143)) and not (layer0_outputs(7876));
    outputs(8088) <= not(layer0_outputs(5702));
    outputs(8089) <= not(layer0_outputs(3568));
    outputs(8090) <= not(layer0_outputs(1065));
    outputs(8091) <= not(layer0_outputs(1275));
    outputs(8092) <= layer0_outputs(6740);
    outputs(8093) <= not(layer0_outputs(2769));
    outputs(8094) <= (layer0_outputs(6040)) and (layer0_outputs(4692));
    outputs(8095) <= not(layer0_outputs(6093));
    outputs(8096) <= not((layer0_outputs(7126)) xor (layer0_outputs(5907)));
    outputs(8097) <= (layer0_outputs(5267)) and (layer0_outputs(6240));
    outputs(8098) <= not(layer0_outputs(1451));
    outputs(8099) <= (layer0_outputs(7947)) and not (layer0_outputs(4068));
    outputs(8100) <= (layer0_outputs(7995)) and not (layer0_outputs(4614));
    outputs(8101) <= not(layer0_outputs(8800));
    outputs(8102) <= not(layer0_outputs(280)) or (layer0_outputs(7644));
    outputs(8103) <= not((layer0_outputs(1199)) or (layer0_outputs(3265)));
    outputs(8104) <= not(layer0_outputs(9719));
    outputs(8105) <= layer0_outputs(4613);
    outputs(8106) <= not(layer0_outputs(6266));
    outputs(8107) <= not(layer0_outputs(7396)) or (layer0_outputs(6967));
    outputs(8108) <= layer0_outputs(1938);
    outputs(8109) <= not(layer0_outputs(6509));
    outputs(8110) <= not((layer0_outputs(8684)) or (layer0_outputs(6859)));
    outputs(8111) <= (layer0_outputs(5072)) xor (layer0_outputs(6981));
    outputs(8112) <= not((layer0_outputs(8486)) xor (layer0_outputs(5145)));
    outputs(8113) <= (layer0_outputs(4040)) and not (layer0_outputs(7777));
    outputs(8114) <= layer0_outputs(8415);
    outputs(8115) <= not(layer0_outputs(4817));
    outputs(8116) <= (layer0_outputs(9596)) xor (layer0_outputs(6499));
    outputs(8117) <= not((layer0_outputs(10225)) xor (layer0_outputs(10144)));
    outputs(8118) <= not((layer0_outputs(9116)) and (layer0_outputs(2973)));
    outputs(8119) <= (layer0_outputs(9523)) and not (layer0_outputs(708));
    outputs(8120) <= not((layer0_outputs(8274)) xor (layer0_outputs(2769)));
    outputs(8121) <= (layer0_outputs(547)) and (layer0_outputs(5382));
    outputs(8122) <= layer0_outputs(3058);
    outputs(8123) <= layer0_outputs(1666);
    outputs(8124) <= layer0_outputs(2339);
    outputs(8125) <= (layer0_outputs(3211)) and not (layer0_outputs(3689));
    outputs(8126) <= (layer0_outputs(9079)) and (layer0_outputs(4563));
    outputs(8127) <= (layer0_outputs(5489)) and (layer0_outputs(4488));
    outputs(8128) <= layer0_outputs(9550);
    outputs(8129) <= not(layer0_outputs(9310));
    outputs(8130) <= layer0_outputs(7997);
    outputs(8131) <= layer0_outputs(1397);
    outputs(8132) <= (layer0_outputs(6334)) xor (layer0_outputs(1948));
    outputs(8133) <= not((layer0_outputs(856)) xor (layer0_outputs(8052)));
    outputs(8134) <= not(layer0_outputs(7304));
    outputs(8135) <= (layer0_outputs(8333)) xor (layer0_outputs(5212));
    outputs(8136) <= layer0_outputs(2893);
    outputs(8137) <= (layer0_outputs(4841)) and (layer0_outputs(6433));
    outputs(8138) <= not(layer0_outputs(6809));
    outputs(8139) <= layer0_outputs(8360);
    outputs(8140) <= not((layer0_outputs(4194)) or (layer0_outputs(5775)));
    outputs(8141) <= not(layer0_outputs(1972)) or (layer0_outputs(5143));
    outputs(8142) <= not(layer0_outputs(5118));
    outputs(8143) <= not((layer0_outputs(9010)) xor (layer0_outputs(2011)));
    outputs(8144) <= not(layer0_outputs(8743));
    outputs(8145) <= (layer0_outputs(5990)) and not (layer0_outputs(2735));
    outputs(8146) <= not(layer0_outputs(2304));
    outputs(8147) <= (layer0_outputs(10135)) and not (layer0_outputs(9537));
    outputs(8148) <= layer0_outputs(5545);
    outputs(8149) <= not(layer0_outputs(9962)) or (layer0_outputs(8312));
    outputs(8150) <= not(layer0_outputs(6105)) or (layer0_outputs(8258));
    outputs(8151) <= not(layer0_outputs(9560));
    outputs(8152) <= not((layer0_outputs(7892)) and (layer0_outputs(3493)));
    outputs(8153) <= layer0_outputs(9621);
    outputs(8154) <= not((layer0_outputs(9198)) or (layer0_outputs(8899)));
    outputs(8155) <= (layer0_outputs(2173)) and not (layer0_outputs(3669));
    outputs(8156) <= (layer0_outputs(9738)) xor (layer0_outputs(3220));
    outputs(8157) <= (layer0_outputs(127)) xor (layer0_outputs(7513));
    outputs(8158) <= not(layer0_outputs(1707));
    outputs(8159) <= layer0_outputs(4692);
    outputs(8160) <= (layer0_outputs(1681)) and not (layer0_outputs(2007));
    outputs(8161) <= not((layer0_outputs(7183)) xor (layer0_outputs(9731)));
    outputs(8162) <= not(layer0_outputs(1868));
    outputs(8163) <= layer0_outputs(10210);
    outputs(8164) <= (layer0_outputs(3489)) and not (layer0_outputs(3923));
    outputs(8165) <= (layer0_outputs(1270)) xor (layer0_outputs(1594));
    outputs(8166) <= not(layer0_outputs(5968));
    outputs(8167) <= not((layer0_outputs(2752)) or (layer0_outputs(9237)));
    outputs(8168) <= layer0_outputs(8710);
    outputs(8169) <= (layer0_outputs(7087)) and not (layer0_outputs(752));
    outputs(8170) <= not(layer0_outputs(8833)) or (layer0_outputs(9183));
    outputs(8171) <= not((layer0_outputs(4487)) or (layer0_outputs(801)));
    outputs(8172) <= (layer0_outputs(5618)) xor (layer0_outputs(7813));
    outputs(8173) <= not(layer0_outputs(3574));
    outputs(8174) <= not((layer0_outputs(7346)) or (layer0_outputs(1447)));
    outputs(8175) <= (layer0_outputs(1408)) and (layer0_outputs(163));
    outputs(8176) <= (layer0_outputs(6523)) xor (layer0_outputs(1485));
    outputs(8177) <= layer0_outputs(7799);
    outputs(8178) <= layer0_outputs(3524);
    outputs(8179) <= layer0_outputs(4904);
    outputs(8180) <= (layer0_outputs(5404)) and not (layer0_outputs(8152));
    outputs(8181) <= layer0_outputs(2533);
    outputs(8182) <= not((layer0_outputs(8977)) or (layer0_outputs(8119)));
    outputs(8183) <= not(layer0_outputs(2361));
    outputs(8184) <= not((layer0_outputs(3949)) xor (layer0_outputs(6249)));
    outputs(8185) <= (layer0_outputs(1007)) and (layer0_outputs(4597));
    outputs(8186) <= (layer0_outputs(148)) and not (layer0_outputs(1508));
    outputs(8187) <= (layer0_outputs(249)) and (layer0_outputs(2792));
    outputs(8188) <= not(layer0_outputs(6933));
    outputs(8189) <= not((layer0_outputs(9876)) or (layer0_outputs(2019)));
    outputs(8190) <= layer0_outputs(9041);
    outputs(8191) <= layer0_outputs(7604);
    outputs(8192) <= (layer0_outputs(3022)) or (layer0_outputs(6829));
    outputs(8193) <= not(layer0_outputs(344)) or (layer0_outputs(2622));
    outputs(8194) <= (layer0_outputs(9439)) and not (layer0_outputs(8944));
    outputs(8195) <= (layer0_outputs(3449)) xor (layer0_outputs(4850));
    outputs(8196) <= not(layer0_outputs(4039));
    outputs(8197) <= layer0_outputs(6790);
    outputs(8198) <= not(layer0_outputs(900));
    outputs(8199) <= not((layer0_outputs(4802)) xor (layer0_outputs(10172)));
    outputs(8200) <= not(layer0_outputs(7433));
    outputs(8201) <= (layer0_outputs(6111)) or (layer0_outputs(7062));
    outputs(8202) <= layer0_outputs(9839);
    outputs(8203) <= not(layer0_outputs(7569)) or (layer0_outputs(6140));
    outputs(8204) <= not((layer0_outputs(5127)) and (layer0_outputs(9755)));
    outputs(8205) <= not(layer0_outputs(9887));
    outputs(8206) <= (layer0_outputs(4831)) and (layer0_outputs(5446));
    outputs(8207) <= (layer0_outputs(4498)) xor (layer0_outputs(10087));
    outputs(8208) <= not((layer0_outputs(1144)) xor (layer0_outputs(1658)));
    outputs(8209) <= not(layer0_outputs(7128)) or (layer0_outputs(4956));
    outputs(8210) <= not(layer0_outputs(3957)) or (layer0_outputs(3777));
    outputs(8211) <= not((layer0_outputs(7531)) xor (layer0_outputs(6574)));
    outputs(8212) <= not((layer0_outputs(1710)) xor (layer0_outputs(438)));
    outputs(8213) <= (layer0_outputs(3077)) xor (layer0_outputs(2911));
    outputs(8214) <= (layer0_outputs(4441)) or (layer0_outputs(7256));
    outputs(8215) <= (layer0_outputs(1076)) xor (layer0_outputs(4892));
    outputs(8216) <= not(layer0_outputs(4458));
    outputs(8217) <= (layer0_outputs(7497)) xor (layer0_outputs(875));
    outputs(8218) <= (layer0_outputs(9186)) and not (layer0_outputs(7883));
    outputs(8219) <= not((layer0_outputs(7020)) xor (layer0_outputs(626)));
    outputs(8220) <= not(layer0_outputs(7358));
    outputs(8221) <= layer0_outputs(7857);
    outputs(8222) <= not(layer0_outputs(2892)) or (layer0_outputs(7059));
    outputs(8223) <= not(layer0_outputs(9871)) or (layer0_outputs(946));
    outputs(8224) <= (layer0_outputs(7167)) or (layer0_outputs(714));
    outputs(8225) <= not(layer0_outputs(8675));
    outputs(8226) <= '1';
    outputs(8227) <= (layer0_outputs(8060)) xor (layer0_outputs(4707));
    outputs(8228) <= not(layer0_outputs(7289));
    outputs(8229) <= not(layer0_outputs(4329)) or (layer0_outputs(602));
    outputs(8230) <= layer0_outputs(2590);
    outputs(8231) <= (layer0_outputs(9246)) or (layer0_outputs(2079));
    outputs(8232) <= not((layer0_outputs(2054)) xor (layer0_outputs(365)));
    outputs(8233) <= not((layer0_outputs(3712)) xor (layer0_outputs(5214)));
    outputs(8234) <= not(layer0_outputs(7874)) or (layer0_outputs(2382));
    outputs(8235) <= (layer0_outputs(8227)) xor (layer0_outputs(174));
    outputs(8236) <= not((layer0_outputs(2852)) xor (layer0_outputs(7418)));
    outputs(8237) <= layer0_outputs(1527);
    outputs(8238) <= layer0_outputs(9383);
    outputs(8239) <= not(layer0_outputs(2773));
    outputs(8240) <= not(layer0_outputs(5463));
    outputs(8241) <= (layer0_outputs(6216)) xor (layer0_outputs(8469));
    outputs(8242) <= (layer0_outputs(3648)) xor (layer0_outputs(7363));
    outputs(8243) <= not(layer0_outputs(7161)) or (layer0_outputs(8287));
    outputs(8244) <= layer0_outputs(9511);
    outputs(8245) <= layer0_outputs(1760);
    outputs(8246) <= not((layer0_outputs(9903)) xor (layer0_outputs(5470)));
    outputs(8247) <= (layer0_outputs(5131)) xor (layer0_outputs(907));
    outputs(8248) <= not(layer0_outputs(8102)) or (layer0_outputs(4229));
    outputs(8249) <= (layer0_outputs(9144)) xor (layer0_outputs(5536));
    outputs(8250) <= (layer0_outputs(9576)) xor (layer0_outputs(20));
    outputs(8251) <= not((layer0_outputs(1302)) and (layer0_outputs(432)));
    outputs(8252) <= (layer0_outputs(3025)) or (layer0_outputs(7403));
    outputs(8253) <= layer0_outputs(9639);
    outputs(8254) <= (layer0_outputs(770)) xor (layer0_outputs(1219));
    outputs(8255) <= layer0_outputs(7120);
    outputs(8256) <= not(layer0_outputs(2882));
    outputs(8257) <= not((layer0_outputs(3575)) xor (layer0_outputs(8952)));
    outputs(8258) <= not((layer0_outputs(8252)) xor (layer0_outputs(6113)));
    outputs(8259) <= not((layer0_outputs(999)) xor (layer0_outputs(9192)));
    outputs(8260) <= layer0_outputs(5554);
    outputs(8261) <= not((layer0_outputs(8689)) xor (layer0_outputs(4320)));
    outputs(8262) <= (layer0_outputs(10053)) xor (layer0_outputs(5594));
    outputs(8263) <= not(layer0_outputs(8761)) or (layer0_outputs(5221));
    outputs(8264) <= layer0_outputs(1003);
    outputs(8265) <= not(layer0_outputs(3938));
    outputs(8266) <= (layer0_outputs(8177)) or (layer0_outputs(3112));
    outputs(8267) <= layer0_outputs(8773);
    outputs(8268) <= not((layer0_outputs(2733)) xor (layer0_outputs(1460)));
    outputs(8269) <= (layer0_outputs(4049)) xor (layer0_outputs(530));
    outputs(8270) <= not(layer0_outputs(1616)) or (layer0_outputs(1352));
    outputs(8271) <= not(layer0_outputs(4772));
    outputs(8272) <= (layer0_outputs(12)) and not (layer0_outputs(6582));
    outputs(8273) <= (layer0_outputs(1523)) and (layer0_outputs(7215));
    outputs(8274) <= layer0_outputs(4491);
    outputs(8275) <= (layer0_outputs(7095)) or (layer0_outputs(10027));
    outputs(8276) <= not((layer0_outputs(5218)) and (layer0_outputs(6260)));
    outputs(8277) <= layer0_outputs(1831);
    outputs(8278) <= (layer0_outputs(441)) xor (layer0_outputs(8936));
    outputs(8279) <= layer0_outputs(9696);
    outputs(8280) <= (layer0_outputs(870)) xor (layer0_outputs(4665));
    outputs(8281) <= layer0_outputs(121);
    outputs(8282) <= (layer0_outputs(408)) xor (layer0_outputs(6925));
    outputs(8283) <= not(layer0_outputs(5999));
    outputs(8284) <= (layer0_outputs(10164)) and (layer0_outputs(2754));
    outputs(8285) <= not(layer0_outputs(9848));
    outputs(8286) <= layer0_outputs(1627);
    outputs(8287) <= (layer0_outputs(10074)) xor (layer0_outputs(3542));
    outputs(8288) <= not((layer0_outputs(9044)) xor (layer0_outputs(4611)));
    outputs(8289) <= (layer0_outputs(6517)) xor (layer0_outputs(6845));
    outputs(8290) <= not(layer0_outputs(7734)) or (layer0_outputs(435));
    outputs(8291) <= (layer0_outputs(3911)) and not (layer0_outputs(4652));
    outputs(8292) <= (layer0_outputs(1442)) xor (layer0_outputs(3409));
    outputs(8293) <= (layer0_outputs(5332)) xor (layer0_outputs(5750));
    outputs(8294) <= (layer0_outputs(6607)) xor (layer0_outputs(6107));
    outputs(8295) <= not((layer0_outputs(10231)) xor (layer0_outputs(264)));
    outputs(8296) <= layer0_outputs(9082);
    outputs(8297) <= not((layer0_outputs(6603)) xor (layer0_outputs(1895)));
    outputs(8298) <= not(layer0_outputs(5346));
    outputs(8299) <= not(layer0_outputs(4303)) or (layer0_outputs(3441));
    outputs(8300) <= not(layer0_outputs(1203));
    outputs(8301) <= layer0_outputs(67);
    outputs(8302) <= not(layer0_outputs(3675)) or (layer0_outputs(7696));
    outputs(8303) <= layer0_outputs(4382);
    outputs(8304) <= not((layer0_outputs(3649)) xor (layer0_outputs(9764)));
    outputs(8305) <= (layer0_outputs(10007)) and (layer0_outputs(4236));
    outputs(8306) <= not(layer0_outputs(1075)) or (layer0_outputs(8531));
    outputs(8307) <= not(layer0_outputs(1660)) or (layer0_outputs(8322));
    outputs(8308) <= (layer0_outputs(7709)) xor (layer0_outputs(3284));
    outputs(8309) <= not(layer0_outputs(3189));
    outputs(8310) <= layer0_outputs(2945);
    outputs(8311) <= (layer0_outputs(7313)) xor (layer0_outputs(6704));
    outputs(8312) <= not((layer0_outputs(5561)) and (layer0_outputs(9888)));
    outputs(8313) <= not((layer0_outputs(7760)) xor (layer0_outputs(4243)));
    outputs(8314) <= not(layer0_outputs(1125));
    outputs(8315) <= layer0_outputs(6620);
    outputs(8316) <= not(layer0_outputs(1243));
    outputs(8317) <= not(layer0_outputs(2579));
    outputs(8318) <= not(layer0_outputs(412));
    outputs(8319) <= not(layer0_outputs(4185));
    outputs(8320) <= (layer0_outputs(7255)) and not (layer0_outputs(5266));
    outputs(8321) <= not((layer0_outputs(1575)) xor (layer0_outputs(2030)));
    outputs(8322) <= not(layer0_outputs(4540));
    outputs(8323) <= not(layer0_outputs(8536));
    outputs(8324) <= not(layer0_outputs(4185));
    outputs(8325) <= (layer0_outputs(96)) xor (layer0_outputs(2498));
    outputs(8326) <= layer0_outputs(1505);
    outputs(8327) <= not((layer0_outputs(826)) and (layer0_outputs(9836)));
    outputs(8328) <= (layer0_outputs(7874)) xor (layer0_outputs(648));
    outputs(8329) <= not((layer0_outputs(973)) xor (layer0_outputs(4279)));
    outputs(8330) <= '1';
    outputs(8331) <= not(layer0_outputs(9316));
    outputs(8332) <= not((layer0_outputs(8593)) xor (layer0_outputs(9903)));
    outputs(8333) <= layer0_outputs(714);
    outputs(8334) <= (layer0_outputs(9045)) xor (layer0_outputs(1434));
    outputs(8335) <= not(layer0_outputs(1749));
    outputs(8336) <= (layer0_outputs(9725)) xor (layer0_outputs(4086));
    outputs(8337) <= (layer0_outputs(3656)) xor (layer0_outputs(7857));
    outputs(8338) <= not(layer0_outputs(7271));
    outputs(8339) <= not(layer0_outputs(5402));
    outputs(8340) <= not((layer0_outputs(5621)) and (layer0_outputs(2582)));
    outputs(8341) <= (layer0_outputs(3717)) xor (layer0_outputs(689));
    outputs(8342) <= not((layer0_outputs(7588)) xor (layer0_outputs(3450)));
    outputs(8343) <= not(layer0_outputs(7952));
    outputs(8344) <= (layer0_outputs(420)) xor (layer0_outputs(7957));
    outputs(8345) <= not(layer0_outputs(7017)) or (layer0_outputs(1149));
    outputs(8346) <= not(layer0_outputs(9405)) or (layer0_outputs(9138));
    outputs(8347) <= layer0_outputs(7643);
    outputs(8348) <= not((layer0_outputs(5220)) xor (layer0_outputs(2427)));
    outputs(8349) <= not(layer0_outputs(5609)) or (layer0_outputs(7275));
    outputs(8350) <= not(layer0_outputs(5770));
    outputs(8351) <= (layer0_outputs(466)) xor (layer0_outputs(3589));
    outputs(8352) <= layer0_outputs(9257);
    outputs(8353) <= layer0_outputs(4849);
    outputs(8354) <= layer0_outputs(3233);
    outputs(8355) <= not(layer0_outputs(7946)) or (layer0_outputs(3762));
    outputs(8356) <= layer0_outputs(8199);
    outputs(8357) <= not((layer0_outputs(5745)) xor (layer0_outputs(3787)));
    outputs(8358) <= not((layer0_outputs(7728)) xor (layer0_outputs(2299)));
    outputs(8359) <= layer0_outputs(3111);
    outputs(8360) <= not(layer0_outputs(1892));
    outputs(8361) <= not((layer0_outputs(138)) xor (layer0_outputs(9055)));
    outputs(8362) <= layer0_outputs(6861);
    outputs(8363) <= layer0_outputs(4347);
    outputs(8364) <= not((layer0_outputs(333)) xor (layer0_outputs(9059)));
    outputs(8365) <= not((layer0_outputs(9424)) xor (layer0_outputs(1927)));
    outputs(8366) <= not((layer0_outputs(7261)) and (layer0_outputs(4099)));
    outputs(8367) <= not(layer0_outputs(6406)) or (layer0_outputs(3685));
    outputs(8368) <= not(layer0_outputs(5742));
    outputs(8369) <= not(layer0_outputs(2538));
    outputs(8370) <= not(layer0_outputs(7309)) or (layer0_outputs(1385));
    outputs(8371) <= (layer0_outputs(9690)) and not (layer0_outputs(7837));
    outputs(8372) <= (layer0_outputs(588)) or (layer0_outputs(6246));
    outputs(8373) <= not((layer0_outputs(1897)) xor (layer0_outputs(3768)));
    outputs(8374) <= layer0_outputs(175);
    outputs(8375) <= (layer0_outputs(5)) and not (layer0_outputs(8529));
    outputs(8376) <= not((layer0_outputs(4448)) xor (layer0_outputs(2169)));
    outputs(8377) <= (layer0_outputs(1727)) and not (layer0_outputs(1251));
    outputs(8378) <= not(layer0_outputs(2076));
    outputs(8379) <= layer0_outputs(7913);
    outputs(8380) <= not(layer0_outputs(5594)) or (layer0_outputs(1001));
    outputs(8381) <= (layer0_outputs(3297)) or (layer0_outputs(1653));
    outputs(8382) <= layer0_outputs(3962);
    outputs(8383) <= layer0_outputs(1229);
    outputs(8384) <= not(layer0_outputs(4343));
    outputs(8385) <= (layer0_outputs(1039)) xor (layer0_outputs(1257));
    outputs(8386) <= not(layer0_outputs(1833)) or (layer0_outputs(6904));
    outputs(8387) <= not((layer0_outputs(5174)) and (layer0_outputs(4232)));
    outputs(8388) <= (layer0_outputs(6868)) or (layer0_outputs(1812));
    outputs(8389) <= layer0_outputs(7123);
    outputs(8390) <= (layer0_outputs(6212)) or (layer0_outputs(8722));
    outputs(8391) <= not(layer0_outputs(3260)) or (layer0_outputs(3025));
    outputs(8392) <= (layer0_outputs(1161)) xor (layer0_outputs(33));
    outputs(8393) <= not(layer0_outputs(4867));
    outputs(8394) <= not(layer0_outputs(4721)) or (layer0_outputs(5270));
    outputs(8395) <= layer0_outputs(7755);
    outputs(8396) <= (layer0_outputs(2644)) xor (layer0_outputs(4104));
    outputs(8397) <= not((layer0_outputs(4648)) xor (layer0_outputs(6845)));
    outputs(8398) <= (layer0_outputs(1071)) and not (layer0_outputs(9545));
    outputs(8399) <= (layer0_outputs(668)) and not (layer0_outputs(9427));
    outputs(8400) <= (layer0_outputs(4708)) xor (layer0_outputs(372));
    outputs(8401) <= layer0_outputs(8015);
    outputs(8402) <= not(layer0_outputs(4509)) or (layer0_outputs(912));
    outputs(8403) <= layer0_outputs(3650);
    outputs(8404) <= (layer0_outputs(4379)) and not (layer0_outputs(3361));
    outputs(8405) <= (layer0_outputs(3291)) and not (layer0_outputs(6190));
    outputs(8406) <= not(layer0_outputs(5345));
    outputs(8407) <= not((layer0_outputs(1328)) xor (layer0_outputs(1910)));
    outputs(8408) <= (layer0_outputs(5619)) xor (layer0_outputs(282));
    outputs(8409) <= not((layer0_outputs(4898)) and (layer0_outputs(1226)));
    outputs(8410) <= (layer0_outputs(2264)) or (layer0_outputs(5213));
    outputs(8411) <= not(layer0_outputs(2668));
    outputs(8412) <= (layer0_outputs(5929)) xor (layer0_outputs(2855));
    outputs(8413) <= not((layer0_outputs(9549)) and (layer0_outputs(5612)));
    outputs(8414) <= not((layer0_outputs(7242)) xor (layer0_outputs(6516)));
    outputs(8415) <= not(layer0_outputs(7553));
    outputs(8416) <= (layer0_outputs(5988)) and not (layer0_outputs(948));
    outputs(8417) <= not((layer0_outputs(7087)) xor (layer0_outputs(9538)));
    outputs(8418) <= layer0_outputs(6305);
    outputs(8419) <= (layer0_outputs(2288)) or (layer0_outputs(9646));
    outputs(8420) <= (layer0_outputs(6483)) xor (layer0_outputs(4107));
    outputs(8421) <= not(layer0_outputs(6630));
    outputs(8422) <= (layer0_outputs(9651)) xor (layer0_outputs(9532));
    outputs(8423) <= not(layer0_outputs(10221));
    outputs(8424) <= not(layer0_outputs(9966));
    outputs(8425) <= not((layer0_outputs(8051)) xor (layer0_outputs(1291)));
    outputs(8426) <= (layer0_outputs(2783)) or (layer0_outputs(1733));
    outputs(8427) <= layer0_outputs(7013);
    outputs(8428) <= not(layer0_outputs(826)) or (layer0_outputs(5541));
    outputs(8429) <= (layer0_outputs(7402)) or (layer0_outputs(1506));
    outputs(8430) <= not(layer0_outputs(9933));
    outputs(8431) <= not((layer0_outputs(2881)) xor (layer0_outputs(2460)));
    outputs(8432) <= not(layer0_outputs(10204)) or (layer0_outputs(564));
    outputs(8433) <= not(layer0_outputs(9897)) or (layer0_outputs(1783));
    outputs(8434) <= not((layer0_outputs(3587)) and (layer0_outputs(3036)));
    outputs(8435) <= not((layer0_outputs(5403)) xor (layer0_outputs(6690)));
    outputs(8436) <= (layer0_outputs(9365)) xor (layer0_outputs(4074));
    outputs(8437) <= (layer0_outputs(1568)) and not (layer0_outputs(5782));
    outputs(8438) <= not((layer0_outputs(9064)) and (layer0_outputs(3525)));
    outputs(8439) <= (layer0_outputs(5925)) xor (layer0_outputs(4260));
    outputs(8440) <= not((layer0_outputs(10139)) or (layer0_outputs(944)));
    outputs(8441) <= not(layer0_outputs(406));
    outputs(8442) <= not((layer0_outputs(3395)) xor (layer0_outputs(8058)));
    outputs(8443) <= not(layer0_outputs(1132));
    outputs(8444) <= not(layer0_outputs(2721)) or (layer0_outputs(7726));
    outputs(8445) <= not((layer0_outputs(4786)) xor (layer0_outputs(5585)));
    outputs(8446) <= not(layer0_outputs(2133));
    outputs(8447) <= (layer0_outputs(6140)) xor (layer0_outputs(8685));
    outputs(8448) <= not(layer0_outputs(2202));
    outputs(8449) <= not(layer0_outputs(3624));
    outputs(8450) <= not(layer0_outputs(7417));
    outputs(8451) <= (layer0_outputs(3042)) xor (layer0_outputs(8921));
    outputs(8452) <= layer0_outputs(7852);
    outputs(8453) <= layer0_outputs(3143);
    outputs(8454) <= not(layer0_outputs(7422)) or (layer0_outputs(1464));
    outputs(8455) <= not(layer0_outputs(9768));
    outputs(8456) <= not((layer0_outputs(7844)) xor (layer0_outputs(3871)));
    outputs(8457) <= (layer0_outputs(972)) and (layer0_outputs(5807));
    outputs(8458) <= (layer0_outputs(3156)) or (layer0_outputs(4789));
    outputs(8459) <= layer0_outputs(3379);
    outputs(8460) <= not(layer0_outputs(1048));
    outputs(8461) <= not((layer0_outputs(10166)) xor (layer0_outputs(1817)));
    outputs(8462) <= (layer0_outputs(4162)) xor (layer0_outputs(9119));
    outputs(8463) <= not(layer0_outputs(4214));
    outputs(8464) <= (layer0_outputs(4769)) xor (layer0_outputs(1487));
    outputs(8465) <= not(layer0_outputs(8980));
    outputs(8466) <= not((layer0_outputs(2415)) xor (layer0_outputs(5288)));
    outputs(8467) <= (layer0_outputs(7605)) xor (layer0_outputs(6664));
    outputs(8468) <= (layer0_outputs(6177)) xor (layer0_outputs(9615));
    outputs(8469) <= not(layer0_outputs(2141));
    outputs(8470) <= not((layer0_outputs(8615)) xor (layer0_outputs(5634)));
    outputs(8471) <= (layer0_outputs(8070)) and not (layer0_outputs(7473));
    outputs(8472) <= (layer0_outputs(7297)) and (layer0_outputs(7707));
    outputs(8473) <= not(layer0_outputs(9597));
    outputs(8474) <= layer0_outputs(3926);
    outputs(8475) <= not(layer0_outputs(2597)) or (layer0_outputs(3738));
    outputs(8476) <= not(layer0_outputs(3380));
    outputs(8477) <= layer0_outputs(7138);
    outputs(8478) <= not(layer0_outputs(7252)) or (layer0_outputs(6079));
    outputs(8479) <= not(layer0_outputs(4345));
    outputs(8480) <= not((layer0_outputs(6133)) and (layer0_outputs(9022)));
    outputs(8481) <= not((layer0_outputs(1636)) xor (layer0_outputs(6045)));
    outputs(8482) <= not(layer0_outputs(9601));
    outputs(8483) <= not(layer0_outputs(9663));
    outputs(8484) <= not(layer0_outputs(2667));
    outputs(8485) <= not((layer0_outputs(2624)) xor (layer0_outputs(9253)));
    outputs(8486) <= (layer0_outputs(7149)) or (layer0_outputs(1918));
    outputs(8487) <= not(layer0_outputs(3668));
    outputs(8488) <= not((layer0_outputs(9710)) or (layer0_outputs(6862)));
    outputs(8489) <= layer0_outputs(1437);
    outputs(8490) <= not(layer0_outputs(8712));
    outputs(8491) <= layer0_outputs(5910);
    outputs(8492) <= layer0_outputs(943);
    outputs(8493) <= (layer0_outputs(5283)) xor (layer0_outputs(4233));
    outputs(8494) <= not((layer0_outputs(1079)) and (layer0_outputs(6049)));
    outputs(8495) <= (layer0_outputs(9609)) xor (layer0_outputs(5086));
    outputs(8496) <= (layer0_outputs(7603)) or (layer0_outputs(1153));
    outputs(8497) <= layer0_outputs(4402);
    outputs(8498) <= (layer0_outputs(1732)) and not (layer0_outputs(7899));
    outputs(8499) <= not((layer0_outputs(9941)) xor (layer0_outputs(9476)));
    outputs(8500) <= not((layer0_outputs(6820)) xor (layer0_outputs(2789)));
    outputs(8501) <= not((layer0_outputs(7914)) xor (layer0_outputs(4592)));
    outputs(8502) <= (layer0_outputs(4826)) or (layer0_outputs(5873));
    outputs(8503) <= not(layer0_outputs(6740));
    outputs(8504) <= layer0_outputs(6696);
    outputs(8505) <= (layer0_outputs(6364)) xor (layer0_outputs(1127));
    outputs(8506) <= '1';
    outputs(8507) <= (layer0_outputs(9712)) or (layer0_outputs(3652));
    outputs(8508) <= not(layer0_outputs(4696));
    outputs(8509) <= (layer0_outputs(6220)) xor (layer0_outputs(5150));
    outputs(8510) <= layer0_outputs(5462);
    outputs(8511) <= layer0_outputs(330);
    outputs(8512) <= not((layer0_outputs(4508)) xor (layer0_outputs(4655)));
    outputs(8513) <= not(layer0_outputs(9108));
    outputs(8514) <= layer0_outputs(9435);
    outputs(8515) <= not((layer0_outputs(8758)) xor (layer0_outputs(3051)));
    outputs(8516) <= not(layer0_outputs(1313));
    outputs(8517) <= not(layer0_outputs(9181)) or (layer0_outputs(5133));
    outputs(8518) <= (layer0_outputs(3543)) and (layer0_outputs(9598));
    outputs(8519) <= (layer0_outputs(6303)) and not (layer0_outputs(2306));
    outputs(8520) <= (layer0_outputs(7419)) or (layer0_outputs(140));
    outputs(8521) <= not(layer0_outputs(6784));
    outputs(8522) <= (layer0_outputs(7328)) xor (layer0_outputs(4588));
    outputs(8523) <= (layer0_outputs(9034)) xor (layer0_outputs(4323));
    outputs(8524) <= not((layer0_outputs(1902)) or (layer0_outputs(1286)));
    outputs(8525) <= not(layer0_outputs(6562)) or (layer0_outputs(1804));
    outputs(8526) <= layer0_outputs(4088);
    outputs(8527) <= layer0_outputs(2147);
    outputs(8528) <= (layer0_outputs(4349)) xor (layer0_outputs(8546));
    outputs(8529) <= not(layer0_outputs(6168));
    outputs(8530) <= not(layer0_outputs(6738)) or (layer0_outputs(9989));
    outputs(8531) <= not((layer0_outputs(555)) xor (layer0_outputs(1654)));
    outputs(8532) <= (layer0_outputs(4599)) and not (layer0_outputs(10169));
    outputs(8533) <= not((layer0_outputs(6694)) xor (layer0_outputs(315)));
    outputs(8534) <= not(layer0_outputs(105));
    outputs(8535) <= layer0_outputs(6469);
    outputs(8536) <= not(layer0_outputs(6665));
    outputs(8537) <= not((layer0_outputs(7604)) xor (layer0_outputs(1737)));
    outputs(8538) <= not(layer0_outputs(6057)) or (layer0_outputs(9355));
    outputs(8539) <= layer0_outputs(576);
    outputs(8540) <= layer0_outputs(8604);
    outputs(8541) <= (layer0_outputs(1472)) xor (layer0_outputs(1879));
    outputs(8542) <= not((layer0_outputs(590)) xor (layer0_outputs(6459)));
    outputs(8543) <= (layer0_outputs(2505)) xor (layer0_outputs(3791));
    outputs(8544) <= not(layer0_outputs(4051));
    outputs(8545) <= (layer0_outputs(5779)) xor (layer0_outputs(1888));
    outputs(8546) <= not((layer0_outputs(9239)) and (layer0_outputs(6299)));
    outputs(8547) <= not((layer0_outputs(3466)) xor (layer0_outputs(6511)));
    outputs(8548) <= not(layer0_outputs(5985)) or (layer0_outputs(8789));
    outputs(8549) <= not((layer0_outputs(8835)) and (layer0_outputs(4595)));
    outputs(8550) <= not(layer0_outputs(2441));
    outputs(8551) <= (layer0_outputs(4155)) xor (layer0_outputs(3135));
    outputs(8552) <= not((layer0_outputs(1124)) xor (layer0_outputs(7972)));
    outputs(8553) <= layer0_outputs(4660);
    outputs(8554) <= (layer0_outputs(443)) xor (layer0_outputs(3024));
    outputs(8555) <= not((layer0_outputs(1961)) xor (layer0_outputs(2486)));
    outputs(8556) <= not((layer0_outputs(783)) xor (layer0_outputs(8630)));
    outputs(8557) <= not(layer0_outputs(559));
    outputs(8558) <= not(layer0_outputs(2658));
    outputs(8559) <= not((layer0_outputs(7497)) and (layer0_outputs(2459)));
    outputs(8560) <= (layer0_outputs(202)) xor (layer0_outputs(1018));
    outputs(8561) <= layer0_outputs(5291);
    outputs(8562) <= layer0_outputs(1678);
    outputs(8563) <= (layer0_outputs(10019)) xor (layer0_outputs(4570));
    outputs(8564) <= not((layer0_outputs(3514)) or (layer0_outputs(2165)));
    outputs(8565) <= layer0_outputs(5037);
    outputs(8566) <= not((layer0_outputs(5637)) and (layer0_outputs(10076)));
    outputs(8567) <= (layer0_outputs(35)) or (layer0_outputs(1437));
    outputs(8568) <= not((layer0_outputs(1775)) xor (layer0_outputs(9588)));
    outputs(8569) <= (layer0_outputs(9384)) or (layer0_outputs(6338));
    outputs(8570) <= not(layer0_outputs(9397)) or (layer0_outputs(5507));
    outputs(8571) <= not((layer0_outputs(2946)) xor (layer0_outputs(2858)));
    outputs(8572) <= (layer0_outputs(3778)) xor (layer0_outputs(2581));
    outputs(8573) <= not((layer0_outputs(451)) or (layer0_outputs(9725)));
    outputs(8574) <= not((layer0_outputs(4094)) and (layer0_outputs(5610)));
    outputs(8575) <= not((layer0_outputs(2752)) xor (layer0_outputs(4657)));
    outputs(8576) <= layer0_outputs(1896);
    outputs(8577) <= layer0_outputs(7039);
    outputs(8578) <= layer0_outputs(8160);
    outputs(8579) <= layer0_outputs(7123);
    outputs(8580) <= not((layer0_outputs(4556)) xor (layer0_outputs(8778)));
    outputs(8581) <= layer0_outputs(4734);
    outputs(8582) <= (layer0_outputs(3113)) and (layer0_outputs(1296));
    outputs(8583) <= not(layer0_outputs(8014));
    outputs(8584) <= not((layer0_outputs(9307)) xor (layer0_outputs(6886)));
    outputs(8585) <= not(layer0_outputs(2877)) or (layer0_outputs(8512));
    outputs(8586) <= not((layer0_outputs(352)) xor (layer0_outputs(5868)));
    outputs(8587) <= layer0_outputs(941);
    outputs(8588) <= not(layer0_outputs(8358)) or (layer0_outputs(6643));
    outputs(8589) <= (layer0_outputs(1439)) and not (layer0_outputs(4549));
    outputs(8590) <= not(layer0_outputs(2677)) or (layer0_outputs(723));
    outputs(8591) <= not(layer0_outputs(552));
    outputs(8592) <= not(layer0_outputs(4511)) or (layer0_outputs(2272));
    outputs(8593) <= not(layer0_outputs(9073));
    outputs(8594) <= not((layer0_outputs(4646)) xor (layer0_outputs(1477)));
    outputs(8595) <= (layer0_outputs(4841)) or (layer0_outputs(9353));
    outputs(8596) <= (layer0_outputs(5950)) or (layer0_outputs(4338));
    outputs(8597) <= layer0_outputs(1390);
    outputs(8598) <= not((layer0_outputs(3406)) and (layer0_outputs(9826)));
    outputs(8599) <= not(layer0_outputs(4915));
    outputs(8600) <= layer0_outputs(121);
    outputs(8601) <= (layer0_outputs(10050)) xor (layer0_outputs(4369));
    outputs(8602) <= not(layer0_outputs(7909));
    outputs(8603) <= layer0_outputs(437);
    outputs(8604) <= (layer0_outputs(3986)) or (layer0_outputs(239));
    outputs(8605) <= not(layer0_outputs(5164));
    outputs(8606) <= not((layer0_outputs(7535)) xor (layer0_outputs(8742)));
    outputs(8607) <= layer0_outputs(6206);
    outputs(8608) <= (layer0_outputs(4830)) or (layer0_outputs(3725));
    outputs(8609) <= not(layer0_outputs(2274));
    outputs(8610) <= not(layer0_outputs(9977));
    outputs(8611) <= not(layer0_outputs(1263));
    outputs(8612) <= (layer0_outputs(9325)) or (layer0_outputs(2186));
    outputs(8613) <= not((layer0_outputs(6987)) xor (layer0_outputs(1311)));
    outputs(8614) <= not(layer0_outputs(8822)) or (layer0_outputs(2266));
    outputs(8615) <= (layer0_outputs(3934)) or (layer0_outputs(6585));
    outputs(8616) <= not(layer0_outputs(5088));
    outputs(8617) <= not(layer0_outputs(7761)) or (layer0_outputs(4236));
    outputs(8618) <= (layer0_outputs(6658)) xor (layer0_outputs(316));
    outputs(8619) <= (layer0_outputs(9107)) and not (layer0_outputs(4463));
    outputs(8620) <= layer0_outputs(7620);
    outputs(8621) <= (layer0_outputs(6485)) xor (layer0_outputs(4298));
    outputs(8622) <= not(layer0_outputs(43)) or (layer0_outputs(6169));
    outputs(8623) <= layer0_outputs(8971);
    outputs(8624) <= layer0_outputs(6563);
    outputs(8625) <= (layer0_outputs(4173)) or (layer0_outputs(8892));
    outputs(8626) <= (layer0_outputs(2491)) and not (layer0_outputs(8825));
    outputs(8627) <= layer0_outputs(1957);
    outputs(8628) <= layer0_outputs(1502);
    outputs(8629) <= not((layer0_outputs(4898)) xor (layer0_outputs(394)));
    outputs(8630) <= (layer0_outputs(8785)) and not (layer0_outputs(2505));
    outputs(8631) <= (layer0_outputs(8870)) or (layer0_outputs(3285));
    outputs(8632) <= (layer0_outputs(9124)) and (layer0_outputs(1495));
    outputs(8633) <= (layer0_outputs(3477)) xor (layer0_outputs(3711));
    outputs(8634) <= (layer0_outputs(10023)) and not (layer0_outputs(4930));
    outputs(8635) <= not((layer0_outputs(8553)) xor (layer0_outputs(9992)));
    outputs(8636) <= not(layer0_outputs(9872));
    outputs(8637) <= layer0_outputs(6464);
    outputs(8638) <= layer0_outputs(5582);
    outputs(8639) <= not(layer0_outputs(6836));
    outputs(8640) <= not((layer0_outputs(15)) and (layer0_outputs(4509)));
    outputs(8641) <= (layer0_outputs(1887)) or (layer0_outputs(9650));
    outputs(8642) <= (layer0_outputs(6594)) and not (layer0_outputs(9412));
    outputs(8643) <= not(layer0_outputs(3027));
    outputs(8644) <= (layer0_outputs(38)) xor (layer0_outputs(3011));
    outputs(8645) <= layer0_outputs(5991);
    outputs(8646) <= not((layer0_outputs(2669)) or (layer0_outputs(4017)));
    outputs(8647) <= not((layer0_outputs(5557)) xor (layer0_outputs(8080)));
    outputs(8648) <= not(layer0_outputs(5680));
    outputs(8649) <= not((layer0_outputs(9631)) xor (layer0_outputs(2660)));
    outputs(8650) <= (layer0_outputs(9895)) and not (layer0_outputs(3273));
    outputs(8651) <= not(layer0_outputs(6680)) or (layer0_outputs(6847));
    outputs(8652) <= not(layer0_outputs(4282)) or (layer0_outputs(6635));
    outputs(8653) <= (layer0_outputs(6090)) xor (layer0_outputs(6453));
    outputs(8654) <= not((layer0_outputs(5891)) or (layer0_outputs(9711)));
    outputs(8655) <= not(layer0_outputs(6517)) or (layer0_outputs(9700));
    outputs(8656) <= not(layer0_outputs(2609)) or (layer0_outputs(4356));
    outputs(8657) <= not(layer0_outputs(3498));
    outputs(8658) <= not(layer0_outputs(34)) or (layer0_outputs(6342));
    outputs(8659) <= layer0_outputs(7113);
    outputs(8660) <= (layer0_outputs(1267)) or (layer0_outputs(497));
    outputs(8661) <= not((layer0_outputs(3344)) xor (layer0_outputs(3010)));
    outputs(8662) <= not(layer0_outputs(8565));
    outputs(8663) <= not(layer0_outputs(926));
    outputs(8664) <= not((layer0_outputs(8856)) xor (layer0_outputs(1261)));
    outputs(8665) <= (layer0_outputs(7651)) or (layer0_outputs(4202));
    outputs(8666) <= layer0_outputs(6246);
    outputs(8667) <= (layer0_outputs(247)) or (layer0_outputs(8538));
    outputs(8668) <= not(layer0_outputs(2273));
    outputs(8669) <= not(layer0_outputs(1951)) or (layer0_outputs(2487));
    outputs(8670) <= (layer0_outputs(4191)) xor (layer0_outputs(3709));
    outputs(8671) <= not((layer0_outputs(10182)) xor (layer0_outputs(6943)));
    outputs(8672) <= not(layer0_outputs(5613));
    outputs(8673) <= (layer0_outputs(820)) and not (layer0_outputs(10171));
    outputs(8674) <= not((layer0_outputs(823)) xor (layer0_outputs(10084)));
    outputs(8675) <= (layer0_outputs(6552)) xor (layer0_outputs(7805));
    outputs(8676) <= not((layer0_outputs(7373)) xor (layer0_outputs(4421)));
    outputs(8677) <= not((layer0_outputs(8537)) xor (layer0_outputs(7545)));
    outputs(8678) <= not((layer0_outputs(4203)) xor (layer0_outputs(1143)));
    outputs(8679) <= (layer0_outputs(3269)) xor (layer0_outputs(4734));
    outputs(8680) <= layer0_outputs(4271);
    outputs(8681) <= not(layer0_outputs(9008));
    outputs(8682) <= (layer0_outputs(2512)) xor (layer0_outputs(1260));
    outputs(8683) <= not(layer0_outputs(614));
    outputs(8684) <= not((layer0_outputs(3047)) xor (layer0_outputs(847)));
    outputs(8685) <= not(layer0_outputs(9004)) or (layer0_outputs(4222));
    outputs(8686) <= (layer0_outputs(3934)) or (layer0_outputs(529));
    outputs(8687) <= not(layer0_outputs(10146));
    outputs(8688) <= not(layer0_outputs(2202));
    outputs(8689) <= (layer0_outputs(716)) xor (layer0_outputs(6720));
    outputs(8690) <= layer0_outputs(3653);
    outputs(8691) <= not((layer0_outputs(1826)) xor (layer0_outputs(5017)));
    outputs(8692) <= not(layer0_outputs(7165)) or (layer0_outputs(9593));
    outputs(8693) <= not((layer0_outputs(2087)) xor (layer0_outputs(9605)));
    outputs(8694) <= not((layer0_outputs(8462)) xor (layer0_outputs(810)));
    outputs(8695) <= (layer0_outputs(3819)) xor (layer0_outputs(3171));
    outputs(8696) <= not((layer0_outputs(9638)) xor (layer0_outputs(4385)));
    outputs(8697) <= not(layer0_outputs(821)) or (layer0_outputs(5398));
    outputs(8698) <= not((layer0_outputs(8004)) xor (layer0_outputs(9892)));
    outputs(8699) <= layer0_outputs(10082);
    outputs(8700) <= layer0_outputs(9115);
    outputs(8701) <= not(layer0_outputs(4058));
    outputs(8702) <= not(layer0_outputs(4722)) or (layer0_outputs(6600));
    outputs(8703) <= not((layer0_outputs(727)) xor (layer0_outputs(359)));
    outputs(8704) <= not((layer0_outputs(9883)) xor (layer0_outputs(2262)));
    outputs(8705) <= not(layer0_outputs(9931));
    outputs(8706) <= not(layer0_outputs(1178)) or (layer0_outputs(5300));
    outputs(8707) <= not((layer0_outputs(166)) xor (layer0_outputs(2426)));
    outputs(8708) <= not((layer0_outputs(8566)) and (layer0_outputs(6452)));
    outputs(8709) <= not((layer0_outputs(3913)) xor (layer0_outputs(9798)));
    outputs(8710) <= not(layer0_outputs(9477));
    outputs(8711) <= (layer0_outputs(8639)) xor (layer0_outputs(2225));
    outputs(8712) <= layer0_outputs(8616);
    outputs(8713) <= not(layer0_outputs(7588)) or (layer0_outputs(9571));
    outputs(8714) <= (layer0_outputs(1979)) and (layer0_outputs(3328));
    outputs(8715) <= not(layer0_outputs(1698)) or (layer0_outputs(339));
    outputs(8716) <= not((layer0_outputs(4264)) xor (layer0_outputs(1550)));
    outputs(8717) <= (layer0_outputs(1074)) and not (layer0_outputs(9539));
    outputs(8718) <= layer0_outputs(3672);
    outputs(8719) <= not(layer0_outputs(6609));
    outputs(8720) <= not((layer0_outputs(8662)) and (layer0_outputs(2903)));
    outputs(8721) <= not(layer0_outputs(9535));
    outputs(8722) <= not((layer0_outputs(8170)) xor (layer0_outputs(4392)));
    outputs(8723) <= not(layer0_outputs(600)) or (layer0_outputs(2631));
    outputs(8724) <= (layer0_outputs(1203)) xor (layer0_outputs(8711));
    outputs(8725) <= layer0_outputs(1216);
    outputs(8726) <= (layer0_outputs(2042)) xor (layer0_outputs(1119));
    outputs(8727) <= not(layer0_outputs(54));
    outputs(8728) <= not(layer0_outputs(10097));
    outputs(8729) <= not((layer0_outputs(238)) xor (layer0_outputs(756)));
    outputs(8730) <= not((layer0_outputs(5423)) xor (layer0_outputs(6929)));
    outputs(8731) <= not(layer0_outputs(3429));
    outputs(8732) <= (layer0_outputs(8979)) xor (layer0_outputs(3692));
    outputs(8733) <= (layer0_outputs(6751)) xor (layer0_outputs(1818));
    outputs(8734) <= layer0_outputs(3037);
    outputs(8735) <= layer0_outputs(9199);
    outputs(8736) <= layer0_outputs(846);
    outputs(8737) <= (layer0_outputs(9123)) xor (layer0_outputs(5235));
    outputs(8738) <= (layer0_outputs(4562)) or (layer0_outputs(7754));
    outputs(8739) <= not(layer0_outputs(5040)) or (layer0_outputs(8128));
    outputs(8740) <= not(layer0_outputs(9007)) or (layer0_outputs(9278));
    outputs(8741) <= (layer0_outputs(10211)) xor (layer0_outputs(8148));
    outputs(8742) <= (layer0_outputs(499)) and not (layer0_outputs(6310));
    outputs(8743) <= not((layer0_outputs(8180)) xor (layer0_outputs(7477)));
    outputs(8744) <= (layer0_outputs(6691)) xor (layer0_outputs(3227));
    outputs(8745) <= not(layer0_outputs(2777));
    outputs(8746) <= not(layer0_outputs(365));
    outputs(8747) <= not((layer0_outputs(1159)) xor (layer0_outputs(8224)));
    outputs(8748) <= not(layer0_outputs(2625)) or (layer0_outputs(8124));
    outputs(8749) <= (layer0_outputs(5252)) xor (layer0_outputs(4919));
    outputs(8750) <= (layer0_outputs(3721)) and (layer0_outputs(4077));
    outputs(8751) <= (layer0_outputs(8535)) xor (layer0_outputs(9482));
    outputs(8752) <= layer0_outputs(6602);
    outputs(8753) <= not(layer0_outputs(4702)) or (layer0_outputs(7626));
    outputs(8754) <= not(layer0_outputs(2506));
    outputs(8755) <= (layer0_outputs(1170)) xor (layer0_outputs(8167));
    outputs(8756) <= not((layer0_outputs(1829)) xor (layer0_outputs(3578)));
    outputs(8757) <= not((layer0_outputs(1740)) xor (layer0_outputs(4658)));
    outputs(8758) <= layer0_outputs(1613);
    outputs(8759) <= not((layer0_outputs(9451)) xor (layer0_outputs(8392)));
    outputs(8760) <= not((layer0_outputs(2122)) and (layer0_outputs(5119)));
    outputs(8761) <= layer0_outputs(3038);
    outputs(8762) <= not((layer0_outputs(8783)) xor (layer0_outputs(1308)));
    outputs(8763) <= not(layer0_outputs(2715));
    outputs(8764) <= not(layer0_outputs(5460)) or (layer0_outputs(3295));
    outputs(8765) <= not(layer0_outputs(3776)) or (layer0_outputs(8620));
    outputs(8766) <= not((layer0_outputs(154)) xor (layer0_outputs(5928)));
    outputs(8767) <= layer0_outputs(2251);
    outputs(8768) <= (layer0_outputs(2371)) xor (layer0_outputs(6365));
    outputs(8769) <= not((layer0_outputs(364)) or (layer0_outputs(7915)));
    outputs(8770) <= (layer0_outputs(9843)) xor (layer0_outputs(8030));
    outputs(8771) <= not(layer0_outputs(2573));
    outputs(8772) <= not((layer0_outputs(6881)) xor (layer0_outputs(1450)));
    outputs(8773) <= layer0_outputs(4080);
    outputs(8774) <= layer0_outputs(1800);
    outputs(8775) <= not(layer0_outputs(1522));
    outputs(8776) <= not(layer0_outputs(6019));
    outputs(8777) <= layer0_outputs(6633);
    outputs(8778) <= not(layer0_outputs(9284));
    outputs(8779) <= not((layer0_outputs(4004)) and (layer0_outputs(6344)));
    outputs(8780) <= (layer0_outputs(7441)) or (layer0_outputs(8308));
    outputs(8781) <= not(layer0_outputs(7706)) or (layer0_outputs(8448));
    outputs(8782) <= not((layer0_outputs(6440)) xor (layer0_outputs(7856)));
    outputs(8783) <= layer0_outputs(9741);
    outputs(8784) <= (layer0_outputs(2969)) xor (layer0_outputs(9142));
    outputs(8785) <= not((layer0_outputs(7740)) xor (layer0_outputs(9746)));
    outputs(8786) <= not((layer0_outputs(5171)) xor (layer0_outputs(8034)));
    outputs(8787) <= not((layer0_outputs(3177)) xor (layer0_outputs(1579)));
    outputs(8788) <= (layer0_outputs(1198)) xor (layer0_outputs(3329));
    outputs(8789) <= not(layer0_outputs(509)) or (layer0_outputs(9808));
    outputs(8790) <= layer0_outputs(2704);
    outputs(8791) <= (layer0_outputs(4486)) and not (layer0_outputs(4322));
    outputs(8792) <= (layer0_outputs(3537)) xor (layer0_outputs(9328));
    outputs(8793) <= layer0_outputs(2793);
    outputs(8794) <= layer0_outputs(4381);
    outputs(8795) <= layer0_outputs(2699);
    outputs(8796) <= (layer0_outputs(3412)) xor (layer0_outputs(79));
    outputs(8797) <= not(layer0_outputs(3282)) or (layer0_outputs(819));
    outputs(8798) <= not(layer0_outputs(383));
    outputs(8799) <= not(layer0_outputs(4906)) or (layer0_outputs(3696));
    outputs(8800) <= layer0_outputs(5726);
    outputs(8801) <= (layer0_outputs(5184)) and (layer0_outputs(2767));
    outputs(8802) <= (layer0_outputs(4707)) and not (layer0_outputs(7418));
    outputs(8803) <= (layer0_outputs(571)) xor (layer0_outputs(2262));
    outputs(8804) <= (layer0_outputs(3272)) xor (layer0_outputs(8729));
    outputs(8805) <= not((layer0_outputs(9236)) xor (layer0_outputs(9788)));
    outputs(8806) <= not(layer0_outputs(88));
    outputs(8807) <= not((layer0_outputs(7860)) and (layer0_outputs(3314)));
    outputs(8808) <= not(layer0_outputs(6871));
    outputs(8809) <= not(layer0_outputs(10019)) or (layer0_outputs(4526));
    outputs(8810) <= not((layer0_outputs(6882)) xor (layer0_outputs(5327)));
    outputs(8811) <= (layer0_outputs(8431)) xor (layer0_outputs(3450));
    outputs(8812) <= not((layer0_outputs(1110)) xor (layer0_outputs(5875)));
    outputs(8813) <= not(layer0_outputs(9264));
    outputs(8814) <= layer0_outputs(3884);
    outputs(8815) <= layer0_outputs(4429);
    outputs(8816) <= (layer0_outputs(6047)) or (layer0_outputs(1593));
    outputs(8817) <= not(layer0_outputs(3506)) or (layer0_outputs(4923));
    outputs(8818) <= not((layer0_outputs(6863)) xor (layer0_outputs(953)));
    outputs(8819) <= not((layer0_outputs(2844)) and (layer0_outputs(9293)));
    outputs(8820) <= layer0_outputs(9959);
    outputs(8821) <= layer0_outputs(1754);
    outputs(8822) <= not((layer0_outputs(5225)) xor (layer0_outputs(9229)));
    outputs(8823) <= (layer0_outputs(7181)) xor (layer0_outputs(6325));
    outputs(8824) <= not(layer0_outputs(3013));
    outputs(8825) <= layer0_outputs(6494);
    outputs(8826) <= (layer0_outputs(8038)) xor (layer0_outputs(4826));
    outputs(8827) <= layer0_outputs(5439);
    outputs(8828) <= not((layer0_outputs(2682)) and (layer0_outputs(7315)));
    outputs(8829) <= not(layer0_outputs(8441));
    outputs(8830) <= not((layer0_outputs(6878)) and (layer0_outputs(8246)));
    outputs(8831) <= not(layer0_outputs(4423)) or (layer0_outputs(4928));
    outputs(8832) <= not(layer0_outputs(3989)) or (layer0_outputs(435));
    outputs(8833) <= not(layer0_outputs(8033));
    outputs(8834) <= not((layer0_outputs(6370)) xor (layer0_outputs(1772)));
    outputs(8835) <= not(layer0_outputs(5064));
    outputs(8836) <= not(layer0_outputs(5466));
    outputs(8837) <= layer0_outputs(1295);
    outputs(8838) <= not((layer0_outputs(3386)) xor (layer0_outputs(2708)));
    outputs(8839) <= not((layer0_outputs(585)) and (layer0_outputs(2709)));
    outputs(8840) <= layer0_outputs(2898);
    outputs(8841) <= not(layer0_outputs(7504));
    outputs(8842) <= (layer0_outputs(10200)) or (layer0_outputs(9851));
    outputs(8843) <= (layer0_outputs(4499)) xor (layer0_outputs(7896));
    outputs(8844) <= (layer0_outputs(9693)) or (layer0_outputs(7815));
    outputs(8845) <= (layer0_outputs(3758)) xor (layer0_outputs(575));
    outputs(8846) <= (layer0_outputs(5732)) and not (layer0_outputs(5537));
    outputs(8847) <= (layer0_outputs(2099)) xor (layer0_outputs(9063));
    outputs(8848) <= (layer0_outputs(3269)) or (layer0_outputs(162));
    outputs(8849) <= (layer0_outputs(6746)) xor (layer0_outputs(1788));
    outputs(8850) <= not(layer0_outputs(2706));
    outputs(8851) <= not((layer0_outputs(711)) xor (layer0_outputs(387)));
    outputs(8852) <= not(layer0_outputs(428));
    outputs(8853) <= not(layer0_outputs(4365)) or (layer0_outputs(7890));
    outputs(8854) <= (layer0_outputs(958)) and not (layer0_outputs(5215));
    outputs(8855) <= not((layer0_outputs(7548)) xor (layer0_outputs(5720)));
    outputs(8856) <= layer0_outputs(449);
    outputs(8857) <= not((layer0_outputs(2729)) xor (layer0_outputs(2227)));
    outputs(8858) <= not(layer0_outputs(10032));
    outputs(8859) <= (layer0_outputs(7057)) xor (layer0_outputs(6742));
    outputs(8860) <= not(layer0_outputs(2076)) or (layer0_outputs(363));
    outputs(8861) <= not(layer0_outputs(622)) or (layer0_outputs(3432));
    outputs(8862) <= not(layer0_outputs(9232));
    outputs(8863) <= not(layer0_outputs(4983));
    outputs(8864) <= not(layer0_outputs(9990));
    outputs(8865) <= layer0_outputs(3240);
    outputs(8866) <= not(layer0_outputs(8191)) or (layer0_outputs(5785));
    outputs(8867) <= layer0_outputs(3459);
    outputs(8868) <= not((layer0_outputs(7750)) or (layer0_outputs(1669)));
    outputs(8869) <= (layer0_outputs(3315)) xor (layer0_outputs(111));
    outputs(8870) <= not(layer0_outputs(6431));
    outputs(8871) <= not(layer0_outputs(6457));
    outputs(8872) <= (layer0_outputs(9415)) and not (layer0_outputs(9407));
    outputs(8873) <= not(layer0_outputs(1959));
    outputs(8874) <= layer0_outputs(4877);
    outputs(8875) <= not((layer0_outputs(3563)) xor (layer0_outputs(4341)));
    outputs(8876) <= layer0_outputs(8901);
    outputs(8877) <= (layer0_outputs(3718)) xor (layer0_outputs(5305));
    outputs(8878) <= not(layer0_outputs(1814));
    outputs(8879) <= (layer0_outputs(3214)) or (layer0_outputs(6741));
    outputs(8880) <= (layer0_outputs(8698)) xor (layer0_outputs(6891));
    outputs(8881) <= not((layer0_outputs(2377)) xor (layer0_outputs(8265)));
    outputs(8882) <= not((layer0_outputs(5715)) xor (layer0_outputs(6945)));
    outputs(8883) <= (layer0_outputs(9436)) or (layer0_outputs(6660));
    outputs(8884) <= layer0_outputs(8651);
    outputs(8885) <= not((layer0_outputs(276)) xor (layer0_outputs(4643)));
    outputs(8886) <= layer0_outputs(577);
    outputs(8887) <= not((layer0_outputs(10202)) xor (layer0_outputs(8551)));
    outputs(8888) <= not(layer0_outputs(8144)) or (layer0_outputs(2727));
    outputs(8889) <= layer0_outputs(1390);
    outputs(8890) <= not(layer0_outputs(8260));
    outputs(8891) <= not(layer0_outputs(8705)) or (layer0_outputs(9822));
    outputs(8892) <= not(layer0_outputs(4332));
    outputs(8893) <= (layer0_outputs(5596)) and not (layer0_outputs(3160));
    outputs(8894) <= not(layer0_outputs(5633));
    outputs(8895) <= layer0_outputs(375);
    outputs(8896) <= not((layer0_outputs(316)) xor (layer0_outputs(884)));
    outputs(8897) <= not(layer0_outputs(7332));
    outputs(8898) <= not(layer0_outputs(4518)) or (layer0_outputs(7085));
    outputs(8899) <= not(layer0_outputs(9412));
    outputs(8900) <= not((layer0_outputs(5766)) xor (layer0_outputs(69)));
    outputs(8901) <= (layer0_outputs(3198)) and not (layer0_outputs(9823));
    outputs(8902) <= not(layer0_outputs(5777)) or (layer0_outputs(2655));
    outputs(8903) <= not((layer0_outputs(7657)) xor (layer0_outputs(2745)));
    outputs(8904) <= (layer0_outputs(4979)) and not (layer0_outputs(7348));
    outputs(8905) <= not(layer0_outputs(1414)) or (layer0_outputs(9776));
    outputs(8906) <= layer0_outputs(402);
    outputs(8907) <= not(layer0_outputs(3347));
    outputs(8908) <= (layer0_outputs(3365)) xor (layer0_outputs(6128));
    outputs(8909) <= not(layer0_outputs(4256)) or (layer0_outputs(3000));
    outputs(8910) <= not(layer0_outputs(5636));
    outputs(8911) <= not((layer0_outputs(806)) xor (layer0_outputs(615)));
    outputs(8912) <= not((layer0_outputs(9743)) xor (layer0_outputs(3753)));
    outputs(8913) <= layer0_outputs(9555);
    outputs(8914) <= not((layer0_outputs(6558)) xor (layer0_outputs(3258)));
    outputs(8915) <= not((layer0_outputs(4917)) xor (layer0_outputs(9939)));
    outputs(8916) <= (layer0_outputs(3245)) or (layer0_outputs(5649));
    outputs(8917) <= layer0_outputs(6402);
    outputs(8918) <= (layer0_outputs(1177)) and not (layer0_outputs(2761));
    outputs(8919) <= not((layer0_outputs(8665)) xor (layer0_outputs(5018)));
    outputs(8920) <= not(layer0_outputs(5593));
    outputs(8921) <= not(layer0_outputs(4078)) or (layer0_outputs(9381));
    outputs(8922) <= (layer0_outputs(3062)) or (layer0_outputs(551));
    outputs(8923) <= not(layer0_outputs(925));
    outputs(8924) <= (layer0_outputs(3366)) or (layer0_outputs(2355));
    outputs(8925) <= not((layer0_outputs(3619)) and (layer0_outputs(7045)));
    outputs(8926) <= not(layer0_outputs(4336)) or (layer0_outputs(1934));
    outputs(8927) <= layer0_outputs(5542);
    outputs(8928) <= (layer0_outputs(7000)) and (layer0_outputs(5650));
    outputs(8929) <= not(layer0_outputs(7203));
    outputs(8930) <= (layer0_outputs(7267)) xor (layer0_outputs(5393));
    outputs(8931) <= (layer0_outputs(63)) or (layer0_outputs(3004));
    outputs(8932) <= not(layer0_outputs(6815));
    outputs(8933) <= (layer0_outputs(9292)) and not (layer0_outputs(3503));
    outputs(8934) <= not((layer0_outputs(5870)) and (layer0_outputs(2400)));
    outputs(8935) <= not((layer0_outputs(1336)) and (layer0_outputs(7970)));
    outputs(8936) <= (layer0_outputs(1604)) or (layer0_outputs(4823));
    outputs(8937) <= (layer0_outputs(2216)) xor (layer0_outputs(4938));
    outputs(8938) <= not(layer0_outputs(7589));
    outputs(8939) <= layer0_outputs(8922);
    outputs(8940) <= not(layer0_outputs(7916));
    outputs(8941) <= (layer0_outputs(9358)) or (layer0_outputs(1414));
    outputs(8942) <= not((layer0_outputs(1233)) or (layer0_outputs(4354)));
    outputs(8943) <= not((layer0_outputs(3125)) xor (layer0_outputs(1929)));
    outputs(8944) <= layer0_outputs(3532);
    outputs(8945) <= not((layer0_outputs(9729)) xor (layer0_outputs(3384)));
    outputs(8946) <= not((layer0_outputs(985)) xor (layer0_outputs(2138)));
    outputs(8947) <= not((layer0_outputs(8275)) xor (layer0_outputs(1180)));
    outputs(8948) <= not((layer0_outputs(8684)) and (layer0_outputs(366)));
    outputs(8949) <= not(layer0_outputs(8924));
    outputs(8950) <= layer0_outputs(3889);
    outputs(8951) <= not(layer0_outputs(1522));
    outputs(8952) <= not((layer0_outputs(410)) xor (layer0_outputs(4573)));
    outputs(8953) <= not(layer0_outputs(1065));
    outputs(8954) <= not((layer0_outputs(1954)) xor (layer0_outputs(8253)));
    outputs(8955) <= (layer0_outputs(143)) or (layer0_outputs(6396));
    outputs(8956) <= not(layer0_outputs(10103));
    outputs(8957) <= layer0_outputs(5144);
    outputs(8958) <= not((layer0_outputs(8499)) xor (layer0_outputs(617)));
    outputs(8959) <= not(layer0_outputs(2492));
    outputs(8960) <= (layer0_outputs(3625)) xor (layer0_outputs(8411));
    outputs(8961) <= (layer0_outputs(6763)) xor (layer0_outputs(4147));
    outputs(8962) <= not(layer0_outputs(6269));
    outputs(8963) <= not(layer0_outputs(3632)) or (layer0_outputs(1971));
    outputs(8964) <= not(layer0_outputs(8146));
    outputs(8965) <= not(layer0_outputs(2940));
    outputs(8966) <= (layer0_outputs(5006)) xor (layer0_outputs(8637));
    outputs(8967) <= (layer0_outputs(9467)) and not (layer0_outputs(8605));
    outputs(8968) <= not((layer0_outputs(9047)) and (layer0_outputs(9672)));
    outputs(8969) <= layer0_outputs(7904);
    outputs(8970) <= not(layer0_outputs(5334)) or (layer0_outputs(5505));
    outputs(8971) <= (layer0_outputs(8540)) xor (layer0_outputs(6200));
    outputs(8972) <= layer0_outputs(5692);
    outputs(8973) <= not((layer0_outputs(4317)) and (layer0_outputs(1312)));
    outputs(8974) <= not(layer0_outputs(1455));
    outputs(8975) <= (layer0_outputs(4478)) xor (layer0_outputs(4903));
    outputs(8976) <= layer0_outputs(6298);
    outputs(8977) <= not((layer0_outputs(406)) and (layer0_outputs(2538)));
    outputs(8978) <= not((layer0_outputs(1046)) xor (layer0_outputs(1382)));
    outputs(8979) <= not((layer0_outputs(4142)) xor (layer0_outputs(9298)));
    outputs(8980) <= not(layer0_outputs(6903)) or (layer0_outputs(2959));
    outputs(8981) <= not(layer0_outputs(2415));
    outputs(8982) <= not((layer0_outputs(7877)) xor (layer0_outputs(783)));
    outputs(8983) <= (layer0_outputs(4201)) xor (layer0_outputs(10106));
    outputs(8984) <= not((layer0_outputs(5205)) and (layer0_outputs(3682)));
    outputs(8985) <= layer0_outputs(760);
    outputs(8986) <= not((layer0_outputs(849)) xor (layer0_outputs(3680)));
    outputs(8987) <= not((layer0_outputs(9134)) or (layer0_outputs(1123)));
    outputs(8988) <= not((layer0_outputs(8976)) and (layer0_outputs(4695)));
    outputs(8989) <= (layer0_outputs(6757)) and not (layer0_outputs(4213));
    outputs(8990) <= (layer0_outputs(9421)) xor (layer0_outputs(5172));
    outputs(8991) <= (layer0_outputs(3866)) xor (layer0_outputs(8428));
    outputs(8992) <= not(layer0_outputs(7898));
    outputs(8993) <= (layer0_outputs(6577)) and (layer0_outputs(7390));
    outputs(8994) <= not((layer0_outputs(1239)) and (layer0_outputs(3146)));
    outputs(8995) <= not(layer0_outputs(5369));
    outputs(8996) <= not(layer0_outputs(5693));
    outputs(8997) <= (layer0_outputs(5480)) xor (layer0_outputs(6405));
    outputs(8998) <= not(layer0_outputs(3988)) or (layer0_outputs(4596));
    outputs(8999) <= (layer0_outputs(6423)) xor (layer0_outputs(9985));
    outputs(9000) <= not(layer0_outputs(5405)) or (layer0_outputs(7179));
    outputs(9001) <= layer0_outputs(35);
    outputs(9002) <= layer0_outputs(8182);
    outputs(9003) <= not((layer0_outputs(4430)) xor (layer0_outputs(3155)));
    outputs(9004) <= not(layer0_outputs(4305));
    outputs(9005) <= not(layer0_outputs(6952));
    outputs(9006) <= (layer0_outputs(6341)) xor (layer0_outputs(3461));
    outputs(9007) <= (layer0_outputs(8909)) and not (layer0_outputs(9396));
    outputs(9008) <= not((layer0_outputs(7152)) xor (layer0_outputs(9226)));
    outputs(9009) <= not(layer0_outputs(7597)) or (layer0_outputs(3286));
    outputs(9010) <= layer0_outputs(6330);
    outputs(9011) <= not(layer0_outputs(3581));
    outputs(9012) <= layer0_outputs(9551);
    outputs(9013) <= not(layer0_outputs(6753)) or (layer0_outputs(4557));
    outputs(9014) <= (layer0_outputs(5347)) and not (layer0_outputs(9708));
    outputs(9015) <= (layer0_outputs(5958)) or (layer0_outputs(1438));
    outputs(9016) <= (layer0_outputs(5242)) xor (layer0_outputs(3640));
    outputs(9017) <= not((layer0_outputs(2561)) xor (layer0_outputs(9907)));
    outputs(9018) <= not((layer0_outputs(9652)) xor (layer0_outputs(8493)));
    outputs(9019) <= layer0_outputs(8740);
    outputs(9020) <= not((layer0_outputs(3158)) xor (layer0_outputs(10055)));
    outputs(9021) <= (layer0_outputs(9128)) or (layer0_outputs(6119));
    outputs(9022) <= not(layer0_outputs(5414));
    outputs(9023) <= (layer0_outputs(3325)) or (layer0_outputs(1843));
    outputs(9024) <= (layer0_outputs(2024)) or (layer0_outputs(4181));
    outputs(9025) <= not(layer0_outputs(7443));
    outputs(9026) <= (layer0_outputs(3150)) and not (layer0_outputs(8063));
    outputs(9027) <= not((layer0_outputs(5074)) xor (layer0_outputs(4672)));
    outputs(9028) <= not(layer0_outputs(8399));
    outputs(9029) <= (layer0_outputs(1566)) or (layer0_outputs(5626));
    outputs(9030) <= not(layer0_outputs(2611)) or (layer0_outputs(9261));
    outputs(9031) <= layer0_outputs(4687);
    outputs(9032) <= (layer0_outputs(705)) xor (layer0_outputs(6692));
    outputs(9033) <= not(layer0_outputs(3218));
    outputs(9034) <= layer0_outputs(7120);
    outputs(9035) <= layer0_outputs(224);
    outputs(9036) <= (layer0_outputs(7119)) or (layer0_outputs(7136));
    outputs(9037) <= not(layer0_outputs(1571));
    outputs(9038) <= layer0_outputs(1281);
    outputs(9039) <= not(layer0_outputs(6380));
    outputs(9040) <= not(layer0_outputs(703));
    outputs(9041) <= not((layer0_outputs(155)) and (layer0_outputs(4806)));
    outputs(9042) <= (layer0_outputs(8389)) xor (layer0_outputs(1431));
    outputs(9043) <= not((layer0_outputs(7894)) and (layer0_outputs(7246)));
    outputs(9044) <= not(layer0_outputs(4805));
    outputs(9045) <= not(layer0_outputs(251));
    outputs(9046) <= not(layer0_outputs(7540)) or (layer0_outputs(680));
    outputs(9047) <= not(layer0_outputs(6343));
    outputs(9048) <= (layer0_outputs(7537)) or (layer0_outputs(3100));
    outputs(9049) <= not(layer0_outputs(2322)) or (layer0_outputs(5530));
    outputs(9050) <= (layer0_outputs(5368)) xor (layer0_outputs(2613));
    outputs(9051) <= not((layer0_outputs(4105)) xor (layer0_outputs(2701)));
    outputs(9052) <= not((layer0_outputs(2128)) or (layer0_outputs(5469)));
    outputs(9053) <= not(layer0_outputs(9601));
    outputs(9054) <= not(layer0_outputs(95)) or (layer0_outputs(5027));
    outputs(9055) <= not((layer0_outputs(4782)) xor (layer0_outputs(5417)));
    outputs(9056) <= layer0_outputs(8743);
    outputs(9057) <= not((layer0_outputs(1872)) xor (layer0_outputs(8294)));
    outputs(9058) <= not((layer0_outputs(6639)) or (layer0_outputs(4490)));
    outputs(9059) <= not((layer0_outputs(5084)) xor (layer0_outputs(1484)));
    outputs(9060) <= (layer0_outputs(6279)) or (layer0_outputs(1846));
    outputs(9061) <= not((layer0_outputs(10088)) xor (layer0_outputs(5354)));
    outputs(9062) <= not((layer0_outputs(569)) xor (layer0_outputs(3010)));
    outputs(9063) <= layer0_outputs(3264);
    outputs(9064) <= not((layer0_outputs(219)) or (layer0_outputs(7097)));
    outputs(9065) <= layer0_outputs(8445);
    outputs(9066) <= layer0_outputs(239);
    outputs(9067) <= not(layer0_outputs(5680));
    outputs(9068) <= (layer0_outputs(7083)) and not (layer0_outputs(3779));
    outputs(9069) <= not((layer0_outputs(9083)) xor (layer0_outputs(6291)));
    outputs(9070) <= not((layer0_outputs(5171)) xor (layer0_outputs(4263)));
    outputs(9071) <= (layer0_outputs(4882)) or (layer0_outputs(4837));
    outputs(9072) <= (layer0_outputs(1628)) xor (layer0_outputs(2596));
    outputs(9073) <= not(layer0_outputs(9442));
    outputs(9074) <= (layer0_outputs(6470)) xor (layer0_outputs(2372));
    outputs(9075) <= (layer0_outputs(3141)) or (layer0_outputs(7506));
    outputs(9076) <= (layer0_outputs(3696)) xor (layer0_outputs(6551));
    outputs(9077) <= not((layer0_outputs(4251)) or (layer0_outputs(6042)));
    outputs(9078) <= not(layer0_outputs(4004)) or (layer0_outputs(453));
    outputs(9079) <= (layer0_outputs(3887)) or (layer0_outputs(2409));
    outputs(9080) <= not(layer0_outputs(2404)) or (layer0_outputs(4685));
    outputs(9081) <= not((layer0_outputs(8277)) xor (layer0_outputs(1212)));
    outputs(9082) <= not((layer0_outputs(619)) xor (layer0_outputs(1066)));
    outputs(9083) <= (layer0_outputs(8756)) xor (layer0_outputs(2671));
    outputs(9084) <= (layer0_outputs(7274)) or (layer0_outputs(4283));
    outputs(9085) <= not(layer0_outputs(5996));
    outputs(9086) <= not(layer0_outputs(9335));
    outputs(9087) <= (layer0_outputs(1299)) xor (layer0_outputs(2916));
    outputs(9088) <= layer0_outputs(9526);
    outputs(9089) <= not(layer0_outputs(9501)) or (layer0_outputs(8563));
    outputs(9090) <= (layer0_outputs(5466)) xor (layer0_outputs(1926));
    outputs(9091) <= (layer0_outputs(425)) or (layer0_outputs(6231));
    outputs(9092) <= not(layer0_outputs(6672));
    outputs(9093) <= not(layer0_outputs(4097));
    outputs(9094) <= (layer0_outputs(546)) xor (layer0_outputs(4694));
    outputs(9095) <= layer0_outputs(1288);
    outputs(9096) <= not(layer0_outputs(5104));
    outputs(9097) <= not((layer0_outputs(3860)) and (layer0_outputs(5088)));
    outputs(9098) <= layer0_outputs(3291);
    outputs(9099) <= not(layer0_outputs(2481));
    outputs(9100) <= layer0_outputs(6810);
    outputs(9101) <= not((layer0_outputs(7737)) xor (layer0_outputs(742)));
    outputs(9102) <= not(layer0_outputs(4361));
    outputs(9103) <= layer0_outputs(3612);
    outputs(9104) <= (layer0_outputs(7695)) xor (layer0_outputs(5930));
    outputs(9105) <= not(layer0_outputs(1661)) or (layer0_outputs(9475));
    outputs(9106) <= not(layer0_outputs(9035)) or (layer0_outputs(2159));
    outputs(9107) <= not(layer0_outputs(7096)) or (layer0_outputs(9789));
    outputs(9108) <= not((layer0_outputs(3841)) xor (layer0_outputs(4862)));
    outputs(9109) <= (layer0_outputs(4454)) xor (layer0_outputs(9143));
    outputs(9110) <= (layer0_outputs(9355)) or (layer0_outputs(8002));
    outputs(9111) <= (layer0_outputs(2725)) xor (layer0_outputs(6950));
    outputs(9112) <= (layer0_outputs(2970)) and (layer0_outputs(170));
    outputs(9113) <= not((layer0_outputs(9178)) xor (layer0_outputs(8661)));
    outputs(9114) <= not(layer0_outputs(3495)) or (layer0_outputs(4277));
    outputs(9115) <= not(layer0_outputs(9517));
    outputs(9116) <= not((layer0_outputs(1055)) and (layer0_outputs(7595)));
    outputs(9117) <= not(layer0_outputs(6553));
    outputs(9118) <= (layer0_outputs(4021)) or (layer0_outputs(5158));
    outputs(9119) <= not((layer0_outputs(628)) xor (layer0_outputs(6551)));
    outputs(9120) <= not(layer0_outputs(329));
    outputs(9121) <= not(layer0_outputs(2657));
    outputs(9122) <= not(layer0_outputs(1075)) or (layer0_outputs(6703));
    outputs(9123) <= not(layer0_outputs(8561)) or (layer0_outputs(5554));
    outputs(9124) <= not(layer0_outputs(335));
    outputs(9125) <= (layer0_outputs(7809)) and not (layer0_outputs(863));
    outputs(9126) <= layer0_outputs(3908);
    outputs(9127) <= layer0_outputs(3381);
    outputs(9128) <= not(layer0_outputs(1905)) or (layer0_outputs(1007));
    outputs(9129) <= (layer0_outputs(8931)) xor (layer0_outputs(1598));
    outputs(9130) <= layer0_outputs(4235);
    outputs(9131) <= not(layer0_outputs(9200));
    outputs(9132) <= (layer0_outputs(9171)) and not (layer0_outputs(3372));
    outputs(9133) <= layer0_outputs(9720);
    outputs(9134) <= not((layer0_outputs(6081)) xor (layer0_outputs(7858)));
    outputs(9135) <= not((layer0_outputs(6247)) xor (layer0_outputs(7199)));
    outputs(9136) <= (layer0_outputs(794)) or (layer0_outputs(2359));
    outputs(9137) <= layer0_outputs(6719);
    outputs(9138) <= layer0_outputs(2783);
    outputs(9139) <= layer0_outputs(9960);
    outputs(9140) <= not((layer0_outputs(8901)) xor (layer0_outputs(8863)));
    outputs(9141) <= (layer0_outputs(984)) xor (layer0_outputs(3016));
    outputs(9142) <= not(layer0_outputs(5660));
    outputs(9143) <= not(layer0_outputs(6573));
    outputs(9144) <= layer0_outputs(7013);
    outputs(9145) <= (layer0_outputs(5072)) or (layer0_outputs(3879));
    outputs(9146) <= not((layer0_outputs(3482)) and (layer0_outputs(7687)));
    outputs(9147) <= not((layer0_outputs(6957)) xor (layer0_outputs(9038)));
    outputs(9148) <= not((layer0_outputs(6282)) xor (layer0_outputs(1303)));
    outputs(9149) <= not(layer0_outputs(8665));
    outputs(9150) <= not((layer0_outputs(2351)) xor (layer0_outputs(593)));
    outputs(9151) <= (layer0_outputs(9692)) xor (layer0_outputs(8568));
    outputs(9152) <= not(layer0_outputs(7861));
    outputs(9153) <= (layer0_outputs(9371)) xor (layer0_outputs(2885));
    outputs(9154) <= not((layer0_outputs(3140)) or (layer0_outputs(8828)));
    outputs(9155) <= not(layer0_outputs(7150));
    outputs(9156) <= not(layer0_outputs(1786)) or (layer0_outputs(1780));
    outputs(9157) <= (layer0_outputs(4129)) xor (layer0_outputs(2823));
    outputs(9158) <= not(layer0_outputs(4179));
    outputs(9159) <= not((layer0_outputs(9879)) or (layer0_outputs(2528)));
    outputs(9160) <= (layer0_outputs(748)) xor (layer0_outputs(10196));
    outputs(9161) <= not(layer0_outputs(6560)) or (layer0_outputs(5914));
    outputs(9162) <= layer0_outputs(7032);
    outputs(9163) <= (layer0_outputs(4197)) xor (layer0_outputs(9009));
    outputs(9164) <= not(layer0_outputs(2539)) or (layer0_outputs(1921));
    outputs(9165) <= (layer0_outputs(6482)) xor (layer0_outputs(1808));
    outputs(9166) <= not((layer0_outputs(8058)) and (layer0_outputs(8869)));
    outputs(9167) <= layer0_outputs(3059);
    outputs(9168) <= not((layer0_outputs(9885)) xor (layer0_outputs(4515)));
    outputs(9169) <= layer0_outputs(4456);
    outputs(9170) <= layer0_outputs(9687);
    outputs(9171) <= not(layer0_outputs(9256)) or (layer0_outputs(558));
    outputs(9172) <= (layer0_outputs(516)) xor (layer0_outputs(9976));
    outputs(9173) <= layer0_outputs(4660);
    outputs(9174) <= not((layer0_outputs(938)) and (layer0_outputs(3235)));
    outputs(9175) <= not((layer0_outputs(480)) xor (layer0_outputs(9847)));
    outputs(9176) <= layer0_outputs(805);
    outputs(9177) <= not(layer0_outputs(9549));
    outputs(9178) <= (layer0_outputs(6890)) and (layer0_outputs(8142));
    outputs(9179) <= not(layer0_outputs(4395)) or (layer0_outputs(6985));
    outputs(9180) <= not(layer0_outputs(6327)) or (layer0_outputs(7603));
    outputs(9181) <= (layer0_outputs(2345)) xor (layer0_outputs(3392));
    outputs(9182) <= not(layer0_outputs(7066));
    outputs(9183) <= not((layer0_outputs(9193)) xor (layer0_outputs(5113)));
    outputs(9184) <= not(layer0_outputs(1284));
    outputs(9185) <= layer0_outputs(8573);
    outputs(9186) <= not(layer0_outputs(7549)) or (layer0_outputs(5061));
    outputs(9187) <= not((layer0_outputs(7500)) xor (layer0_outputs(181)));
    outputs(9188) <= (layer0_outputs(250)) xor (layer0_outputs(4347));
    outputs(9189) <= (layer0_outputs(3533)) and (layer0_outputs(5328));
    outputs(9190) <= not((layer0_outputs(6705)) xor (layer0_outputs(3927)));
    outputs(9191) <= layer0_outputs(2183);
    outputs(9192) <= not((layer0_outputs(1238)) xor (layer0_outputs(8185)));
    outputs(9193) <= (layer0_outputs(2436)) xor (layer0_outputs(414));
    outputs(9194) <= (layer0_outputs(1119)) or (layer0_outputs(2418));
    outputs(9195) <= not(layer0_outputs(5109)) or (layer0_outputs(923));
    outputs(9196) <= not((layer0_outputs(8018)) and (layer0_outputs(5359)));
    outputs(9197) <= not(layer0_outputs(1944)) or (layer0_outputs(3479));
    outputs(9198) <= (layer0_outputs(10224)) xor (layer0_outputs(3857));
    outputs(9199) <= not((layer0_outputs(8297)) xor (layer0_outputs(3311)));
    outputs(9200) <= layer0_outputs(7696);
    outputs(9201) <= not(layer0_outputs(7575));
    outputs(9202) <= (layer0_outputs(4607)) xor (layer0_outputs(622));
    outputs(9203) <= not((layer0_outputs(1240)) and (layer0_outputs(4087)));
    outputs(9204) <= not(layer0_outputs(1657)) or (layer0_outputs(4400));
    outputs(9205) <= not(layer0_outputs(9659));
    outputs(9206) <= (layer0_outputs(10201)) xor (layer0_outputs(1234));
    outputs(9207) <= not(layer0_outputs(7894));
    outputs(9208) <= not(layer0_outputs(3873)) or (layer0_outputs(8490));
    outputs(9209) <= layer0_outputs(2091);
    outputs(9210) <= not(layer0_outputs(5279));
    outputs(9211) <= (layer0_outputs(5233)) xor (layer0_outputs(6631));
    outputs(9212) <= not(layer0_outputs(9806)) or (layer0_outputs(2802));
    outputs(9213) <= not(layer0_outputs(3054));
    outputs(9214) <= not(layer0_outputs(1654));
    outputs(9215) <= not(layer0_outputs(6217)) or (layer0_outputs(5471));
    outputs(9216) <= not(layer0_outputs(7106));
    outputs(9217) <= not(layer0_outputs(3166));
    outputs(9218) <= (layer0_outputs(8831)) and (layer0_outputs(9190));
    outputs(9219) <= (layer0_outputs(24)) and (layer0_outputs(4124));
    outputs(9220) <= not(layer0_outputs(4225));
    outputs(9221) <= not((layer0_outputs(9702)) xor (layer0_outputs(2285)));
    outputs(9222) <= (layer0_outputs(9146)) xor (layer0_outputs(6735));
    outputs(9223) <= (layer0_outputs(6841)) and not (layer0_outputs(3308));
    outputs(9224) <= layer0_outputs(6387);
    outputs(9225) <= not(layer0_outputs(9514));
    outputs(9226) <= layer0_outputs(8413);
    outputs(9227) <= layer0_outputs(3230);
    outputs(9228) <= not(layer0_outputs(2721)) or (layer0_outputs(1399));
    outputs(9229) <= not((layer0_outputs(5344)) or (layer0_outputs(8653)));
    outputs(9230) <= not((layer0_outputs(8725)) xor (layer0_outputs(8292)));
    outputs(9231) <= not(layer0_outputs(6892));
    outputs(9232) <= (layer0_outputs(6545)) xor (layer0_outputs(405));
    outputs(9233) <= not((layer0_outputs(61)) xor (layer0_outputs(1083)));
    outputs(9234) <= (layer0_outputs(9457)) xor (layer0_outputs(3119));
    outputs(9235) <= (layer0_outputs(4205)) xor (layer0_outputs(5700));
    outputs(9236) <= (layer0_outputs(918)) and not (layer0_outputs(2927));
    outputs(9237) <= (layer0_outputs(9103)) and (layer0_outputs(5576));
    outputs(9238) <= not(layer0_outputs(355));
    outputs(9239) <= not((layer0_outputs(5849)) and (layer0_outputs(10232)));
    outputs(9240) <= layer0_outputs(8387);
    outputs(9241) <= not((layer0_outputs(9685)) xor (layer0_outputs(9226)));
    outputs(9242) <= (layer0_outputs(7428)) xor (layer0_outputs(9757));
    outputs(9243) <= (layer0_outputs(3340)) xor (layer0_outputs(2305));
    outputs(9244) <= layer0_outputs(9904);
    outputs(9245) <= not((layer0_outputs(8104)) xor (layer0_outputs(8830)));
    outputs(9246) <= not(layer0_outputs(1848));
    outputs(9247) <= layer0_outputs(2474);
    outputs(9248) <= (layer0_outputs(3082)) and (layer0_outputs(5816));
    outputs(9249) <= (layer0_outputs(2467)) and (layer0_outputs(800));
    outputs(9250) <= not((layer0_outputs(2050)) or (layer0_outputs(5590)));
    outputs(9251) <= not(layer0_outputs(1130));
    outputs(9252) <= not(layer0_outputs(315)) or (layer0_outputs(6666));
    outputs(9253) <= (layer0_outputs(7488)) and not (layer0_outputs(2256));
    outputs(9254) <= '0';
    outputs(9255) <= (layer0_outputs(8868)) and not (layer0_outputs(5641));
    outputs(9256) <= not(layer0_outputs(5322));
    outputs(9257) <= (layer0_outputs(8209)) xor (layer0_outputs(5050));
    outputs(9258) <= layer0_outputs(4688);
    outputs(9259) <= not((layer0_outputs(1008)) or (layer0_outputs(8382)));
    outputs(9260) <= layer0_outputs(6662);
    outputs(9261) <= (layer0_outputs(5428)) xor (layer0_outputs(5802));
    outputs(9262) <= (layer0_outputs(2226)) and not (layer0_outputs(9413));
    outputs(9263) <= (layer0_outputs(10042)) and not (layer0_outputs(9484));
    outputs(9264) <= layer0_outputs(6752);
    outputs(9265) <= (layer0_outputs(9505)) xor (layer0_outputs(8829));
    outputs(9266) <= not(layer0_outputs(2063));
    outputs(9267) <= (layer0_outputs(3883)) and not (layer0_outputs(6743));
    outputs(9268) <= (layer0_outputs(5832)) xor (layer0_outputs(6311));
    outputs(9269) <= not(layer0_outputs(8633)) or (layer0_outputs(8571));
    outputs(9270) <= not(layer0_outputs(5946));
    outputs(9271) <= not(layer0_outputs(2511));
    outputs(9272) <= not((layer0_outputs(1365)) xor (layer0_outputs(2286)));
    outputs(9273) <= not(layer0_outputs(8637));
    outputs(9274) <= (layer0_outputs(3662)) xor (layer0_outputs(6614));
    outputs(9275) <= not((layer0_outputs(2890)) xor (layer0_outputs(3334)));
    outputs(9276) <= not(layer0_outputs(1960));
    outputs(9277) <= layer0_outputs(1846);
    outputs(9278) <= not(layer0_outputs(3700));
    outputs(9279) <= not((layer0_outputs(7374)) xor (layer0_outputs(6769)));
    outputs(9280) <= not(layer0_outputs(2529));
    outputs(9281) <= not((layer0_outputs(6826)) xor (layer0_outputs(9677)));
    outputs(9282) <= (layer0_outputs(4855)) or (layer0_outputs(6464));
    outputs(9283) <= layer0_outputs(8368);
    outputs(9284) <= layer0_outputs(7927);
    outputs(9285) <= not(layer0_outputs(5944));
    outputs(9286) <= (layer0_outputs(5975)) and (layer0_outputs(4314));
    outputs(9287) <= not((layer0_outputs(6403)) or (layer0_outputs(1754)));
    outputs(9288) <= not(layer0_outputs(426));
    outputs(9289) <= (layer0_outputs(3354)) xor (layer0_outputs(7241));
    outputs(9290) <= not((layer0_outputs(1857)) and (layer0_outputs(444)));
    outputs(9291) <= (layer0_outputs(537)) xor (layer0_outputs(6099));
    outputs(9292) <= (layer0_outputs(9541)) and not (layer0_outputs(2747));
    outputs(9293) <= not(layer0_outputs(3918));
    outputs(9294) <= (layer0_outputs(5614)) xor (layer0_outputs(3062));
    outputs(9295) <= layer0_outputs(6788);
    outputs(9296) <= (layer0_outputs(8594)) xor (layer0_outputs(9473));
    outputs(9297) <= (layer0_outputs(3948)) and not (layer0_outputs(749));
    outputs(9298) <= (layer0_outputs(4325)) xor (layer0_outputs(4678));
    outputs(9299) <= not(layer0_outputs(2403));
    outputs(9300) <= (layer0_outputs(927)) xor (layer0_outputs(9774));
    outputs(9301) <= not((layer0_outputs(2477)) xor (layer0_outputs(6656)));
    outputs(9302) <= (layer0_outputs(7681)) xor (layer0_outputs(3562));
    outputs(9303) <= not(layer0_outputs(5158));
    outputs(9304) <= (layer0_outputs(7700)) and (layer0_outputs(7102));
    outputs(9305) <= layer0_outputs(5284);
    outputs(9306) <= layer0_outputs(8688);
    outputs(9307) <= layer0_outputs(2015);
    outputs(9308) <= not(layer0_outputs(6579));
    outputs(9309) <= not((layer0_outputs(1307)) xor (layer0_outputs(9901)));
    outputs(9310) <= (layer0_outputs(109)) and not (layer0_outputs(1093));
    outputs(9311) <= (layer0_outputs(8675)) xor (layer0_outputs(472));
    outputs(9312) <= not((layer0_outputs(10000)) and (layer0_outputs(934)));
    outputs(9313) <= layer0_outputs(5488);
    outputs(9314) <= not(layer0_outputs(6130));
    outputs(9315) <= not((layer0_outputs(5960)) xor (layer0_outputs(2710)));
    outputs(9316) <= layer0_outputs(7137);
    outputs(9317) <= (layer0_outputs(2228)) xor (layer0_outputs(16));
    outputs(9318) <= not((layer0_outputs(6125)) xor (layer0_outputs(847)));
    outputs(9319) <= layer0_outputs(2571);
    outputs(9320) <= not((layer0_outputs(329)) or (layer0_outputs(9160)));
    outputs(9321) <= not((layer0_outputs(4128)) xor (layer0_outputs(198)));
    outputs(9322) <= (layer0_outputs(6069)) xor (layer0_outputs(4144));
    outputs(9323) <= not((layer0_outputs(3901)) xor (layer0_outputs(7303)));
    outputs(9324) <= not(layer0_outputs(7453)) or (layer0_outputs(145));
    outputs(9325) <= not(layer0_outputs(9665));
    outputs(9326) <= layer0_outputs(5036);
    outputs(9327) <= not((layer0_outputs(9305)) xor (layer0_outputs(8750)));
    outputs(9328) <= layer0_outputs(10128);
    outputs(9329) <= (layer0_outputs(2032)) xor (layer0_outputs(2818));
    outputs(9330) <= not(layer0_outputs(7001)) or (layer0_outputs(1997));
    outputs(9331) <= not(layer0_outputs(7878)) or (layer0_outputs(8190));
    outputs(9332) <= (layer0_outputs(5186)) xor (layer0_outputs(17));
    outputs(9333) <= (layer0_outputs(4047)) xor (layer0_outputs(2290));
    outputs(9334) <= layer0_outputs(5338);
    outputs(9335) <= (layer0_outputs(4544)) xor (layer0_outputs(5667));
    outputs(9336) <= not(layer0_outputs(3043));
    outputs(9337) <= (layer0_outputs(6688)) and not (layer0_outputs(5575));
    outputs(9338) <= not((layer0_outputs(5161)) xor (layer0_outputs(1228)));
    outputs(9339) <= not(layer0_outputs(7464));
    outputs(9340) <= layer0_outputs(2574);
    outputs(9341) <= layer0_outputs(5626);
    outputs(9342) <= not((layer0_outputs(5752)) xor (layer0_outputs(6963)));
    outputs(9343) <= layer0_outputs(748);
    outputs(9344) <= not(layer0_outputs(3455));
    outputs(9345) <= not(layer0_outputs(7994));
    outputs(9346) <= layer0_outputs(7024);
    outputs(9347) <= not(layer0_outputs(9804));
    outputs(9348) <= layer0_outputs(9048);
    outputs(9349) <= (layer0_outputs(9702)) xor (layer0_outputs(3270));
    outputs(9350) <= not(layer0_outputs(6340));
    outputs(9351) <= (layer0_outputs(1222)) and (layer0_outputs(5907));
    outputs(9352) <= not((layer0_outputs(5387)) xor (layer0_outputs(4374)));
    outputs(9353) <= (layer0_outputs(7033)) xor (layer0_outputs(7226));
    outputs(9354) <= not(layer0_outputs(8846));
    outputs(9355) <= layer0_outputs(8807);
    outputs(9356) <= (layer0_outputs(7160)) and (layer0_outputs(31));
    outputs(9357) <= layer0_outputs(1213);
    outputs(9358) <= layer0_outputs(4269);
    outputs(9359) <= (layer0_outputs(5721)) and not (layer0_outputs(7186));
    outputs(9360) <= not((layer0_outputs(9637)) and (layer0_outputs(5943)));
    outputs(9361) <= (layer0_outputs(7652)) and not (layer0_outputs(9154));
    outputs(9362) <= layer0_outputs(3401);
    outputs(9363) <= not(layer0_outputs(3101));
    outputs(9364) <= (layer0_outputs(1983)) and not (layer0_outputs(3034));
    outputs(9365) <= (layer0_outputs(5477)) and not (layer0_outputs(1294));
    outputs(9366) <= not(layer0_outputs(5506));
    outputs(9367) <= not((layer0_outputs(5995)) xor (layer0_outputs(7833)));
    outputs(9368) <= (layer0_outputs(7996)) xor (layer0_outputs(401));
    outputs(9369) <= (layer0_outputs(10120)) and (layer0_outputs(931));
    outputs(9370) <= layer0_outputs(1048);
    outputs(9371) <= layer0_outputs(7508);
    outputs(9372) <= not(layer0_outputs(5407)) or (layer0_outputs(6640));
    outputs(9373) <= not((layer0_outputs(9694)) and (layer0_outputs(6288)));
    outputs(9374) <= not(layer0_outputs(2712));
    outputs(9375) <= layer0_outputs(4493);
    outputs(9376) <= layer0_outputs(7205);
    outputs(9377) <= (layer0_outputs(4768)) xor (layer0_outputs(8440));
    outputs(9378) <= (layer0_outputs(7607)) and (layer0_outputs(3856));
    outputs(9379) <= not((layer0_outputs(8924)) xor (layer0_outputs(548)));
    outputs(9380) <= (layer0_outputs(2871)) xor (layer0_outputs(5276));
    outputs(9381) <= not((layer0_outputs(6366)) xor (layer0_outputs(1020)));
    outputs(9382) <= (layer0_outputs(3853)) and not (layer0_outputs(8300));
    outputs(9383) <= not(layer0_outputs(6659));
    outputs(9384) <= layer0_outputs(1967);
    outputs(9385) <= not(layer0_outputs(2577));
    outputs(9386) <= not(layer0_outputs(8338));
    outputs(9387) <= (layer0_outputs(4769)) and not (layer0_outputs(2842));
    outputs(9388) <= not((layer0_outputs(3086)) xor (layer0_outputs(9289)));
    outputs(9389) <= layer0_outputs(831);
    outputs(9390) <= (layer0_outputs(1316)) xor (layer0_outputs(752));
    outputs(9391) <= not(layer0_outputs(5976));
    outputs(9392) <= (layer0_outputs(9878)) xor (layer0_outputs(6270));
    outputs(9393) <= (layer0_outputs(1689)) xor (layer0_outputs(84));
    outputs(9394) <= (layer0_outputs(734)) and not (layer0_outputs(1840));
    outputs(9395) <= (layer0_outputs(9775)) xor (layer0_outputs(1683));
    outputs(9396) <= not((layer0_outputs(6363)) or (layer0_outputs(1525)));
    outputs(9397) <= (layer0_outputs(1562)) xor (layer0_outputs(2901));
    outputs(9398) <= not((layer0_outputs(8808)) xor (layer0_outputs(591)));
    outputs(9399) <= (layer0_outputs(6767)) and not (layer0_outputs(8927));
    outputs(9400) <= layer0_outputs(4565);
    outputs(9401) <= (layer0_outputs(50)) xor (layer0_outputs(8400));
    outputs(9402) <= (layer0_outputs(7888)) xor (layer0_outputs(4133));
    outputs(9403) <= layer0_outputs(883);
    outputs(9404) <= (layer0_outputs(8702)) and not (layer0_outputs(2233));
    outputs(9405) <= (layer0_outputs(3153)) xor (layer0_outputs(4741));
    outputs(9406) <= layer0_outputs(10098);
    outputs(9407) <= layer0_outputs(8748);
    outputs(9408) <= (layer0_outputs(1330)) and (layer0_outputs(5390));
    outputs(9409) <= (layer0_outputs(3186)) and (layer0_outputs(2961));
    outputs(9410) <= layer0_outputs(3065);
    outputs(9411) <= not(layer0_outputs(1013));
    outputs(9412) <= (layer0_outputs(4728)) and not (layer0_outputs(3646));
    outputs(9413) <= not(layer0_outputs(5492));
    outputs(9414) <= not((layer0_outputs(8903)) xor (layer0_outputs(2595)));
    outputs(9415) <= not(layer0_outputs(10087));
    outputs(9416) <= not(layer0_outputs(1614));
    outputs(9417) <= (layer0_outputs(2090)) and (layer0_outputs(4964));
    outputs(9418) <= not((layer0_outputs(5965)) xor (layer0_outputs(10049)));
    outputs(9419) <= not(layer0_outputs(203));
    outputs(9420) <= (layer0_outputs(2241)) xor (layer0_outputs(2321));
    outputs(9421) <= layer0_outputs(7063);
    outputs(9422) <= layer0_outputs(3142);
    outputs(9423) <= not(layer0_outputs(2410));
    outputs(9424) <= layer0_outputs(8351);
    outputs(9425) <= layer0_outputs(7986);
    outputs(9426) <= (layer0_outputs(7174)) xor (layer0_outputs(1903));
    outputs(9427) <= not(layer0_outputs(1282)) or (layer0_outputs(6791));
    outputs(9428) <= layer0_outputs(7172);
    outputs(9429) <= (layer0_outputs(7642)) and not (layer0_outputs(1393));
    outputs(9430) <= not(layer0_outputs(9002));
    outputs(9431) <= (layer0_outputs(8634)) and not (layer0_outputs(6627));
    outputs(9432) <= not(layer0_outputs(5124));
    outputs(9433) <= not(layer0_outputs(5319)) or (layer0_outputs(966));
    outputs(9434) <= (layer0_outputs(9731)) and not (layer0_outputs(1826));
    outputs(9435) <= layer0_outputs(692);
    outputs(9436) <= not((layer0_outputs(4832)) xor (layer0_outputs(6922)));
    outputs(9437) <= not((layer0_outputs(7353)) xor (layer0_outputs(4373)));
    outputs(9438) <= (layer0_outputs(9254)) and (layer0_outputs(7871));
    outputs(9439) <= not(layer0_outputs(6307));
    outputs(9440) <= layer0_outputs(7358);
    outputs(9441) <= not((layer0_outputs(1498)) xor (layer0_outputs(3239)));
    outputs(9442) <= (layer0_outputs(6385)) or (layer0_outputs(10134));
    outputs(9443) <= layer0_outputs(4075);
    outputs(9444) <= not(layer0_outputs(3656));
    outputs(9445) <= not((layer0_outputs(2083)) xor (layer0_outputs(9153)));
    outputs(9446) <= not(layer0_outputs(9428));
    outputs(9447) <= not(layer0_outputs(2316));
    outputs(9448) <= layer0_outputs(5106);
    outputs(9449) <= not((layer0_outputs(868)) xor (layer0_outputs(7900)));
    outputs(9450) <= layer0_outputs(3692);
    outputs(9451) <= not(layer0_outputs(4207));
    outputs(9452) <= layer0_outputs(7218);
    outputs(9453) <= not(layer0_outputs(1646));
    outputs(9454) <= layer0_outputs(1714);
    outputs(9455) <= (layer0_outputs(4531)) xor (layer0_outputs(8465));
    outputs(9456) <= (layer0_outputs(9309)) and (layer0_outputs(6538));
    outputs(9457) <= (layer0_outputs(2812)) and not (layer0_outputs(9896));
    outputs(9458) <= not((layer0_outputs(9599)) xor (layer0_outputs(903)));
    outputs(9459) <= not(layer0_outputs(8915));
    outputs(9460) <= layer0_outputs(2308);
    outputs(9461) <= not(layer0_outputs(6561));
    outputs(9462) <= (layer0_outputs(1041)) and (layer0_outputs(4749));
    outputs(9463) <= (layer0_outputs(1397)) and not (layer0_outputs(4344));
    outputs(9464) <= not(layer0_outputs(4118)) or (layer0_outputs(1890));
    outputs(9465) <= layer0_outputs(9848);
    outputs(9466) <= (layer0_outputs(2991)) and not (layer0_outputs(6593));
    outputs(9467) <= not((layer0_outputs(9497)) or (layer0_outputs(3780)));
    outputs(9468) <= not((layer0_outputs(4497)) or (layer0_outputs(1137)));
    outputs(9469) <= layer0_outputs(4616);
    outputs(9470) <= layer0_outputs(7811);
    outputs(9471) <= (layer0_outputs(5734)) xor (layer0_outputs(2873));
    outputs(9472) <= (layer0_outputs(6518)) and not (layer0_outputs(861));
    outputs(9473) <= (layer0_outputs(6022)) and not (layer0_outputs(7632));
    outputs(9474) <= not(layer0_outputs(8619));
    outputs(9475) <= (layer0_outputs(5321)) xor (layer0_outputs(5396));
    outputs(9476) <= layer0_outputs(7084);
    outputs(9477) <= (layer0_outputs(7749)) xor (layer0_outputs(6800));
    outputs(9478) <= layer0_outputs(4028);
    outputs(9479) <= not((layer0_outputs(6016)) or (layer0_outputs(2193)));
    outputs(9480) <= not((layer0_outputs(9096)) or (layer0_outputs(9667)));
    outputs(9481) <= layer0_outputs(9179);
    outputs(9482) <= layer0_outputs(9216);
    outputs(9483) <= not(layer0_outputs(641)) or (layer0_outputs(1027));
    outputs(9484) <= (layer0_outputs(6726)) and not (layer0_outputs(9083));
    outputs(9485) <= layer0_outputs(1461);
    outputs(9486) <= not(layer0_outputs(5116));
    outputs(9487) <= layer0_outputs(7595);
    outputs(9488) <= not(layer0_outputs(3203)) or (layer0_outputs(1022));
    outputs(9489) <= (layer0_outputs(1948)) and not (layer0_outputs(9372));
    outputs(9490) <= layer0_outputs(6994);
    outputs(9491) <= layer0_outputs(3659);
    outputs(9492) <= not((layer0_outputs(6887)) and (layer0_outputs(6862)));
    outputs(9493) <= not(layer0_outputs(2347));
    outputs(9494) <= (layer0_outputs(3724)) and not (layer0_outputs(5502));
    outputs(9495) <= not(layer0_outputs(7196)) or (layer0_outputs(8941));
    outputs(9496) <= (layer0_outputs(4487)) xor (layer0_outputs(4821));
    outputs(9497) <= layer0_outputs(2907);
    outputs(9498) <= layer0_outputs(3346);
    outputs(9499) <= not(layer0_outputs(6185));
    outputs(9500) <= (layer0_outputs(386)) xor (layer0_outputs(2578));
    outputs(9501) <= (layer0_outputs(5193)) xor (layer0_outputs(737));
    outputs(9502) <= not((layer0_outputs(5161)) xor (layer0_outputs(632)));
    outputs(9503) <= not((layer0_outputs(9260)) xor (layer0_outputs(5620)));
    outputs(9504) <= not(layer0_outputs(5142)) or (layer0_outputs(6162));
    outputs(9505) <= layer0_outputs(2912);
    outputs(9506) <= (layer0_outputs(2323)) xor (layer0_outputs(8417));
    outputs(9507) <= not(layer0_outputs(1768));
    outputs(9508) <= layer0_outputs(7530);
    outputs(9509) <= layer0_outputs(2086);
    outputs(9510) <= not((layer0_outputs(418)) or (layer0_outputs(1582)));
    outputs(9511) <= not((layer0_outputs(5071)) xor (layer0_outputs(7028)));
    outputs(9512) <= (layer0_outputs(5073)) and (layer0_outputs(567));
    outputs(9513) <= layer0_outputs(9850);
    outputs(9514) <= not(layer0_outputs(2414));
    outputs(9515) <= not(layer0_outputs(8535));
    outputs(9516) <= not((layer0_outputs(6209)) xor (layer0_outputs(8603)));
    outputs(9517) <= layer0_outputs(6772);
    outputs(9518) <= not(layer0_outputs(6439)) or (layer0_outputs(9270));
    outputs(9519) <= not(layer0_outputs(5809));
    outputs(9520) <= layer0_outputs(6015);
    outputs(9521) <= (layer0_outputs(9031)) and (layer0_outputs(4059));
    outputs(9522) <= layer0_outputs(1031);
    outputs(9523) <= not(layer0_outputs(3917));
    outputs(9524) <= layer0_outputs(5038);
    outputs(9525) <= not(layer0_outputs(5750));
    outputs(9526) <= layer0_outputs(7214);
    outputs(9527) <= (layer0_outputs(3932)) xor (layer0_outputs(3618));
    outputs(9528) <= (layer0_outputs(9628)) and not (layer0_outputs(8589));
    outputs(9529) <= not(layer0_outputs(7321));
    outputs(9530) <= not((layer0_outputs(1640)) or (layer0_outputs(1151)));
    outputs(9531) <= layer0_outputs(7850);
    outputs(9532) <= (layer0_outputs(5423)) xor (layer0_outputs(431));
    outputs(9533) <= layer0_outputs(2816);
    outputs(9534) <= not(layer0_outputs(1354));
    outputs(9535) <= layer0_outputs(8362);
    outputs(9536) <= (layer0_outputs(8847)) and (layer0_outputs(1357));
    outputs(9537) <= not(layer0_outputs(4308));
    outputs(9538) <= (layer0_outputs(6867)) and (layer0_outputs(6980));
    outputs(9539) <= layer0_outputs(5961);
    outputs(9540) <= layer0_outputs(5893);
    outputs(9541) <= not(layer0_outputs(8140));
    outputs(9542) <= (layer0_outputs(9588)) and not (layer0_outputs(9091));
    outputs(9543) <= not((layer0_outputs(5046)) xor (layer0_outputs(1370)));
    outputs(9544) <= layer0_outputs(7697);
    outputs(9545) <= not((layer0_outputs(9052)) and (layer0_outputs(2834)));
    outputs(9546) <= not((layer0_outputs(4904)) xor (layer0_outputs(9088)));
    outputs(9547) <= (layer0_outputs(6775)) and not (layer0_outputs(8843));
    outputs(9548) <= (layer0_outputs(8493)) and (layer0_outputs(1976));
    outputs(9549) <= not(layer0_outputs(5239));
    outputs(9550) <= not((layer0_outputs(1659)) or (layer0_outputs(1986)));
    outputs(9551) <= (layer0_outputs(6310)) and not (layer0_outputs(2410));
    outputs(9552) <= layer0_outputs(2259);
    outputs(9553) <= not(layer0_outputs(3329));
    outputs(9554) <= (layer0_outputs(4355)) and (layer0_outputs(9129));
    outputs(9555) <= layer0_outputs(7194);
    outputs(9556) <= not((layer0_outputs(8843)) or (layer0_outputs(2802)));
    outputs(9557) <= (layer0_outputs(9533)) and not (layer0_outputs(4276));
    outputs(9558) <= layer0_outputs(8601);
    outputs(9559) <= layer0_outputs(2247);
    outputs(9560) <= not((layer0_outputs(5079)) xor (layer0_outputs(4055)));
    outputs(9561) <= layer0_outputs(5646);
    outputs(9562) <= (layer0_outputs(3411)) xor (layer0_outputs(7266));
    outputs(9563) <= not((layer0_outputs(5751)) xor (layer0_outputs(8059)));
    outputs(9564) <= layer0_outputs(3635);
    outputs(9565) <= not(layer0_outputs(6678));
    outputs(9566) <= not((layer0_outputs(3931)) xor (layer0_outputs(7158)));
    outputs(9567) <= layer0_outputs(8780);
    outputs(9568) <= (layer0_outputs(4044)) and not (layer0_outputs(1855));
    outputs(9569) <= (layer0_outputs(6631)) and (layer0_outputs(3781));
    outputs(9570) <= not(layer0_outputs(10112));
    outputs(9571) <= not((layer0_outputs(2049)) xor (layer0_outputs(7006)));
    outputs(9572) <= not(layer0_outputs(3704));
    outputs(9573) <= (layer0_outputs(5090)) and not (layer0_outputs(9085));
    outputs(9574) <= (layer0_outputs(3941)) and not (layer0_outputs(352));
    outputs(9575) <= not(layer0_outputs(7679)) or (layer0_outputs(7335));
    outputs(9576) <= layer0_outputs(6255);
    outputs(9577) <= (layer0_outputs(1140)) xor (layer0_outputs(7799));
    outputs(9578) <= (layer0_outputs(122)) xor (layer0_outputs(8294));
    outputs(9579) <= layer0_outputs(5166);
    outputs(9580) <= not((layer0_outputs(4238)) xor (layer0_outputs(7233)));
    outputs(9581) <= (layer0_outputs(1098)) xor (layer0_outputs(3244));
    outputs(9582) <= not(layer0_outputs(5181)) or (layer0_outputs(8287));
    outputs(9583) <= layer0_outputs(8975);
    outputs(9584) <= (layer0_outputs(1513)) and not (layer0_outputs(631));
    outputs(9585) <= layer0_outputs(945);
    outputs(9586) <= (layer0_outputs(3408)) xor (layer0_outputs(4567));
    outputs(9587) <= not((layer0_outputs(8520)) xor (layer0_outputs(5468)));
    outputs(9588) <= not((layer0_outputs(4551)) or (layer0_outputs(789)));
    outputs(9589) <= not(layer0_outputs(5850));
    outputs(9590) <= not(layer0_outputs(2658));
    outputs(9591) <= layer0_outputs(10033);
    outputs(9592) <= layer0_outputs(3341);
    outputs(9593) <= not((layer0_outputs(1262)) and (layer0_outputs(3335)));
    outputs(9594) <= (layer0_outputs(488)) and not (layer0_outputs(9449));
    outputs(9595) <= not(layer0_outputs(412));
    outputs(9596) <= not(layer0_outputs(3435));
    outputs(9597) <= (layer0_outputs(3886)) xor (layer0_outputs(8508));
    outputs(9598) <= (layer0_outputs(5808)) xor (layer0_outputs(1231));
    outputs(9599) <= (layer0_outputs(10006)) or (layer0_outputs(152));
    outputs(9600) <= not(layer0_outputs(1067));
    outputs(9601) <= (layer0_outputs(4093)) and not (layer0_outputs(2501));
    outputs(9602) <= not((layer0_outputs(5819)) xor (layer0_outputs(2762)));
    outputs(9603) <= not(layer0_outputs(3733));
    outputs(9604) <= not((layer0_outputs(9127)) xor (layer0_outputs(5964)));
    outputs(9605) <= not((layer0_outputs(9058)) xor (layer0_outputs(1193)));
    outputs(9606) <= not((layer0_outputs(7691)) xor (layer0_outputs(3640)));
    outputs(9607) <= not(layer0_outputs(8502)) or (layer0_outputs(10132));
    outputs(9608) <= not(layer0_outputs(7869)) or (layer0_outputs(3630));
    outputs(9609) <= not((layer0_outputs(9443)) or (layer0_outputs(1378)));
    outputs(9610) <= (layer0_outputs(5946)) xor (layer0_outputs(992));
    outputs(9611) <= not((layer0_outputs(4884)) and (layer0_outputs(5412)));
    outputs(9612) <= (layer0_outputs(7617)) xor (layer0_outputs(7269));
    outputs(9613) <= not((layer0_outputs(6318)) or (layer0_outputs(4999)));
    outputs(9614) <= not((layer0_outputs(9378)) xor (layer0_outputs(4843)));
    outputs(9615) <= not(layer0_outputs(7492)) or (layer0_outputs(4682));
    outputs(9616) <= (layer0_outputs(8069)) xor (layer0_outputs(61));
    outputs(9617) <= not((layer0_outputs(2178)) and (layer0_outputs(5222)));
    outputs(9618) <= not(layer0_outputs(695));
    outputs(9619) <= not((layer0_outputs(2020)) xor (layer0_outputs(5637)));
    outputs(9620) <= (layer0_outputs(4760)) and not (layer0_outputs(7949));
    outputs(9621) <= layer0_outputs(9632);
    outputs(9622) <= layer0_outputs(9222);
    outputs(9623) <= (layer0_outputs(1822)) xor (layer0_outputs(5569));
    outputs(9624) <= (layer0_outputs(620)) xor (layer0_outputs(2687));
    outputs(9625) <= not((layer0_outputs(1268)) xor (layer0_outputs(9485)));
    outputs(9626) <= (layer0_outputs(2800)) or (layer0_outputs(2568));
    outputs(9627) <= (layer0_outputs(2345)) xor (layer0_outputs(2589));
    outputs(9628) <= not(layer0_outputs(8179));
    outputs(9629) <= not((layer0_outputs(4107)) xor (layer0_outputs(3748)));
    outputs(9630) <= not((layer0_outputs(1435)) xor (layer0_outputs(6124)));
    outputs(9631) <= not((layer0_outputs(8776)) xor (layer0_outputs(2557)));
    outputs(9632) <= layer0_outputs(2245);
    outputs(9633) <= (layer0_outputs(5696)) and not (layer0_outputs(8510));
    outputs(9634) <= (layer0_outputs(5360)) and not (layer0_outputs(4084));
    outputs(9635) <= (layer0_outputs(8116)) xor (layer0_outputs(6800));
    outputs(9636) <= (layer0_outputs(9616)) or (layer0_outputs(4020));
    outputs(9637) <= not((layer0_outputs(5749)) and (layer0_outputs(3698)));
    outputs(9638) <= not((layer0_outputs(4913)) xor (layer0_outputs(624)));
    outputs(9639) <= not(layer0_outputs(6094));
    outputs(9640) <= not(layer0_outputs(5926));
    outputs(9641) <= not(layer0_outputs(9096));
    outputs(9642) <= (layer0_outputs(8160)) and not (layer0_outputs(2301));
    outputs(9643) <= layer0_outputs(5216);
    outputs(9644) <= (layer0_outputs(3711)) and not (layer0_outputs(4798));
    outputs(9645) <= not((layer0_outputs(5876)) xor (layer0_outputs(2958)));
    outputs(9646) <= not(layer0_outputs(4029)) or (layer0_outputs(4449));
    outputs(9647) <= (layer0_outputs(4142)) and not (layer0_outputs(6297));
    outputs(9648) <= layer0_outputs(5755);
    outputs(9649) <= (layer0_outputs(8788)) or (layer0_outputs(8380));
    outputs(9650) <= not((layer0_outputs(580)) xor (layer0_outputs(5226)));
    outputs(9651) <= not(layer0_outputs(1898));
    outputs(9652) <= not(layer0_outputs(9357)) or (layer0_outputs(2599));
    outputs(9653) <= not((layer0_outputs(6681)) or (layer0_outputs(2954)));
    outputs(9654) <= (layer0_outputs(8290)) and not (layer0_outputs(9164));
    outputs(9655) <= layer0_outputs(4457);
    outputs(9656) <= (layer0_outputs(2664)) and not (layer0_outputs(4240));
    outputs(9657) <= not(layer0_outputs(5200));
    outputs(9658) <= (layer0_outputs(53)) and (layer0_outputs(4931));
    outputs(9659) <= not(layer0_outputs(7783));
    outputs(9660) <= not(layer0_outputs(649));
    outputs(9661) <= not(layer0_outputs(9813));
    outputs(9662) <= not((layer0_outputs(6428)) and (layer0_outputs(4865)));
    outputs(9663) <= not(layer0_outputs(125));
    outputs(9664) <= layer0_outputs(5548);
    outputs(9665) <= not((layer0_outputs(8634)) xor (layer0_outputs(6700)));
    outputs(9666) <= not(layer0_outputs(1462));
    outputs(9667) <= not((layer0_outputs(8599)) or (layer0_outputs(6913)));
    outputs(9668) <= (layer0_outputs(2909)) and not (layer0_outputs(8027));
    outputs(9669) <= not((layer0_outputs(10066)) xor (layer0_outputs(4018)));
    outputs(9670) <= not(layer0_outputs(1695));
    outputs(9671) <= not((layer0_outputs(539)) xor (layer0_outputs(5579)));
    outputs(9672) <= not(layer0_outputs(3486));
    outputs(9673) <= not((layer0_outputs(7253)) or (layer0_outputs(8099)));
    outputs(9674) <= not((layer0_outputs(6139)) or (layer0_outputs(2554)));
    outputs(9675) <= not((layer0_outputs(2772)) xor (layer0_outputs(9569)));
    outputs(9676) <= (layer0_outputs(5093)) and (layer0_outputs(5903));
    outputs(9677) <= not(layer0_outputs(9548));
    outputs(9678) <= layer0_outputs(5981);
    outputs(9679) <= (layer0_outputs(7779)) and not (layer0_outputs(8343));
    outputs(9680) <= not((layer0_outputs(8329)) xor (layer0_outputs(7617)));
    outputs(9681) <= (layer0_outputs(5689)) and not (layer0_outputs(3501));
    outputs(9682) <= not(layer0_outputs(5886));
    outputs(9683) <= not((layer0_outputs(7321)) or (layer0_outputs(6967)));
    outputs(9684) <= layer0_outputs(9138);
    outputs(9685) <= not((layer0_outputs(9502)) and (layer0_outputs(5658)));
    outputs(9686) <= not(layer0_outputs(99));
    outputs(9687) <= not(layer0_outputs(9307));
    outputs(9688) <= layer0_outputs(10218);
    outputs(9689) <= layer0_outputs(4937);
    outputs(9690) <= not(layer0_outputs(3395));
    outputs(9691) <= (layer0_outputs(9457)) xor (layer0_outputs(18));
    outputs(9692) <= not(layer0_outputs(2717));
    outputs(9693) <= layer0_outputs(7231);
    outputs(9694) <= not(layer0_outputs(5068));
    outputs(9695) <= (layer0_outputs(9195)) and not (layer0_outputs(4694));
    outputs(9696) <= (layer0_outputs(8162)) and not (layer0_outputs(3526));
    outputs(9697) <= not((layer0_outputs(433)) xor (layer0_outputs(4304)));
    outputs(9698) <= layer0_outputs(9186);
    outputs(9699) <= not(layer0_outputs(8356));
    outputs(9700) <= not(layer0_outputs(6360));
    outputs(9701) <= not((layer0_outputs(4834)) or (layer0_outputs(2514)));
    outputs(9702) <= not((layer0_outputs(290)) xor (layer0_outputs(429)));
    outputs(9703) <= layer0_outputs(9817);
    outputs(9704) <= not((layer0_outputs(7989)) xor (layer0_outputs(2804)));
    outputs(9705) <= not(layer0_outputs(8192));
    outputs(9706) <= not((layer0_outputs(4568)) and (layer0_outputs(6356)));
    outputs(9707) <= (layer0_outputs(8075)) and not (layer0_outputs(6843));
    outputs(9708) <= layer0_outputs(7420);
    outputs(9709) <= (layer0_outputs(5523)) and not (layer0_outputs(3610));
    outputs(9710) <= layer0_outputs(9447);
    outputs(9711) <= not((layer0_outputs(3197)) xor (layer0_outputs(2720)));
    outputs(9712) <= (layer0_outputs(9456)) or (layer0_outputs(6309));
    outputs(9713) <= not(layer0_outputs(6803));
    outputs(9714) <= not((layer0_outputs(8311)) xor (layer0_outputs(8106)));
    outputs(9715) <= not(layer0_outputs(6617));
    outputs(9716) <= not(layer0_outputs(3571));
    outputs(9717) <= (layer0_outputs(6378)) xor (layer0_outputs(5904));
    outputs(9718) <= not(layer0_outputs(4495)) or (layer0_outputs(6760));
    outputs(9719) <= (layer0_outputs(9553)) and not (layer0_outputs(7065));
    outputs(9720) <= layer0_outputs(4457);
    outputs(9721) <= layer0_outputs(1064);
    outputs(9722) <= (layer0_outputs(779)) xor (layer0_outputs(5878));
    outputs(9723) <= layer0_outputs(7902);
    outputs(9724) <= (layer0_outputs(10124)) xor (layer0_outputs(3141));
    outputs(9725) <= layer0_outputs(8096);
    outputs(9726) <= not(layer0_outputs(2936));
    outputs(9727) <= layer0_outputs(464);
    outputs(9728) <= layer0_outputs(1229);
    outputs(9729) <= (layer0_outputs(9420)) xor (layer0_outputs(816));
    outputs(9730) <= not(layer0_outputs(9718));
    outputs(9731) <= (layer0_outputs(724)) and not (layer0_outputs(2194));
    outputs(9732) <= (layer0_outputs(3811)) and not (layer0_outputs(4942));
    outputs(9733) <= not(layer0_outputs(26)) or (layer0_outputs(7184));
    outputs(9734) <= layer0_outputs(9532);
    outputs(9735) <= (layer0_outputs(3419)) xor (layer0_outputs(2871));
    outputs(9736) <= (layer0_outputs(8623)) xor (layer0_outputs(2103));
    outputs(9737) <= layer0_outputs(5483);
    outputs(9738) <= not((layer0_outputs(8106)) xor (layer0_outputs(8703)));
    outputs(9739) <= layer0_outputs(2537);
    outputs(9740) <= (layer0_outputs(8244)) xor (layer0_outputs(2890));
    outputs(9741) <= layer0_outputs(6734);
    outputs(9742) <= (layer0_outputs(2091)) and not (layer0_outputs(541));
    outputs(9743) <= layer0_outputs(150);
    outputs(9744) <= (layer0_outputs(4414)) and not (layer0_outputs(3737));
    outputs(9745) <= not(layer0_outputs(4420));
    outputs(9746) <= (layer0_outputs(7277)) and (layer0_outputs(7207));
    outputs(9747) <= not(layer0_outputs(9664));
    outputs(9748) <= (layer0_outputs(1699)) xor (layer0_outputs(4362));
    outputs(9749) <= (layer0_outputs(1496)) xor (layer0_outputs(9569));
    outputs(9750) <= not((layer0_outputs(2344)) xor (layer0_outputs(1204)));
    outputs(9751) <= not(layer0_outputs(1946));
    outputs(9752) <= (layer0_outputs(7364)) and (layer0_outputs(6925));
    outputs(9753) <= (layer0_outputs(9441)) xor (layer0_outputs(2634));
    outputs(9754) <= (layer0_outputs(3665)) and (layer0_outputs(6322));
    outputs(9755) <= not(layer0_outputs(8614));
    outputs(9756) <= layer0_outputs(7371);
    outputs(9757) <= (layer0_outputs(10171)) and not (layer0_outputs(5677));
    outputs(9758) <= layer0_outputs(1091);
    outputs(9759) <= not(layer0_outputs(1643));
    outputs(9760) <= not(layer0_outputs(3115));
    outputs(9761) <= layer0_outputs(1574);
    outputs(9762) <= (layer0_outputs(6103)) xor (layer0_outputs(8150));
    outputs(9763) <= not(layer0_outputs(2565));
    outputs(9764) <= (layer0_outputs(4759)) and not (layer0_outputs(6875));
    outputs(9765) <= not(layer0_outputs(4140));
    outputs(9766) <= not(layer0_outputs(9944));
    outputs(9767) <= not(layer0_outputs(6007));
    outputs(9768) <= layer0_outputs(100);
    outputs(9769) <= layer0_outputs(6229);
    outputs(9770) <= not(layer0_outputs(7621));
    outputs(9771) <= (layer0_outputs(7355)) and (layer0_outputs(8764));
    outputs(9772) <= (layer0_outputs(5460)) xor (layer0_outputs(9102));
    outputs(9773) <= layer0_outputs(6629);
    outputs(9774) <= not(layer0_outputs(5918));
    outputs(9775) <= layer0_outputs(7646);
    outputs(9776) <= layer0_outputs(10017);
    outputs(9777) <= not(layer0_outputs(5480));
    outputs(9778) <= (layer0_outputs(8364)) xor (layer0_outputs(8354));
    outputs(9779) <= not(layer0_outputs(6394));
    outputs(9780) <= layer0_outputs(5328);
    outputs(9781) <= not((layer0_outputs(3090)) or (layer0_outputs(2706)));
    outputs(9782) <= not((layer0_outputs(7156)) or (layer0_outputs(1793)));
    outputs(9783) <= not(layer0_outputs(5800)) or (layer0_outputs(4130));
    outputs(9784) <= (layer0_outputs(8436)) xor (layer0_outputs(4431));
    outputs(9785) <= (layer0_outputs(136)) xor (layer0_outputs(8327));
    outputs(9786) <= not((layer0_outputs(1920)) or (layer0_outputs(8020)));
    outputs(9787) <= not((layer0_outputs(9137)) xor (layer0_outputs(4247)));
    outputs(9788) <= not(layer0_outputs(3617)) or (layer0_outputs(4629));
    outputs(9789) <= not(layer0_outputs(2177));
    outputs(9790) <= not(layer0_outputs(5131));
    outputs(9791) <= (layer0_outputs(9976)) and not (layer0_outputs(6384));
    outputs(9792) <= (layer0_outputs(3551)) and (layer0_outputs(3159));
    outputs(9793) <= layer0_outputs(7017);
    outputs(9794) <= (layer0_outputs(4825)) xor (layer0_outputs(647));
    outputs(9795) <= not((layer0_outputs(1649)) xor (layer0_outputs(6376)));
    outputs(9796) <= (layer0_outputs(10158)) xor (layer0_outputs(8207));
    outputs(9797) <= not((layer0_outputs(1834)) xor (layer0_outputs(3828)));
    outputs(9798) <= (layer0_outputs(1046)) and not (layer0_outputs(2320));
    outputs(9799) <= not((layer0_outputs(1381)) xor (layer0_outputs(3784)));
    outputs(9800) <= (layer0_outputs(9269)) and not (layer0_outputs(6009));
    outputs(9801) <= layer0_outputs(7890);
    outputs(9802) <= not((layer0_outputs(2056)) xor (layer0_outputs(9367)));
    outputs(9803) <= (layer0_outputs(3417)) and not (layer0_outputs(5590));
    outputs(9804) <= not((layer0_outputs(3612)) xor (layer0_outputs(6441)));
    outputs(9805) <= (layer0_outputs(7118)) and (layer0_outputs(7889));
    outputs(9806) <= layer0_outputs(7695);
    outputs(9807) <= not(layer0_outputs(3275));
    outputs(9808) <= (layer0_outputs(2370)) and not (layer0_outputs(8638));
    outputs(9809) <= (layer0_outputs(7042)) xor (layer0_outputs(6811));
    outputs(9810) <= not((layer0_outputs(2712)) xor (layer0_outputs(6693)));
    outputs(9811) <= not(layer0_outputs(10014));
    outputs(9812) <= not(layer0_outputs(9448));
    outputs(9813) <= layer0_outputs(759);
    outputs(9814) <= layer0_outputs(640);
    outputs(9815) <= not((layer0_outputs(9082)) or (layer0_outputs(2761)));
    outputs(9816) <= not(layer0_outputs(69)) or (layer0_outputs(4704));
    outputs(9817) <= layer0_outputs(7877);
    outputs(9818) <= (layer0_outputs(8267)) or (layer0_outputs(6991));
    outputs(9819) <= not((layer0_outputs(2065)) xor (layer0_outputs(1739)));
    outputs(9820) <= not((layer0_outputs(6555)) xor (layer0_outputs(5518)));
    outputs(9821) <= (layer0_outputs(6065)) and not (layer0_outputs(893));
    outputs(9822) <= not(layer0_outputs(3839));
    outputs(9823) <= layer0_outputs(8465);
    outputs(9824) <= (layer0_outputs(2522)) and not (layer0_outputs(4858));
    outputs(9825) <= not((layer0_outputs(2562)) or (layer0_outputs(1860)));
    outputs(9826) <= not(layer0_outputs(8687));
    outputs(9827) <= layer0_outputs(7247);
    outputs(9828) <= not(layer0_outputs(9586));
    outputs(9829) <= not((layer0_outputs(9149)) xor (layer0_outputs(8875)));
    outputs(9830) <= not(layer0_outputs(7648));
    outputs(9831) <= not(layer0_outputs(5938));
    outputs(9832) <= layer0_outputs(6446);
    outputs(9833) <= (layer0_outputs(6126)) and not (layer0_outputs(5050));
    outputs(9834) <= layer0_outputs(8512);
    outputs(9835) <= not(layer0_outputs(10219));
    outputs(9836) <= not((layer0_outputs(7206)) or (layer0_outputs(4824)));
    outputs(9837) <= (layer0_outputs(409)) xor (layer0_outputs(4731));
    outputs(9838) <= layer0_outputs(1187);
    outputs(9839) <= layer0_outputs(7278);
    outputs(9840) <= not(layer0_outputs(5371));
    outputs(9841) <= (layer0_outputs(4417)) xor (layer0_outputs(1368));
    outputs(9842) <= not((layer0_outputs(6261)) xor (layer0_outputs(980)));
    outputs(9843) <= not(layer0_outputs(1153));
    outputs(9844) <= layer0_outputs(5596);
    outputs(9845) <= (layer0_outputs(1345)) and (layer0_outputs(3808));
    outputs(9846) <= (layer0_outputs(6890)) xor (layer0_outputs(3931));
    outputs(9847) <= not((layer0_outputs(9301)) xor (layer0_outputs(2931)));
    outputs(9848) <= not(layer0_outputs(4732));
    outputs(9849) <= layer0_outputs(2828);
    outputs(9850) <= not((layer0_outputs(5500)) xor (layer0_outputs(2846)));
    outputs(9851) <= (layer0_outputs(6358)) xor (layer0_outputs(7810));
    outputs(9852) <= (layer0_outputs(6148)) and (layer0_outputs(852));
    outputs(9853) <= layer0_outputs(5209);
    outputs(9854) <= (layer0_outputs(4056)) and not (layer0_outputs(5741));
    outputs(9855) <= not(layer0_outputs(2833)) or (layer0_outputs(8850));
    outputs(9856) <= not(layer0_outputs(2854));
    outputs(9857) <= not(layer0_outputs(3298));
    outputs(9858) <= (layer0_outputs(1347)) and not (layer0_outputs(2610));
    outputs(9859) <= (layer0_outputs(4318)) and not (layer0_outputs(7154));
    outputs(9860) <= not((layer0_outputs(1294)) xor (layer0_outputs(6218)));
    outputs(9861) <= not(layer0_outputs(913));
    outputs(9862) <= not(layer0_outputs(6305));
    outputs(9863) <= not(layer0_outputs(2008));
    outputs(9864) <= not((layer0_outputs(1430)) or (layer0_outputs(6765)));
    outputs(9865) <= layer0_outputs(549);
    outputs(9866) <= layer0_outputs(1120);
    outputs(9867) <= not((layer0_outputs(886)) xor (layer0_outputs(5031)));
    outputs(9868) <= not(layer0_outputs(7829));
    outputs(9869) <= (layer0_outputs(4941)) and not (layer0_outputs(2389));
    outputs(9870) <= not(layer0_outputs(8653));
    outputs(9871) <= not((layer0_outputs(7571)) xor (layer0_outputs(4312)));
    outputs(9872) <= (layer0_outputs(5727)) xor (layer0_outputs(8739));
    outputs(9873) <= (layer0_outputs(551)) xor (layer0_outputs(6033));
    outputs(9874) <= layer0_outputs(1494);
    outputs(9875) <= not(layer0_outputs(3952));
    outputs(9876) <= layer0_outputs(3215);
    outputs(9877) <= not(layer0_outputs(1662));
    outputs(9878) <= not(layer0_outputs(9937));
    outputs(9879) <= (layer0_outputs(8406)) and not (layer0_outputs(6300));
    outputs(9880) <= not(layer0_outputs(2210));
    outputs(9881) <= (layer0_outputs(5318)) xor (layer0_outputs(1432));
    outputs(9882) <= (layer0_outputs(5651)) and (layer0_outputs(5174));
    outputs(9883) <= (layer0_outputs(5730)) xor (layer0_outputs(5008));
    outputs(9884) <= layer0_outputs(4645);
    outputs(9885) <= not(layer0_outputs(7036)) or (layer0_outputs(7226));
    outputs(9886) <= not(layer0_outputs(3914));
    outputs(9887) <= (layer0_outputs(6844)) xor (layer0_outputs(9884));
    outputs(9888) <= (layer0_outputs(2548)) and not (layer0_outputs(1719));
    outputs(9889) <= layer0_outputs(441);
    outputs(9890) <= not(layer0_outputs(1713));
    outputs(9891) <= not((layer0_outputs(2820)) xor (layer0_outputs(917)));
    outputs(9892) <= not(layer0_outputs(6380)) or (layer0_outputs(8269));
    outputs(9893) <= not(layer0_outputs(70));
    outputs(9894) <= not(layer0_outputs(3110));
    outputs(9895) <= (layer0_outputs(345)) xor (layer0_outputs(7143));
    outputs(9896) <= not((layer0_outputs(2696)) xor (layer0_outputs(817)));
    outputs(9897) <= not((layer0_outputs(1042)) xor (layer0_outputs(3991)));
    outputs(9898) <= layer0_outputs(9989);
    outputs(9899) <= not((layer0_outputs(1988)) xor (layer0_outputs(8577)));
    outputs(9900) <= not(layer0_outputs(2406));
    outputs(9901) <= layer0_outputs(408);
    outputs(9902) <= layer0_outputs(7727);
    outputs(9903) <= (layer0_outputs(4186)) xor (layer0_outputs(1002));
    outputs(9904) <= not((layer0_outputs(745)) or (layer0_outputs(3249)));
    outputs(9905) <= not(layer0_outputs(8123));
    outputs(9906) <= (layer0_outputs(1393)) xor (layer0_outputs(3888));
    outputs(9907) <= not((layer0_outputs(4936)) or (layer0_outputs(1300)));
    outputs(9908) <= layer0_outputs(1720);
    outputs(9909) <= layer0_outputs(1004);
    outputs(9910) <= not(layer0_outputs(2110));
    outputs(9911) <= (layer0_outputs(5983)) and not (layer0_outputs(9167));
    outputs(9912) <= not(layer0_outputs(7555));
    outputs(9913) <= not((layer0_outputs(1561)) and (layer0_outputs(4605)));
    outputs(9914) <= not(layer0_outputs(1175));
    outputs(9915) <= not(layer0_outputs(7451));
    outputs(9916) <= not(layer0_outputs(2736)) or (layer0_outputs(3251));
    outputs(9917) <= (layer0_outputs(9006)) or (layer0_outputs(1185));
    outputs(9918) <= (layer0_outputs(3714)) and not (layer0_outputs(6054));
    outputs(9919) <= not((layer0_outputs(3511)) xor (layer0_outputs(5847)));
    outputs(9920) <= layer0_outputs(2416);
    outputs(9921) <= not(layer0_outputs(3885));
    outputs(9922) <= not(layer0_outputs(1342));
    outputs(9923) <= not(layer0_outputs(6654));
    outputs(9924) <= not((layer0_outputs(445)) xor (layer0_outputs(1424)));
    outputs(9925) <= (layer0_outputs(9068)) and (layer0_outputs(7213));
    outputs(9926) <= not(layer0_outputs(2191));
    outputs(9927) <= layer0_outputs(486);
    outputs(9928) <= layer0_outputs(5085);
    outputs(9929) <= (layer0_outputs(2891)) xor (layer0_outputs(6106));
    outputs(9930) <= layer0_outputs(5275);
    outputs(9931) <= not(layer0_outputs(3006));
    outputs(9932) <= layer0_outputs(1592);
    outputs(9933) <= (layer0_outputs(9570)) xor (layer0_outputs(3600));
    outputs(9934) <= not(layer0_outputs(368));
    outputs(9935) <= not((layer0_outputs(7230)) xor (layer0_outputs(10123)));
    outputs(9936) <= not(layer0_outputs(6810)) or (layer0_outputs(1805));
    outputs(9937) <= layer0_outputs(3899);
    outputs(9938) <= not(layer0_outputs(9022));
    outputs(9939) <= (layer0_outputs(6864)) xor (layer0_outputs(2127));
    outputs(9940) <= (layer0_outputs(6463)) xor (layer0_outputs(917));
    outputs(9941) <= (layer0_outputs(3041)) and not (layer0_outputs(9423));
    outputs(9942) <= not(layer0_outputs(7302));
    outputs(9943) <= (layer0_outputs(5138)) and (layer0_outputs(985));
    outputs(9944) <= layer0_outputs(6759);
    outputs(9945) <= not(layer0_outputs(1000));
    outputs(9946) <= (layer0_outputs(2516)) xor (layer0_outputs(8969));
    outputs(9947) <= (layer0_outputs(4455)) xor (layer0_outputs(9358));
    outputs(9948) <= (layer0_outputs(8400)) and not (layer0_outputs(8944));
    outputs(9949) <= layer0_outputs(2066);
    outputs(9950) <= layer0_outputs(103);
    outputs(9951) <= not(layer0_outputs(1644));
    outputs(9952) <= (layer0_outputs(7572)) and not (layer0_outputs(7458));
    outputs(9953) <= (layer0_outputs(8771)) and not (layer0_outputs(1163));
    outputs(9954) <= not(layer0_outputs(4475));
    outputs(9955) <= (layer0_outputs(5409)) and (layer0_outputs(10223));
    outputs(9956) <= not((layer0_outputs(179)) or (layer0_outputs(539)));
    outputs(9957) <= not(layer0_outputs(672));
    outputs(9958) <= not((layer0_outputs(10140)) and (layer0_outputs(9869)));
    outputs(9959) <= not(layer0_outputs(4659));
    outputs(9960) <= not(layer0_outputs(7365));
    outputs(9961) <= (layer0_outputs(9978)) xor (layer0_outputs(4900));
    outputs(9962) <= not(layer0_outputs(744));
    outputs(9963) <= not((layer0_outputs(1452)) xor (layer0_outputs(6434)));
    outputs(9964) <= (layer0_outputs(1045)) xor (layer0_outputs(7338));
    outputs(9965) <= not(layer0_outputs(2437));
    outputs(9966) <= layer0_outputs(8096);
    outputs(9967) <= layer0_outputs(4700);
    outputs(9968) <= not((layer0_outputs(6798)) xor (layer0_outputs(389)));
    outputs(9969) <= not((layer0_outputs(2987)) xor (layer0_outputs(6255)));
    outputs(9970) <= not(layer0_outputs(5972)) or (layer0_outputs(4061));
    outputs(9971) <= not(layer0_outputs(9153)) or (layer0_outputs(3362));
    outputs(9972) <= (layer0_outputs(5444)) and not (layer0_outputs(1050));
    outputs(9973) <= not((layer0_outputs(2807)) or (layer0_outputs(6005)));
    outputs(9974) <= not(layer0_outputs(3287));
    outputs(9975) <= layer0_outputs(6402);
    outputs(9976) <= not(layer0_outputs(4954));
    outputs(9977) <= not((layer0_outputs(4601)) or (layer0_outputs(10115)));
    outputs(9978) <= not(layer0_outputs(2691));
    outputs(9979) <= layer0_outputs(8973);
    outputs(9980) <= (layer0_outputs(3987)) and not (layer0_outputs(3935));
    outputs(9981) <= layer0_outputs(3475);
    outputs(9982) <= layer0_outputs(7568);
    outputs(9983) <= not((layer0_outputs(9567)) xor (layer0_outputs(3895)));
    outputs(9984) <= (layer0_outputs(5223)) xor (layer0_outputs(1097));
    outputs(9985) <= not(layer0_outputs(2649));
    outputs(9986) <= not(layer0_outputs(3908));
    outputs(9987) <= not(layer0_outputs(8405));
    outputs(9988) <= (layer0_outputs(4600)) and not (layer0_outputs(10229));
    outputs(9989) <= not(layer0_outputs(4865));
    outputs(9990) <= (layer0_outputs(8153)) and (layer0_outputs(6001));
    outputs(9991) <= (layer0_outputs(3029)) or (layer0_outputs(2307));
    outputs(9992) <= layer0_outputs(82);
    outputs(9993) <= (layer0_outputs(9160)) xor (layer0_outputs(7631));
    outputs(9994) <= not((layer0_outputs(3881)) xor (layer0_outputs(8184)));
    outputs(9995) <= (layer0_outputs(655)) or (layer0_outputs(5553));
    outputs(9996) <= (layer0_outputs(1771)) and (layer0_outputs(5511));
    outputs(9997) <= not((layer0_outputs(1764)) xor (layer0_outputs(4634)));
    outputs(9998) <= not(layer0_outputs(7743));
    outputs(9999) <= not(layer0_outputs(8103));
    outputs(10000) <= not(layer0_outputs(3499));
    outputs(10001) <= (layer0_outputs(5525)) and not (layer0_outputs(5291));
    outputs(10002) <= not((layer0_outputs(5341)) and (layer0_outputs(545)));
    outputs(10003) <= not((layer0_outputs(8761)) xor (layer0_outputs(8541)));
    outputs(10004) <= not(layer0_outputs(3914));
    outputs(10005) <= (layer0_outputs(6747)) and not (layer0_outputs(4702));
    outputs(10006) <= not((layer0_outputs(5909)) or (layer0_outputs(6204)));
    outputs(10007) <= layer0_outputs(555);
    outputs(10008) <= not((layer0_outputs(4340)) xor (layer0_outputs(3457)));
    outputs(10009) <= not(layer0_outputs(7556));
    outputs(10010) <= layer0_outputs(385);
    outputs(10011) <= not(layer0_outputs(574));
    outputs(10012) <= layer0_outputs(2343);
    outputs(10013) <= (layer0_outputs(6721)) xor (layer0_outputs(8857));
    outputs(10014) <= not((layer0_outputs(8655)) or (layer0_outputs(5628)));
    outputs(10015) <= (layer0_outputs(8131)) xor (layer0_outputs(3854));
    outputs(10016) <= not((layer0_outputs(9658)) xor (layer0_outputs(3351)));
    outputs(10017) <= not(layer0_outputs(9238));
    outputs(10018) <= not(layer0_outputs(499));
    outputs(10019) <= (layer0_outputs(9232)) and not (layer0_outputs(6685));
    outputs(10020) <= (layer0_outputs(4221)) and not (layer0_outputs(5835));
    outputs(10021) <= not((layer0_outputs(10022)) or (layer0_outputs(7004)));
    outputs(10022) <= not((layer0_outputs(6234)) xor (layer0_outputs(8021)));
    outputs(10023) <= not((layer0_outputs(2134)) or (layer0_outputs(5924)));
    outputs(10024) <= layer0_outputs(6998);
    outputs(10025) <= (layer0_outputs(2424)) and (layer0_outputs(8456));
    outputs(10026) <= not(layer0_outputs(5363));
    outputs(10027) <= (layer0_outputs(2713)) xor (layer0_outputs(5649));
    outputs(10028) <= not(layer0_outputs(7943));
    outputs(10029) <= not((layer0_outputs(829)) xor (layer0_outputs(6391)));
    outputs(10030) <= layer0_outputs(2108);
    outputs(10031) <= (layer0_outputs(4775)) and not (layer0_outputs(9833));
    outputs(10032) <= (layer0_outputs(7907)) xor (layer0_outputs(461));
    outputs(10033) <= not((layer0_outputs(4777)) xor (layer0_outputs(9446)));
    outputs(10034) <= layer0_outputs(3188);
    outputs(10035) <= not(layer0_outputs(8302));
    outputs(10036) <= (layer0_outputs(7867)) xor (layer0_outputs(4428));
    outputs(10037) <= (layer0_outputs(5607)) and not (layer0_outputs(919));
    outputs(10038) <= (layer0_outputs(5469)) and not (layer0_outputs(9870));
    outputs(10039) <= not(layer0_outputs(5527));
    outputs(10040) <= layer0_outputs(3221);
    outputs(10041) <= (layer0_outputs(9760)) or (layer0_outputs(10062));
    outputs(10042) <= (layer0_outputs(6559)) and not (layer0_outputs(6429));
    outputs(10043) <= (layer0_outputs(7212)) and not (layer0_outputs(1999));
    outputs(10044) <= not((layer0_outputs(7801)) xor (layer0_outputs(7524)));
    outputs(10045) <= layer0_outputs(5154);
    outputs(10046) <= not(layer0_outputs(3952));
    outputs(10047) <= not(layer0_outputs(8706));
    outputs(10048) <= (layer0_outputs(4285)) xor (layer0_outputs(1059));
    outputs(10049) <= not(layer0_outputs(8143)) or (layer0_outputs(4186));
    outputs(10050) <= (layer0_outputs(9247)) and (layer0_outputs(10092));
    outputs(10051) <= not((layer0_outputs(7843)) xor (layer0_outputs(8856)));
    outputs(10052) <= (layer0_outputs(8206)) xor (layer0_outputs(9577));
    outputs(10053) <= not((layer0_outputs(9623)) xor (layer0_outputs(5033)));
    outputs(10054) <= not((layer0_outputs(738)) xor (layer0_outputs(4721)));
    outputs(10055) <= not(layer0_outputs(6035)) or (layer0_outputs(8742));
    outputs(10056) <= not(layer0_outputs(9176));
    outputs(10057) <= (layer0_outputs(2387)) and not (layer0_outputs(3879));
    outputs(10058) <= not((layer0_outputs(7057)) xor (layer0_outputs(5846)));
    outputs(10059) <= (layer0_outputs(7670)) xor (layer0_outputs(10057));
    outputs(10060) <= (layer0_outputs(5415)) xor (layer0_outputs(9527));
    outputs(10061) <= (layer0_outputs(3396)) xor (layer0_outputs(4819));
    outputs(10062) <= not(layer0_outputs(4217));
    outputs(10063) <= layer0_outputs(107);
    outputs(10064) <= not(layer0_outputs(5936));
    outputs(10065) <= not(layer0_outputs(1130));
    outputs(10066) <= (layer0_outputs(2718)) xor (layer0_outputs(9889));
    outputs(10067) <= not((layer0_outputs(9861)) or (layer0_outputs(2697)));
    outputs(10068) <= not((layer0_outputs(6175)) and (layer0_outputs(2963)));
    outputs(10069) <= (layer0_outputs(7768)) and not (layer0_outputs(4434));
    outputs(10070) <= not(layer0_outputs(2591));
    outputs(10071) <= not((layer0_outputs(9718)) or (layer0_outputs(552)));
    outputs(10072) <= (layer0_outputs(8909)) and not (layer0_outputs(6272));
    outputs(10073) <= not(layer0_outputs(4452));
    outputs(10074) <= (layer0_outputs(2522)) and (layer0_outputs(3137));
    outputs(10075) <= (layer0_outputs(9343)) and not (layer0_outputs(5259));
    outputs(10076) <= not((layer0_outputs(6408)) or (layer0_outputs(1812)));
    outputs(10077) <= layer0_outputs(779);
    outputs(10078) <= layer0_outputs(4394);
    outputs(10079) <= (layer0_outputs(6244)) and (layer0_outputs(3855));
    outputs(10080) <= (layer0_outputs(1282)) xor (layer0_outputs(4988));
    outputs(10081) <= not((layer0_outputs(3364)) xor (layer0_outputs(3697)));
    outputs(10082) <= not((layer0_outputs(3040)) xor (layer0_outputs(4547)));
    outputs(10083) <= not(layer0_outputs(6895));
    outputs(10084) <= not((layer0_outputs(3549)) or (layer0_outputs(7962)));
    outputs(10085) <= (layer0_outputs(4642)) and not (layer0_outputs(9061));
    outputs(10086) <= layer0_outputs(189);
    outputs(10087) <= (layer0_outputs(4164)) or (layer0_outputs(2282));
    outputs(10088) <= (layer0_outputs(6493)) xor (layer0_outputs(6121));
    outputs(10089) <= not(layer0_outputs(7558));
    outputs(10090) <= (layer0_outputs(8518)) and not (layer0_outputs(99));
    outputs(10091) <= (layer0_outputs(3172)) xor (layer0_outputs(6999));
    outputs(10092) <= not((layer0_outputs(3045)) xor (layer0_outputs(3316)));
    outputs(10093) <= not(layer0_outputs(5419));
    outputs(10094) <= (layer0_outputs(6244)) and not (layer0_outputs(8466));
    outputs(10095) <= not((layer0_outputs(10199)) xor (layer0_outputs(2121)));
    outputs(10096) <= layer0_outputs(1597);
    outputs(10097) <= not((layer0_outputs(6644)) xor (layer0_outputs(5714)));
    outputs(10098) <= (layer0_outputs(8334)) and not (layer0_outputs(5132));
    outputs(10099) <= not(layer0_outputs(9244));
    outputs(10100) <= not(layer0_outputs(3113));
    outputs(10101) <= not((layer0_outputs(6419)) xor (layer0_outputs(5020)));
    outputs(10102) <= (layer0_outputs(1273)) and not (layer0_outputs(3886));
    outputs(10103) <= (layer0_outputs(5644)) and not (layer0_outputs(3367));
    outputs(10104) <= not(layer0_outputs(3306));
    outputs(10105) <= (layer0_outputs(8731)) xor (layer0_outputs(3107));
    outputs(10106) <= not(layer0_outputs(2286));
    outputs(10107) <= (layer0_outputs(1024)) xor (layer0_outputs(7314));
    outputs(10108) <= layer0_outputs(5442);
    outputs(10109) <= (layer0_outputs(6638)) xor (layer0_outputs(4459));
    outputs(10110) <= layer0_outputs(3086);
    outputs(10111) <= not(layer0_outputs(7923)) or (layer0_outputs(448));
    outputs(10112) <= not((layer0_outputs(1526)) xor (layer0_outputs(9308)));
    outputs(10113) <= (layer0_outputs(6135)) and not (layer0_outputs(8033));
    outputs(10114) <= (layer0_outputs(3057)) and (layer0_outputs(9057));
    outputs(10115) <= (layer0_outputs(703)) and not (layer0_outputs(3756));
    outputs(10116) <= not(layer0_outputs(915));
    outputs(10117) <= not(layer0_outputs(4638));
    outputs(10118) <= (layer0_outputs(840)) xor (layer0_outputs(8028));
    outputs(10119) <= not(layer0_outputs(7931));
    outputs(10120) <= not((layer0_outputs(4384)) or (layer0_outputs(2794)));
    outputs(10121) <= not(layer0_outputs(1838));
    outputs(10122) <= not((layer0_outputs(9167)) or (layer0_outputs(3323)));
    outputs(10123) <= (layer0_outputs(9915)) and not (layer0_outputs(5139));
    outputs(10124) <= not((layer0_outputs(3248)) or (layer0_outputs(1857)));
    outputs(10125) <= (layer0_outputs(5525)) xor (layer0_outputs(4138));
    outputs(10126) <= layer0_outputs(5589);
    outputs(10127) <= not(layer0_outputs(7682));
    outputs(10128) <= not(layer0_outputs(8899));
    outputs(10129) <= layer0_outputs(8847);
    outputs(10130) <= not(layer0_outputs(9338));
    outputs(10131) <= not(layer0_outputs(9356));
    outputs(10132) <= layer0_outputs(5041);
    outputs(10133) <= layer0_outputs(8872);
    outputs(10134) <= not(layer0_outputs(4241)) or (layer0_outputs(674));
    outputs(10135) <= not((layer0_outputs(5211)) xor (layer0_outputs(5081)));
    outputs(10136) <= not(layer0_outputs(8766)) or (layer0_outputs(8035));
    outputs(10137) <= (layer0_outputs(4260)) and (layer0_outputs(3151));
    outputs(10138) <= layer0_outputs(7910);
    outputs(10139) <= layer0_outputs(2275);
    outputs(10140) <= (layer0_outputs(6052)) and not (layer0_outputs(7342));
    outputs(10141) <= not((layer0_outputs(982)) xor (layer0_outputs(6522)));
    outputs(10142) <= (layer0_outputs(9275)) xor (layer0_outputs(6926));
    outputs(10143) <= not((layer0_outputs(4452)) or (layer0_outputs(6882)));
    outputs(10144) <= not(layer0_outputs(9334));
    outputs(10145) <= not((layer0_outputs(7012)) xor (layer0_outputs(4915)));
    outputs(10146) <= (layer0_outputs(2498)) and (layer0_outputs(9081));
    outputs(10147) <= layer0_outputs(8149);
    outputs(10148) <= (layer0_outputs(9846)) and not (layer0_outputs(754));
    outputs(10149) <= not((layer0_outputs(9801)) or (layer0_outputs(4756)));
    outputs(10150) <= not(layer0_outputs(8804)) or (layer0_outputs(3375));
    outputs(10151) <= not((layer0_outputs(6043)) xor (layer0_outputs(1256)));
    outputs(10152) <= not(layer0_outputs(5217));
    outputs(10153) <= not((layer0_outputs(6062)) or (layer0_outputs(9510)));
    outputs(10154) <= not(layer0_outputs(9952)) or (layer0_outputs(4639));
    outputs(10155) <= layer0_outputs(3289);
    outputs(10156) <= not((layer0_outputs(2509)) xor (layer0_outputs(1290)));
    outputs(10157) <= (layer0_outputs(7054)) and not (layer0_outputs(8697));
    outputs(10158) <= layer0_outputs(7708);
    outputs(10159) <= not((layer0_outputs(3368)) xor (layer0_outputs(8326)));
    outputs(10160) <= not(layer0_outputs(7693));
    outputs(10161) <= (layer0_outputs(6853)) and not (layer0_outputs(5934));
    outputs(10162) <= layer0_outputs(3454);
    outputs(10163) <= layer0_outputs(4971);
    outputs(10164) <= not(layer0_outputs(2825));
    outputs(10165) <= layer0_outputs(5858);
    outputs(10166) <= layer0_outputs(5535);
    outputs(10167) <= layer0_outputs(6048);
    outputs(10168) <= not(layer0_outputs(1584));
    outputs(10169) <= layer0_outputs(98);
    outputs(10170) <= not((layer0_outputs(3805)) or (layer0_outputs(4169)));
    outputs(10171) <= not((layer0_outputs(8671)) or (layer0_outputs(1758)));
    outputs(10172) <= layer0_outputs(6022);
    outputs(10173) <= not((layer0_outputs(6799)) and (layer0_outputs(345)));
    outputs(10174) <= not(layer0_outputs(9177));
    outputs(10175) <= layer0_outputs(1995);
    outputs(10176) <= not((layer0_outputs(9918)) xor (layer0_outputs(8514)));
    outputs(10177) <= not(layer0_outputs(3219));
    outputs(10178) <= (layer0_outputs(3325)) xor (layer0_outputs(6383));
    outputs(10179) <= not(layer0_outputs(2559));
    outputs(10180) <= not((layer0_outputs(7959)) or (layer0_outputs(6235)));
    outputs(10181) <= not((layer0_outputs(3431)) xor (layer0_outputs(1345)));
    outputs(10182) <= (layer0_outputs(6121)) and not (layer0_outputs(6242));
    outputs(10183) <= layer0_outputs(3451);
    outputs(10184) <= (layer0_outputs(1094)) and not (layer0_outputs(4092));
    outputs(10185) <= (layer0_outputs(7108)) and (layer0_outputs(7060));
    outputs(10186) <= not((layer0_outputs(3356)) xor (layer0_outputs(5111)));
    outputs(10187) <= layer0_outputs(4830);
    outputs(10188) <= (layer0_outputs(1477)) xor (layer0_outputs(5399));
    outputs(10189) <= not(layer0_outputs(1270));
    outputs(10190) <= not((layer0_outputs(9866)) xor (layer0_outputs(6389)));
    outputs(10191) <= layer0_outputs(8596);
    outputs(10192) <= not(layer0_outputs(6745));
    outputs(10193) <= not((layer0_outputs(4358)) xor (layer0_outputs(2195)));
    outputs(10194) <= (layer0_outputs(7904)) xor (layer0_outputs(6068));
    outputs(10195) <= (layer0_outputs(3898)) or (layer0_outputs(2728));
    outputs(10196) <= (layer0_outputs(3185)) and (layer0_outputs(10002));
    outputs(10197) <= layer0_outputs(5956);
    outputs(10198) <= (layer0_outputs(7493)) and (layer0_outputs(3856));
    outputs(10199) <= not((layer0_outputs(3942)) xor (layer0_outputs(4341)));
    outputs(10200) <= not(layer0_outputs(1235));
    outputs(10201) <= (layer0_outputs(5664)) and not (layer0_outputs(4073));
    outputs(10202) <= (layer0_outputs(3699)) and not (layer0_outputs(4291));
    outputs(10203) <= (layer0_outputs(9508)) xor (layer0_outputs(712));
    outputs(10204) <= (layer0_outputs(3370)) and not (layer0_outputs(9323));
    outputs(10205) <= (layer0_outputs(7808)) xor (layer0_outputs(8695));
    outputs(10206) <= not(layer0_outputs(10205));
    outputs(10207) <= not(layer0_outputs(360));
    outputs(10208) <= (layer0_outputs(6924)) and not (layer0_outputs(6249));
    outputs(10209) <= not((layer0_outputs(6701)) xor (layer0_outputs(8066)));
    outputs(10210) <= not((layer0_outputs(7798)) xor (layer0_outputs(1494)));
    outputs(10211) <= (layer0_outputs(966)) or (layer0_outputs(4272));
    outputs(10212) <= (layer0_outputs(2247)) or (layer0_outputs(4103));
    outputs(10213) <= not((layer0_outputs(7004)) xor (layer0_outputs(470)));
    outputs(10214) <= not(layer0_outputs(2300));
    outputs(10215) <= not(layer0_outputs(587));
    outputs(10216) <= (layer0_outputs(8055)) and not (layer0_outputs(3592));
    outputs(10217) <= not(layer0_outputs(979));
    outputs(10218) <= (layer0_outputs(7640)) xor (layer0_outputs(7574));
    outputs(10219) <= (layer0_outputs(6342)) and not (layer0_outputs(1543));
    outputs(10220) <= not(layer0_outputs(5396));
    outputs(10221) <= not(layer0_outputs(3023));
    outputs(10222) <= not(layer0_outputs(6422));
    outputs(10223) <= not((layer0_outputs(3299)) xor (layer0_outputs(543)));
    outputs(10224) <= (layer0_outputs(4550)) and not (layer0_outputs(4549));
    outputs(10225) <= layer0_outputs(4759);
    outputs(10226) <= not((layer0_outputs(7482)) xor (layer0_outputs(1580)));
    outputs(10227) <= layer0_outputs(728);
    outputs(10228) <= not((layer0_outputs(3049)) or (layer0_outputs(6855)));
    outputs(10229) <= layer0_outputs(4589);
    outputs(10230) <= (layer0_outputs(2745)) xor (layer0_outputs(6610));
    outputs(10231) <= layer0_outputs(3458);
    outputs(10232) <= layer0_outputs(8368);
    outputs(10233) <= (layer0_outputs(8591)) xor (layer0_outputs(9586));
    outputs(10234) <= not(layer0_outputs(9932));
    outputs(10235) <= layer0_outputs(194);
    outputs(10236) <= (layer0_outputs(1680)) xor (layer0_outputs(3924));
    outputs(10237) <= (layer0_outputs(5346)) xor (layer0_outputs(9536));
    outputs(10238) <= layer0_outputs(77);
    outputs(10239) <= (layer0_outputs(7660)) xor (layer0_outputs(1599));

end Behavioral;
