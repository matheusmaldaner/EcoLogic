library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(9 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= (inputs(68)) and not (inputs(17));
    layer0_outputs(1) <= (inputs(232)) xor (inputs(239));
    layer0_outputs(2) <= not(inputs(243));
    layer0_outputs(3) <= not(inputs(41));
    layer0_outputs(4) <= not(inputs(78)) or (inputs(142));
    layer0_outputs(5) <= not(inputs(19));
    layer0_outputs(6) <= not(inputs(90)) or (inputs(47));
    layer0_outputs(7) <= not((inputs(233)) or (inputs(90)));
    layer0_outputs(8) <= (inputs(197)) xor (inputs(51));
    layer0_outputs(9) <= not((inputs(101)) xor (inputs(8)));
    layer0_outputs(10) <= (inputs(92)) and not (inputs(51));
    layer0_outputs(11) <= (inputs(196)) or (inputs(99));
    layer0_outputs(12) <= not((inputs(8)) xor (inputs(131)));
    layer0_outputs(13) <= (inputs(201)) or (inputs(37));
    layer0_outputs(14) <= (inputs(252)) xor (inputs(22));
    layer0_outputs(15) <= inputs(237);
    layer0_outputs(16) <= (inputs(161)) and (inputs(59));
    layer0_outputs(17) <= inputs(67);
    layer0_outputs(18) <= (inputs(157)) and not (inputs(35));
    layer0_outputs(19) <= not(inputs(69)) or (inputs(209));
    layer0_outputs(20) <= (inputs(50)) xor (inputs(177));
    layer0_outputs(21) <= inputs(246);
    layer0_outputs(22) <= (inputs(160)) and not (inputs(1));
    layer0_outputs(23) <= not(inputs(37));
    layer0_outputs(24) <= (inputs(158)) or (inputs(141));
    layer0_outputs(25) <= not(inputs(100));
    layer0_outputs(26) <= inputs(157);
    layer0_outputs(27) <= '0';
    layer0_outputs(28) <= inputs(69);
    layer0_outputs(29) <= not((inputs(247)) xor (inputs(218)));
    layer0_outputs(30) <= not((inputs(149)) xor (inputs(19)));
    layer0_outputs(31) <= inputs(72);
    layer0_outputs(32) <= not(inputs(27)) or (inputs(209));
    layer0_outputs(33) <= not(inputs(174)) or (inputs(47));
    layer0_outputs(34) <= not(inputs(235));
    layer0_outputs(35) <= not((inputs(184)) or (inputs(250)));
    layer0_outputs(36) <= inputs(20);
    layer0_outputs(37) <= '1';
    layer0_outputs(38) <= inputs(221);
    layer0_outputs(39) <= not((inputs(124)) or (inputs(189)));
    layer0_outputs(40) <= not((inputs(166)) xor (inputs(4)));
    layer0_outputs(41) <= not((inputs(100)) or (inputs(12)));
    layer0_outputs(42) <= not(inputs(232)) or (inputs(171));
    layer0_outputs(43) <= not(inputs(68));
    layer0_outputs(44) <= not((inputs(250)) or (inputs(215)));
    layer0_outputs(45) <= (inputs(157)) or (inputs(194));
    layer0_outputs(46) <= (inputs(140)) xor (inputs(14));
    layer0_outputs(47) <= not((inputs(202)) or (inputs(189)));
    layer0_outputs(48) <= (inputs(219)) or (inputs(84));
    layer0_outputs(49) <= (inputs(178)) or (inputs(65));
    layer0_outputs(50) <= (inputs(217)) and not (inputs(208));
    layer0_outputs(51) <= (inputs(106)) or (inputs(5));
    layer0_outputs(52) <= (inputs(92)) or (inputs(122));
    layer0_outputs(53) <= not((inputs(59)) or (inputs(162)));
    layer0_outputs(54) <= not((inputs(40)) or (inputs(174)));
    layer0_outputs(55) <= not((inputs(227)) xor (inputs(243)));
    layer0_outputs(56) <= not(inputs(92));
    layer0_outputs(57) <= not((inputs(44)) or (inputs(99)));
    layer0_outputs(58) <= (inputs(70)) or (inputs(251));
    layer0_outputs(59) <= not(inputs(185)) or (inputs(240));
    layer0_outputs(60) <= not((inputs(7)) or (inputs(234)));
    layer0_outputs(61) <= (inputs(143)) and not (inputs(178));
    layer0_outputs(62) <= '0';
    layer0_outputs(63) <= (inputs(186)) xor (inputs(52));
    layer0_outputs(64) <= (inputs(23)) xor (inputs(29));
    layer0_outputs(65) <= inputs(143);
    layer0_outputs(66) <= not(inputs(21));
    layer0_outputs(67) <= not(inputs(152)) or (inputs(73));
    layer0_outputs(68) <= (inputs(48)) and (inputs(223));
    layer0_outputs(69) <= inputs(202);
    layer0_outputs(70) <= inputs(229);
    layer0_outputs(71) <= (inputs(237)) or (inputs(56));
    layer0_outputs(72) <= (inputs(193)) and not (inputs(31));
    layer0_outputs(73) <= not(inputs(111)) or (inputs(235));
    layer0_outputs(74) <= not((inputs(47)) or (inputs(253)));
    layer0_outputs(75) <= (inputs(97)) and (inputs(89));
    layer0_outputs(76) <= (inputs(178)) and (inputs(244));
    layer0_outputs(77) <= '0';
    layer0_outputs(78) <= (inputs(181)) or (inputs(59));
    layer0_outputs(79) <= not((inputs(2)) and (inputs(20)));
    layer0_outputs(80) <= not((inputs(135)) or (inputs(197)));
    layer0_outputs(81) <= (inputs(240)) and not (inputs(101));
    layer0_outputs(82) <= not(inputs(103));
    layer0_outputs(83) <= (inputs(234)) xor (inputs(82));
    layer0_outputs(84) <= (inputs(153)) or (inputs(132));
    layer0_outputs(85) <= (inputs(47)) or (inputs(84));
    layer0_outputs(86) <= (inputs(206)) xor (inputs(102));
    layer0_outputs(87) <= (inputs(70)) and not (inputs(242));
    layer0_outputs(88) <= (inputs(83)) xor (inputs(174));
    layer0_outputs(89) <= not((inputs(39)) or (inputs(40)));
    layer0_outputs(90) <= not((inputs(7)) xor (inputs(181)));
    layer0_outputs(91) <= (inputs(98)) or (inputs(166));
    layer0_outputs(92) <= (inputs(225)) and not (inputs(248));
    layer0_outputs(93) <= not((inputs(58)) or (inputs(150)));
    layer0_outputs(94) <= not((inputs(243)) xor (inputs(242)));
    layer0_outputs(95) <= (inputs(114)) xor (inputs(174));
    layer0_outputs(96) <= not((inputs(237)) or (inputs(236)));
    layer0_outputs(97) <= inputs(199);
    layer0_outputs(98) <= (inputs(236)) xor (inputs(185));
    layer0_outputs(99) <= not(inputs(20));
    layer0_outputs(100) <= (inputs(104)) and not (inputs(224));
    layer0_outputs(101) <= not((inputs(180)) or (inputs(60)));
    layer0_outputs(102) <= not((inputs(247)) xor (inputs(218)));
    layer0_outputs(103) <= inputs(69);
    layer0_outputs(104) <= not(inputs(95));
    layer0_outputs(105) <= not((inputs(62)) xor (inputs(16)));
    layer0_outputs(106) <= not(inputs(104)) or (inputs(137));
    layer0_outputs(107) <= (inputs(153)) and not (inputs(11));
    layer0_outputs(108) <= (inputs(101)) or (inputs(86));
    layer0_outputs(109) <= not((inputs(227)) and (inputs(248)));
    layer0_outputs(110) <= (inputs(163)) xor (inputs(191));
    layer0_outputs(111) <= inputs(228);
    layer0_outputs(112) <= not((inputs(199)) or (inputs(15)));
    layer0_outputs(113) <= '1';
    layer0_outputs(114) <= (inputs(159)) or (inputs(107));
    layer0_outputs(115) <= not((inputs(102)) xor (inputs(167)));
    layer0_outputs(116) <= not((inputs(170)) or (inputs(236)));
    layer0_outputs(117) <= (inputs(4)) and not (inputs(21));
    layer0_outputs(118) <= (inputs(168)) xor (inputs(239));
    layer0_outputs(119) <= not(inputs(106));
    layer0_outputs(120) <= not(inputs(102));
    layer0_outputs(121) <= (inputs(234)) and not (inputs(141));
    layer0_outputs(122) <= (inputs(28)) and (inputs(65));
    layer0_outputs(123) <= (inputs(161)) xor (inputs(6));
    layer0_outputs(124) <= not(inputs(121)) or (inputs(69));
    layer0_outputs(125) <= inputs(151);
    layer0_outputs(126) <= (inputs(222)) or (inputs(58));
    layer0_outputs(127) <= not(inputs(88)) or (inputs(82));
    layer0_outputs(128) <= (inputs(122)) or (inputs(0));
    layer0_outputs(129) <= not((inputs(253)) xor (inputs(123)));
    layer0_outputs(130) <= inputs(77);
    layer0_outputs(131) <= not((inputs(147)) or (inputs(164)));
    layer0_outputs(132) <= not(inputs(200));
    layer0_outputs(133) <= not(inputs(198));
    layer0_outputs(134) <= not((inputs(188)) or (inputs(59)));
    layer0_outputs(135) <= not((inputs(247)) xor (inputs(181)));
    layer0_outputs(136) <= inputs(25);
    layer0_outputs(137) <= '1';
    layer0_outputs(138) <= (inputs(102)) and not (inputs(28));
    layer0_outputs(139) <= not(inputs(102)) or (inputs(161));
    layer0_outputs(140) <= not(inputs(202)) or (inputs(29));
    layer0_outputs(141) <= not(inputs(173));
    layer0_outputs(142) <= not(inputs(131)) or (inputs(24));
    layer0_outputs(143) <= '1';
    layer0_outputs(144) <= (inputs(33)) and not (inputs(218));
    layer0_outputs(145) <= (inputs(14)) or (inputs(139));
    layer0_outputs(146) <= (inputs(196)) and not (inputs(114));
    layer0_outputs(147) <= (inputs(57)) or (inputs(77));
    layer0_outputs(148) <= inputs(122);
    layer0_outputs(149) <= inputs(183);
    layer0_outputs(150) <= not((inputs(39)) xor (inputs(81)));
    layer0_outputs(151) <= (inputs(53)) and not (inputs(38));
    layer0_outputs(152) <= not(inputs(193));
    layer0_outputs(153) <= not(inputs(85));
    layer0_outputs(154) <= (inputs(71)) or (inputs(95));
    layer0_outputs(155) <= not(inputs(87)) or (inputs(205));
    layer0_outputs(156) <= not(inputs(190)) or (inputs(30));
    layer0_outputs(157) <= inputs(56);
    layer0_outputs(158) <= (inputs(48)) xor (inputs(210));
    layer0_outputs(159) <= not(inputs(21)) or (inputs(82));
    layer0_outputs(160) <= (inputs(199)) and not (inputs(177));
    layer0_outputs(161) <= (inputs(10)) and not (inputs(128));
    layer0_outputs(162) <= not(inputs(151)) or (inputs(248));
    layer0_outputs(163) <= not((inputs(93)) or (inputs(197)));
    layer0_outputs(164) <= (inputs(225)) xor (inputs(166));
    layer0_outputs(165) <= (inputs(29)) and not (inputs(4));
    layer0_outputs(166) <= not(inputs(181)) or (inputs(29));
    layer0_outputs(167) <= not((inputs(205)) xor (inputs(231)));
    layer0_outputs(168) <= not((inputs(251)) or (inputs(101)));
    layer0_outputs(169) <= not(inputs(181));
    layer0_outputs(170) <= (inputs(96)) xor (inputs(58));
    layer0_outputs(171) <= not((inputs(37)) or (inputs(158)));
    layer0_outputs(172) <= not(inputs(215));
    layer0_outputs(173) <= (inputs(153)) and not (inputs(116));
    layer0_outputs(174) <= (inputs(41)) xor (inputs(254));
    layer0_outputs(175) <= (inputs(118)) and not (inputs(240));
    layer0_outputs(176) <= not((inputs(218)) or (inputs(204)));
    layer0_outputs(177) <= (inputs(237)) and (inputs(241));
    layer0_outputs(178) <= (inputs(33)) xor (inputs(251));
    layer0_outputs(179) <= inputs(66);
    layer0_outputs(180) <= not((inputs(251)) or (inputs(242)));
    layer0_outputs(181) <= inputs(10);
    layer0_outputs(182) <= (inputs(181)) and not (inputs(78));
    layer0_outputs(183) <= inputs(121);
    layer0_outputs(184) <= (inputs(52)) or (inputs(8));
    layer0_outputs(185) <= (inputs(104)) and not (inputs(186));
    layer0_outputs(186) <= (inputs(2)) and not (inputs(124));
    layer0_outputs(187) <= not(inputs(108));
    layer0_outputs(188) <= (inputs(126)) and not (inputs(19));
    layer0_outputs(189) <= (inputs(16)) xor (inputs(229));
    layer0_outputs(190) <= inputs(179);
    layer0_outputs(191) <= not(inputs(118)) or (inputs(18));
    layer0_outputs(192) <= not((inputs(156)) xor (inputs(127)));
    layer0_outputs(193) <= not(inputs(220));
    layer0_outputs(194) <= (inputs(240)) or (inputs(159));
    layer0_outputs(195) <= (inputs(62)) or (inputs(78));
    layer0_outputs(196) <= not(inputs(136));
    layer0_outputs(197) <= not(inputs(64)) or (inputs(11));
    layer0_outputs(198) <= (inputs(255)) and (inputs(32));
    layer0_outputs(199) <= (inputs(43)) xor (inputs(34));
    layer0_outputs(200) <= not(inputs(183));
    layer0_outputs(201) <= (inputs(213)) and not (inputs(13));
    layer0_outputs(202) <= not(inputs(214)) or (inputs(211));
    layer0_outputs(203) <= not(inputs(66));
    layer0_outputs(204) <= not(inputs(220)) or (inputs(226));
    layer0_outputs(205) <= not(inputs(151));
    layer0_outputs(206) <= not(inputs(132)) or (inputs(79));
    layer0_outputs(207) <= (inputs(203)) and not (inputs(10));
    layer0_outputs(208) <= (inputs(101)) or (inputs(225));
    layer0_outputs(209) <= inputs(198);
    layer0_outputs(210) <= not((inputs(102)) or (inputs(141)));
    layer0_outputs(211) <= (inputs(27)) or (inputs(200));
    layer0_outputs(212) <= not(inputs(37)) or (inputs(125));
    layer0_outputs(213) <= not((inputs(194)) or (inputs(170)));
    layer0_outputs(214) <= not(inputs(237));
    layer0_outputs(215) <= inputs(165);
    layer0_outputs(216) <= not((inputs(165)) or (inputs(97)));
    layer0_outputs(217) <= inputs(119);
    layer0_outputs(218) <= inputs(230);
    layer0_outputs(219) <= inputs(56);
    layer0_outputs(220) <= not(inputs(66));
    layer0_outputs(221) <= not((inputs(151)) or (inputs(228)));
    layer0_outputs(222) <= (inputs(61)) or (inputs(139));
    layer0_outputs(223) <= not((inputs(174)) or (inputs(247)));
    layer0_outputs(224) <= not(inputs(88)) or (inputs(16));
    layer0_outputs(225) <= inputs(246);
    layer0_outputs(226) <= inputs(118);
    layer0_outputs(227) <= not(inputs(180)) or (inputs(127));
    layer0_outputs(228) <= (inputs(166)) and not (inputs(94));
    layer0_outputs(229) <= (inputs(41)) xor (inputs(73));
    layer0_outputs(230) <= not((inputs(82)) or (inputs(150)));
    layer0_outputs(231) <= not(inputs(82));
    layer0_outputs(232) <= not(inputs(197));
    layer0_outputs(233) <= not(inputs(27));
    layer0_outputs(234) <= '1';
    layer0_outputs(235) <= (inputs(14)) xor (inputs(135));
    layer0_outputs(236) <= not((inputs(220)) xor (inputs(31)));
    layer0_outputs(237) <= inputs(153);
    layer0_outputs(238) <= not(inputs(184)) or (inputs(231));
    layer0_outputs(239) <= (inputs(64)) or (inputs(153));
    layer0_outputs(240) <= not(inputs(166)) or (inputs(249));
    layer0_outputs(241) <= not(inputs(99)) or (inputs(66));
    layer0_outputs(242) <= not(inputs(99)) or (inputs(253));
    layer0_outputs(243) <= (inputs(244)) or (inputs(225));
    layer0_outputs(244) <= inputs(218);
    layer0_outputs(245) <= not(inputs(7)) or (inputs(238));
    layer0_outputs(246) <= not(inputs(150)) or (inputs(66));
    layer0_outputs(247) <= not((inputs(218)) or (inputs(190)));
    layer0_outputs(248) <= inputs(38);
    layer0_outputs(249) <= not(inputs(204));
    layer0_outputs(250) <= (inputs(187)) and not (inputs(114));
    layer0_outputs(251) <= not(inputs(173));
    layer0_outputs(252) <= (inputs(57)) or (inputs(147));
    layer0_outputs(253) <= not(inputs(203)) or (inputs(19));
    layer0_outputs(254) <= not(inputs(70));
    layer0_outputs(255) <= not((inputs(51)) or (inputs(220)));
    layer0_outputs(256) <= not(inputs(157));
    layer0_outputs(257) <= not(inputs(232)) or (inputs(69));
    layer0_outputs(258) <= not((inputs(139)) or (inputs(39)));
    layer0_outputs(259) <= not(inputs(88));
    layer0_outputs(260) <= inputs(131);
    layer0_outputs(261) <= not((inputs(118)) xor (inputs(174)));
    layer0_outputs(262) <= not(inputs(126));
    layer0_outputs(263) <= inputs(12);
    layer0_outputs(264) <= not((inputs(93)) or (inputs(222)));
    layer0_outputs(265) <= not((inputs(214)) and (inputs(234)));
    layer0_outputs(266) <= not((inputs(42)) or (inputs(38)));
    layer0_outputs(267) <= not(inputs(207));
    layer0_outputs(268) <= (inputs(28)) and (inputs(5));
    layer0_outputs(269) <= (inputs(196)) xor (inputs(26));
    layer0_outputs(270) <= not(inputs(150));
    layer0_outputs(271) <= (inputs(210)) xor (inputs(178));
    layer0_outputs(272) <= not(inputs(28));
    layer0_outputs(273) <= not(inputs(163));
    layer0_outputs(274) <= not(inputs(126));
    layer0_outputs(275) <= (inputs(89)) and not (inputs(233));
    layer0_outputs(276) <= (inputs(94)) or (inputs(96));
    layer0_outputs(277) <= not((inputs(27)) or (inputs(103)));
    layer0_outputs(278) <= inputs(1);
    layer0_outputs(279) <= (inputs(34)) or (inputs(68));
    layer0_outputs(280) <= not((inputs(117)) or (inputs(45)));
    layer0_outputs(281) <= not(inputs(194)) or (inputs(205));
    layer0_outputs(282) <= not(inputs(175));
    layer0_outputs(283) <= not(inputs(165));
    layer0_outputs(284) <= not((inputs(157)) or (inputs(169)));
    layer0_outputs(285) <= not(inputs(68)) or (inputs(158));
    layer0_outputs(286) <= not((inputs(92)) or (inputs(235)));
    layer0_outputs(287) <= not((inputs(100)) xor (inputs(57)));
    layer0_outputs(288) <= inputs(121);
    layer0_outputs(289) <= inputs(150);
    layer0_outputs(290) <= '1';
    layer0_outputs(291) <= not((inputs(240)) xor (inputs(174)));
    layer0_outputs(292) <= not(inputs(137)) or (inputs(95));
    layer0_outputs(293) <= (inputs(221)) or (inputs(147));
    layer0_outputs(294) <= not(inputs(199)) or (inputs(137));
    layer0_outputs(295) <= (inputs(197)) or (inputs(198));
    layer0_outputs(296) <= not(inputs(38));
    layer0_outputs(297) <= inputs(151);
    layer0_outputs(298) <= not(inputs(172)) or (inputs(98));
    layer0_outputs(299) <= not(inputs(93));
    layer0_outputs(300) <= not((inputs(61)) or (inputs(115)));
    layer0_outputs(301) <= (inputs(75)) and not (inputs(80));
    layer0_outputs(302) <= not((inputs(207)) or (inputs(92)));
    layer0_outputs(303) <= (inputs(16)) xor (inputs(157));
    layer0_outputs(304) <= not(inputs(229)) or (inputs(220));
    layer0_outputs(305) <= not(inputs(166));
    layer0_outputs(306) <= (inputs(170)) and (inputs(88));
    layer0_outputs(307) <= inputs(130);
    layer0_outputs(308) <= (inputs(211)) or (inputs(214));
    layer0_outputs(309) <= not((inputs(148)) or (inputs(134)));
    layer0_outputs(310) <= not((inputs(132)) or (inputs(76)));
    layer0_outputs(311) <= inputs(124);
    layer0_outputs(312) <= (inputs(233)) or (inputs(97));
    layer0_outputs(313) <= not((inputs(177)) or (inputs(73)));
    layer0_outputs(314) <= (inputs(133)) and not (inputs(239));
    layer0_outputs(315) <= inputs(91);
    layer0_outputs(316) <= (inputs(201)) xor (inputs(252));
    layer0_outputs(317) <= not((inputs(6)) or (inputs(84)));
    layer0_outputs(318) <= not((inputs(171)) xor (inputs(10)));
    layer0_outputs(319) <= (inputs(246)) or (inputs(107));
    layer0_outputs(320) <= (inputs(160)) and not (inputs(105));
    layer0_outputs(321) <= inputs(152);
    layer0_outputs(322) <= not((inputs(234)) or (inputs(70)));
    layer0_outputs(323) <= not(inputs(90)) or (inputs(45));
    layer0_outputs(324) <= not((inputs(223)) or (inputs(56)));
    layer0_outputs(325) <= not((inputs(150)) or (inputs(39)));
    layer0_outputs(326) <= not(inputs(216));
    layer0_outputs(327) <= '1';
    layer0_outputs(328) <= (inputs(153)) or (inputs(68));
    layer0_outputs(329) <= (inputs(180)) xor (inputs(9));
    layer0_outputs(330) <= (inputs(138)) and not (inputs(45));
    layer0_outputs(331) <= inputs(58);
    layer0_outputs(332) <= not(inputs(232));
    layer0_outputs(333) <= inputs(180);
    layer0_outputs(334) <= (inputs(179)) or (inputs(203));
    layer0_outputs(335) <= (inputs(245)) and not (inputs(129));
    layer0_outputs(336) <= (inputs(180)) and not (inputs(214));
    layer0_outputs(337) <= '0';
    layer0_outputs(338) <= not(inputs(136)) or (inputs(31));
    layer0_outputs(339) <= (inputs(211)) and not (inputs(49));
    layer0_outputs(340) <= (inputs(153)) or (inputs(203));
    layer0_outputs(341) <= not(inputs(142));
    layer0_outputs(342) <= not(inputs(236));
    layer0_outputs(343) <= (inputs(7)) or (inputs(207));
    layer0_outputs(344) <= not(inputs(150)) or (inputs(222));
    layer0_outputs(345) <= (inputs(32)) and (inputs(169));
    layer0_outputs(346) <= (inputs(34)) xor (inputs(191));
    layer0_outputs(347) <= inputs(252);
    layer0_outputs(348) <= (inputs(235)) and not (inputs(227));
    layer0_outputs(349) <= (inputs(97)) or (inputs(107));
    layer0_outputs(350) <= (inputs(116)) and not (inputs(234));
    layer0_outputs(351) <= not(inputs(139)) or (inputs(76));
    layer0_outputs(352) <= not((inputs(94)) or (inputs(199)));
    layer0_outputs(353) <= (inputs(155)) and not (inputs(22));
    layer0_outputs(354) <= not((inputs(208)) or (inputs(170)));
    layer0_outputs(355) <= not((inputs(24)) or (inputs(190)));
    layer0_outputs(356) <= (inputs(72)) and (inputs(212));
    layer0_outputs(357) <= not((inputs(143)) and (inputs(54)));
    layer0_outputs(358) <= not((inputs(64)) xor (inputs(106)));
    layer0_outputs(359) <= (inputs(13)) or (inputs(75));
    layer0_outputs(360) <= not(inputs(102));
    layer0_outputs(361) <= not((inputs(236)) or (inputs(218)));
    layer0_outputs(362) <= not(inputs(178));
    layer0_outputs(363) <= (inputs(221)) and not (inputs(226));
    layer0_outputs(364) <= (inputs(102)) and not (inputs(244));
    layer0_outputs(365) <= not(inputs(141)) or (inputs(205));
    layer0_outputs(366) <= not(inputs(162));
    layer0_outputs(367) <= inputs(135);
    layer0_outputs(368) <= not((inputs(138)) or (inputs(250)));
    layer0_outputs(369) <= not(inputs(135));
    layer0_outputs(370) <= not((inputs(61)) and (inputs(171)));
    layer0_outputs(371) <= not((inputs(7)) xor (inputs(233)));
    layer0_outputs(372) <= not(inputs(3)) or (inputs(241));
    layer0_outputs(373) <= not((inputs(202)) or (inputs(218)));
    layer0_outputs(374) <= not((inputs(147)) xor (inputs(252)));
    layer0_outputs(375) <= not(inputs(84)) or (inputs(221));
    layer0_outputs(376) <= not(inputs(90)) or (inputs(204));
    layer0_outputs(377) <= '0';
    layer0_outputs(378) <= inputs(102);
    layer0_outputs(379) <= not((inputs(114)) xor (inputs(147)));
    layer0_outputs(380) <= not(inputs(167));
    layer0_outputs(381) <= (inputs(77)) or (inputs(63));
    layer0_outputs(382) <= not((inputs(58)) xor (inputs(141)));
    layer0_outputs(383) <= (inputs(54)) xor (inputs(236));
    layer0_outputs(384) <= not(inputs(118));
    layer0_outputs(385) <= not((inputs(228)) or (inputs(223)));
    layer0_outputs(386) <= (inputs(0)) xor (inputs(219));
    layer0_outputs(387) <= (inputs(65)) and not (inputs(37));
    layer0_outputs(388) <= not((inputs(93)) or (inputs(253)));
    layer0_outputs(389) <= (inputs(155)) and not (inputs(114));
    layer0_outputs(390) <= not((inputs(152)) and (inputs(152)));
    layer0_outputs(391) <= not(inputs(101)) or (inputs(64));
    layer0_outputs(392) <= (inputs(27)) xor (inputs(20));
    layer0_outputs(393) <= inputs(130);
    layer0_outputs(394) <= (inputs(211)) or (inputs(51));
    layer0_outputs(395) <= not(inputs(164));
    layer0_outputs(396) <= not(inputs(91)) or (inputs(128));
    layer0_outputs(397) <= (inputs(246)) or (inputs(251));
    layer0_outputs(398) <= (inputs(160)) and not (inputs(62));
    layer0_outputs(399) <= (inputs(23)) or (inputs(170));
    layer0_outputs(400) <= (inputs(185)) and not (inputs(234));
    layer0_outputs(401) <= not(inputs(152));
    layer0_outputs(402) <= (inputs(237)) and (inputs(8));
    layer0_outputs(403) <= not(inputs(235)) or (inputs(213));
    layer0_outputs(404) <= inputs(228);
    layer0_outputs(405) <= (inputs(168)) and not (inputs(92));
    layer0_outputs(406) <= not(inputs(253)) or (inputs(209));
    layer0_outputs(407) <= (inputs(20)) and not (inputs(165));
    layer0_outputs(408) <= (inputs(127)) xor (inputs(55));
    layer0_outputs(409) <= (inputs(168)) and not (inputs(13));
    layer0_outputs(410) <= not(inputs(200)) or (inputs(53));
    layer0_outputs(411) <= (inputs(52)) xor (inputs(193));
    layer0_outputs(412) <= inputs(182);
    layer0_outputs(413) <= (inputs(123)) and not (inputs(94));
    layer0_outputs(414) <= not(inputs(51)) or (inputs(133));
    layer0_outputs(415) <= inputs(120);
    layer0_outputs(416) <= not((inputs(81)) or (inputs(136)));
    layer0_outputs(417) <= not((inputs(2)) or (inputs(172)));
    layer0_outputs(418) <= inputs(92);
    layer0_outputs(419) <= (inputs(147)) and not (inputs(189));
    layer0_outputs(420) <= inputs(89);
    layer0_outputs(421) <= (inputs(119)) and not (inputs(221));
    layer0_outputs(422) <= inputs(249);
    layer0_outputs(423) <= (inputs(157)) or (inputs(23));
    layer0_outputs(424) <= not((inputs(81)) xor (inputs(46)));
    layer0_outputs(425) <= not((inputs(62)) or (inputs(109)));
    layer0_outputs(426) <= (inputs(94)) xor (inputs(113));
    layer0_outputs(427) <= not((inputs(124)) or (inputs(26)));
    layer0_outputs(428) <= inputs(165);
    layer0_outputs(429) <= not((inputs(4)) or (inputs(37)));
    layer0_outputs(430) <= (inputs(200)) and (inputs(171));
    layer0_outputs(431) <= (inputs(142)) xor (inputs(201));
    layer0_outputs(432) <= (inputs(94)) or (inputs(181));
    layer0_outputs(433) <= (inputs(22)) or (inputs(162));
    layer0_outputs(434) <= (inputs(227)) and not (inputs(115));
    layer0_outputs(435) <= not(inputs(41)) or (inputs(4));
    layer0_outputs(436) <= not((inputs(194)) xor (inputs(205)));
    layer0_outputs(437) <= (inputs(136)) and not (inputs(213));
    layer0_outputs(438) <= (inputs(76)) and not (inputs(202));
    layer0_outputs(439) <= not((inputs(201)) xor (inputs(11)));
    layer0_outputs(440) <= not(inputs(56));
    layer0_outputs(441) <= (inputs(191)) or (inputs(82));
    layer0_outputs(442) <= inputs(60);
    layer0_outputs(443) <= (inputs(200)) xor (inputs(63));
    layer0_outputs(444) <= (inputs(123)) and (inputs(252));
    layer0_outputs(445) <= not(inputs(87));
    layer0_outputs(446) <= (inputs(55)) xor (inputs(7));
    layer0_outputs(447) <= (inputs(101)) xor (inputs(131));
    layer0_outputs(448) <= not((inputs(27)) or (inputs(43)));
    layer0_outputs(449) <= not((inputs(104)) or (inputs(63)));
    layer0_outputs(450) <= not(inputs(54)) or (inputs(249));
    layer0_outputs(451) <= (inputs(107)) and not (inputs(61));
    layer0_outputs(452) <= (inputs(173)) or (inputs(78));
    layer0_outputs(453) <= not((inputs(199)) or (inputs(131)));
    layer0_outputs(454) <= (inputs(137)) xor (inputs(170));
    layer0_outputs(455) <= (inputs(178)) and not (inputs(112));
    layer0_outputs(456) <= not((inputs(96)) xor (inputs(200)));
    layer0_outputs(457) <= not(inputs(137)) or (inputs(250));
    layer0_outputs(458) <= (inputs(72)) and not (inputs(167));
    layer0_outputs(459) <= not((inputs(44)) or (inputs(127)));
    layer0_outputs(460) <= not((inputs(164)) or (inputs(50)));
    layer0_outputs(461) <= not((inputs(218)) or (inputs(188)));
    layer0_outputs(462) <= (inputs(127)) and not (inputs(238));
    layer0_outputs(463) <= (inputs(125)) or (inputs(109));
    layer0_outputs(464) <= (inputs(33)) and (inputs(145));
    layer0_outputs(465) <= (inputs(24)) and (inputs(129));
    layer0_outputs(466) <= inputs(251);
    layer0_outputs(467) <= not(inputs(102)) or (inputs(53));
    layer0_outputs(468) <= (inputs(228)) or (inputs(149));
    layer0_outputs(469) <= (inputs(224)) xor (inputs(212));
    layer0_outputs(470) <= not(inputs(57)) or (inputs(172));
    layer0_outputs(471) <= '1';
    layer0_outputs(472) <= inputs(215);
    layer0_outputs(473) <= not(inputs(91));
    layer0_outputs(474) <= (inputs(240)) and (inputs(193));
    layer0_outputs(475) <= (inputs(98)) xor (inputs(117));
    layer0_outputs(476) <= (inputs(92)) xor (inputs(90));
    layer0_outputs(477) <= (inputs(200)) or (inputs(163));
    layer0_outputs(478) <= '0';
    layer0_outputs(479) <= not(inputs(122));
    layer0_outputs(480) <= not((inputs(18)) or (inputs(144)));
    layer0_outputs(481) <= not((inputs(33)) or (inputs(120)));
    layer0_outputs(482) <= (inputs(251)) and (inputs(79));
    layer0_outputs(483) <= not(inputs(215)) or (inputs(61));
    layer0_outputs(484) <= (inputs(250)) and (inputs(168));
    layer0_outputs(485) <= not(inputs(97));
    layer0_outputs(486) <= (inputs(214)) and not (inputs(147));
    layer0_outputs(487) <= not((inputs(23)) or (inputs(109)));
    layer0_outputs(488) <= not((inputs(89)) or (inputs(189)));
    layer0_outputs(489) <= (inputs(123)) and not (inputs(82));
    layer0_outputs(490) <= (inputs(183)) and not (inputs(114));
    layer0_outputs(491) <= not(inputs(155)) or (inputs(13));
    layer0_outputs(492) <= not(inputs(39)) or (inputs(13));
    layer0_outputs(493) <= not(inputs(40)) or (inputs(48));
    layer0_outputs(494) <= inputs(59);
    layer0_outputs(495) <= not((inputs(249)) or (inputs(233)));
    layer0_outputs(496) <= not(inputs(155)) or (inputs(49));
    layer0_outputs(497) <= inputs(80);
    layer0_outputs(498) <= (inputs(187)) and not (inputs(95));
    layer0_outputs(499) <= (inputs(235)) xor (inputs(230));
    layer0_outputs(500) <= (inputs(32)) or (inputs(23));
    layer0_outputs(501) <= not(inputs(120)) or (inputs(12));
    layer0_outputs(502) <= inputs(122);
    layer0_outputs(503) <= inputs(221);
    layer0_outputs(504) <= inputs(189);
    layer0_outputs(505) <= (inputs(156)) and not (inputs(98));
    layer0_outputs(506) <= (inputs(160)) xor (inputs(248));
    layer0_outputs(507) <= inputs(120);
    layer0_outputs(508) <= (inputs(99)) and not (inputs(59));
    layer0_outputs(509) <= not(inputs(76));
    layer0_outputs(510) <= not(inputs(39)) or (inputs(228));
    layer0_outputs(511) <= (inputs(128)) or (inputs(114));
    layer0_outputs(512) <= not((inputs(159)) xor (inputs(217)));
    layer0_outputs(513) <= not(inputs(106)) or (inputs(13));
    layer0_outputs(514) <= not((inputs(176)) and (inputs(17)));
    layer0_outputs(515) <= not((inputs(205)) or (inputs(189)));
    layer0_outputs(516) <= not(inputs(231));
    layer0_outputs(517) <= not((inputs(230)) and (inputs(1)));
    layer0_outputs(518) <= not((inputs(49)) xor (inputs(105)));
    layer0_outputs(519) <= inputs(153);
    layer0_outputs(520) <= inputs(92);
    layer0_outputs(521) <= (inputs(196)) and not (inputs(246));
    layer0_outputs(522) <= '1';
    layer0_outputs(523) <= inputs(107);
    layer0_outputs(524) <= (inputs(102)) and not (inputs(254));
    layer0_outputs(525) <= (inputs(71)) or (inputs(242));
    layer0_outputs(526) <= (inputs(130)) xor (inputs(195));
    layer0_outputs(527) <= not((inputs(79)) xor (inputs(120)));
    layer0_outputs(528) <= not(inputs(27)) or (inputs(18));
    layer0_outputs(529) <= not(inputs(105));
    layer0_outputs(530) <= (inputs(148)) xor (inputs(224));
    layer0_outputs(531) <= not((inputs(153)) or (inputs(34)));
    layer0_outputs(532) <= not((inputs(46)) and (inputs(163)));
    layer0_outputs(533) <= (inputs(238)) and (inputs(216));
    layer0_outputs(534) <= not(inputs(130)) or (inputs(74));
    layer0_outputs(535) <= (inputs(14)) and (inputs(33));
    layer0_outputs(536) <= (inputs(115)) or (inputs(138));
    layer0_outputs(537) <= not(inputs(154));
    layer0_outputs(538) <= not((inputs(151)) or (inputs(233)));
    layer0_outputs(539) <= not((inputs(165)) or (inputs(37)));
    layer0_outputs(540) <= not(inputs(107));
    layer0_outputs(541) <= inputs(40);
    layer0_outputs(542) <= inputs(240);
    layer0_outputs(543) <= (inputs(48)) or (inputs(157));
    layer0_outputs(544) <= not((inputs(3)) or (inputs(148)));
    layer0_outputs(545) <= inputs(173);
    layer0_outputs(546) <= inputs(56);
    layer0_outputs(547) <= (inputs(29)) xor (inputs(67));
    layer0_outputs(548) <= not((inputs(249)) or (inputs(135)));
    layer0_outputs(549) <= (inputs(114)) xor (inputs(67));
    layer0_outputs(550) <= not(inputs(112));
    layer0_outputs(551) <= not(inputs(70));
    layer0_outputs(552) <= (inputs(3)) or (inputs(122));
    layer0_outputs(553) <= (inputs(194)) xor (inputs(230));
    layer0_outputs(554) <= (inputs(149)) and not (inputs(211));
    layer0_outputs(555) <= (inputs(235)) and not (inputs(17));
    layer0_outputs(556) <= inputs(124);
    layer0_outputs(557) <= (inputs(163)) and not (inputs(247));
    layer0_outputs(558) <= (inputs(156)) or (inputs(232));
    layer0_outputs(559) <= not(inputs(165));
    layer0_outputs(560) <= (inputs(234)) xor (inputs(116));
    layer0_outputs(561) <= (inputs(231)) and not (inputs(196));
    layer0_outputs(562) <= not((inputs(74)) xor (inputs(11)));
    layer0_outputs(563) <= (inputs(32)) or (inputs(16));
    layer0_outputs(564) <= (inputs(214)) or (inputs(222));
    layer0_outputs(565) <= not((inputs(139)) xor (inputs(134)));
    layer0_outputs(566) <= (inputs(175)) xor (inputs(226));
    layer0_outputs(567) <= not(inputs(39));
    layer0_outputs(568) <= not((inputs(109)) xor (inputs(87)));
    layer0_outputs(569) <= (inputs(190)) or (inputs(75));
    layer0_outputs(570) <= (inputs(220)) or (inputs(201));
    layer0_outputs(571) <= (inputs(69)) or (inputs(172));
    layer0_outputs(572) <= not(inputs(250)) or (inputs(154));
    layer0_outputs(573) <= not((inputs(72)) or (inputs(2)));
    layer0_outputs(574) <= not((inputs(88)) or (inputs(13)));
    layer0_outputs(575) <= not((inputs(133)) or (inputs(220)));
    layer0_outputs(576) <= not(inputs(77)) or (inputs(246));
    layer0_outputs(577) <= not(inputs(121)) or (inputs(13));
    layer0_outputs(578) <= (inputs(29)) or (inputs(152));
    layer0_outputs(579) <= not(inputs(130)) or (inputs(145));
    layer0_outputs(580) <= (inputs(72)) and not (inputs(11));
    layer0_outputs(581) <= (inputs(102)) and not (inputs(32));
    layer0_outputs(582) <= not((inputs(91)) or (inputs(237)));
    layer0_outputs(583) <= not(inputs(125)) or (inputs(20));
    layer0_outputs(584) <= (inputs(119)) or (inputs(250));
    layer0_outputs(585) <= not((inputs(143)) and (inputs(30)));
    layer0_outputs(586) <= not(inputs(76));
    layer0_outputs(587) <= (inputs(54)) xor (inputs(30));
    layer0_outputs(588) <= (inputs(89)) or (inputs(111));
    layer0_outputs(589) <= (inputs(246)) xor (inputs(1));
    layer0_outputs(590) <= '0';
    layer0_outputs(591) <= not((inputs(77)) xor (inputs(44)));
    layer0_outputs(592) <= not(inputs(185)) or (inputs(117));
    layer0_outputs(593) <= not(inputs(50));
    layer0_outputs(594) <= not(inputs(216)) or (inputs(146));
    layer0_outputs(595) <= (inputs(173)) xor (inputs(140));
    layer0_outputs(596) <= (inputs(135)) or (inputs(79));
    layer0_outputs(597) <= not(inputs(204));
    layer0_outputs(598) <= (inputs(30)) or (inputs(147));
    layer0_outputs(599) <= (inputs(5)) or (inputs(178));
    layer0_outputs(600) <= (inputs(26)) and not (inputs(7));
    layer0_outputs(601) <= not((inputs(132)) xor (inputs(241)));
    layer0_outputs(602) <= (inputs(19)) and (inputs(50));
    layer0_outputs(603) <= not((inputs(70)) or (inputs(147)));
    layer0_outputs(604) <= '1';
    layer0_outputs(605) <= not(inputs(101));
    layer0_outputs(606) <= not(inputs(167)) or (inputs(10));
    layer0_outputs(607) <= (inputs(251)) or (inputs(21));
    layer0_outputs(608) <= not(inputs(115));
    layer0_outputs(609) <= (inputs(106)) or (inputs(6));
    layer0_outputs(610) <= (inputs(112)) or (inputs(54));
    layer0_outputs(611) <= not(inputs(170));
    layer0_outputs(612) <= (inputs(205)) or (inputs(101));
    layer0_outputs(613) <= (inputs(192)) or (inputs(207));
    layer0_outputs(614) <= not(inputs(134)) or (inputs(245));
    layer0_outputs(615) <= inputs(94);
    layer0_outputs(616) <= (inputs(53)) xor (inputs(112));
    layer0_outputs(617) <= not((inputs(190)) or (inputs(178)));
    layer0_outputs(618) <= not(inputs(105));
    layer0_outputs(619) <= not((inputs(202)) and (inputs(113)));
    layer0_outputs(620) <= inputs(101);
    layer0_outputs(621) <= (inputs(38)) or (inputs(183));
    layer0_outputs(622) <= not(inputs(119)) or (inputs(149));
    layer0_outputs(623) <= (inputs(184)) or (inputs(211));
    layer0_outputs(624) <= (inputs(223)) or (inputs(165));
    layer0_outputs(625) <= '0';
    layer0_outputs(626) <= (inputs(19)) and not (inputs(163));
    layer0_outputs(627) <= (inputs(98)) or (inputs(233));
    layer0_outputs(628) <= (inputs(222)) or (inputs(126));
    layer0_outputs(629) <= (inputs(155)) and not (inputs(235));
    layer0_outputs(630) <= inputs(51);
    layer0_outputs(631) <= not(inputs(104));
    layer0_outputs(632) <= (inputs(231)) xor (inputs(227));
    layer0_outputs(633) <= (inputs(21)) or (inputs(187));
    layer0_outputs(634) <= not((inputs(164)) xor (inputs(186)));
    layer0_outputs(635) <= not((inputs(253)) xor (inputs(193)));
    layer0_outputs(636) <= (inputs(150)) and (inputs(237));
    layer0_outputs(637) <= (inputs(230)) and not (inputs(202));
    layer0_outputs(638) <= not(inputs(201)) or (inputs(32));
    layer0_outputs(639) <= not(inputs(152));
    layer0_outputs(640) <= not(inputs(85)) or (inputs(24));
    layer0_outputs(641) <= inputs(233);
    layer0_outputs(642) <= not(inputs(210));
    layer0_outputs(643) <= not(inputs(229)) or (inputs(176));
    layer0_outputs(644) <= (inputs(98)) or (inputs(122));
    layer0_outputs(645) <= not(inputs(158));
    layer0_outputs(646) <= not(inputs(76));
    layer0_outputs(647) <= not((inputs(101)) or (inputs(70)));
    layer0_outputs(648) <= (inputs(252)) and (inputs(17));
    layer0_outputs(649) <= '1';
    layer0_outputs(650) <= not(inputs(43)) or (inputs(6));
    layer0_outputs(651) <= not(inputs(58));
    layer0_outputs(652) <= not((inputs(28)) and (inputs(161)));
    layer0_outputs(653) <= (inputs(64)) or (inputs(99));
    layer0_outputs(654) <= (inputs(132)) and not (inputs(112));
    layer0_outputs(655) <= not(inputs(79)) or (inputs(25));
    layer0_outputs(656) <= not(inputs(195)) or (inputs(177));
    layer0_outputs(657) <= not(inputs(90)) or (inputs(0));
    layer0_outputs(658) <= (inputs(209)) or (inputs(171));
    layer0_outputs(659) <= not(inputs(227)) or (inputs(6));
    layer0_outputs(660) <= (inputs(245)) and not (inputs(175));
    layer0_outputs(661) <= (inputs(31)) or (inputs(7));
    layer0_outputs(662) <= (inputs(201)) and not (inputs(131));
    layer0_outputs(663) <= (inputs(211)) and (inputs(143));
    layer0_outputs(664) <= inputs(188);
    layer0_outputs(665) <= (inputs(86)) and not (inputs(43));
    layer0_outputs(666) <= not((inputs(232)) or (inputs(66)));
    layer0_outputs(667) <= inputs(107);
    layer0_outputs(668) <= (inputs(71)) and not (inputs(30));
    layer0_outputs(669) <= not((inputs(196)) or (inputs(218)));
    layer0_outputs(670) <= (inputs(213)) xor (inputs(244));
    layer0_outputs(671) <= (inputs(44)) xor (inputs(219));
    layer0_outputs(672) <= not(inputs(103)) or (inputs(220));
    layer0_outputs(673) <= inputs(61);
    layer0_outputs(674) <= not(inputs(178)) or (inputs(26));
    layer0_outputs(675) <= not(inputs(49));
    layer0_outputs(676) <= (inputs(210)) and (inputs(250));
    layer0_outputs(677) <= not(inputs(134));
    layer0_outputs(678) <= not((inputs(92)) and (inputs(74)));
    layer0_outputs(679) <= not(inputs(112)) or (inputs(20));
    layer0_outputs(680) <= not((inputs(249)) or (inputs(45)));
    layer0_outputs(681) <= not((inputs(20)) xor (inputs(238)));
    layer0_outputs(682) <= not((inputs(87)) xor (inputs(224)));
    layer0_outputs(683) <= not(inputs(149));
    layer0_outputs(684) <= not(inputs(112));
    layer0_outputs(685) <= not(inputs(119));
    layer0_outputs(686) <= not((inputs(50)) xor (inputs(0)));
    layer0_outputs(687) <= not((inputs(96)) xor (inputs(67)));
    layer0_outputs(688) <= (inputs(67)) and not (inputs(1));
    layer0_outputs(689) <= inputs(104);
    layer0_outputs(690) <= not(inputs(72));
    layer0_outputs(691) <= not((inputs(188)) xor (inputs(225)));
    layer0_outputs(692) <= not(inputs(180));
    layer0_outputs(693) <= not(inputs(88));
    layer0_outputs(694) <= (inputs(127)) or (inputs(1));
    layer0_outputs(695) <= not((inputs(113)) xor (inputs(67)));
    layer0_outputs(696) <= inputs(182);
    layer0_outputs(697) <= inputs(227);
    layer0_outputs(698) <= not((inputs(224)) or (inputs(149)));
    layer0_outputs(699) <= inputs(202);
    layer0_outputs(700) <= (inputs(229)) and not (inputs(11));
    layer0_outputs(701) <= (inputs(238)) or (inputs(195));
    layer0_outputs(702) <= not(inputs(137));
    layer0_outputs(703) <= (inputs(177)) and (inputs(42));
    layer0_outputs(704) <= not(inputs(171)) or (inputs(27));
    layer0_outputs(705) <= (inputs(147)) and (inputs(127));
    layer0_outputs(706) <= not(inputs(162));
    layer0_outputs(707) <= (inputs(230)) and not (inputs(16));
    layer0_outputs(708) <= not(inputs(159));
    layer0_outputs(709) <= not((inputs(239)) or (inputs(56)));
    layer0_outputs(710) <= (inputs(39)) xor (inputs(139));
    layer0_outputs(711) <= not(inputs(134)) or (inputs(214));
    layer0_outputs(712) <= (inputs(118)) and not (inputs(161));
    layer0_outputs(713) <= not((inputs(181)) and (inputs(179)));
    layer0_outputs(714) <= '1';
    layer0_outputs(715) <= (inputs(33)) xor (inputs(3));
    layer0_outputs(716) <= '1';
    layer0_outputs(717) <= (inputs(58)) and (inputs(154));
    layer0_outputs(718) <= not(inputs(200)) or (inputs(78));
    layer0_outputs(719) <= not((inputs(190)) and (inputs(251)));
    layer0_outputs(720) <= not(inputs(104));
    layer0_outputs(721) <= not((inputs(61)) xor (inputs(158)));
    layer0_outputs(722) <= (inputs(51)) and not (inputs(241));
    layer0_outputs(723) <= '0';
    layer0_outputs(724) <= not(inputs(201)) or (inputs(20));
    layer0_outputs(725) <= inputs(74);
    layer0_outputs(726) <= (inputs(155)) or (inputs(207));
    layer0_outputs(727) <= (inputs(5)) or (inputs(137));
    layer0_outputs(728) <= inputs(8);
    layer0_outputs(729) <= (inputs(144)) or (inputs(201));
    layer0_outputs(730) <= inputs(96);
    layer0_outputs(731) <= (inputs(230)) or (inputs(105));
    layer0_outputs(732) <= not(inputs(188)) or (inputs(108));
    layer0_outputs(733) <= inputs(219);
    layer0_outputs(734) <= not(inputs(129));
    layer0_outputs(735) <= not((inputs(171)) xor (inputs(52)));
    layer0_outputs(736) <= '1';
    layer0_outputs(737) <= not((inputs(251)) or (inputs(90)));
    layer0_outputs(738) <= not(inputs(119));
    layer0_outputs(739) <= (inputs(47)) and not (inputs(226));
    layer0_outputs(740) <= (inputs(130)) and (inputs(21));
    layer0_outputs(741) <= not(inputs(196));
    layer0_outputs(742) <= (inputs(10)) and not (inputs(26));
    layer0_outputs(743) <= not((inputs(207)) xor (inputs(171)));
    layer0_outputs(744) <= not((inputs(42)) or (inputs(181)));
    layer0_outputs(745) <= not(inputs(242)) or (inputs(190));
    layer0_outputs(746) <= (inputs(179)) and not (inputs(13));
    layer0_outputs(747) <= not(inputs(116)) or (inputs(228));
    layer0_outputs(748) <= inputs(168);
    layer0_outputs(749) <= not((inputs(232)) xor (inputs(6)));
    layer0_outputs(750) <= inputs(57);
    layer0_outputs(751) <= (inputs(13)) or (inputs(18));
    layer0_outputs(752) <= not((inputs(35)) or (inputs(215)));
    layer0_outputs(753) <= (inputs(31)) or (inputs(103));
    layer0_outputs(754) <= (inputs(254)) or (inputs(50));
    layer0_outputs(755) <= not((inputs(10)) xor (inputs(132)));
    layer0_outputs(756) <= (inputs(44)) xor (inputs(9));
    layer0_outputs(757) <= not(inputs(0)) or (inputs(11));
    layer0_outputs(758) <= (inputs(248)) and (inputs(185));
    layer0_outputs(759) <= (inputs(20)) or (inputs(20));
    layer0_outputs(760) <= not((inputs(249)) or (inputs(218)));
    layer0_outputs(761) <= inputs(105);
    layer0_outputs(762) <= (inputs(77)) or (inputs(138));
    layer0_outputs(763) <= '0';
    layer0_outputs(764) <= not(inputs(143)) or (inputs(242));
    layer0_outputs(765) <= not((inputs(238)) xor (inputs(102)));
    layer0_outputs(766) <= not((inputs(218)) xor (inputs(45)));
    layer0_outputs(767) <= (inputs(216)) or (inputs(30));
    layer0_outputs(768) <= not((inputs(145)) xor (inputs(190)));
    layer0_outputs(769) <= not(inputs(216)) or (inputs(18));
    layer0_outputs(770) <= inputs(140);
    layer0_outputs(771) <= not((inputs(181)) or (inputs(128)));
    layer0_outputs(772) <= '0';
    layer0_outputs(773) <= (inputs(180)) xor (inputs(115));
    layer0_outputs(774) <= inputs(135);
    layer0_outputs(775) <= inputs(61);
    layer0_outputs(776) <= '1';
    layer0_outputs(777) <= not((inputs(128)) xor (inputs(78)));
    layer0_outputs(778) <= not((inputs(129)) or (inputs(137)));
    layer0_outputs(779) <= not((inputs(166)) or (inputs(194)));
    layer0_outputs(780) <= inputs(43);
    layer0_outputs(781) <= (inputs(116)) or (inputs(0));
    layer0_outputs(782) <= not((inputs(81)) xor (inputs(60)));
    layer0_outputs(783) <= not(inputs(118));
    layer0_outputs(784) <= (inputs(95)) and not (inputs(247));
    layer0_outputs(785) <= (inputs(63)) xor (inputs(56));
    layer0_outputs(786) <= not((inputs(206)) or (inputs(77)));
    layer0_outputs(787) <= (inputs(168)) and not (inputs(201));
    layer0_outputs(788) <= inputs(68);
    layer0_outputs(789) <= not((inputs(156)) xor (inputs(223)));
    layer0_outputs(790) <= not(inputs(24));
    layer0_outputs(791) <= (inputs(119)) or (inputs(146));
    layer0_outputs(792) <= (inputs(4)) xor (inputs(17));
    layer0_outputs(793) <= (inputs(230)) or (inputs(229));
    layer0_outputs(794) <= (inputs(154)) and not (inputs(3));
    layer0_outputs(795) <= not((inputs(239)) xor (inputs(163)));
    layer0_outputs(796) <= not((inputs(194)) or (inputs(235)));
    layer0_outputs(797) <= not(inputs(34));
    layer0_outputs(798) <= not(inputs(155));
    layer0_outputs(799) <= (inputs(173)) and not (inputs(31));
    layer0_outputs(800) <= not((inputs(119)) or (inputs(132)));
    layer0_outputs(801) <= not(inputs(55));
    layer0_outputs(802) <= (inputs(1)) xor (inputs(100));
    layer0_outputs(803) <= (inputs(232)) and not (inputs(188));
    layer0_outputs(804) <= not(inputs(28)) or (inputs(109));
    layer0_outputs(805) <= inputs(118);
    layer0_outputs(806) <= (inputs(61)) or (inputs(68));
    layer0_outputs(807) <= (inputs(60)) xor (inputs(93));
    layer0_outputs(808) <= (inputs(74)) and not (inputs(23));
    layer0_outputs(809) <= not(inputs(145)) or (inputs(208));
    layer0_outputs(810) <= (inputs(183)) and not (inputs(189));
    layer0_outputs(811) <= not(inputs(0)) or (inputs(185));
    layer0_outputs(812) <= (inputs(27)) xor (inputs(12));
    layer0_outputs(813) <= not((inputs(232)) xor (inputs(22)));
    layer0_outputs(814) <= not((inputs(219)) xor (inputs(199)));
    layer0_outputs(815) <= (inputs(184)) or (inputs(162));
    layer0_outputs(816) <= inputs(39);
    layer0_outputs(817) <= not(inputs(79)) or (inputs(5));
    layer0_outputs(818) <= not(inputs(106));
    layer0_outputs(819) <= inputs(119);
    layer0_outputs(820) <= inputs(229);
    layer0_outputs(821) <= not((inputs(255)) or (inputs(36)));
    layer0_outputs(822) <= (inputs(162)) xor (inputs(84));
    layer0_outputs(823) <= '0';
    layer0_outputs(824) <= (inputs(12)) or (inputs(221));
    layer0_outputs(825) <= not(inputs(250)) or (inputs(50));
    layer0_outputs(826) <= not(inputs(11)) or (inputs(17));
    layer0_outputs(827) <= not((inputs(96)) xor (inputs(80)));
    layer0_outputs(828) <= (inputs(201)) and not (inputs(162));
    layer0_outputs(829) <= not(inputs(46)) or (inputs(190));
    layer0_outputs(830) <= not(inputs(136)) or (inputs(21));
    layer0_outputs(831) <= not((inputs(255)) xor (inputs(52)));
    layer0_outputs(832) <= not((inputs(218)) xor (inputs(32)));
    layer0_outputs(833) <= not(inputs(156)) or (inputs(66));
    layer0_outputs(834) <= not((inputs(48)) xor (inputs(152)));
    layer0_outputs(835) <= (inputs(205)) or (inputs(26));
    layer0_outputs(836) <= not(inputs(121));
    layer0_outputs(837) <= (inputs(81)) xor (inputs(140));
    layer0_outputs(838) <= inputs(115);
    layer0_outputs(839) <= (inputs(153)) and not (inputs(40));
    layer0_outputs(840) <= (inputs(64)) or (inputs(251));
    layer0_outputs(841) <= not(inputs(245));
    layer0_outputs(842) <= (inputs(141)) or (inputs(237));
    layer0_outputs(843) <= '1';
    layer0_outputs(844) <= not((inputs(168)) xor (inputs(60)));
    layer0_outputs(845) <= not(inputs(212));
    layer0_outputs(846) <= (inputs(185)) or (inputs(206));
    layer0_outputs(847) <= (inputs(208)) and not (inputs(47));
    layer0_outputs(848) <= not(inputs(100));
    layer0_outputs(849) <= not((inputs(11)) xor (inputs(108)));
    layer0_outputs(850) <= (inputs(23)) and (inputs(241));
    layer0_outputs(851) <= not((inputs(168)) xor (inputs(215)));
    layer0_outputs(852) <= (inputs(98)) and (inputs(53));
    layer0_outputs(853) <= not(inputs(101));
    layer0_outputs(854) <= not(inputs(220)) or (inputs(160));
    layer0_outputs(855) <= '0';
    layer0_outputs(856) <= not(inputs(153)) or (inputs(180));
    layer0_outputs(857) <= (inputs(3)) and not (inputs(163));
    layer0_outputs(858) <= (inputs(215)) and not (inputs(44));
    layer0_outputs(859) <= '1';
    layer0_outputs(860) <= inputs(154);
    layer0_outputs(861) <= inputs(251);
    layer0_outputs(862) <= not((inputs(106)) or (inputs(153)));
    layer0_outputs(863) <= (inputs(36)) and (inputs(252));
    layer0_outputs(864) <= (inputs(228)) xor (inputs(161));
    layer0_outputs(865) <= (inputs(246)) and not (inputs(243));
    layer0_outputs(866) <= not(inputs(14)) or (inputs(114));
    layer0_outputs(867) <= not(inputs(220));
    layer0_outputs(868) <= (inputs(166)) or (inputs(141));
    layer0_outputs(869) <= not((inputs(249)) and (inputs(111)));
    layer0_outputs(870) <= not((inputs(99)) or (inputs(106)));
    layer0_outputs(871) <= (inputs(88)) and not (inputs(134));
    layer0_outputs(872) <= (inputs(167)) and not (inputs(244));
    layer0_outputs(873) <= not((inputs(160)) or (inputs(166)));
    layer0_outputs(874) <= not((inputs(162)) or (inputs(164)));
    layer0_outputs(875) <= inputs(155);
    layer0_outputs(876) <= (inputs(132)) and not (inputs(193));
    layer0_outputs(877) <= (inputs(73)) and not (inputs(127));
    layer0_outputs(878) <= not(inputs(204));
    layer0_outputs(879) <= inputs(25);
    layer0_outputs(880) <= not((inputs(205)) or (inputs(249)));
    layer0_outputs(881) <= '1';
    layer0_outputs(882) <= inputs(132);
    layer0_outputs(883) <= (inputs(192)) and not (inputs(160));
    layer0_outputs(884) <= not((inputs(60)) xor (inputs(236)));
    layer0_outputs(885) <= not(inputs(102)) or (inputs(195));
    layer0_outputs(886) <= (inputs(115)) and not (inputs(22));
    layer0_outputs(887) <= '0';
    layer0_outputs(888) <= inputs(39);
    layer0_outputs(889) <= not((inputs(128)) or (inputs(208)));
    layer0_outputs(890) <= inputs(65);
    layer0_outputs(891) <= not((inputs(90)) or (inputs(229)));
    layer0_outputs(892) <= not(inputs(36));
    layer0_outputs(893) <= not((inputs(58)) and (inputs(223)));
    layer0_outputs(894) <= not(inputs(124));
    layer0_outputs(895) <= not((inputs(234)) or (inputs(54)));
    layer0_outputs(896) <= not((inputs(60)) or (inputs(220)));
    layer0_outputs(897) <= inputs(12);
    layer0_outputs(898) <= not((inputs(70)) or (inputs(75)));
    layer0_outputs(899) <= inputs(47);
    layer0_outputs(900) <= (inputs(199)) and not (inputs(215));
    layer0_outputs(901) <= not((inputs(85)) xor (inputs(159)));
    layer0_outputs(902) <= (inputs(206)) xor (inputs(59));
    layer0_outputs(903) <= '0';
    layer0_outputs(904) <= (inputs(28)) and not (inputs(247));
    layer0_outputs(905) <= (inputs(230)) xor (inputs(29));
    layer0_outputs(906) <= not((inputs(232)) xor (inputs(168)));
    layer0_outputs(907) <= (inputs(60)) or (inputs(8));
    layer0_outputs(908) <= inputs(155);
    layer0_outputs(909) <= not((inputs(192)) xor (inputs(68)));
    layer0_outputs(910) <= not(inputs(152)) or (inputs(52));
    layer0_outputs(911) <= not(inputs(196));
    layer0_outputs(912) <= (inputs(25)) xor (inputs(219));
    layer0_outputs(913) <= not((inputs(226)) xor (inputs(84)));
    layer0_outputs(914) <= not(inputs(101));
    layer0_outputs(915) <= (inputs(125)) and not (inputs(13));
    layer0_outputs(916) <= (inputs(72)) and not (inputs(103));
    layer0_outputs(917) <= not(inputs(26)) or (inputs(250));
    layer0_outputs(918) <= not((inputs(255)) or (inputs(159)));
    layer0_outputs(919) <= not(inputs(121)) or (inputs(204));
    layer0_outputs(920) <= not((inputs(113)) or (inputs(246)));
    layer0_outputs(921) <= '1';
    layer0_outputs(922) <= not((inputs(104)) or (inputs(255)));
    layer0_outputs(923) <= (inputs(49)) or (inputs(121));
    layer0_outputs(924) <= not((inputs(255)) or (inputs(183)));
    layer0_outputs(925) <= inputs(67);
    layer0_outputs(926) <= inputs(56);
    layer0_outputs(927) <= (inputs(42)) or (inputs(197));
    layer0_outputs(928) <= not((inputs(164)) or (inputs(185)));
    layer0_outputs(929) <= inputs(197);
    layer0_outputs(930) <= not((inputs(197)) or (inputs(76)));
    layer0_outputs(931) <= (inputs(155)) and not (inputs(75));
    layer0_outputs(932) <= (inputs(23)) or (inputs(7));
    layer0_outputs(933) <= not((inputs(149)) xor (inputs(112)));
    layer0_outputs(934) <= (inputs(183)) and not (inputs(241));
    layer0_outputs(935) <= not(inputs(101)) or (inputs(244));
    layer0_outputs(936) <= (inputs(39)) and (inputs(185));
    layer0_outputs(937) <= (inputs(250)) and not (inputs(242));
    layer0_outputs(938) <= not(inputs(243));
    layer0_outputs(939) <= (inputs(243)) and not (inputs(53));
    layer0_outputs(940) <= (inputs(87)) or (inputs(235));
    layer0_outputs(941) <= not((inputs(217)) xor (inputs(168)));
    layer0_outputs(942) <= not(inputs(168));
    layer0_outputs(943) <= not((inputs(37)) and (inputs(227)));
    layer0_outputs(944) <= inputs(118);
    layer0_outputs(945) <= inputs(7);
    layer0_outputs(946) <= inputs(106);
    layer0_outputs(947) <= not(inputs(248)) or (inputs(36));
    layer0_outputs(948) <= not(inputs(60)) or (inputs(119));
    layer0_outputs(949) <= not(inputs(207)) or (inputs(207));
    layer0_outputs(950) <= (inputs(113)) xor (inputs(30));
    layer0_outputs(951) <= not((inputs(65)) xor (inputs(221)));
    layer0_outputs(952) <= (inputs(103)) or (inputs(139));
    layer0_outputs(953) <= '0';
    layer0_outputs(954) <= not(inputs(85));
    layer0_outputs(955) <= (inputs(222)) or (inputs(42));
    layer0_outputs(956) <= inputs(149);
    layer0_outputs(957) <= (inputs(254)) or (inputs(240));
    layer0_outputs(958) <= (inputs(148)) and not (inputs(254));
    layer0_outputs(959) <= (inputs(156)) and not (inputs(161));
    layer0_outputs(960) <= not(inputs(109)) or (inputs(227));
    layer0_outputs(961) <= (inputs(181)) and not (inputs(8));
    layer0_outputs(962) <= inputs(71);
    layer0_outputs(963) <= not((inputs(217)) or (inputs(228)));
    layer0_outputs(964) <= not(inputs(39));
    layer0_outputs(965) <= not(inputs(102)) or (inputs(65));
    layer0_outputs(966) <= not((inputs(141)) or (inputs(96)));
    layer0_outputs(967) <= inputs(202);
    layer0_outputs(968) <= (inputs(123)) and not (inputs(66));
    layer0_outputs(969) <= (inputs(219)) and (inputs(33));
    layer0_outputs(970) <= not(inputs(13)) or (inputs(37));
    layer0_outputs(971) <= '1';
    layer0_outputs(972) <= (inputs(79)) xor (inputs(165));
    layer0_outputs(973) <= (inputs(128)) and not (inputs(94));
    layer0_outputs(974) <= (inputs(161)) and not (inputs(231));
    layer0_outputs(975) <= inputs(164);
    layer0_outputs(976) <= (inputs(141)) and not (inputs(251));
    layer0_outputs(977) <= not(inputs(71));
    layer0_outputs(978) <= not(inputs(137)) or (inputs(158));
    layer0_outputs(979) <= not((inputs(104)) xor (inputs(20)));
    layer0_outputs(980) <= not(inputs(58)) or (inputs(114));
    layer0_outputs(981) <= not((inputs(84)) or (inputs(110)));
    layer0_outputs(982) <= (inputs(142)) and (inputs(112));
    layer0_outputs(983) <= not(inputs(117)) or (inputs(249));
    layer0_outputs(984) <= not(inputs(58));
    layer0_outputs(985) <= inputs(41);
    layer0_outputs(986) <= inputs(215);
    layer0_outputs(987) <= (inputs(83)) or (inputs(105));
    layer0_outputs(988) <= inputs(107);
    layer0_outputs(989) <= (inputs(246)) and (inputs(31));
    layer0_outputs(990) <= not(inputs(46));
    layer0_outputs(991) <= not((inputs(60)) or (inputs(76)));
    layer0_outputs(992) <= not((inputs(210)) or (inputs(142)));
    layer0_outputs(993) <= not((inputs(39)) or (inputs(158)));
    layer0_outputs(994) <= (inputs(55)) and not (inputs(244));
    layer0_outputs(995) <= (inputs(214)) xor (inputs(32));
    layer0_outputs(996) <= not((inputs(128)) xor (inputs(135)));
    layer0_outputs(997) <= (inputs(146)) and not (inputs(252));
    layer0_outputs(998) <= not(inputs(153)) or (inputs(245));
    layer0_outputs(999) <= (inputs(238)) and not (inputs(71));
    layer0_outputs(1000) <= inputs(118);
    layer0_outputs(1001) <= not((inputs(138)) xor (inputs(209)));
    layer0_outputs(1002) <= inputs(137);
    layer0_outputs(1003) <= (inputs(96)) xor (inputs(216));
    layer0_outputs(1004) <= not(inputs(198));
    layer0_outputs(1005) <= inputs(55);
    layer0_outputs(1006) <= inputs(89);
    layer0_outputs(1007) <= not((inputs(103)) or (inputs(94)));
    layer0_outputs(1008) <= not(inputs(127)) or (inputs(8));
    layer0_outputs(1009) <= not((inputs(31)) or (inputs(240)));
    layer0_outputs(1010) <= not((inputs(190)) xor (inputs(178)));
    layer0_outputs(1011) <= (inputs(72)) or (inputs(67));
    layer0_outputs(1012) <= not(inputs(243));
    layer0_outputs(1013) <= (inputs(197)) and not (inputs(210));
    layer0_outputs(1014) <= not(inputs(66));
    layer0_outputs(1015) <= not(inputs(145));
    layer0_outputs(1016) <= '0';
    layer0_outputs(1017) <= not(inputs(27));
    layer0_outputs(1018) <= not((inputs(120)) xor (inputs(129)));
    layer0_outputs(1019) <= not(inputs(103)) or (inputs(29));
    layer0_outputs(1020) <= not(inputs(55)) or (inputs(167));
    layer0_outputs(1021) <= (inputs(77)) or (inputs(40));
    layer0_outputs(1022) <= (inputs(58)) xor (inputs(11));
    layer0_outputs(1023) <= '1';
    layer0_outputs(1024) <= inputs(106);
    layer0_outputs(1025) <= inputs(100);
    layer0_outputs(1026) <= inputs(140);
    layer0_outputs(1027) <= not(inputs(93)) or (inputs(194));
    layer0_outputs(1028) <= inputs(119);
    layer0_outputs(1029) <= not((inputs(154)) or (inputs(8)));
    layer0_outputs(1030) <= not(inputs(150)) or (inputs(215));
    layer0_outputs(1031) <= (inputs(84)) and not (inputs(208));
    layer0_outputs(1032) <= (inputs(84)) or (inputs(180));
    layer0_outputs(1033) <= not((inputs(49)) xor (inputs(171)));
    layer0_outputs(1034) <= not(inputs(119));
    layer0_outputs(1035) <= (inputs(152)) and not (inputs(27));
    layer0_outputs(1036) <= (inputs(55)) or (inputs(54));
    layer0_outputs(1037) <= not(inputs(39));
    layer0_outputs(1038) <= inputs(172);
    layer0_outputs(1039) <= not((inputs(228)) or (inputs(154)));
    layer0_outputs(1040) <= (inputs(151)) xor (inputs(95));
    layer0_outputs(1041) <= (inputs(248)) xor (inputs(250));
    layer0_outputs(1042) <= (inputs(15)) xor (inputs(198));
    layer0_outputs(1043) <= not(inputs(73)) or (inputs(27));
    layer0_outputs(1044) <= (inputs(8)) xor (inputs(120));
    layer0_outputs(1045) <= '0';
    layer0_outputs(1046) <= not(inputs(136)) or (inputs(171));
    layer0_outputs(1047) <= not((inputs(179)) xor (inputs(24)));
    layer0_outputs(1048) <= not(inputs(221));
    layer0_outputs(1049) <= not((inputs(153)) xor (inputs(19)));
    layer0_outputs(1050) <= (inputs(141)) xor (inputs(206));
    layer0_outputs(1051) <= (inputs(115)) and not (inputs(242));
    layer0_outputs(1052) <= '1';
    layer0_outputs(1053) <= (inputs(125)) and not (inputs(210));
    layer0_outputs(1054) <= inputs(47);
    layer0_outputs(1055) <= not((inputs(141)) or (inputs(147)));
    layer0_outputs(1056) <= not(inputs(106)) or (inputs(195));
    layer0_outputs(1057) <= not(inputs(69)) or (inputs(8));
    layer0_outputs(1058) <= not((inputs(39)) or (inputs(123)));
    layer0_outputs(1059) <= not((inputs(254)) or (inputs(163)));
    layer0_outputs(1060) <= (inputs(106)) and not (inputs(177));
    layer0_outputs(1061) <= inputs(112);
    layer0_outputs(1062) <= (inputs(158)) and not (inputs(177));
    layer0_outputs(1063) <= inputs(121);
    layer0_outputs(1064) <= not((inputs(78)) xor (inputs(164)));
    layer0_outputs(1065) <= not(inputs(120)) or (inputs(202));
    layer0_outputs(1066) <= (inputs(67)) and not (inputs(191));
    layer0_outputs(1067) <= (inputs(73)) or (inputs(144));
    layer0_outputs(1068) <= inputs(112);
    layer0_outputs(1069) <= (inputs(165)) or (inputs(223));
    layer0_outputs(1070) <= not((inputs(195)) or (inputs(191)));
    layer0_outputs(1071) <= inputs(49);
    layer0_outputs(1072) <= not(inputs(119)) or (inputs(7));
    layer0_outputs(1073) <= not(inputs(197));
    layer0_outputs(1074) <= inputs(249);
    layer0_outputs(1075) <= not((inputs(65)) and (inputs(61)));
    layer0_outputs(1076) <= not(inputs(112)) or (inputs(210));
    layer0_outputs(1077) <= inputs(200);
    layer0_outputs(1078) <= not(inputs(100));
    layer0_outputs(1079) <= (inputs(139)) and not (inputs(194));
    layer0_outputs(1080) <= inputs(104);
    layer0_outputs(1081) <= (inputs(109)) or (inputs(109));
    layer0_outputs(1082) <= (inputs(3)) or (inputs(237));
    layer0_outputs(1083) <= not(inputs(210)) or (inputs(66));
    layer0_outputs(1084) <= (inputs(9)) or (inputs(63));
    layer0_outputs(1085) <= (inputs(152)) xor (inputs(248));
    layer0_outputs(1086) <= (inputs(158)) and (inputs(104));
    layer0_outputs(1087) <= (inputs(9)) xor (inputs(186));
    layer0_outputs(1088) <= not((inputs(32)) xor (inputs(214)));
    layer0_outputs(1089) <= (inputs(229)) and not (inputs(84));
    layer0_outputs(1090) <= not(inputs(53));
    layer0_outputs(1091) <= (inputs(103)) or (inputs(118));
    layer0_outputs(1092) <= (inputs(222)) xor (inputs(91));
    layer0_outputs(1093) <= (inputs(52)) or (inputs(199));
    layer0_outputs(1094) <= '1';
    layer0_outputs(1095) <= (inputs(237)) xor (inputs(166));
    layer0_outputs(1096) <= not((inputs(90)) or (inputs(228)));
    layer0_outputs(1097) <= inputs(103);
    layer0_outputs(1098) <= not(inputs(187));
    layer0_outputs(1099) <= inputs(96);
    layer0_outputs(1100) <= inputs(241);
    layer0_outputs(1101) <= not((inputs(60)) xor (inputs(78)));
    layer0_outputs(1102) <= not(inputs(238)) or (inputs(14));
    layer0_outputs(1103) <= (inputs(18)) xor (inputs(163));
    layer0_outputs(1104) <= (inputs(96)) or (inputs(212));
    layer0_outputs(1105) <= (inputs(196)) and (inputs(42));
    layer0_outputs(1106) <= (inputs(117)) and not (inputs(52));
    layer0_outputs(1107) <= (inputs(30)) xor (inputs(148));
    layer0_outputs(1108) <= not(inputs(74));
    layer0_outputs(1109) <= (inputs(63)) and not (inputs(110));
    layer0_outputs(1110) <= not(inputs(236));
    layer0_outputs(1111) <= (inputs(21)) or (inputs(5));
    layer0_outputs(1112) <= (inputs(94)) or (inputs(140));
    layer0_outputs(1113) <= not((inputs(243)) or (inputs(110)));
    layer0_outputs(1114) <= not((inputs(17)) xor (inputs(159)));
    layer0_outputs(1115) <= inputs(186);
    layer0_outputs(1116) <= (inputs(98)) or (inputs(59));
    layer0_outputs(1117) <= not((inputs(40)) xor (inputs(8)));
    layer0_outputs(1118) <= inputs(59);
    layer0_outputs(1119) <= not(inputs(226));
    layer0_outputs(1120) <= (inputs(243)) and not (inputs(53));
    layer0_outputs(1121) <= not((inputs(211)) or (inputs(114)));
    layer0_outputs(1122) <= not((inputs(48)) or (inputs(140)));
    layer0_outputs(1123) <= not((inputs(144)) and (inputs(110)));
    layer0_outputs(1124) <= '1';
    layer0_outputs(1125) <= (inputs(238)) or (inputs(40));
    layer0_outputs(1126) <= inputs(111);
    layer0_outputs(1127) <= '0';
    layer0_outputs(1128) <= inputs(90);
    layer0_outputs(1129) <= (inputs(153)) or (inputs(119));
    layer0_outputs(1130) <= not((inputs(31)) or (inputs(206)));
    layer0_outputs(1131) <= inputs(221);
    layer0_outputs(1132) <= not((inputs(160)) or (inputs(167)));
    layer0_outputs(1133) <= not(inputs(195)) or (inputs(29));
    layer0_outputs(1134) <= not(inputs(121)) or (inputs(50));
    layer0_outputs(1135) <= (inputs(11)) and not (inputs(50));
    layer0_outputs(1136) <= inputs(94);
    layer0_outputs(1137) <= (inputs(160)) or (inputs(90));
    layer0_outputs(1138) <= not((inputs(161)) or (inputs(197)));
    layer0_outputs(1139) <= '1';
    layer0_outputs(1140) <= (inputs(23)) and not (inputs(202));
    layer0_outputs(1141) <= not(inputs(29)) or (inputs(224));
    layer0_outputs(1142) <= not((inputs(172)) and (inputs(132)));
    layer0_outputs(1143) <= (inputs(119)) and not (inputs(235));
    layer0_outputs(1144) <= not(inputs(111));
    layer0_outputs(1145) <= not((inputs(188)) or (inputs(6)));
    layer0_outputs(1146) <= inputs(160);
    layer0_outputs(1147) <= inputs(94);
    layer0_outputs(1148) <= (inputs(180)) and not (inputs(226));
    layer0_outputs(1149) <= not((inputs(226)) xor (inputs(158)));
    layer0_outputs(1150) <= '1';
    layer0_outputs(1151) <= not((inputs(14)) or (inputs(51)));
    layer0_outputs(1152) <= not((inputs(172)) or (inputs(171)));
    layer0_outputs(1153) <= (inputs(110)) xor (inputs(193));
    layer0_outputs(1154) <= inputs(209);
    layer0_outputs(1155) <= inputs(136);
    layer0_outputs(1156) <= (inputs(176)) and not (inputs(245));
    layer0_outputs(1157) <= (inputs(204)) or (inputs(194));
    layer0_outputs(1158) <= not(inputs(117));
    layer0_outputs(1159) <= '0';
    layer0_outputs(1160) <= (inputs(214)) or (inputs(13));
    layer0_outputs(1161) <= not(inputs(63)) or (inputs(43));
    layer0_outputs(1162) <= not(inputs(148));
    layer0_outputs(1163) <= (inputs(136)) and not (inputs(50));
    layer0_outputs(1164) <= inputs(88);
    layer0_outputs(1165) <= not(inputs(187)) or (inputs(169));
    layer0_outputs(1166) <= not((inputs(27)) xor (inputs(247)));
    layer0_outputs(1167) <= inputs(158);
    layer0_outputs(1168) <= (inputs(115)) or (inputs(124));
    layer0_outputs(1169) <= inputs(254);
    layer0_outputs(1170) <= '1';
    layer0_outputs(1171) <= not((inputs(143)) and (inputs(43)));
    layer0_outputs(1172) <= inputs(77);
    layer0_outputs(1173) <= not(inputs(18)) or (inputs(97));
    layer0_outputs(1174) <= (inputs(147)) xor (inputs(32));
    layer0_outputs(1175) <= not((inputs(243)) xor (inputs(115)));
    layer0_outputs(1176) <= (inputs(239)) or (inputs(205));
    layer0_outputs(1177) <= not(inputs(158));
    layer0_outputs(1178) <= (inputs(241)) xor (inputs(217));
    layer0_outputs(1179) <= (inputs(241)) xor (inputs(69));
    layer0_outputs(1180) <= (inputs(199)) and not (inputs(189));
    layer0_outputs(1181) <= not((inputs(201)) or (inputs(128)));
    layer0_outputs(1182) <= not(inputs(44)) or (inputs(110));
    layer0_outputs(1183) <= (inputs(127)) and not (inputs(52));
    layer0_outputs(1184) <= not(inputs(69));
    layer0_outputs(1185) <= (inputs(189)) or (inputs(36));
    layer0_outputs(1186) <= (inputs(198)) and not (inputs(43));
    layer0_outputs(1187) <= not(inputs(162));
    layer0_outputs(1188) <= not((inputs(44)) xor (inputs(190)));
    layer0_outputs(1189) <= not((inputs(38)) or (inputs(118)));
    layer0_outputs(1190) <= not(inputs(137));
    layer0_outputs(1191) <= not((inputs(166)) xor (inputs(97)));
    layer0_outputs(1192) <= (inputs(117)) and not (inputs(65));
    layer0_outputs(1193) <= not(inputs(79)) or (inputs(238));
    layer0_outputs(1194) <= not(inputs(153));
    layer0_outputs(1195) <= inputs(70);
    layer0_outputs(1196) <= inputs(141);
    layer0_outputs(1197) <= inputs(42);
    layer0_outputs(1198) <= not(inputs(87));
    layer0_outputs(1199) <= (inputs(82)) and not (inputs(62));
    layer0_outputs(1200) <= (inputs(250)) xor (inputs(68));
    layer0_outputs(1201) <= not(inputs(166)) or (inputs(209));
    layer0_outputs(1202) <= '0';
    layer0_outputs(1203) <= not(inputs(42));
    layer0_outputs(1204) <= not((inputs(158)) xor (inputs(81)));
    layer0_outputs(1205) <= (inputs(146)) or (inputs(94));
    layer0_outputs(1206) <= (inputs(153)) and not (inputs(103));
    layer0_outputs(1207) <= not(inputs(117));
    layer0_outputs(1208) <= not(inputs(168)) or (inputs(79));
    layer0_outputs(1209) <= not(inputs(202));
    layer0_outputs(1210) <= not(inputs(154));
    layer0_outputs(1211) <= (inputs(159)) or (inputs(151));
    layer0_outputs(1212) <= (inputs(182)) xor (inputs(195));
    layer0_outputs(1213) <= '1';
    layer0_outputs(1214) <= (inputs(90)) and not (inputs(26));
    layer0_outputs(1215) <= not(inputs(187)) or (inputs(146));
    layer0_outputs(1216) <= (inputs(240)) xor (inputs(237));
    layer0_outputs(1217) <= inputs(72);
    layer0_outputs(1218) <= (inputs(183)) xor (inputs(89));
    layer0_outputs(1219) <= not(inputs(247));
    layer0_outputs(1220) <= (inputs(7)) and not (inputs(239));
    layer0_outputs(1221) <= inputs(156);
    layer0_outputs(1222) <= (inputs(137)) and not (inputs(188));
    layer0_outputs(1223) <= inputs(103);
    layer0_outputs(1224) <= not(inputs(59)) or (inputs(210));
    layer0_outputs(1225) <= not(inputs(77)) or (inputs(248));
    layer0_outputs(1226) <= not(inputs(245)) or (inputs(95));
    layer0_outputs(1227) <= '0';
    layer0_outputs(1228) <= not(inputs(56));
    layer0_outputs(1229) <= inputs(17);
    layer0_outputs(1230) <= (inputs(73)) and not (inputs(11));
    layer0_outputs(1231) <= not(inputs(237)) or (inputs(67));
    layer0_outputs(1232) <= '0';
    layer0_outputs(1233) <= not((inputs(44)) or (inputs(20)));
    layer0_outputs(1234) <= (inputs(70)) or (inputs(208));
    layer0_outputs(1235) <= not(inputs(26)) or (inputs(243));
    layer0_outputs(1236) <= not((inputs(90)) xor (inputs(253)));
    layer0_outputs(1237) <= not((inputs(234)) or (inputs(109)));
    layer0_outputs(1238) <= not((inputs(25)) xor (inputs(122)));
    layer0_outputs(1239) <= not((inputs(31)) or (inputs(24)));
    layer0_outputs(1240) <= not(inputs(229));
    layer0_outputs(1241) <= (inputs(7)) and not (inputs(145));
    layer0_outputs(1242) <= inputs(159);
    layer0_outputs(1243) <= not((inputs(201)) xor (inputs(222)));
    layer0_outputs(1244) <= not((inputs(251)) xor (inputs(25)));
    layer0_outputs(1245) <= inputs(149);
    layer0_outputs(1246) <= (inputs(197)) or (inputs(189));
    layer0_outputs(1247) <= (inputs(26)) and not (inputs(245));
    layer0_outputs(1248) <= (inputs(113)) and not (inputs(240));
    layer0_outputs(1249) <= inputs(82);
    layer0_outputs(1250) <= inputs(253);
    layer0_outputs(1251) <= inputs(167);
    layer0_outputs(1252) <= not(inputs(90));
    layer0_outputs(1253) <= not(inputs(136));
    layer0_outputs(1254) <= inputs(121);
    layer0_outputs(1255) <= inputs(144);
    layer0_outputs(1256) <= not((inputs(144)) xor (inputs(53)));
    layer0_outputs(1257) <= not((inputs(36)) xor (inputs(162)));
    layer0_outputs(1258) <= not(inputs(181));
    layer0_outputs(1259) <= not(inputs(150));
    layer0_outputs(1260) <= inputs(87);
    layer0_outputs(1261) <= not(inputs(88)) or (inputs(148));
    layer0_outputs(1262) <= not((inputs(72)) or (inputs(178)));
    layer0_outputs(1263) <= (inputs(72)) and not (inputs(53));
    layer0_outputs(1264) <= inputs(222);
    layer0_outputs(1265) <= not((inputs(218)) xor (inputs(94)));
    layer0_outputs(1266) <= (inputs(110)) or (inputs(58));
    layer0_outputs(1267) <= (inputs(63)) and not (inputs(239));
    layer0_outputs(1268) <= not(inputs(68));
    layer0_outputs(1269) <= '0';
    layer0_outputs(1270) <= (inputs(238)) and not (inputs(177));
    layer0_outputs(1271) <= '1';
    layer0_outputs(1272) <= (inputs(11)) xor (inputs(253));
    layer0_outputs(1273) <= (inputs(153)) and not (inputs(119));
    layer0_outputs(1274) <= (inputs(34)) and not (inputs(118));
    layer0_outputs(1275) <= not((inputs(187)) or (inputs(215)));
    layer0_outputs(1276) <= (inputs(154)) or (inputs(36));
    layer0_outputs(1277) <= not(inputs(119)) or (inputs(131));
    layer0_outputs(1278) <= not(inputs(113));
    layer0_outputs(1279) <= not((inputs(224)) xor (inputs(102)));
    layer0_outputs(1280) <= not(inputs(128));
    layer0_outputs(1281) <= inputs(182);
    layer0_outputs(1282) <= not(inputs(136)) or (inputs(29));
    layer0_outputs(1283) <= not((inputs(144)) xor (inputs(188)));
    layer0_outputs(1284) <= (inputs(99)) or (inputs(217));
    layer0_outputs(1285) <= not((inputs(82)) or (inputs(104)));
    layer0_outputs(1286) <= not(inputs(165));
    layer0_outputs(1287) <= (inputs(108)) or (inputs(25));
    layer0_outputs(1288) <= inputs(244);
    layer0_outputs(1289) <= not(inputs(159));
    layer0_outputs(1290) <= not((inputs(72)) and (inputs(67)));
    layer0_outputs(1291) <= not((inputs(246)) xor (inputs(74)));
    layer0_outputs(1292) <= (inputs(217)) and (inputs(251));
    layer0_outputs(1293) <= (inputs(122)) and not (inputs(251));
    layer0_outputs(1294) <= not(inputs(133));
    layer0_outputs(1295) <= (inputs(38)) and not (inputs(204));
    layer0_outputs(1296) <= not(inputs(171));
    layer0_outputs(1297) <= not((inputs(188)) or (inputs(194)));
    layer0_outputs(1298) <= not(inputs(224)) or (inputs(191));
    layer0_outputs(1299) <= (inputs(131)) and not (inputs(49));
    layer0_outputs(1300) <= (inputs(153)) or (inputs(116));
    layer0_outputs(1301) <= not((inputs(169)) xor (inputs(128)));
    layer0_outputs(1302) <= inputs(230);
    layer0_outputs(1303) <= not(inputs(198)) or (inputs(45));
    layer0_outputs(1304) <= (inputs(124)) and not (inputs(145));
    layer0_outputs(1305) <= not(inputs(91));
    layer0_outputs(1306) <= (inputs(231)) xor (inputs(241));
    layer0_outputs(1307) <= not(inputs(101)) or (inputs(126));
    layer0_outputs(1308) <= inputs(71);
    layer0_outputs(1309) <= not(inputs(194));
    layer0_outputs(1310) <= (inputs(43)) and not (inputs(35));
    layer0_outputs(1311) <= not((inputs(129)) xor (inputs(106)));
    layer0_outputs(1312) <= (inputs(166)) or (inputs(193));
    layer0_outputs(1313) <= not(inputs(209));
    layer0_outputs(1314) <= inputs(90);
    layer0_outputs(1315) <= not(inputs(216));
    layer0_outputs(1316) <= not((inputs(80)) and (inputs(13)));
    layer0_outputs(1317) <= (inputs(210)) or (inputs(212));
    layer0_outputs(1318) <= (inputs(0)) and not (inputs(111));
    layer0_outputs(1319) <= not(inputs(197)) or (inputs(208));
    layer0_outputs(1320) <= not((inputs(99)) xor (inputs(241)));
    layer0_outputs(1321) <= inputs(59);
    layer0_outputs(1322) <= not((inputs(97)) or (inputs(168)));
    layer0_outputs(1323) <= not(inputs(122));
    layer0_outputs(1324) <= inputs(152);
    layer0_outputs(1325) <= not(inputs(167)) or (inputs(108));
    layer0_outputs(1326) <= (inputs(60)) and not (inputs(14));
    layer0_outputs(1327) <= '1';
    layer0_outputs(1328) <= not((inputs(87)) xor (inputs(85)));
    layer0_outputs(1329) <= not((inputs(147)) or (inputs(80)));
    layer0_outputs(1330) <= (inputs(169)) and not (inputs(78));
    layer0_outputs(1331) <= not(inputs(251)) or (inputs(145));
    layer0_outputs(1332) <= inputs(151);
    layer0_outputs(1333) <= (inputs(118)) and not (inputs(163));
    layer0_outputs(1334) <= inputs(165);
    layer0_outputs(1335) <= (inputs(189)) and not (inputs(22));
    layer0_outputs(1336) <= (inputs(52)) or (inputs(4));
    layer0_outputs(1337) <= (inputs(81)) and (inputs(176));
    layer0_outputs(1338) <= inputs(197);
    layer0_outputs(1339) <= not((inputs(239)) or (inputs(34)));
    layer0_outputs(1340) <= inputs(113);
    layer0_outputs(1341) <= not(inputs(149));
    layer0_outputs(1342) <= (inputs(205)) and not (inputs(66));
    layer0_outputs(1343) <= inputs(159);
    layer0_outputs(1344) <= not(inputs(160));
    layer0_outputs(1345) <= (inputs(165)) and not (inputs(238));
    layer0_outputs(1346) <= inputs(69);
    layer0_outputs(1347) <= not(inputs(101));
    layer0_outputs(1348) <= not(inputs(104));
    layer0_outputs(1349) <= inputs(166);
    layer0_outputs(1350) <= not((inputs(21)) and (inputs(10)));
    layer0_outputs(1351) <= '1';
    layer0_outputs(1352) <= not(inputs(165)) or (inputs(234));
    layer0_outputs(1353) <= not((inputs(137)) xor (inputs(63)));
    layer0_outputs(1354) <= (inputs(75)) xor (inputs(242));
    layer0_outputs(1355) <= not((inputs(4)) or (inputs(147)));
    layer0_outputs(1356) <= not(inputs(99));
    layer0_outputs(1357) <= (inputs(234)) and not (inputs(48));
    layer0_outputs(1358) <= (inputs(131)) or (inputs(136));
    layer0_outputs(1359) <= not((inputs(130)) xor (inputs(81)));
    layer0_outputs(1360) <= not(inputs(110)) or (inputs(7));
    layer0_outputs(1361) <= not((inputs(44)) xor (inputs(181)));
    layer0_outputs(1362) <= not((inputs(221)) xor (inputs(154)));
    layer0_outputs(1363) <= not((inputs(54)) or (inputs(172)));
    layer0_outputs(1364) <= not(inputs(7)) or (inputs(212));
    layer0_outputs(1365) <= inputs(39);
    layer0_outputs(1366) <= (inputs(221)) and not (inputs(85));
    layer0_outputs(1367) <= not(inputs(73)) or (inputs(4));
    layer0_outputs(1368) <= (inputs(100)) and not (inputs(194));
    layer0_outputs(1369) <= (inputs(149)) xor (inputs(175));
    layer0_outputs(1370) <= (inputs(15)) and not (inputs(234));
    layer0_outputs(1371) <= not((inputs(39)) or (inputs(162)));
    layer0_outputs(1372) <= (inputs(19)) or (inputs(123));
    layer0_outputs(1373) <= not(inputs(125)) or (inputs(245));
    layer0_outputs(1374) <= not((inputs(24)) or (inputs(210)));
    layer0_outputs(1375) <= inputs(81);
    layer0_outputs(1376) <= (inputs(44)) and (inputs(118));
    layer0_outputs(1377) <= not((inputs(179)) xor (inputs(238)));
    layer0_outputs(1378) <= (inputs(108)) xor (inputs(205));
    layer0_outputs(1379) <= '1';
    layer0_outputs(1380) <= (inputs(154)) xor (inputs(106));
    layer0_outputs(1381) <= not(inputs(51)) or (inputs(220));
    layer0_outputs(1382) <= not((inputs(158)) xor (inputs(249)));
    layer0_outputs(1383) <= (inputs(126)) and not (inputs(167));
    layer0_outputs(1384) <= (inputs(218)) or (inputs(79));
    layer0_outputs(1385) <= not(inputs(254));
    layer0_outputs(1386) <= not(inputs(211)) or (inputs(46));
    layer0_outputs(1387) <= (inputs(52)) xor (inputs(149));
    layer0_outputs(1388) <= inputs(34);
    layer0_outputs(1389) <= not(inputs(213)) or (inputs(125));
    layer0_outputs(1390) <= not(inputs(19));
    layer0_outputs(1391) <= not((inputs(194)) or (inputs(15)));
    layer0_outputs(1392) <= not((inputs(21)) or (inputs(131)));
    layer0_outputs(1393) <= inputs(137);
    layer0_outputs(1394) <= not(inputs(231)) or (inputs(163));
    layer0_outputs(1395) <= not(inputs(21));
    layer0_outputs(1396) <= (inputs(247)) and (inputs(175));
    layer0_outputs(1397) <= not((inputs(252)) or (inputs(225)));
    layer0_outputs(1398) <= not((inputs(248)) xor (inputs(57)));
    layer0_outputs(1399) <= not((inputs(56)) or (inputs(231)));
    layer0_outputs(1400) <= inputs(179);
    layer0_outputs(1401) <= not(inputs(152));
    layer0_outputs(1402) <= inputs(189);
    layer0_outputs(1403) <= '1';
    layer0_outputs(1404) <= (inputs(253)) or (inputs(91));
    layer0_outputs(1405) <= (inputs(16)) and (inputs(130));
    layer0_outputs(1406) <= not((inputs(246)) xor (inputs(41)));
    layer0_outputs(1407) <= (inputs(82)) and not (inputs(115));
    layer0_outputs(1408) <= (inputs(28)) and not (inputs(112));
    layer0_outputs(1409) <= (inputs(193)) xor (inputs(208));
    layer0_outputs(1410) <= inputs(182);
    layer0_outputs(1411) <= not((inputs(92)) or (inputs(126)));
    layer0_outputs(1412) <= not((inputs(2)) or (inputs(59)));
    layer0_outputs(1413) <= '1';
    layer0_outputs(1414) <= (inputs(216)) or (inputs(128));
    layer0_outputs(1415) <= inputs(186);
    layer0_outputs(1416) <= '1';
    layer0_outputs(1417) <= not((inputs(71)) xor (inputs(95)));
    layer0_outputs(1418) <= (inputs(174)) and not (inputs(244));
    layer0_outputs(1419) <= (inputs(172)) and not (inputs(14));
    layer0_outputs(1420) <= (inputs(198)) or (inputs(213));
    layer0_outputs(1421) <= (inputs(186)) or (inputs(243));
    layer0_outputs(1422) <= not((inputs(229)) xor (inputs(210)));
    layer0_outputs(1423) <= not(inputs(129));
    layer0_outputs(1424) <= not(inputs(42));
    layer0_outputs(1425) <= not(inputs(198));
    layer0_outputs(1426) <= not((inputs(247)) or (inputs(182)));
    layer0_outputs(1427) <= not(inputs(216)) or (inputs(26));
    layer0_outputs(1428) <= (inputs(89)) and not (inputs(9));
    layer0_outputs(1429) <= (inputs(87)) and not (inputs(236));
    layer0_outputs(1430) <= inputs(54);
    layer0_outputs(1431) <= not(inputs(132));
    layer0_outputs(1432) <= inputs(203);
    layer0_outputs(1433) <= (inputs(120)) and not (inputs(82));
    layer0_outputs(1434) <= (inputs(141)) and not (inputs(6));
    layer0_outputs(1435) <= not(inputs(102)) or (inputs(210));
    layer0_outputs(1436) <= not((inputs(126)) xor (inputs(176)));
    layer0_outputs(1437) <= (inputs(75)) and (inputs(16));
    layer0_outputs(1438) <= not((inputs(110)) or (inputs(237)));
    layer0_outputs(1439) <= (inputs(138)) or (inputs(122));
    layer0_outputs(1440) <= (inputs(104)) or (inputs(234));
    layer0_outputs(1441) <= inputs(10);
    layer0_outputs(1442) <= not((inputs(117)) xor (inputs(236)));
    layer0_outputs(1443) <= not(inputs(131));
    layer0_outputs(1444) <= (inputs(145)) or (inputs(8));
    layer0_outputs(1445) <= not((inputs(169)) and (inputs(172)));
    layer0_outputs(1446) <= (inputs(42)) or (inputs(206));
    layer0_outputs(1447) <= inputs(182);
    layer0_outputs(1448) <= inputs(72);
    layer0_outputs(1449) <= '0';
    layer0_outputs(1450) <= (inputs(133)) and not (inputs(16));
    layer0_outputs(1451) <= (inputs(192)) xor (inputs(74));
    layer0_outputs(1452) <= inputs(33);
    layer0_outputs(1453) <= (inputs(4)) or (inputs(44));
    layer0_outputs(1454) <= '0';
    layer0_outputs(1455) <= (inputs(191)) or (inputs(52));
    layer0_outputs(1456) <= not((inputs(162)) xor (inputs(168)));
    layer0_outputs(1457) <= not(inputs(223));
    layer0_outputs(1458) <= (inputs(196)) or (inputs(188));
    layer0_outputs(1459) <= not(inputs(47)) or (inputs(234));
    layer0_outputs(1460) <= inputs(82);
    layer0_outputs(1461) <= (inputs(131)) xor (inputs(68));
    layer0_outputs(1462) <= (inputs(247)) xor (inputs(83));
    layer0_outputs(1463) <= (inputs(230)) and not (inputs(93));
    layer0_outputs(1464) <= not((inputs(215)) or (inputs(73)));
    layer0_outputs(1465) <= (inputs(214)) and not (inputs(147));
    layer0_outputs(1466) <= (inputs(209)) xor (inputs(26));
    layer0_outputs(1467) <= (inputs(172)) or (inputs(69));
    layer0_outputs(1468) <= '1';
    layer0_outputs(1469) <= (inputs(195)) and not (inputs(81));
    layer0_outputs(1470) <= not(inputs(54));
    layer0_outputs(1471) <= (inputs(180)) or (inputs(125));
    layer0_outputs(1472) <= inputs(124);
    layer0_outputs(1473) <= (inputs(145)) xor (inputs(109));
    layer0_outputs(1474) <= (inputs(7)) xor (inputs(116));
    layer0_outputs(1475) <= (inputs(79)) or (inputs(71));
    layer0_outputs(1476) <= inputs(138);
    layer0_outputs(1477) <= (inputs(236)) and not (inputs(206));
    layer0_outputs(1478) <= not(inputs(124));
    layer0_outputs(1479) <= (inputs(229)) or (inputs(53));
    layer0_outputs(1480) <= inputs(135);
    layer0_outputs(1481) <= not((inputs(222)) xor (inputs(126)));
    layer0_outputs(1482) <= (inputs(9)) or (inputs(166));
    layer0_outputs(1483) <= (inputs(124)) or (inputs(135));
    layer0_outputs(1484) <= (inputs(96)) xor (inputs(118));
    layer0_outputs(1485) <= not(inputs(108));
    layer0_outputs(1486) <= (inputs(186)) or (inputs(186));
    layer0_outputs(1487) <= (inputs(114)) or (inputs(250));
    layer0_outputs(1488) <= (inputs(131)) and not (inputs(31));
    layer0_outputs(1489) <= not((inputs(170)) or (inputs(228)));
    layer0_outputs(1490) <= not((inputs(40)) or (inputs(57)));
    layer0_outputs(1491) <= not(inputs(202)) or (inputs(225));
    layer0_outputs(1492) <= inputs(138);
    layer0_outputs(1493) <= inputs(246);
    layer0_outputs(1494) <= (inputs(177)) and (inputs(209));
    layer0_outputs(1495) <= not(inputs(220)) or (inputs(135));
    layer0_outputs(1496) <= (inputs(142)) or (inputs(91));
    layer0_outputs(1497) <= inputs(120);
    layer0_outputs(1498) <= not(inputs(136)) or (inputs(44));
    layer0_outputs(1499) <= not(inputs(87)) or (inputs(29));
    layer0_outputs(1500) <= (inputs(147)) xor (inputs(9));
    layer0_outputs(1501) <= not(inputs(216)) or (inputs(225));
    layer0_outputs(1502) <= not((inputs(72)) xor (inputs(211)));
    layer0_outputs(1503) <= (inputs(129)) xor (inputs(187));
    layer0_outputs(1504) <= inputs(215);
    layer0_outputs(1505) <= inputs(99);
    layer0_outputs(1506) <= (inputs(5)) and not (inputs(72));
    layer0_outputs(1507) <= not(inputs(151));
    layer0_outputs(1508) <= not(inputs(105));
    layer0_outputs(1509) <= inputs(50);
    layer0_outputs(1510) <= not((inputs(174)) or (inputs(164)));
    layer0_outputs(1511) <= inputs(118);
    layer0_outputs(1512) <= (inputs(47)) and not (inputs(216));
    layer0_outputs(1513) <= not((inputs(177)) xor (inputs(231)));
    layer0_outputs(1514) <= not(inputs(59)) or (inputs(255));
    layer0_outputs(1515) <= not((inputs(89)) xor (inputs(31)));
    layer0_outputs(1516) <= '0';
    layer0_outputs(1517) <= inputs(100);
    layer0_outputs(1518) <= not(inputs(143));
    layer0_outputs(1519) <= not((inputs(6)) xor (inputs(71)));
    layer0_outputs(1520) <= inputs(119);
    layer0_outputs(1521) <= not((inputs(239)) xor (inputs(11)));
    layer0_outputs(1522) <= not(inputs(181)) or (inputs(33));
    layer0_outputs(1523) <= not(inputs(148)) or (inputs(223));
    layer0_outputs(1524) <= not(inputs(116));
    layer0_outputs(1525) <= '1';
    layer0_outputs(1526) <= (inputs(86)) and (inputs(201));
    layer0_outputs(1527) <= not(inputs(22));
    layer0_outputs(1528) <= (inputs(31)) xor (inputs(96));
    layer0_outputs(1529) <= not((inputs(85)) and (inputs(143)));
    layer0_outputs(1530) <= inputs(107);
    layer0_outputs(1531) <= not(inputs(53)) or (inputs(157));
    layer0_outputs(1532) <= inputs(90);
    layer0_outputs(1533) <= not(inputs(155)) or (inputs(179));
    layer0_outputs(1534) <= '0';
    layer0_outputs(1535) <= (inputs(174)) and not (inputs(100));
    layer0_outputs(1536) <= (inputs(143)) xor (inputs(25));
    layer0_outputs(1537) <= inputs(172);
    layer0_outputs(1538) <= not(inputs(20));
    layer0_outputs(1539) <= not(inputs(190));
    layer0_outputs(1540) <= not((inputs(171)) xor (inputs(62)));
    layer0_outputs(1541) <= not((inputs(114)) or (inputs(232)));
    layer0_outputs(1542) <= (inputs(102)) and not (inputs(146));
    layer0_outputs(1543) <= not((inputs(129)) or (inputs(103)));
    layer0_outputs(1544) <= not(inputs(100)) or (inputs(141));
    layer0_outputs(1545) <= (inputs(191)) xor (inputs(70));
    layer0_outputs(1546) <= not((inputs(128)) or (inputs(109)));
    layer0_outputs(1547) <= not(inputs(27));
    layer0_outputs(1548) <= (inputs(105)) and not (inputs(9));
    layer0_outputs(1549) <= not((inputs(216)) or (inputs(185)));
    layer0_outputs(1550) <= not((inputs(183)) xor (inputs(214)));
    layer0_outputs(1551) <= not(inputs(104));
    layer0_outputs(1552) <= (inputs(207)) xor (inputs(143));
    layer0_outputs(1553) <= not(inputs(82));
    layer0_outputs(1554) <= not((inputs(25)) or (inputs(53)));
    layer0_outputs(1555) <= not(inputs(102));
    layer0_outputs(1556) <= not((inputs(96)) or (inputs(50)));
    layer0_outputs(1557) <= not((inputs(161)) xor (inputs(124)));
    layer0_outputs(1558) <= not((inputs(48)) xor (inputs(115)));
    layer0_outputs(1559) <= not(inputs(183));
    layer0_outputs(1560) <= not((inputs(144)) and (inputs(5)));
    layer0_outputs(1561) <= not((inputs(145)) or (inputs(150)));
    layer0_outputs(1562) <= inputs(187);
    layer0_outputs(1563) <= not(inputs(56)) or (inputs(100));
    layer0_outputs(1564) <= not((inputs(62)) or (inputs(33)));
    layer0_outputs(1565) <= not(inputs(183)) or (inputs(134));
    layer0_outputs(1566) <= not((inputs(83)) or (inputs(150)));
    layer0_outputs(1567) <= (inputs(106)) and not (inputs(249));
    layer0_outputs(1568) <= not(inputs(211)) or (inputs(114));
    layer0_outputs(1569) <= inputs(156);
    layer0_outputs(1570) <= not((inputs(179)) or (inputs(6)));
    layer0_outputs(1571) <= (inputs(162)) or (inputs(229));
    layer0_outputs(1572) <= '0';
    layer0_outputs(1573) <= not((inputs(222)) and (inputs(43)));
    layer0_outputs(1574) <= (inputs(177)) xor (inputs(73));
    layer0_outputs(1575) <= (inputs(131)) or (inputs(14));
    layer0_outputs(1576) <= (inputs(226)) or (inputs(197));
    layer0_outputs(1577) <= inputs(69);
    layer0_outputs(1578) <= (inputs(197)) or (inputs(195));
    layer0_outputs(1579) <= (inputs(167)) and not (inputs(132));
    layer0_outputs(1580) <= not((inputs(56)) or (inputs(125)));
    layer0_outputs(1581) <= (inputs(238)) and not (inputs(144));
    layer0_outputs(1582) <= inputs(91);
    layer0_outputs(1583) <= (inputs(74)) xor (inputs(126));
    layer0_outputs(1584) <= not(inputs(196));
    layer0_outputs(1585) <= (inputs(104)) or (inputs(232));
    layer0_outputs(1586) <= '1';
    layer0_outputs(1587) <= not((inputs(90)) or (inputs(146)));
    layer0_outputs(1588) <= not(inputs(116)) or (inputs(128));
    layer0_outputs(1589) <= (inputs(32)) xor (inputs(40));
    layer0_outputs(1590) <= (inputs(120)) and not (inputs(132));
    layer0_outputs(1591) <= (inputs(4)) and not (inputs(33));
    layer0_outputs(1592) <= not(inputs(169));
    layer0_outputs(1593) <= inputs(111);
    layer0_outputs(1594) <= (inputs(209)) and (inputs(18));
    layer0_outputs(1595) <= not(inputs(41));
    layer0_outputs(1596) <= not((inputs(69)) or (inputs(24)));
    layer0_outputs(1597) <= (inputs(132)) or (inputs(26));
    layer0_outputs(1598) <= '1';
    layer0_outputs(1599) <= (inputs(249)) and not (inputs(23));
    layer0_outputs(1600) <= not((inputs(93)) xor (inputs(16)));
    layer0_outputs(1601) <= not((inputs(46)) xor (inputs(171)));
    layer0_outputs(1602) <= not(inputs(182));
    layer0_outputs(1603) <= not(inputs(151)) or (inputs(52));
    layer0_outputs(1604) <= (inputs(117)) xor (inputs(97));
    layer0_outputs(1605) <= (inputs(30)) xor (inputs(74));
    layer0_outputs(1606) <= not((inputs(233)) or (inputs(109)));
    layer0_outputs(1607) <= not(inputs(228));
    layer0_outputs(1608) <= not(inputs(149));
    layer0_outputs(1609) <= (inputs(178)) and not (inputs(189));
    layer0_outputs(1610) <= not((inputs(10)) xor (inputs(63)));
    layer0_outputs(1611) <= (inputs(117)) and not (inputs(57));
    layer0_outputs(1612) <= (inputs(136)) or (inputs(233));
    layer0_outputs(1613) <= (inputs(109)) xor (inputs(17));
    layer0_outputs(1614) <= not(inputs(165));
    layer0_outputs(1615) <= not(inputs(180)) or (inputs(39));
    layer0_outputs(1616) <= not((inputs(5)) and (inputs(211)));
    layer0_outputs(1617) <= (inputs(218)) and not (inputs(171));
    layer0_outputs(1618) <= not((inputs(178)) or (inputs(72)));
    layer0_outputs(1619) <= inputs(206);
    layer0_outputs(1620) <= not((inputs(237)) and (inputs(30)));
    layer0_outputs(1621) <= not(inputs(28)) or (inputs(208));
    layer0_outputs(1622) <= (inputs(133)) and not (inputs(58));
    layer0_outputs(1623) <= not(inputs(0));
    layer0_outputs(1624) <= (inputs(196)) xor (inputs(254));
    layer0_outputs(1625) <= inputs(53);
    layer0_outputs(1626) <= not(inputs(46));
    layer0_outputs(1627) <= (inputs(216)) and not (inputs(208));
    layer0_outputs(1628) <= not((inputs(132)) xor (inputs(12)));
    layer0_outputs(1629) <= not(inputs(213));
    layer0_outputs(1630) <= not(inputs(119));
    layer0_outputs(1631) <= (inputs(193)) and (inputs(96));
    layer0_outputs(1632) <= (inputs(82)) and not (inputs(157));
    layer0_outputs(1633) <= not((inputs(78)) or (inputs(229)));
    layer0_outputs(1634) <= (inputs(131)) and not (inputs(119));
    layer0_outputs(1635) <= (inputs(232)) and not (inputs(126));
    layer0_outputs(1636) <= not(inputs(132));
    layer0_outputs(1637) <= not(inputs(92)) or (inputs(161));
    layer0_outputs(1638) <= (inputs(87)) xor (inputs(130));
    layer0_outputs(1639) <= (inputs(151)) and not (inputs(229));
    layer0_outputs(1640) <= (inputs(194)) xor (inputs(110));
    layer0_outputs(1641) <= (inputs(101)) and not (inputs(178));
    layer0_outputs(1642) <= not(inputs(180)) or (inputs(159));
    layer0_outputs(1643) <= inputs(184);
    layer0_outputs(1644) <= (inputs(75)) and not (inputs(153));
    layer0_outputs(1645) <= not(inputs(240));
    layer0_outputs(1646) <= not((inputs(235)) or (inputs(200)));
    layer0_outputs(1647) <= (inputs(4)) and not (inputs(37));
    layer0_outputs(1648) <= (inputs(141)) and not (inputs(212));
    layer0_outputs(1649) <= (inputs(104)) or (inputs(163));
    layer0_outputs(1650) <= not((inputs(34)) or (inputs(120)));
    layer0_outputs(1651) <= (inputs(86)) or (inputs(140));
    layer0_outputs(1652) <= not(inputs(248));
    layer0_outputs(1653) <= inputs(138);
    layer0_outputs(1654) <= not((inputs(39)) xor (inputs(29)));
    layer0_outputs(1655) <= (inputs(178)) and not (inputs(63));
    layer0_outputs(1656) <= (inputs(149)) or (inputs(252));
    layer0_outputs(1657) <= (inputs(1)) or (inputs(41));
    layer0_outputs(1658) <= not(inputs(205));
    layer0_outputs(1659) <= inputs(214);
    layer0_outputs(1660) <= inputs(130);
    layer0_outputs(1661) <= not((inputs(19)) or (inputs(104)));
    layer0_outputs(1662) <= (inputs(139)) xor (inputs(44));
    layer0_outputs(1663) <= (inputs(131)) and not (inputs(252));
    layer0_outputs(1664) <= inputs(34);
    layer0_outputs(1665) <= (inputs(124)) or (inputs(74));
    layer0_outputs(1666) <= (inputs(164)) or (inputs(44));
    layer0_outputs(1667) <= (inputs(209)) and not (inputs(85));
    layer0_outputs(1668) <= not(inputs(155)) or (inputs(0));
    layer0_outputs(1669) <= '1';
    layer0_outputs(1670) <= (inputs(55)) and not (inputs(22));
    layer0_outputs(1671) <= (inputs(181)) xor (inputs(158));
    layer0_outputs(1672) <= not(inputs(215)) or (inputs(245));
    layer0_outputs(1673) <= not((inputs(23)) xor (inputs(144)));
    layer0_outputs(1674) <= (inputs(135)) and not (inputs(65));
    layer0_outputs(1675) <= not(inputs(107));
    layer0_outputs(1676) <= not(inputs(212)) or (inputs(14));
    layer0_outputs(1677) <= '1';
    layer0_outputs(1678) <= not((inputs(85)) or (inputs(142)));
    layer0_outputs(1679) <= not(inputs(126));
    layer0_outputs(1680) <= not(inputs(73)) or (inputs(243));
    layer0_outputs(1681) <= not((inputs(69)) and (inputs(87)));
    layer0_outputs(1682) <= not((inputs(181)) or (inputs(53)));
    layer0_outputs(1683) <= not(inputs(234)) or (inputs(74));
    layer0_outputs(1684) <= not(inputs(135)) or (inputs(38));
    layer0_outputs(1685) <= (inputs(59)) xor (inputs(103));
    layer0_outputs(1686) <= (inputs(122)) and (inputs(73));
    layer0_outputs(1687) <= not(inputs(68));
    layer0_outputs(1688) <= not((inputs(123)) or (inputs(153)));
    layer0_outputs(1689) <= inputs(142);
    layer0_outputs(1690) <= (inputs(229)) xor (inputs(25));
    layer0_outputs(1691) <= (inputs(217)) and not (inputs(80));
    layer0_outputs(1692) <= (inputs(107)) and not (inputs(0));
    layer0_outputs(1693) <= not((inputs(173)) or (inputs(239)));
    layer0_outputs(1694) <= '0';
    layer0_outputs(1695) <= (inputs(183)) xor (inputs(16));
    layer0_outputs(1696) <= (inputs(125)) and not (inputs(242));
    layer0_outputs(1697) <= (inputs(239)) or (inputs(209));
    layer0_outputs(1698) <= not((inputs(127)) xor (inputs(221)));
    layer0_outputs(1699) <= not(inputs(134));
    layer0_outputs(1700) <= not((inputs(56)) xor (inputs(63)));
    layer0_outputs(1701) <= '1';
    layer0_outputs(1702) <= not(inputs(91));
    layer0_outputs(1703) <= not((inputs(139)) or (inputs(50)));
    layer0_outputs(1704) <= (inputs(157)) and not (inputs(129));
    layer0_outputs(1705) <= '0';
    layer0_outputs(1706) <= not((inputs(26)) or (inputs(214)));
    layer0_outputs(1707) <= (inputs(43)) and not (inputs(62));
    layer0_outputs(1708) <= (inputs(200)) or (inputs(230));
    layer0_outputs(1709) <= not((inputs(25)) or (inputs(107)));
    layer0_outputs(1710) <= not(inputs(179));
    layer0_outputs(1711) <= (inputs(234)) and not (inputs(94));
    layer0_outputs(1712) <= not(inputs(37));
    layer0_outputs(1713) <= not(inputs(255)) or (inputs(255));
    layer0_outputs(1714) <= inputs(76);
    layer0_outputs(1715) <= not((inputs(244)) xor (inputs(238)));
    layer0_outputs(1716) <= not((inputs(182)) or (inputs(21)));
    layer0_outputs(1717) <= inputs(133);
    layer0_outputs(1718) <= not(inputs(205)) or (inputs(18));
    layer0_outputs(1719) <= '0';
    layer0_outputs(1720) <= not(inputs(39));
    layer0_outputs(1721) <= inputs(167);
    layer0_outputs(1722) <= not((inputs(41)) or (inputs(140)));
    layer0_outputs(1723) <= (inputs(218)) or (inputs(235));
    layer0_outputs(1724) <= '1';
    layer0_outputs(1725) <= inputs(94);
    layer0_outputs(1726) <= not(inputs(103)) or (inputs(2));
    layer0_outputs(1727) <= (inputs(138)) xor (inputs(246));
    layer0_outputs(1728) <= inputs(191);
    layer0_outputs(1729) <= not((inputs(111)) or (inputs(179)));
    layer0_outputs(1730) <= not((inputs(6)) xor (inputs(124)));
    layer0_outputs(1731) <= not((inputs(255)) or (inputs(97)));
    layer0_outputs(1732) <= not(inputs(213));
    layer0_outputs(1733) <= inputs(42);
    layer0_outputs(1734) <= not(inputs(102)) or (inputs(192));
    layer0_outputs(1735) <= (inputs(120)) and not (inputs(239));
    layer0_outputs(1736) <= (inputs(242)) or (inputs(78));
    layer0_outputs(1737) <= '0';
    layer0_outputs(1738) <= (inputs(180)) and not (inputs(248));
    layer0_outputs(1739) <= not(inputs(173));
    layer0_outputs(1740) <= (inputs(100)) and not (inputs(27));
    layer0_outputs(1741) <= (inputs(62)) and not (inputs(65));
    layer0_outputs(1742) <= (inputs(121)) and not (inputs(190));
    layer0_outputs(1743) <= (inputs(46)) and not (inputs(89));
    layer0_outputs(1744) <= not(inputs(85)) or (inputs(32));
    layer0_outputs(1745) <= not(inputs(69)) or (inputs(43));
    layer0_outputs(1746) <= not(inputs(179)) or (inputs(142));
    layer0_outputs(1747) <= not(inputs(249)) or (inputs(47));
    layer0_outputs(1748) <= inputs(203);
    layer0_outputs(1749) <= (inputs(47)) and (inputs(244));
    layer0_outputs(1750) <= (inputs(110)) and not (inputs(96));
    layer0_outputs(1751) <= not((inputs(74)) or (inputs(13)));
    layer0_outputs(1752) <= not((inputs(203)) or (inputs(23)));
    layer0_outputs(1753) <= not(inputs(61)) or (inputs(174));
    layer0_outputs(1754) <= (inputs(83)) xor (inputs(32));
    layer0_outputs(1755) <= inputs(154);
    layer0_outputs(1756) <= (inputs(49)) or (inputs(191));
    layer0_outputs(1757) <= not(inputs(118)) or (inputs(190));
    layer0_outputs(1758) <= inputs(85);
    layer0_outputs(1759) <= not((inputs(104)) xor (inputs(253)));
    layer0_outputs(1760) <= (inputs(150)) and not (inputs(93));
    layer0_outputs(1761) <= (inputs(39)) or (inputs(54));
    layer0_outputs(1762) <= (inputs(228)) or (inputs(105));
    layer0_outputs(1763) <= inputs(137);
    layer0_outputs(1764) <= (inputs(188)) and not (inputs(129));
    layer0_outputs(1765) <= not(inputs(27)) or (inputs(208));
    layer0_outputs(1766) <= (inputs(34)) or (inputs(190));
    layer0_outputs(1767) <= not((inputs(252)) xor (inputs(222)));
    layer0_outputs(1768) <= not(inputs(254)) or (inputs(51));
    layer0_outputs(1769) <= not((inputs(10)) xor (inputs(22)));
    layer0_outputs(1770) <= not((inputs(121)) or (inputs(85)));
    layer0_outputs(1771) <= (inputs(23)) and not (inputs(227));
    layer0_outputs(1772) <= (inputs(175)) and (inputs(70));
    layer0_outputs(1773) <= (inputs(201)) and not (inputs(131));
    layer0_outputs(1774) <= not(inputs(157)) or (inputs(128));
    layer0_outputs(1775) <= (inputs(68)) or (inputs(54));
    layer0_outputs(1776) <= not((inputs(6)) xor (inputs(208)));
    layer0_outputs(1777) <= (inputs(127)) or (inputs(23));
    layer0_outputs(1778) <= '0';
    layer0_outputs(1779) <= not(inputs(163));
    layer0_outputs(1780) <= inputs(9);
    layer0_outputs(1781) <= not(inputs(181)) or (inputs(208));
    layer0_outputs(1782) <= not(inputs(23));
    layer0_outputs(1783) <= (inputs(61)) and (inputs(15));
    layer0_outputs(1784) <= not((inputs(80)) xor (inputs(155)));
    layer0_outputs(1785) <= not(inputs(182));
    layer0_outputs(1786) <= inputs(151);
    layer0_outputs(1787) <= inputs(135);
    layer0_outputs(1788) <= not((inputs(87)) xor (inputs(5)));
    layer0_outputs(1789) <= not((inputs(62)) or (inputs(220)));
    layer0_outputs(1790) <= not(inputs(212));
    layer0_outputs(1791) <= not((inputs(236)) or (inputs(30)));
    layer0_outputs(1792) <= not((inputs(42)) or (inputs(172)));
    layer0_outputs(1793) <= inputs(206);
    layer0_outputs(1794) <= not(inputs(220)) or (inputs(161));
    layer0_outputs(1795) <= (inputs(6)) and not (inputs(184));
    layer0_outputs(1796) <= not(inputs(106));
    layer0_outputs(1797) <= (inputs(18)) xor (inputs(32));
    layer0_outputs(1798) <= (inputs(121)) and not (inputs(53));
    layer0_outputs(1799) <= not(inputs(239));
    layer0_outputs(1800) <= inputs(157);
    layer0_outputs(1801) <= not(inputs(138)) or (inputs(19));
    layer0_outputs(1802) <= (inputs(13)) and not (inputs(62));
    layer0_outputs(1803) <= not((inputs(16)) xor (inputs(68)));
    layer0_outputs(1804) <= (inputs(233)) xor (inputs(19));
    layer0_outputs(1805) <= not((inputs(132)) xor (inputs(12)));
    layer0_outputs(1806) <= (inputs(54)) or (inputs(170));
    layer0_outputs(1807) <= not(inputs(101)) or (inputs(226));
    layer0_outputs(1808) <= (inputs(87)) and not (inputs(156));
    layer0_outputs(1809) <= (inputs(30)) and not (inputs(187));
    layer0_outputs(1810) <= not((inputs(184)) or (inputs(232)));
    layer0_outputs(1811) <= (inputs(202)) xor (inputs(218));
    layer0_outputs(1812) <= not(inputs(91));
    layer0_outputs(1813) <= not((inputs(255)) and (inputs(46)));
    layer0_outputs(1814) <= not(inputs(85));
    layer0_outputs(1815) <= (inputs(58)) and not (inputs(252));
    layer0_outputs(1816) <= not(inputs(157));
    layer0_outputs(1817) <= (inputs(137)) and not (inputs(204));
    layer0_outputs(1818) <= (inputs(169)) and not (inputs(47));
    layer0_outputs(1819) <= not((inputs(152)) or (inputs(126)));
    layer0_outputs(1820) <= (inputs(196)) and not (inputs(232));
    layer0_outputs(1821) <= inputs(39);
    layer0_outputs(1822) <= not(inputs(210)) or (inputs(35));
    layer0_outputs(1823) <= inputs(3);
    layer0_outputs(1824) <= (inputs(219)) or (inputs(163));
    layer0_outputs(1825) <= not(inputs(171)) or (inputs(208));
    layer0_outputs(1826) <= (inputs(83)) or (inputs(98));
    layer0_outputs(1827) <= (inputs(170)) and not (inputs(159));
    layer0_outputs(1828) <= inputs(255);
    layer0_outputs(1829) <= inputs(64);
    layer0_outputs(1830) <= inputs(194);
    layer0_outputs(1831) <= (inputs(175)) xor (inputs(163));
    layer0_outputs(1832) <= '1';
    layer0_outputs(1833) <= not(inputs(168));
    layer0_outputs(1834) <= (inputs(28)) or (inputs(1));
    layer0_outputs(1835) <= (inputs(78)) or (inputs(209));
    layer0_outputs(1836) <= not(inputs(251));
    layer0_outputs(1837) <= not(inputs(185)) or (inputs(145));
    layer0_outputs(1838) <= not(inputs(219));
    layer0_outputs(1839) <= not((inputs(113)) or (inputs(97)));
    layer0_outputs(1840) <= not((inputs(244)) xor (inputs(109)));
    layer0_outputs(1841) <= (inputs(218)) or (inputs(55));
    layer0_outputs(1842) <= not(inputs(221)) or (inputs(9));
    layer0_outputs(1843) <= not(inputs(187)) or (inputs(125));
    layer0_outputs(1844) <= not((inputs(170)) xor (inputs(204)));
    layer0_outputs(1845) <= inputs(172);
    layer0_outputs(1846) <= (inputs(155)) and not (inputs(249));
    layer0_outputs(1847) <= not((inputs(212)) xor (inputs(56)));
    layer0_outputs(1848) <= (inputs(63)) and not (inputs(91));
    layer0_outputs(1849) <= not(inputs(54)) or (inputs(115));
    layer0_outputs(1850) <= not((inputs(90)) or (inputs(206)));
    layer0_outputs(1851) <= '1';
    layer0_outputs(1852) <= not(inputs(102)) or (inputs(207));
    layer0_outputs(1853) <= not(inputs(254)) or (inputs(45));
    layer0_outputs(1854) <= not((inputs(250)) and (inputs(84)));
    layer0_outputs(1855) <= not(inputs(88)) or (inputs(126));
    layer0_outputs(1856) <= (inputs(76)) or (inputs(200));
    layer0_outputs(1857) <= not((inputs(161)) or (inputs(67)));
    layer0_outputs(1858) <= not((inputs(114)) xor (inputs(145)));
    layer0_outputs(1859) <= (inputs(156)) xor (inputs(78));
    layer0_outputs(1860) <= not(inputs(230));
    layer0_outputs(1861) <= not((inputs(151)) or (inputs(216)));
    layer0_outputs(1862) <= not(inputs(82));
    layer0_outputs(1863) <= (inputs(26)) and (inputs(129));
    layer0_outputs(1864) <= '0';
    layer0_outputs(1865) <= (inputs(87)) and not (inputs(178));
    layer0_outputs(1866) <= inputs(72);
    layer0_outputs(1867) <= not(inputs(60));
    layer0_outputs(1868) <= not(inputs(67));
    layer0_outputs(1869) <= (inputs(65)) or (inputs(234));
    layer0_outputs(1870) <= inputs(42);
    layer0_outputs(1871) <= not(inputs(184)) or (inputs(73));
    layer0_outputs(1872) <= not((inputs(134)) xor (inputs(162)));
    layer0_outputs(1873) <= (inputs(184)) xor (inputs(45));
    layer0_outputs(1874) <= (inputs(129)) or (inputs(165));
    layer0_outputs(1875) <= not(inputs(2));
    layer0_outputs(1876) <= '1';
    layer0_outputs(1877) <= (inputs(119)) or (inputs(234));
    layer0_outputs(1878) <= not(inputs(163));
    layer0_outputs(1879) <= not(inputs(92));
    layer0_outputs(1880) <= not((inputs(4)) xor (inputs(105)));
    layer0_outputs(1881) <= not(inputs(89));
    layer0_outputs(1882) <= not((inputs(180)) or (inputs(36)));
    layer0_outputs(1883) <= not(inputs(60));
    layer0_outputs(1884) <= (inputs(86)) or (inputs(229));
    layer0_outputs(1885) <= (inputs(40)) and not (inputs(93));
    layer0_outputs(1886) <= not((inputs(159)) and (inputs(191)));
    layer0_outputs(1887) <= (inputs(220)) or (inputs(132));
    layer0_outputs(1888) <= (inputs(130)) or (inputs(223));
    layer0_outputs(1889) <= not(inputs(182)) or (inputs(205));
    layer0_outputs(1890) <= not(inputs(23));
    layer0_outputs(1891) <= not((inputs(32)) xor (inputs(19)));
    layer0_outputs(1892) <= not((inputs(180)) or (inputs(239)));
    layer0_outputs(1893) <= not(inputs(138));
    layer0_outputs(1894) <= not(inputs(231));
    layer0_outputs(1895) <= (inputs(210)) and not (inputs(237));
    layer0_outputs(1896) <= inputs(144);
    layer0_outputs(1897) <= (inputs(10)) xor (inputs(98));
    layer0_outputs(1898) <= not(inputs(140));
    layer0_outputs(1899) <= not(inputs(45)) or (inputs(174));
    layer0_outputs(1900) <= not((inputs(185)) or (inputs(134)));
    layer0_outputs(1901) <= not(inputs(149));
    layer0_outputs(1902) <= inputs(180);
    layer0_outputs(1903) <= (inputs(80)) xor (inputs(186));
    layer0_outputs(1904) <= not(inputs(32));
    layer0_outputs(1905) <= not((inputs(22)) or (inputs(29)));
    layer0_outputs(1906) <= '0';
    layer0_outputs(1907) <= not((inputs(94)) xor (inputs(18)));
    layer0_outputs(1908) <= (inputs(74)) and not (inputs(236));
    layer0_outputs(1909) <= (inputs(128)) and not (inputs(241));
    layer0_outputs(1910) <= (inputs(39)) and not (inputs(27));
    layer0_outputs(1911) <= not(inputs(52));
    layer0_outputs(1912) <= (inputs(117)) and not (inputs(97));
    layer0_outputs(1913) <= not((inputs(37)) xor (inputs(154)));
    layer0_outputs(1914) <= not(inputs(99));
    layer0_outputs(1915) <= inputs(108);
    layer0_outputs(1916) <= not((inputs(60)) or (inputs(59)));
    layer0_outputs(1917) <= not(inputs(175));
    layer0_outputs(1918) <= not(inputs(88)) or (inputs(170));
    layer0_outputs(1919) <= not((inputs(241)) xor (inputs(167)));
    layer0_outputs(1920) <= (inputs(66)) or (inputs(227));
    layer0_outputs(1921) <= (inputs(78)) and not (inputs(97));
    layer0_outputs(1922) <= inputs(106);
    layer0_outputs(1923) <= (inputs(203)) and not (inputs(97));
    layer0_outputs(1924) <= (inputs(151)) and not (inputs(175));
    layer0_outputs(1925) <= (inputs(84)) xor (inputs(188));
    layer0_outputs(1926) <= not((inputs(220)) or (inputs(247)));
    layer0_outputs(1927) <= not((inputs(178)) or (inputs(69)));
    layer0_outputs(1928) <= inputs(92);
    layer0_outputs(1929) <= not(inputs(86));
    layer0_outputs(1930) <= not(inputs(87)) or (inputs(162));
    layer0_outputs(1931) <= not(inputs(209)) or (inputs(17));
    layer0_outputs(1932) <= not((inputs(172)) or (inputs(9)));
    layer0_outputs(1933) <= not(inputs(53)) or (inputs(129));
    layer0_outputs(1934) <= not((inputs(134)) or (inputs(156)));
    layer0_outputs(1935) <= not((inputs(34)) xor (inputs(179)));
    layer0_outputs(1936) <= inputs(120);
    layer0_outputs(1937) <= not((inputs(76)) or (inputs(160)));
    layer0_outputs(1938) <= (inputs(15)) and not (inputs(28));
    layer0_outputs(1939) <= inputs(210);
    layer0_outputs(1940) <= inputs(55);
    layer0_outputs(1941) <= not((inputs(239)) xor (inputs(5)));
    layer0_outputs(1942) <= not((inputs(101)) xor (inputs(237)));
    layer0_outputs(1943) <= not(inputs(181));
    layer0_outputs(1944) <= (inputs(5)) xor (inputs(208));
    layer0_outputs(1945) <= not(inputs(6)) or (inputs(227));
    layer0_outputs(1946) <= not((inputs(155)) or (inputs(179)));
    layer0_outputs(1947) <= not((inputs(199)) xor (inputs(191)));
    layer0_outputs(1948) <= (inputs(46)) xor (inputs(67));
    layer0_outputs(1949) <= not((inputs(210)) and (inputs(21)));
    layer0_outputs(1950) <= not(inputs(171));
    layer0_outputs(1951) <= (inputs(222)) or (inputs(252));
    layer0_outputs(1952) <= not(inputs(232)) or (inputs(202));
    layer0_outputs(1953) <= (inputs(167)) and not (inputs(18));
    layer0_outputs(1954) <= not(inputs(133)) or (inputs(228));
    layer0_outputs(1955) <= inputs(189);
    layer0_outputs(1956) <= not(inputs(95)) or (inputs(194));
    layer0_outputs(1957) <= not((inputs(15)) and (inputs(199)));
    layer0_outputs(1958) <= not(inputs(214));
    layer0_outputs(1959) <= inputs(201);
    layer0_outputs(1960) <= (inputs(153)) xor (inputs(5));
    layer0_outputs(1961) <= (inputs(123)) and not (inputs(36));
    layer0_outputs(1962) <= '1';
    layer0_outputs(1963) <= not((inputs(147)) or (inputs(122)));
    layer0_outputs(1964) <= not((inputs(4)) and (inputs(31)));
    layer0_outputs(1965) <= not((inputs(228)) or (inputs(70)));
    layer0_outputs(1966) <= not(inputs(25));
    layer0_outputs(1967) <= '1';
    layer0_outputs(1968) <= not(inputs(148)) or (inputs(193));
    layer0_outputs(1969) <= not((inputs(245)) and (inputs(79)));
    layer0_outputs(1970) <= (inputs(218)) and not (inputs(174));
    layer0_outputs(1971) <= not((inputs(87)) xor (inputs(145)));
    layer0_outputs(1972) <= (inputs(33)) xor (inputs(106));
    layer0_outputs(1973) <= inputs(183);
    layer0_outputs(1974) <= (inputs(25)) and not (inputs(93));
    layer0_outputs(1975) <= not(inputs(186)) or (inputs(99));
    layer0_outputs(1976) <= not((inputs(77)) or (inputs(94)));
    layer0_outputs(1977) <= not((inputs(16)) or (inputs(144)));
    layer0_outputs(1978) <= (inputs(63)) or (inputs(231));
    layer0_outputs(1979) <= (inputs(11)) or (inputs(81));
    layer0_outputs(1980) <= not((inputs(125)) or (inputs(47)));
    layer0_outputs(1981) <= inputs(140);
    layer0_outputs(1982) <= not((inputs(194)) or (inputs(157)));
    layer0_outputs(1983) <= inputs(77);
    layer0_outputs(1984) <= not((inputs(125)) xor (inputs(139)));
    layer0_outputs(1985) <= not(inputs(193));
    layer0_outputs(1986) <= (inputs(22)) and (inputs(35));
    layer0_outputs(1987) <= (inputs(153)) and not (inputs(18));
    layer0_outputs(1988) <= not(inputs(111));
    layer0_outputs(1989) <= (inputs(49)) and (inputs(44));
    layer0_outputs(1990) <= not(inputs(95));
    layer0_outputs(1991) <= not(inputs(255));
    layer0_outputs(1992) <= not(inputs(136));
    layer0_outputs(1993) <= not(inputs(239));
    layer0_outputs(1994) <= not((inputs(252)) xor (inputs(148)));
    layer0_outputs(1995) <= (inputs(252)) or (inputs(89));
    layer0_outputs(1996) <= not(inputs(87)) or (inputs(43));
    layer0_outputs(1997) <= (inputs(42)) xor (inputs(229));
    layer0_outputs(1998) <= not((inputs(65)) or (inputs(148)));
    layer0_outputs(1999) <= (inputs(82)) xor (inputs(255));
    layer0_outputs(2000) <= (inputs(182)) xor (inputs(41));
    layer0_outputs(2001) <= (inputs(216)) and not (inputs(49));
    layer0_outputs(2002) <= inputs(166);
    layer0_outputs(2003) <= not(inputs(81)) or (inputs(24));
    layer0_outputs(2004) <= not(inputs(104)) or (inputs(67));
    layer0_outputs(2005) <= not(inputs(167));
    layer0_outputs(2006) <= (inputs(196)) and not (inputs(253));
    layer0_outputs(2007) <= not(inputs(253));
    layer0_outputs(2008) <= not(inputs(239)) or (inputs(216));
    layer0_outputs(2009) <= (inputs(38)) or (inputs(239));
    layer0_outputs(2010) <= inputs(100);
    layer0_outputs(2011) <= (inputs(227)) and not (inputs(161));
    layer0_outputs(2012) <= inputs(153);
    layer0_outputs(2013) <= inputs(152);
    layer0_outputs(2014) <= not(inputs(216)) or (inputs(111));
    layer0_outputs(2015) <= inputs(203);
    layer0_outputs(2016) <= not(inputs(186));
    layer0_outputs(2017) <= not((inputs(163)) or (inputs(187)));
    layer0_outputs(2018) <= not((inputs(153)) or (inputs(25)));
    layer0_outputs(2019) <= not(inputs(38)) or (inputs(13));
    layer0_outputs(2020) <= (inputs(91)) or (inputs(238));
    layer0_outputs(2021) <= not(inputs(188));
    layer0_outputs(2022) <= inputs(6);
    layer0_outputs(2023) <= inputs(217);
    layer0_outputs(2024) <= not(inputs(189)) or (inputs(45));
    layer0_outputs(2025) <= (inputs(71)) or (inputs(204));
    layer0_outputs(2026) <= inputs(154);
    layer0_outputs(2027) <= not((inputs(140)) or (inputs(115)));
    layer0_outputs(2028) <= inputs(100);
    layer0_outputs(2029) <= '0';
    layer0_outputs(2030) <= not(inputs(231)) or (inputs(13));
    layer0_outputs(2031) <= not(inputs(132));
    layer0_outputs(2032) <= not((inputs(245)) or (inputs(83)));
    layer0_outputs(2033) <= not(inputs(141));
    layer0_outputs(2034) <= (inputs(238)) xor (inputs(212));
    layer0_outputs(2035) <= '1';
    layer0_outputs(2036) <= not((inputs(160)) and (inputs(82)));
    layer0_outputs(2037) <= not(inputs(22));
    layer0_outputs(2038) <= (inputs(253)) and not (inputs(207));
    layer0_outputs(2039) <= not((inputs(194)) or (inputs(5)));
    layer0_outputs(2040) <= not(inputs(8)) or (inputs(220));
    layer0_outputs(2041) <= (inputs(165)) and not (inputs(228));
    layer0_outputs(2042) <= (inputs(53)) or (inputs(65));
    layer0_outputs(2043) <= (inputs(142)) and (inputs(146));
    layer0_outputs(2044) <= inputs(203);
    layer0_outputs(2045) <= not((inputs(236)) or (inputs(61)));
    layer0_outputs(2046) <= not((inputs(57)) xor (inputs(208)));
    layer0_outputs(2047) <= (inputs(223)) xor (inputs(105));
    layer0_outputs(2048) <= '1';
    layer0_outputs(2049) <= not((inputs(143)) or (inputs(215)));
    layer0_outputs(2050) <= (inputs(199)) or (inputs(127));
    layer0_outputs(2051) <= (inputs(105)) and not (inputs(0));
    layer0_outputs(2052) <= not((inputs(217)) or (inputs(104)));
    layer0_outputs(2053) <= (inputs(106)) and not (inputs(254));
    layer0_outputs(2054) <= not((inputs(92)) or (inputs(93)));
    layer0_outputs(2055) <= not(inputs(34));
    layer0_outputs(2056) <= '0';
    layer0_outputs(2057) <= not(inputs(107));
    layer0_outputs(2058) <= (inputs(86)) and not (inputs(32));
    layer0_outputs(2059) <= not(inputs(42)) or (inputs(94));
    layer0_outputs(2060) <= (inputs(131)) or (inputs(59));
    layer0_outputs(2061) <= not(inputs(252)) or (inputs(49));
    layer0_outputs(2062) <= inputs(234);
    layer0_outputs(2063) <= (inputs(146)) or (inputs(169));
    layer0_outputs(2064) <= (inputs(43)) and not (inputs(254));
    layer0_outputs(2065) <= (inputs(189)) or (inputs(252));
    layer0_outputs(2066) <= (inputs(175)) and not (inputs(245));
    layer0_outputs(2067) <= (inputs(158)) or (inputs(180));
    layer0_outputs(2068) <= (inputs(190)) or (inputs(250));
    layer0_outputs(2069) <= not(inputs(96)) or (inputs(23));
    layer0_outputs(2070) <= not((inputs(18)) or (inputs(103)));
    layer0_outputs(2071) <= (inputs(170)) or (inputs(38));
    layer0_outputs(2072) <= not(inputs(65));
    layer0_outputs(2073) <= not((inputs(138)) or (inputs(81)));
    layer0_outputs(2074) <= not(inputs(123));
    layer0_outputs(2075) <= inputs(150);
    layer0_outputs(2076) <= inputs(124);
    layer0_outputs(2077) <= (inputs(86)) and not (inputs(62));
    layer0_outputs(2078) <= (inputs(18)) or (inputs(182));
    layer0_outputs(2079) <= '0';
    layer0_outputs(2080) <= not(inputs(247)) or (inputs(207));
    layer0_outputs(2081) <= '1';
    layer0_outputs(2082) <= inputs(68);
    layer0_outputs(2083) <= not(inputs(26)) or (inputs(62));
    layer0_outputs(2084) <= inputs(156);
    layer0_outputs(2085) <= (inputs(198)) and not (inputs(206));
    layer0_outputs(2086) <= (inputs(198)) or (inputs(80));
    layer0_outputs(2087) <= not((inputs(34)) or (inputs(231)));
    layer0_outputs(2088) <= not((inputs(21)) or (inputs(14)));
    layer0_outputs(2089) <= (inputs(84)) xor (inputs(41));
    layer0_outputs(2090) <= not((inputs(157)) or (inputs(132)));
    layer0_outputs(2091) <= inputs(231);
    layer0_outputs(2092) <= (inputs(219)) and not (inputs(206));
    layer0_outputs(2093) <= (inputs(153)) and not (inputs(182));
    layer0_outputs(2094) <= (inputs(128)) or (inputs(86));
    layer0_outputs(2095) <= (inputs(9)) or (inputs(194));
    layer0_outputs(2096) <= (inputs(18)) or (inputs(130));
    layer0_outputs(2097) <= (inputs(117)) and not (inputs(80));
    layer0_outputs(2098) <= not((inputs(54)) xor (inputs(144)));
    layer0_outputs(2099) <= not((inputs(239)) xor (inputs(228)));
    layer0_outputs(2100) <= inputs(57);
    layer0_outputs(2101) <= inputs(84);
    layer0_outputs(2102) <= not((inputs(211)) or (inputs(188)));
    layer0_outputs(2103) <= (inputs(145)) xor (inputs(166));
    layer0_outputs(2104) <= not(inputs(179));
    layer0_outputs(2105) <= inputs(57);
    layer0_outputs(2106) <= not(inputs(242));
    layer0_outputs(2107) <= not(inputs(100)) or (inputs(13));
    layer0_outputs(2108) <= not((inputs(87)) xor (inputs(70)));
    layer0_outputs(2109) <= not((inputs(35)) xor (inputs(196)));
    layer0_outputs(2110) <= inputs(41);
    layer0_outputs(2111) <= not(inputs(92));
    layer0_outputs(2112) <= (inputs(118)) and not (inputs(38));
    layer0_outputs(2113) <= (inputs(25)) xor (inputs(76));
    layer0_outputs(2114) <= '0';
    layer0_outputs(2115) <= not((inputs(106)) or (inputs(150)));
    layer0_outputs(2116) <= inputs(254);
    layer0_outputs(2117) <= not((inputs(206)) or (inputs(68)));
    layer0_outputs(2118) <= (inputs(57)) or (inputs(37));
    layer0_outputs(2119) <= not(inputs(47));
    layer0_outputs(2120) <= not(inputs(182));
    layer0_outputs(2121) <= (inputs(107)) and not (inputs(22));
    layer0_outputs(2122) <= not((inputs(228)) and (inputs(7)));
    layer0_outputs(2123) <= (inputs(71)) and not (inputs(204));
    layer0_outputs(2124) <= '0';
    layer0_outputs(2125) <= inputs(182);
    layer0_outputs(2126) <= inputs(207);
    layer0_outputs(2127) <= inputs(214);
    layer0_outputs(2128) <= inputs(40);
    layer0_outputs(2129) <= (inputs(180)) or (inputs(251));
    layer0_outputs(2130) <= not((inputs(91)) or (inputs(122)));
    layer0_outputs(2131) <= not(inputs(193));
    layer0_outputs(2132) <= '1';
    layer0_outputs(2133) <= not(inputs(201)) or (inputs(32));
    layer0_outputs(2134) <= inputs(214);
    layer0_outputs(2135) <= not(inputs(52)) or (inputs(144));
    layer0_outputs(2136) <= (inputs(192)) and not (inputs(2));
    layer0_outputs(2137) <= (inputs(179)) and not (inputs(6));
    layer0_outputs(2138) <= '0';
    layer0_outputs(2139) <= (inputs(255)) and not (inputs(143));
    layer0_outputs(2140) <= inputs(59);
    layer0_outputs(2141) <= not((inputs(76)) xor (inputs(75)));
    layer0_outputs(2142) <= inputs(82);
    layer0_outputs(2143) <= not(inputs(229));
    layer0_outputs(2144) <= inputs(118);
    layer0_outputs(2145) <= '1';
    layer0_outputs(2146) <= (inputs(40)) and not (inputs(90));
    layer0_outputs(2147) <= '0';
    layer0_outputs(2148) <= (inputs(203)) and not (inputs(7));
    layer0_outputs(2149) <= not(inputs(114));
    layer0_outputs(2150) <= not((inputs(216)) xor (inputs(240)));
    layer0_outputs(2151) <= not((inputs(158)) and (inputs(243)));
    layer0_outputs(2152) <= not((inputs(172)) or (inputs(187)));
    layer0_outputs(2153) <= not(inputs(217));
    layer0_outputs(2154) <= (inputs(106)) xor (inputs(210));
    layer0_outputs(2155) <= not(inputs(202));
    layer0_outputs(2156) <= not((inputs(148)) xor (inputs(4)));
    layer0_outputs(2157) <= not(inputs(151)) or (inputs(127));
    layer0_outputs(2158) <= not((inputs(150)) or (inputs(220)));
    layer0_outputs(2159) <= '1';
    layer0_outputs(2160) <= not(inputs(132));
    layer0_outputs(2161) <= not((inputs(108)) xor (inputs(233)));
    layer0_outputs(2162) <= not((inputs(15)) xor (inputs(150)));
    layer0_outputs(2163) <= inputs(255);
    layer0_outputs(2164) <= (inputs(116)) and not (inputs(84));
    layer0_outputs(2165) <= (inputs(200)) and not (inputs(31));
    layer0_outputs(2166) <= (inputs(12)) and (inputs(12));
    layer0_outputs(2167) <= not(inputs(179)) or (inputs(64));
    layer0_outputs(2168) <= not((inputs(84)) or (inputs(42)));
    layer0_outputs(2169) <= (inputs(178)) and not (inputs(15));
    layer0_outputs(2170) <= not(inputs(188)) or (inputs(253));
    layer0_outputs(2171) <= (inputs(230)) or (inputs(106));
    layer0_outputs(2172) <= (inputs(198)) and not (inputs(110));
    layer0_outputs(2173) <= not((inputs(96)) or (inputs(221)));
    layer0_outputs(2174) <= (inputs(167)) and not (inputs(251));
    layer0_outputs(2175) <= not((inputs(64)) or (inputs(234)));
    layer0_outputs(2176) <= not(inputs(186)) or (inputs(65));
    layer0_outputs(2177) <= not((inputs(10)) or (inputs(110)));
    layer0_outputs(2178) <= not((inputs(96)) or (inputs(101)));
    layer0_outputs(2179) <= inputs(119);
    layer0_outputs(2180) <= '0';
    layer0_outputs(2181) <= not(inputs(124));
    layer0_outputs(2182) <= (inputs(176)) and not (inputs(245));
    layer0_outputs(2183) <= (inputs(23)) and not (inputs(91));
    layer0_outputs(2184) <= '0';
    layer0_outputs(2185) <= (inputs(65)) or (inputs(177));
    layer0_outputs(2186) <= not(inputs(158)) or (inputs(236));
    layer0_outputs(2187) <= (inputs(133)) and not (inputs(38));
    layer0_outputs(2188) <= (inputs(193)) and not (inputs(34));
    layer0_outputs(2189) <= not(inputs(84)) or (inputs(194));
    layer0_outputs(2190) <= not((inputs(173)) xor (inputs(4)));
    layer0_outputs(2191) <= not(inputs(120)) or (inputs(62));
    layer0_outputs(2192) <= not(inputs(164)) or (inputs(45));
    layer0_outputs(2193) <= not(inputs(80));
    layer0_outputs(2194) <= not(inputs(30)) or (inputs(240));
    layer0_outputs(2195) <= not(inputs(44));
    layer0_outputs(2196) <= (inputs(250)) and not (inputs(141));
    layer0_outputs(2197) <= not((inputs(162)) xor (inputs(190)));
    layer0_outputs(2198) <= (inputs(186)) and not (inputs(206));
    layer0_outputs(2199) <= '1';
    layer0_outputs(2200) <= (inputs(102)) and not (inputs(251));
    layer0_outputs(2201) <= (inputs(239)) and (inputs(239));
    layer0_outputs(2202) <= (inputs(25)) xor (inputs(114));
    layer0_outputs(2203) <= not((inputs(184)) or (inputs(222)));
    layer0_outputs(2204) <= (inputs(50)) and (inputs(110));
    layer0_outputs(2205) <= not((inputs(214)) or (inputs(98)));
    layer0_outputs(2206) <= (inputs(84)) or (inputs(250));
    layer0_outputs(2207) <= (inputs(254)) xor (inputs(121));
    layer0_outputs(2208) <= not((inputs(91)) xor (inputs(12)));
    layer0_outputs(2209) <= not(inputs(123));
    layer0_outputs(2210) <= not((inputs(110)) or (inputs(133)));
    layer0_outputs(2211) <= not((inputs(8)) xor (inputs(169)));
    layer0_outputs(2212) <= not(inputs(183));
    layer0_outputs(2213) <= inputs(87);
    layer0_outputs(2214) <= (inputs(170)) or (inputs(96));
    layer0_outputs(2215) <= not(inputs(122));
    layer0_outputs(2216) <= inputs(182);
    layer0_outputs(2217) <= not(inputs(54)) or (inputs(117));
    layer0_outputs(2218) <= not(inputs(177)) or (inputs(254));
    layer0_outputs(2219) <= (inputs(12)) or (inputs(183));
    layer0_outputs(2220) <= not(inputs(74));
    layer0_outputs(2221) <= not(inputs(40)) or (inputs(88));
    layer0_outputs(2222) <= '0';
    layer0_outputs(2223) <= not(inputs(112)) or (inputs(21));
    layer0_outputs(2224) <= (inputs(3)) xor (inputs(241));
    layer0_outputs(2225) <= (inputs(9)) and (inputs(144));
    layer0_outputs(2226) <= not(inputs(51)) or (inputs(96));
    layer0_outputs(2227) <= (inputs(219)) or (inputs(178));
    layer0_outputs(2228) <= inputs(167);
    layer0_outputs(2229) <= not(inputs(71));
    layer0_outputs(2230) <= (inputs(143)) or (inputs(125));
    layer0_outputs(2231) <= (inputs(47)) and not (inputs(31));
    layer0_outputs(2232) <= (inputs(251)) xor (inputs(158));
    layer0_outputs(2233) <= '0';
    layer0_outputs(2234) <= (inputs(171)) and not (inputs(175));
    layer0_outputs(2235) <= inputs(235);
    layer0_outputs(2236) <= not((inputs(87)) or (inputs(247)));
    layer0_outputs(2237) <= (inputs(167)) and not (inputs(196));
    layer0_outputs(2238) <= (inputs(7)) or (inputs(39));
    layer0_outputs(2239) <= not(inputs(181));
    layer0_outputs(2240) <= not(inputs(214));
    layer0_outputs(2241) <= (inputs(116)) and not (inputs(44));
    layer0_outputs(2242) <= (inputs(138)) xor (inputs(57));
    layer0_outputs(2243) <= (inputs(138)) and not (inputs(210));
    layer0_outputs(2244) <= not((inputs(22)) xor (inputs(41)));
    layer0_outputs(2245) <= (inputs(8)) or (inputs(31));
    layer0_outputs(2246) <= (inputs(251)) xor (inputs(232));
    layer0_outputs(2247) <= (inputs(133)) and not (inputs(14));
    layer0_outputs(2248) <= (inputs(244)) or (inputs(48));
    layer0_outputs(2249) <= not(inputs(152));
    layer0_outputs(2250) <= inputs(166);
    layer0_outputs(2251) <= not(inputs(199));
    layer0_outputs(2252) <= (inputs(161)) and not (inputs(111));
    layer0_outputs(2253) <= (inputs(16)) xor (inputs(100));
    layer0_outputs(2254) <= not((inputs(47)) and (inputs(81)));
    layer0_outputs(2255) <= not((inputs(181)) or (inputs(29)));
    layer0_outputs(2256) <= (inputs(96)) or (inputs(42));
    layer0_outputs(2257) <= not(inputs(207));
    layer0_outputs(2258) <= not(inputs(89));
    layer0_outputs(2259) <= not((inputs(38)) and (inputs(85)));
    layer0_outputs(2260) <= inputs(104);
    layer0_outputs(2261) <= inputs(131);
    layer0_outputs(2262) <= (inputs(235)) or (inputs(137));
    layer0_outputs(2263) <= (inputs(122)) or (inputs(54));
    layer0_outputs(2264) <= not((inputs(173)) or (inputs(219)));
    layer0_outputs(2265) <= not((inputs(197)) or (inputs(100)));
    layer0_outputs(2266) <= not((inputs(44)) or (inputs(180)));
    layer0_outputs(2267) <= inputs(213);
    layer0_outputs(2268) <= (inputs(54)) or (inputs(162));
    layer0_outputs(2269) <= (inputs(181)) or (inputs(149));
    layer0_outputs(2270) <= (inputs(70)) and not (inputs(123));
    layer0_outputs(2271) <= not((inputs(239)) or (inputs(176)));
    layer0_outputs(2272) <= not(inputs(195));
    layer0_outputs(2273) <= inputs(86);
    layer0_outputs(2274) <= (inputs(153)) or (inputs(149));
    layer0_outputs(2275) <= (inputs(18)) xor (inputs(187));
    layer0_outputs(2276) <= not((inputs(125)) or (inputs(117)));
    layer0_outputs(2277) <= not((inputs(21)) or (inputs(95)));
    layer0_outputs(2278) <= not(inputs(215)) or (inputs(182));
    layer0_outputs(2279) <= not((inputs(226)) xor (inputs(52)));
    layer0_outputs(2280) <= not(inputs(73));
    layer0_outputs(2281) <= not(inputs(246));
    layer0_outputs(2282) <= (inputs(34)) xor (inputs(128));
    layer0_outputs(2283) <= not(inputs(188));
    layer0_outputs(2284) <= not((inputs(57)) xor (inputs(247)));
    layer0_outputs(2285) <= not((inputs(43)) xor (inputs(17)));
    layer0_outputs(2286) <= not(inputs(136)) or (inputs(108));
    layer0_outputs(2287) <= (inputs(169)) and not (inputs(46));
    layer0_outputs(2288) <= not((inputs(198)) or (inputs(53)));
    layer0_outputs(2289) <= (inputs(87)) and not (inputs(145));
    layer0_outputs(2290) <= (inputs(146)) and not (inputs(112));
    layer0_outputs(2291) <= not(inputs(131)) or (inputs(35));
    layer0_outputs(2292) <= not((inputs(139)) xor (inputs(71)));
    layer0_outputs(2293) <= inputs(203);
    layer0_outputs(2294) <= (inputs(131)) or (inputs(229));
    layer0_outputs(2295) <= not((inputs(9)) or (inputs(100)));
    layer0_outputs(2296) <= inputs(68);
    layer0_outputs(2297) <= inputs(153);
    layer0_outputs(2298) <= inputs(117);
    layer0_outputs(2299) <= not(inputs(158));
    layer0_outputs(2300) <= (inputs(54)) and not (inputs(227));
    layer0_outputs(2301) <= (inputs(233)) or (inputs(9));
    layer0_outputs(2302) <= not(inputs(167));
    layer0_outputs(2303) <= (inputs(242)) or (inputs(116));
    layer0_outputs(2304) <= (inputs(222)) or (inputs(184));
    layer0_outputs(2305) <= (inputs(217)) xor (inputs(208));
    layer0_outputs(2306) <= not(inputs(226));
    layer0_outputs(2307) <= not(inputs(45));
    layer0_outputs(2308) <= not((inputs(244)) or (inputs(123)));
    layer0_outputs(2309) <= (inputs(151)) and not (inputs(83));
    layer0_outputs(2310) <= not(inputs(117));
    layer0_outputs(2311) <= (inputs(211)) and not (inputs(44));
    layer0_outputs(2312) <= not((inputs(53)) and (inputs(5)));
    layer0_outputs(2313) <= (inputs(28)) xor (inputs(217));
    layer0_outputs(2314) <= not(inputs(79)) or (inputs(167));
    layer0_outputs(2315) <= not(inputs(190)) or (inputs(9));
    layer0_outputs(2316) <= not((inputs(208)) or (inputs(125)));
    layer0_outputs(2317) <= not((inputs(155)) or (inputs(140)));
    layer0_outputs(2318) <= (inputs(20)) and (inputs(99));
    layer0_outputs(2319) <= not((inputs(108)) or (inputs(56)));
    layer0_outputs(2320) <= not(inputs(199));
    layer0_outputs(2321) <= not((inputs(1)) and (inputs(160)));
    layer0_outputs(2322) <= not(inputs(24)) or (inputs(17));
    layer0_outputs(2323) <= (inputs(142)) or (inputs(210));
    layer0_outputs(2324) <= not(inputs(148));
    layer0_outputs(2325) <= not(inputs(135)) or (inputs(233));
    layer0_outputs(2326) <= inputs(252);
    layer0_outputs(2327) <= not(inputs(229)) or (inputs(48));
    layer0_outputs(2328) <= (inputs(21)) and not (inputs(41));
    layer0_outputs(2329) <= (inputs(118)) xor (inputs(247));
    layer0_outputs(2330) <= (inputs(102)) and not (inputs(198));
    layer0_outputs(2331) <= (inputs(4)) xor (inputs(234));
    layer0_outputs(2332) <= not(inputs(134)) or (inputs(41));
    layer0_outputs(2333) <= inputs(189);
    layer0_outputs(2334) <= (inputs(98)) or (inputs(108));
    layer0_outputs(2335) <= inputs(194);
    layer0_outputs(2336) <= not(inputs(215)) or (inputs(16));
    layer0_outputs(2337) <= not(inputs(86));
    layer0_outputs(2338) <= not(inputs(96));
    layer0_outputs(2339) <= (inputs(189)) or (inputs(191));
    layer0_outputs(2340) <= not((inputs(245)) xor (inputs(85)));
    layer0_outputs(2341) <= not((inputs(57)) xor (inputs(252)));
    layer0_outputs(2342) <= inputs(58);
    layer0_outputs(2343) <= not((inputs(146)) xor (inputs(134)));
    layer0_outputs(2344) <= (inputs(78)) and not (inputs(54));
    layer0_outputs(2345) <= (inputs(152)) or (inputs(151));
    layer0_outputs(2346) <= not(inputs(69));
    layer0_outputs(2347) <= (inputs(127)) and not (inputs(80));
    layer0_outputs(2348) <= not(inputs(101));
    layer0_outputs(2349) <= (inputs(45)) and (inputs(12));
    layer0_outputs(2350) <= not((inputs(34)) xor (inputs(85)));
    layer0_outputs(2351) <= not(inputs(38)) or (inputs(227));
    layer0_outputs(2352) <= not((inputs(144)) or (inputs(221)));
    layer0_outputs(2353) <= (inputs(78)) xor (inputs(99));
    layer0_outputs(2354) <= inputs(181);
    layer0_outputs(2355) <= not((inputs(44)) or (inputs(191)));
    layer0_outputs(2356) <= (inputs(189)) or (inputs(187));
    layer0_outputs(2357) <= not(inputs(150));
    layer0_outputs(2358) <= (inputs(206)) xor (inputs(189));
    layer0_outputs(2359) <= inputs(98);
    layer0_outputs(2360) <= inputs(234);
    layer0_outputs(2361) <= (inputs(215)) or (inputs(61));
    layer0_outputs(2362) <= inputs(216);
    layer0_outputs(2363) <= (inputs(78)) and not (inputs(248));
    layer0_outputs(2364) <= inputs(164);
    layer0_outputs(2365) <= not(inputs(161)) or (inputs(158));
    layer0_outputs(2366) <= (inputs(95)) xor (inputs(146));
    layer0_outputs(2367) <= not(inputs(125));
    layer0_outputs(2368) <= inputs(165);
    layer0_outputs(2369) <= not((inputs(137)) or (inputs(99)));
    layer0_outputs(2370) <= not((inputs(8)) xor (inputs(242)));
    layer0_outputs(2371) <= (inputs(199)) and not (inputs(224));
    layer0_outputs(2372) <= inputs(30);
    layer0_outputs(2373) <= (inputs(1)) xor (inputs(122));
    layer0_outputs(2374) <= not(inputs(161)) or (inputs(12));
    layer0_outputs(2375) <= not(inputs(142)) or (inputs(46));
    layer0_outputs(2376) <= not((inputs(193)) or (inputs(201)));
    layer0_outputs(2377) <= '1';
    layer0_outputs(2378) <= '1';
    layer0_outputs(2379) <= not((inputs(253)) or (inputs(75)));
    layer0_outputs(2380) <= not(inputs(144));
    layer0_outputs(2381) <= not(inputs(115)) or (inputs(192));
    layer0_outputs(2382) <= (inputs(139)) or (inputs(211));
    layer0_outputs(2383) <= inputs(206);
    layer0_outputs(2384) <= not((inputs(173)) and (inputs(227)));
    layer0_outputs(2385) <= (inputs(165)) or (inputs(203));
    layer0_outputs(2386) <= inputs(66);
    layer0_outputs(2387) <= (inputs(86)) and not (inputs(197));
    layer0_outputs(2388) <= not(inputs(90)) or (inputs(114));
    layer0_outputs(2389) <= not((inputs(83)) xor (inputs(40)));
    layer0_outputs(2390) <= not((inputs(106)) xor (inputs(60)));
    layer0_outputs(2391) <= (inputs(162)) and not (inputs(158));
    layer0_outputs(2392) <= (inputs(70)) and not (inputs(7));
    layer0_outputs(2393) <= not(inputs(38));
    layer0_outputs(2394) <= not((inputs(32)) xor (inputs(130)));
    layer0_outputs(2395) <= not((inputs(238)) or (inputs(92)));
    layer0_outputs(2396) <= not((inputs(187)) or (inputs(160)));
    layer0_outputs(2397) <= (inputs(249)) or (inputs(212));
    layer0_outputs(2398) <= inputs(180);
    layer0_outputs(2399) <= (inputs(17)) and not (inputs(127));
    layer0_outputs(2400) <= (inputs(203)) and not (inputs(231));
    layer0_outputs(2401) <= not((inputs(208)) xor (inputs(206)));
    layer0_outputs(2402) <= inputs(137);
    layer0_outputs(2403) <= not((inputs(251)) xor (inputs(58)));
    layer0_outputs(2404) <= not(inputs(65));
    layer0_outputs(2405) <= inputs(253);
    layer0_outputs(2406) <= inputs(99);
    layer0_outputs(2407) <= (inputs(108)) or (inputs(221));
    layer0_outputs(2408) <= (inputs(205)) xor (inputs(1));
    layer0_outputs(2409) <= not(inputs(171)) or (inputs(147));
    layer0_outputs(2410) <= inputs(13);
    layer0_outputs(2411) <= (inputs(45)) xor (inputs(55));
    layer0_outputs(2412) <= (inputs(136)) and not (inputs(142));
    layer0_outputs(2413) <= (inputs(126)) xor (inputs(147));
    layer0_outputs(2414) <= (inputs(99)) and not (inputs(236));
    layer0_outputs(2415) <= (inputs(53)) xor (inputs(200));
    layer0_outputs(2416) <= (inputs(109)) and not (inputs(21));
    layer0_outputs(2417) <= (inputs(110)) and (inputs(28));
    layer0_outputs(2418) <= inputs(219);
    layer0_outputs(2419) <= '0';
    layer0_outputs(2420) <= (inputs(234)) xor (inputs(18));
    layer0_outputs(2421) <= inputs(216);
    layer0_outputs(2422) <= not(inputs(102));
    layer0_outputs(2423) <= not(inputs(9)) or (inputs(157));
    layer0_outputs(2424) <= (inputs(204)) or (inputs(71));
    layer0_outputs(2425) <= inputs(88);
    layer0_outputs(2426) <= not(inputs(170));
    layer0_outputs(2427) <= inputs(38);
    layer0_outputs(2428) <= (inputs(110)) and not (inputs(109));
    layer0_outputs(2429) <= not((inputs(134)) xor (inputs(32)));
    layer0_outputs(2430) <= inputs(34);
    layer0_outputs(2431) <= '1';
    layer0_outputs(2432) <= not(inputs(154)) or (inputs(209));
    layer0_outputs(2433) <= not(inputs(207)) or (inputs(175));
    layer0_outputs(2434) <= inputs(140);
    layer0_outputs(2435) <= (inputs(182)) or (inputs(165));
    layer0_outputs(2436) <= not((inputs(43)) and (inputs(81)));
    layer0_outputs(2437) <= not((inputs(56)) xor (inputs(251)));
    layer0_outputs(2438) <= (inputs(138)) and not (inputs(42));
    layer0_outputs(2439) <= (inputs(50)) or (inputs(138));
    layer0_outputs(2440) <= not((inputs(110)) and (inputs(41)));
    layer0_outputs(2441) <= not(inputs(217)) or (inputs(19));
    layer0_outputs(2442) <= not((inputs(172)) or (inputs(171)));
    layer0_outputs(2443) <= not((inputs(63)) or (inputs(200)));
    layer0_outputs(2444) <= inputs(137);
    layer0_outputs(2445) <= not(inputs(120));
    layer0_outputs(2446) <= not(inputs(212)) or (inputs(62));
    layer0_outputs(2447) <= (inputs(155)) xor (inputs(225));
    layer0_outputs(2448) <= (inputs(95)) and not (inputs(1));
    layer0_outputs(2449) <= (inputs(23)) and not (inputs(83));
    layer0_outputs(2450) <= not((inputs(253)) or (inputs(91)));
    layer0_outputs(2451) <= (inputs(63)) and (inputs(14));
    layer0_outputs(2452) <= (inputs(52)) and not (inputs(246));
    layer0_outputs(2453) <= not((inputs(201)) and (inputs(72)));
    layer0_outputs(2454) <= (inputs(37)) xor (inputs(169));
    layer0_outputs(2455) <= (inputs(220)) xor (inputs(188));
    layer0_outputs(2456) <= not((inputs(212)) xor (inputs(75)));
    layer0_outputs(2457) <= not((inputs(45)) or (inputs(223)));
    layer0_outputs(2458) <= (inputs(72)) and not (inputs(220));
    layer0_outputs(2459) <= not(inputs(233));
    layer0_outputs(2460) <= (inputs(86)) and not (inputs(230));
    layer0_outputs(2461) <= (inputs(155)) and not (inputs(46));
    layer0_outputs(2462) <= (inputs(181)) xor (inputs(161));
    layer0_outputs(2463) <= not(inputs(128));
    layer0_outputs(2464) <= not((inputs(116)) or (inputs(24)));
    layer0_outputs(2465) <= inputs(198);
    layer0_outputs(2466) <= (inputs(48)) and not (inputs(133));
    layer0_outputs(2467) <= (inputs(33)) and (inputs(3));
    layer0_outputs(2468) <= (inputs(88)) and not (inputs(150));
    layer0_outputs(2469) <= inputs(164);
    layer0_outputs(2470) <= '1';
    layer0_outputs(2471) <= not(inputs(208)) or (inputs(205));
    layer0_outputs(2472) <= (inputs(184)) and not (inputs(130));
    layer0_outputs(2473) <= (inputs(149)) or (inputs(167));
    layer0_outputs(2474) <= (inputs(26)) or (inputs(110));
    layer0_outputs(2475) <= (inputs(196)) xor (inputs(34));
    layer0_outputs(2476) <= (inputs(45)) and (inputs(223));
    layer0_outputs(2477) <= not(inputs(40)) or (inputs(231));
    layer0_outputs(2478) <= inputs(66);
    layer0_outputs(2479) <= not(inputs(217)) or (inputs(250));
    layer0_outputs(2480) <= (inputs(193)) and not (inputs(142));
    layer0_outputs(2481) <= inputs(186);
    layer0_outputs(2482) <= (inputs(146)) or (inputs(118));
    layer0_outputs(2483) <= not((inputs(108)) xor (inputs(68)));
    layer0_outputs(2484) <= not(inputs(71)) or (inputs(14));
    layer0_outputs(2485) <= (inputs(135)) or (inputs(143));
    layer0_outputs(2486) <= not((inputs(208)) xor (inputs(25)));
    layer0_outputs(2487) <= (inputs(194)) or (inputs(166));
    layer0_outputs(2488) <= not(inputs(155)) or (inputs(174));
    layer0_outputs(2489) <= not(inputs(145)) or (inputs(7));
    layer0_outputs(2490) <= not(inputs(42)) or (inputs(225));
    layer0_outputs(2491) <= inputs(41);
    layer0_outputs(2492) <= (inputs(206)) xor (inputs(6));
    layer0_outputs(2493) <= (inputs(167)) and not (inputs(39));
    layer0_outputs(2494) <= inputs(40);
    layer0_outputs(2495) <= not((inputs(172)) or (inputs(23)));
    layer0_outputs(2496) <= (inputs(243)) and (inputs(128));
    layer0_outputs(2497) <= not(inputs(35)) or (inputs(81));
    layer0_outputs(2498) <= (inputs(116)) and not (inputs(10));
    layer0_outputs(2499) <= not((inputs(61)) or (inputs(133)));
    layer0_outputs(2500) <= inputs(212);
    layer0_outputs(2501) <= not((inputs(99)) xor (inputs(148)));
    layer0_outputs(2502) <= not(inputs(230)) or (inputs(145));
    layer0_outputs(2503) <= not(inputs(123));
    layer0_outputs(2504) <= not(inputs(76)) or (inputs(35));
    layer0_outputs(2505) <= not((inputs(122)) xor (inputs(249)));
    layer0_outputs(2506) <= not((inputs(204)) xor (inputs(147)));
    layer0_outputs(2507) <= (inputs(164)) and not (inputs(177));
    layer0_outputs(2508) <= (inputs(192)) xor (inputs(86));
    layer0_outputs(2509) <= inputs(128);
    layer0_outputs(2510) <= '0';
    layer0_outputs(2511) <= inputs(1);
    layer0_outputs(2512) <= (inputs(212)) and not (inputs(79));
    layer0_outputs(2513) <= (inputs(228)) or (inputs(197));
    layer0_outputs(2514) <= inputs(173);
    layer0_outputs(2515) <= not((inputs(233)) or (inputs(209)));
    layer0_outputs(2516) <= not(inputs(200)) or (inputs(44));
    layer0_outputs(2517) <= not((inputs(28)) or (inputs(138)));
    layer0_outputs(2518) <= '1';
    layer0_outputs(2519) <= not((inputs(235)) xor (inputs(35)));
    layer0_outputs(2520) <= not(inputs(143));
    layer0_outputs(2521) <= not(inputs(165)) or (inputs(6));
    layer0_outputs(2522) <= not(inputs(122)) or (inputs(156));
    layer0_outputs(2523) <= not((inputs(45)) and (inputs(244)));
    layer0_outputs(2524) <= (inputs(131)) and not (inputs(1));
    layer0_outputs(2525) <= inputs(147);
    layer0_outputs(2526) <= (inputs(247)) and (inputs(235));
    layer0_outputs(2527) <= not(inputs(227));
    layer0_outputs(2528) <= not((inputs(34)) xor (inputs(167)));
    layer0_outputs(2529) <= (inputs(108)) or (inputs(172));
    layer0_outputs(2530) <= not(inputs(116));
    layer0_outputs(2531) <= not(inputs(50)) or (inputs(11));
    layer0_outputs(2532) <= inputs(214);
    layer0_outputs(2533) <= not(inputs(60)) or (inputs(15));
    layer0_outputs(2534) <= not(inputs(33)) or (inputs(157));
    layer0_outputs(2535) <= (inputs(40)) or (inputs(253));
    layer0_outputs(2536) <= not((inputs(123)) or (inputs(194)));
    layer0_outputs(2537) <= (inputs(178)) or (inputs(224));
    layer0_outputs(2538) <= not(inputs(174));
    layer0_outputs(2539) <= '0';
    layer0_outputs(2540) <= (inputs(114)) and not (inputs(5));
    layer0_outputs(2541) <= (inputs(130)) xor (inputs(47));
    layer0_outputs(2542) <= inputs(183);
    layer0_outputs(2543) <= (inputs(222)) xor (inputs(255));
    layer0_outputs(2544) <= not((inputs(86)) or (inputs(28)));
    layer0_outputs(2545) <= inputs(164);
    layer0_outputs(2546) <= not((inputs(174)) xor (inputs(245)));
    layer0_outputs(2547) <= not(inputs(88));
    layer0_outputs(2548) <= (inputs(109)) or (inputs(4));
    layer0_outputs(2549) <= inputs(93);
    layer0_outputs(2550) <= not((inputs(0)) xor (inputs(196)));
    layer0_outputs(2551) <= (inputs(192)) and (inputs(156));
    layer0_outputs(2552) <= not((inputs(191)) xor (inputs(148)));
    layer0_outputs(2553) <= not((inputs(216)) or (inputs(211)));
    layer0_outputs(2554) <= inputs(105);
    layer0_outputs(2555) <= not(inputs(71)) or (inputs(51));
    layer0_outputs(2556) <= '1';
    layer0_outputs(2557) <= (inputs(5)) xor (inputs(68));
    layer0_outputs(2558) <= (inputs(123)) and not (inputs(25));
    layer0_outputs(2559) <= (inputs(244)) and not (inputs(65));
    layer0_outputs(2560) <= not((inputs(217)) or (inputs(11)));
    layer0_outputs(2561) <= (inputs(245)) or (inputs(58));
    layer0_outputs(2562) <= inputs(24);
    layer0_outputs(2563) <= (inputs(169)) and not (inputs(130));
    layer0_outputs(2564) <= (inputs(38)) and not (inputs(20));
    layer0_outputs(2565) <= (inputs(230)) and not (inputs(61));
    layer0_outputs(2566) <= inputs(109);
    layer0_outputs(2567) <= inputs(35);
    layer0_outputs(2568) <= (inputs(157)) and not (inputs(19));
    layer0_outputs(2569) <= not(inputs(250));
    layer0_outputs(2570) <= (inputs(107)) and not (inputs(172));
    layer0_outputs(2571) <= not(inputs(136));
    layer0_outputs(2572) <= not(inputs(173));
    layer0_outputs(2573) <= (inputs(56)) and not (inputs(125));
    layer0_outputs(2574) <= not(inputs(139)) or (inputs(96));
    layer0_outputs(2575) <= (inputs(117)) and not (inputs(89));
    layer0_outputs(2576) <= '1';
    layer0_outputs(2577) <= (inputs(90)) and not (inputs(62));
    layer0_outputs(2578) <= not((inputs(143)) xor (inputs(46)));
    layer0_outputs(2579) <= (inputs(114)) and not (inputs(30));
    layer0_outputs(2580) <= not((inputs(191)) xor (inputs(211)));
    layer0_outputs(2581) <= not((inputs(115)) xor (inputs(52)));
    layer0_outputs(2582) <= not((inputs(17)) and (inputs(0)));
    layer0_outputs(2583) <= (inputs(49)) and (inputs(144));
    layer0_outputs(2584) <= (inputs(203)) and not (inputs(200));
    layer0_outputs(2585) <= inputs(138);
    layer0_outputs(2586) <= (inputs(34)) xor (inputs(150));
    layer0_outputs(2587) <= (inputs(205)) or (inputs(22));
    layer0_outputs(2588) <= (inputs(71)) and not (inputs(223));
    layer0_outputs(2589) <= not((inputs(181)) or (inputs(190)));
    layer0_outputs(2590) <= (inputs(83)) xor (inputs(35));
    layer0_outputs(2591) <= (inputs(61)) and not (inputs(75));
    layer0_outputs(2592) <= (inputs(91)) xor (inputs(192));
    layer0_outputs(2593) <= (inputs(226)) and not (inputs(203));
    layer0_outputs(2594) <= not(inputs(246)) or (inputs(13));
    layer0_outputs(2595) <= not((inputs(212)) and (inputs(158)));
    layer0_outputs(2596) <= (inputs(130)) or (inputs(93));
    layer0_outputs(2597) <= inputs(55);
    layer0_outputs(2598) <= not((inputs(156)) or (inputs(94)));
    layer0_outputs(2599) <= (inputs(151)) or (inputs(165));
    layer0_outputs(2600) <= (inputs(235)) and (inputs(235));
    layer0_outputs(2601) <= '0';
    layer0_outputs(2602) <= not(inputs(248));
    layer0_outputs(2603) <= not((inputs(240)) or (inputs(98)));
    layer0_outputs(2604) <= not((inputs(158)) xor (inputs(40)));
    layer0_outputs(2605) <= (inputs(139)) and not (inputs(13));
    layer0_outputs(2606) <= not(inputs(93)) or (inputs(28));
    layer0_outputs(2607) <= not((inputs(78)) and (inputs(252)));
    layer0_outputs(2608) <= (inputs(165)) and not (inputs(116));
    layer0_outputs(2609) <= not(inputs(207));
    layer0_outputs(2610) <= (inputs(167)) and not (inputs(94));
    layer0_outputs(2611) <= not(inputs(66));
    layer0_outputs(2612) <= not((inputs(154)) or (inputs(129)));
    layer0_outputs(2613) <= (inputs(118)) and not (inputs(179));
    layer0_outputs(2614) <= inputs(195);
    layer0_outputs(2615) <= (inputs(76)) xor (inputs(178));
    layer0_outputs(2616) <= not((inputs(116)) or (inputs(21)));
    layer0_outputs(2617) <= (inputs(174)) xor (inputs(241));
    layer0_outputs(2618) <= not(inputs(248));
    layer0_outputs(2619) <= not(inputs(189));
    layer0_outputs(2620) <= not(inputs(108)) or (inputs(95));
    layer0_outputs(2621) <= not(inputs(69));
    layer0_outputs(2622) <= (inputs(219)) xor (inputs(229));
    layer0_outputs(2623) <= not((inputs(244)) xor (inputs(149)));
    layer0_outputs(2624) <= '0';
    layer0_outputs(2625) <= not(inputs(143));
    layer0_outputs(2626) <= inputs(30);
    layer0_outputs(2627) <= (inputs(214)) or (inputs(103));
    layer0_outputs(2628) <= not((inputs(182)) xor (inputs(104)));
    layer0_outputs(2629) <= not((inputs(55)) or (inputs(214)));
    layer0_outputs(2630) <= '1';
    layer0_outputs(2631) <= not((inputs(157)) xor (inputs(9)));
    layer0_outputs(2632) <= (inputs(139)) and (inputs(177));
    layer0_outputs(2633) <= inputs(148);
    layer0_outputs(2634) <= not((inputs(238)) or (inputs(106)));
    layer0_outputs(2635) <= '1';
    layer0_outputs(2636) <= inputs(251);
    layer0_outputs(2637) <= (inputs(204)) and not (inputs(146));
    layer0_outputs(2638) <= (inputs(103)) xor (inputs(64));
    layer0_outputs(2639) <= (inputs(182)) or (inputs(234));
    layer0_outputs(2640) <= '0';
    layer0_outputs(2641) <= (inputs(87)) xor (inputs(85));
    layer0_outputs(2642) <= not((inputs(88)) or (inputs(78)));
    layer0_outputs(2643) <= not(inputs(151));
    layer0_outputs(2644) <= (inputs(1)) or (inputs(109));
    layer0_outputs(2645) <= (inputs(58)) xor (inputs(192));
    layer0_outputs(2646) <= not(inputs(93));
    layer0_outputs(2647) <= (inputs(106)) or (inputs(206));
    layer0_outputs(2648) <= (inputs(66)) xor (inputs(181));
    layer0_outputs(2649) <= (inputs(47)) and not (inputs(134));
    layer0_outputs(2650) <= inputs(148);
    layer0_outputs(2651) <= (inputs(98)) and not (inputs(82));
    layer0_outputs(2652) <= inputs(150);
    layer0_outputs(2653) <= inputs(73);
    layer0_outputs(2654) <= not(inputs(93));
    layer0_outputs(2655) <= (inputs(72)) or (inputs(196));
    layer0_outputs(2656) <= (inputs(53)) and not (inputs(11));
    layer0_outputs(2657) <= not((inputs(84)) xor (inputs(133)));
    layer0_outputs(2658) <= not(inputs(113));
    layer0_outputs(2659) <= (inputs(188)) or (inputs(75));
    layer0_outputs(2660) <= (inputs(162)) or (inputs(38));
    layer0_outputs(2661) <= (inputs(123)) or (inputs(82));
    layer0_outputs(2662) <= inputs(115);
    layer0_outputs(2663) <= '1';
    layer0_outputs(2664) <= not(inputs(218));
    layer0_outputs(2665) <= (inputs(152)) and (inputs(249));
    layer0_outputs(2666) <= not((inputs(248)) or (inputs(10)));
    layer0_outputs(2667) <= (inputs(64)) or (inputs(97));
    layer0_outputs(2668) <= not((inputs(120)) xor (inputs(43)));
    layer0_outputs(2669) <= not(inputs(152));
    layer0_outputs(2670) <= not(inputs(33)) or (inputs(72));
    layer0_outputs(2671) <= not((inputs(41)) or (inputs(244)));
    layer0_outputs(2672) <= (inputs(74)) xor (inputs(170));
    layer0_outputs(2673) <= (inputs(169)) and not (inputs(253));
    layer0_outputs(2674) <= not(inputs(95));
    layer0_outputs(2675) <= (inputs(9)) or (inputs(168));
    layer0_outputs(2676) <= '0';
    layer0_outputs(2677) <= not(inputs(176));
    layer0_outputs(2678) <= '0';
    layer0_outputs(2679) <= (inputs(145)) xor (inputs(170));
    layer0_outputs(2680) <= not(inputs(37)) or (inputs(124));
    layer0_outputs(2681) <= not(inputs(36));
    layer0_outputs(2682) <= not(inputs(241)) or (inputs(19));
    layer0_outputs(2683) <= not((inputs(74)) or (inputs(51)));
    layer0_outputs(2684) <= not((inputs(50)) xor (inputs(99)));
    layer0_outputs(2685) <= inputs(101);
    layer0_outputs(2686) <= not(inputs(61));
    layer0_outputs(2687) <= (inputs(29)) or (inputs(57));
    layer0_outputs(2688) <= (inputs(7)) or (inputs(197));
    layer0_outputs(2689) <= '0';
    layer0_outputs(2690) <= not((inputs(224)) xor (inputs(244)));
    layer0_outputs(2691) <= not(inputs(155)) or (inputs(219));
    layer0_outputs(2692) <= not(inputs(133)) or (inputs(127));
    layer0_outputs(2693) <= inputs(120);
    layer0_outputs(2694) <= (inputs(113)) or (inputs(54));
    layer0_outputs(2695) <= (inputs(202)) and not (inputs(103));
    layer0_outputs(2696) <= inputs(86);
    layer0_outputs(2697) <= '0';
    layer0_outputs(2698) <= (inputs(70)) and not (inputs(216));
    layer0_outputs(2699) <= not((inputs(70)) or (inputs(35)));
    layer0_outputs(2700) <= not((inputs(75)) xor (inputs(45)));
    layer0_outputs(2701) <= not(inputs(141)) or (inputs(48));
    layer0_outputs(2702) <= (inputs(254)) and not (inputs(228));
    layer0_outputs(2703) <= '0';
    layer0_outputs(2704) <= inputs(196);
    layer0_outputs(2705) <= not(inputs(225));
    layer0_outputs(2706) <= inputs(173);
    layer0_outputs(2707) <= (inputs(13)) and not (inputs(148));
    layer0_outputs(2708) <= not((inputs(118)) xor (inputs(70)));
    layer0_outputs(2709) <= not((inputs(220)) or (inputs(250)));
    layer0_outputs(2710) <= not(inputs(246)) or (inputs(144));
    layer0_outputs(2711) <= inputs(91);
    layer0_outputs(2712) <= not((inputs(232)) or (inputs(53)));
    layer0_outputs(2713) <= not((inputs(210)) or (inputs(147)));
    layer0_outputs(2714) <= (inputs(146)) and not (inputs(205));
    layer0_outputs(2715) <= (inputs(50)) or (inputs(223));
    layer0_outputs(2716) <= (inputs(54)) and not (inputs(115));
    layer0_outputs(2717) <= not(inputs(12));
    layer0_outputs(2718) <= not((inputs(105)) or (inputs(243)));
    layer0_outputs(2719) <= not((inputs(164)) or (inputs(213)));
    layer0_outputs(2720) <= not((inputs(123)) and (inputs(124)));
    layer0_outputs(2721) <= (inputs(250)) xor (inputs(187));
    layer0_outputs(2722) <= not((inputs(143)) xor (inputs(59)));
    layer0_outputs(2723) <= inputs(69);
    layer0_outputs(2724) <= not((inputs(188)) xor (inputs(195)));
    layer0_outputs(2725) <= not(inputs(54));
    layer0_outputs(2726) <= not((inputs(13)) or (inputs(171)));
    layer0_outputs(2727) <= not((inputs(28)) xor (inputs(132)));
    layer0_outputs(2728) <= not(inputs(217));
    layer0_outputs(2729) <= (inputs(148)) or (inputs(247));
    layer0_outputs(2730) <= not(inputs(12));
    layer0_outputs(2731) <= not(inputs(166));
    layer0_outputs(2732) <= inputs(53);
    layer0_outputs(2733) <= '0';
    layer0_outputs(2734) <= not((inputs(149)) and (inputs(29)));
    layer0_outputs(2735) <= (inputs(0)) xor (inputs(245));
    layer0_outputs(2736) <= inputs(102);
    layer0_outputs(2737) <= (inputs(70)) xor (inputs(242));
    layer0_outputs(2738) <= (inputs(38)) or (inputs(156));
    layer0_outputs(2739) <= not((inputs(240)) xor (inputs(92)));
    layer0_outputs(2740) <= not((inputs(5)) xor (inputs(131)));
    layer0_outputs(2741) <= (inputs(132)) xor (inputs(52));
    layer0_outputs(2742) <= inputs(246);
    layer0_outputs(2743) <= not((inputs(87)) or (inputs(132)));
    layer0_outputs(2744) <= (inputs(35)) xor (inputs(180));
    layer0_outputs(2745) <= not((inputs(203)) and (inputs(38)));
    layer0_outputs(2746) <= (inputs(115)) and not (inputs(207));
    layer0_outputs(2747) <= inputs(206);
    layer0_outputs(2748) <= not(inputs(154));
    layer0_outputs(2749) <= inputs(121);
    layer0_outputs(2750) <= not((inputs(14)) and (inputs(60)));
    layer0_outputs(2751) <= not(inputs(207));
    layer0_outputs(2752) <= inputs(100);
    layer0_outputs(2753) <= not(inputs(184)) or (inputs(195));
    layer0_outputs(2754) <= not(inputs(63)) or (inputs(65));
    layer0_outputs(2755) <= not(inputs(184));
    layer0_outputs(2756) <= (inputs(8)) or (inputs(150));
    layer0_outputs(2757) <= (inputs(92)) or (inputs(225));
    layer0_outputs(2758) <= inputs(56);
    layer0_outputs(2759) <= (inputs(86)) and not (inputs(128));
    layer0_outputs(2760) <= inputs(173);
    layer0_outputs(2761) <= '0';
    layer0_outputs(2762) <= not((inputs(156)) or (inputs(170)));
    layer0_outputs(2763) <= '0';
    layer0_outputs(2764) <= not((inputs(137)) or (inputs(251)));
    layer0_outputs(2765) <= not(inputs(168));
    layer0_outputs(2766) <= (inputs(85)) or (inputs(137));
    layer0_outputs(2767) <= not((inputs(200)) or (inputs(82)));
    layer0_outputs(2768) <= (inputs(201)) and not (inputs(190));
    layer0_outputs(2769) <= not(inputs(103)) or (inputs(149));
    layer0_outputs(2770) <= not((inputs(161)) or (inputs(216)));
    layer0_outputs(2771) <= not(inputs(121)) or (inputs(190));
    layer0_outputs(2772) <= '0';
    layer0_outputs(2773) <= inputs(161);
    layer0_outputs(2774) <= inputs(168);
    layer0_outputs(2775) <= not(inputs(115)) or (inputs(200));
    layer0_outputs(2776) <= inputs(230);
    layer0_outputs(2777) <= not(inputs(37));
    layer0_outputs(2778) <= not((inputs(163)) or (inputs(53)));
    layer0_outputs(2779) <= (inputs(83)) xor (inputs(79));
    layer0_outputs(2780) <= (inputs(179)) or (inputs(222));
    layer0_outputs(2781) <= not(inputs(137));
    layer0_outputs(2782) <= (inputs(6)) and not (inputs(25));
    layer0_outputs(2783) <= (inputs(67)) and (inputs(159));
    layer0_outputs(2784) <= not(inputs(148));
    layer0_outputs(2785) <= not((inputs(149)) xor (inputs(254)));
    layer0_outputs(2786) <= (inputs(27)) and not (inputs(242));
    layer0_outputs(2787) <= not(inputs(11)) or (inputs(15));
    layer0_outputs(2788) <= not(inputs(164)) or (inputs(159));
    layer0_outputs(2789) <= (inputs(95)) or (inputs(148));
    layer0_outputs(2790) <= not(inputs(164));
    layer0_outputs(2791) <= inputs(98);
    layer0_outputs(2792) <= inputs(168);
    layer0_outputs(2793) <= (inputs(253)) or (inputs(103));
    layer0_outputs(2794) <= not((inputs(2)) and (inputs(75)));
    layer0_outputs(2795) <= not(inputs(134)) or (inputs(41));
    layer0_outputs(2796) <= (inputs(150)) xor (inputs(159));
    layer0_outputs(2797) <= '1';
    layer0_outputs(2798) <= (inputs(136)) and not (inputs(62));
    layer0_outputs(2799) <= inputs(109);
    layer0_outputs(2800) <= (inputs(139)) xor (inputs(109));
    layer0_outputs(2801) <= (inputs(92)) and not (inputs(160));
    layer0_outputs(2802) <= (inputs(156)) xor (inputs(6));
    layer0_outputs(2803) <= inputs(44);
    layer0_outputs(2804) <= (inputs(223)) or (inputs(242));
    layer0_outputs(2805) <= not((inputs(76)) or (inputs(75)));
    layer0_outputs(2806) <= inputs(58);
    layer0_outputs(2807) <= not((inputs(116)) or (inputs(52)));
    layer0_outputs(2808) <= not(inputs(110)) or (inputs(175));
    layer0_outputs(2809) <= '1';
    layer0_outputs(2810) <= inputs(66);
    layer0_outputs(2811) <= not(inputs(203)) or (inputs(236));
    layer0_outputs(2812) <= (inputs(64)) and not (inputs(7));
    layer0_outputs(2813) <= (inputs(78)) and not (inputs(159));
    layer0_outputs(2814) <= (inputs(215)) and not (inputs(242));
    layer0_outputs(2815) <= not((inputs(40)) or (inputs(55)));
    layer0_outputs(2816) <= inputs(133);
    layer0_outputs(2817) <= not((inputs(83)) or (inputs(249)));
    layer0_outputs(2818) <= inputs(212);
    layer0_outputs(2819) <= not(inputs(60));
    layer0_outputs(2820) <= not(inputs(6)) or (inputs(188));
    layer0_outputs(2821) <= (inputs(116)) and not (inputs(9));
    layer0_outputs(2822) <= not((inputs(177)) xor (inputs(82)));
    layer0_outputs(2823) <= inputs(119);
    layer0_outputs(2824) <= not(inputs(152)) or (inputs(84));
    layer0_outputs(2825) <= not((inputs(245)) xor (inputs(34)));
    layer0_outputs(2826) <= inputs(167);
    layer0_outputs(2827) <= (inputs(81)) and not (inputs(35));
    layer0_outputs(2828) <= (inputs(216)) or (inputs(99));
    layer0_outputs(2829) <= not((inputs(179)) xor (inputs(244)));
    layer0_outputs(2830) <= inputs(118);
    layer0_outputs(2831) <= (inputs(88)) and not (inputs(6));
    layer0_outputs(2832) <= inputs(250);
    layer0_outputs(2833) <= (inputs(163)) or (inputs(78));
    layer0_outputs(2834) <= not((inputs(233)) or (inputs(118)));
    layer0_outputs(2835) <= inputs(224);
    layer0_outputs(2836) <= not(inputs(159));
    layer0_outputs(2837) <= (inputs(83)) and not (inputs(64));
    layer0_outputs(2838) <= (inputs(146)) and not (inputs(121));
    layer0_outputs(2839) <= not(inputs(38));
    layer0_outputs(2840) <= inputs(100);
    layer0_outputs(2841) <= (inputs(134)) and not (inputs(30));
    layer0_outputs(2842) <= not(inputs(95)) or (inputs(80));
    layer0_outputs(2843) <= (inputs(195)) or (inputs(177));
    layer0_outputs(2844) <= inputs(168);
    layer0_outputs(2845) <= not((inputs(31)) xor (inputs(93)));
    layer0_outputs(2846) <= not(inputs(199)) or (inputs(37));
    layer0_outputs(2847) <= not((inputs(159)) or (inputs(154)));
    layer0_outputs(2848) <= (inputs(23)) or (inputs(116));
    layer0_outputs(2849) <= (inputs(180)) and not (inputs(190));
    layer0_outputs(2850) <= '1';
    layer0_outputs(2851) <= (inputs(93)) and not (inputs(241));
    layer0_outputs(2852) <= not((inputs(161)) or (inputs(170)));
    layer0_outputs(2853) <= inputs(55);
    layer0_outputs(2854) <= not((inputs(141)) or (inputs(105)));
    layer0_outputs(2855) <= not((inputs(223)) or (inputs(211)));
    layer0_outputs(2856) <= not(inputs(221)) or (inputs(31));
    layer0_outputs(2857) <= not(inputs(70));
    layer0_outputs(2858) <= (inputs(70)) and not (inputs(227));
    layer0_outputs(2859) <= (inputs(45)) or (inputs(118));
    layer0_outputs(2860) <= not(inputs(108));
    layer0_outputs(2861) <= not(inputs(205));
    layer0_outputs(2862) <= not(inputs(56)) or (inputs(131));
    layer0_outputs(2863) <= not((inputs(98)) xor (inputs(64)));
    layer0_outputs(2864) <= not((inputs(81)) or (inputs(62)));
    layer0_outputs(2865) <= not((inputs(254)) or (inputs(15)));
    layer0_outputs(2866) <= not(inputs(112));
    layer0_outputs(2867) <= inputs(42);
    layer0_outputs(2868) <= not(inputs(71)) or (inputs(27));
    layer0_outputs(2869) <= inputs(219);
    layer0_outputs(2870) <= not(inputs(166)) or (inputs(98));
    layer0_outputs(2871) <= not(inputs(134)) or (inputs(191));
    layer0_outputs(2872) <= not(inputs(129));
    layer0_outputs(2873) <= not((inputs(92)) or (inputs(202)));
    layer0_outputs(2874) <= (inputs(101)) and (inputs(152));
    layer0_outputs(2875) <= (inputs(124)) or (inputs(34));
    layer0_outputs(2876) <= inputs(59);
    layer0_outputs(2877) <= inputs(191);
    layer0_outputs(2878) <= not(inputs(226));
    layer0_outputs(2879) <= (inputs(165)) xor (inputs(182));
    layer0_outputs(2880) <= not(inputs(241)) or (inputs(24));
    layer0_outputs(2881) <= not((inputs(115)) xor (inputs(38)));
    layer0_outputs(2882) <= (inputs(122)) and not (inputs(169));
    layer0_outputs(2883) <= (inputs(203)) xor (inputs(19));
    layer0_outputs(2884) <= not((inputs(13)) or (inputs(164)));
    layer0_outputs(2885) <= not((inputs(67)) or (inputs(137)));
    layer0_outputs(2886) <= not((inputs(202)) and (inputs(252)));
    layer0_outputs(2887) <= (inputs(207)) or (inputs(85));
    layer0_outputs(2888) <= (inputs(59)) or (inputs(161));
    layer0_outputs(2889) <= not((inputs(206)) and (inputs(62)));
    layer0_outputs(2890) <= not((inputs(227)) and (inputs(193)));
    layer0_outputs(2891) <= inputs(96);
    layer0_outputs(2892) <= (inputs(140)) or (inputs(189));
    layer0_outputs(2893) <= not(inputs(107)) or (inputs(244));
    layer0_outputs(2894) <= (inputs(76)) or (inputs(15));
    layer0_outputs(2895) <= not((inputs(79)) and (inputs(221)));
    layer0_outputs(2896) <= not((inputs(248)) and (inputs(141)));
    layer0_outputs(2897) <= not(inputs(156));
    layer0_outputs(2898) <= '1';
    layer0_outputs(2899) <= (inputs(32)) xor (inputs(42));
    layer0_outputs(2900) <= not((inputs(127)) xor (inputs(47)));
    layer0_outputs(2901) <= not(inputs(140));
    layer0_outputs(2902) <= (inputs(133)) or (inputs(62));
    layer0_outputs(2903) <= not(inputs(230)) or (inputs(159));
    layer0_outputs(2904) <= (inputs(231)) and not (inputs(219));
    layer0_outputs(2905) <= inputs(84);
    layer0_outputs(2906) <= not(inputs(65)) or (inputs(55));
    layer0_outputs(2907) <= not((inputs(140)) or (inputs(170)));
    layer0_outputs(2908) <= inputs(251);
    layer0_outputs(2909) <= inputs(214);
    layer0_outputs(2910) <= (inputs(154)) and not (inputs(3));
    layer0_outputs(2911) <= not((inputs(47)) and (inputs(130)));
    layer0_outputs(2912) <= not(inputs(119));
    layer0_outputs(2913) <= not((inputs(210)) xor (inputs(74)));
    layer0_outputs(2914) <= not((inputs(88)) or (inputs(227)));
    layer0_outputs(2915) <= not(inputs(97));
    layer0_outputs(2916) <= inputs(101);
    layer0_outputs(2917) <= (inputs(211)) and not (inputs(56));
    layer0_outputs(2918) <= not(inputs(88));
    layer0_outputs(2919) <= not(inputs(107)) or (inputs(8));
    layer0_outputs(2920) <= (inputs(182)) and not (inputs(83));
    layer0_outputs(2921) <= (inputs(140)) or (inputs(25));
    layer0_outputs(2922) <= (inputs(42)) and not (inputs(213));
    layer0_outputs(2923) <= inputs(177);
    layer0_outputs(2924) <= not((inputs(243)) xor (inputs(108)));
    layer0_outputs(2925) <= not(inputs(196));
    layer0_outputs(2926) <= not(inputs(43)) or (inputs(243));
    layer0_outputs(2927) <= (inputs(190)) or (inputs(253));
    layer0_outputs(2928) <= not((inputs(39)) or (inputs(91)));
    layer0_outputs(2929) <= not((inputs(171)) or (inputs(123)));
    layer0_outputs(2930) <= '0';
    layer0_outputs(2931) <= not((inputs(184)) or (inputs(235)));
    layer0_outputs(2932) <= (inputs(126)) xor (inputs(159));
    layer0_outputs(2933) <= not(inputs(148));
    layer0_outputs(2934) <= not(inputs(42));
    layer0_outputs(2935) <= not((inputs(155)) xor (inputs(112)));
    layer0_outputs(2936) <= not((inputs(30)) or (inputs(117)));
    layer0_outputs(2937) <= not(inputs(70));
    layer0_outputs(2938) <= (inputs(8)) and (inputs(98));
    layer0_outputs(2939) <= not(inputs(204));
    layer0_outputs(2940) <= not(inputs(9)) or (inputs(18));
    layer0_outputs(2941) <= not((inputs(177)) xor (inputs(129)));
    layer0_outputs(2942) <= not((inputs(218)) xor (inputs(212)));
    layer0_outputs(2943) <= not(inputs(105)) or (inputs(155));
    layer0_outputs(2944) <= not((inputs(104)) xor (inputs(254)));
    layer0_outputs(2945) <= (inputs(149)) and not (inputs(67));
    layer0_outputs(2946) <= (inputs(160)) and not (inputs(174));
    layer0_outputs(2947) <= (inputs(195)) or (inputs(124));
    layer0_outputs(2948) <= not(inputs(157)) or (inputs(229));
    layer0_outputs(2949) <= not(inputs(14));
    layer0_outputs(2950) <= (inputs(154)) xor (inputs(53));
    layer0_outputs(2951) <= not((inputs(140)) and (inputs(189)));
    layer0_outputs(2952) <= not(inputs(118)) or (inputs(100));
    layer0_outputs(2953) <= (inputs(142)) xor (inputs(60));
    layer0_outputs(2954) <= not((inputs(126)) or (inputs(75)));
    layer0_outputs(2955) <= (inputs(225)) xor (inputs(210));
    layer0_outputs(2956) <= not(inputs(97));
    layer0_outputs(2957) <= not((inputs(66)) or (inputs(40)));
    layer0_outputs(2958) <= not(inputs(238));
    layer0_outputs(2959) <= (inputs(89)) or (inputs(36));
    layer0_outputs(2960) <= (inputs(66)) or (inputs(205));
    layer0_outputs(2961) <= inputs(136);
    layer0_outputs(2962) <= inputs(64);
    layer0_outputs(2963) <= inputs(184);
    layer0_outputs(2964) <= not(inputs(230));
    layer0_outputs(2965) <= (inputs(36)) and not (inputs(131));
    layer0_outputs(2966) <= not(inputs(86));
    layer0_outputs(2967) <= (inputs(238)) or (inputs(20));
    layer0_outputs(2968) <= (inputs(248)) and not (inputs(208));
    layer0_outputs(2969) <= (inputs(245)) and (inputs(70));
    layer0_outputs(2970) <= (inputs(218)) or (inputs(100));
    layer0_outputs(2971) <= (inputs(170)) xor (inputs(239));
    layer0_outputs(2972) <= (inputs(229)) or (inputs(74));
    layer0_outputs(2973) <= not(inputs(184)) or (inputs(229));
    layer0_outputs(2974) <= (inputs(182)) xor (inputs(164));
    layer0_outputs(2975) <= not((inputs(173)) or (inputs(24)));
    layer0_outputs(2976) <= not(inputs(52));
    layer0_outputs(2977) <= not((inputs(180)) and (inputs(91)));
    layer0_outputs(2978) <= '0';
    layer0_outputs(2979) <= (inputs(135)) or (inputs(150));
    layer0_outputs(2980) <= (inputs(79)) or (inputs(145));
    layer0_outputs(2981) <= '0';
    layer0_outputs(2982) <= (inputs(95)) and not (inputs(248));
    layer0_outputs(2983) <= inputs(213);
    layer0_outputs(2984) <= '0';
    layer0_outputs(2985) <= '1';
    layer0_outputs(2986) <= (inputs(132)) and not (inputs(191));
    layer0_outputs(2987) <= not(inputs(201)) or (inputs(36));
    layer0_outputs(2988) <= not((inputs(73)) xor (inputs(128)));
    layer0_outputs(2989) <= not(inputs(195));
    layer0_outputs(2990) <= (inputs(184)) xor (inputs(90));
    layer0_outputs(2991) <= not((inputs(227)) xor (inputs(9)));
    layer0_outputs(2992) <= (inputs(103)) or (inputs(62));
    layer0_outputs(2993) <= '0';
    layer0_outputs(2994) <= not((inputs(37)) xor (inputs(4)));
    layer0_outputs(2995) <= (inputs(185)) or (inputs(11));
    layer0_outputs(2996) <= (inputs(187)) xor (inputs(24));
    layer0_outputs(2997) <= (inputs(163)) or (inputs(77));
    layer0_outputs(2998) <= (inputs(226)) xor (inputs(86));
    layer0_outputs(2999) <= (inputs(152)) or (inputs(8));
    layer0_outputs(3000) <= not(inputs(86));
    layer0_outputs(3001) <= not((inputs(155)) or (inputs(65)));
    layer0_outputs(3002) <= not((inputs(243)) and (inputs(193)));
    layer0_outputs(3003) <= (inputs(142)) xor (inputs(41));
    layer0_outputs(3004) <= (inputs(229)) and not (inputs(25));
    layer0_outputs(3005) <= not(inputs(120));
    layer0_outputs(3006) <= inputs(173);
    layer0_outputs(3007) <= (inputs(156)) and not (inputs(149));
    layer0_outputs(3008) <= not(inputs(217)) or (inputs(33));
    layer0_outputs(3009) <= not(inputs(233)) or (inputs(191));
    layer0_outputs(3010) <= not(inputs(125)) or (inputs(239));
    layer0_outputs(3011) <= (inputs(29)) or (inputs(123));
    layer0_outputs(3012) <= not((inputs(31)) xor (inputs(218)));
    layer0_outputs(3013) <= not(inputs(198));
    layer0_outputs(3014) <= (inputs(231)) xor (inputs(33));
    layer0_outputs(3015) <= (inputs(36)) or (inputs(132));
    layer0_outputs(3016) <= inputs(203);
    layer0_outputs(3017) <= not((inputs(181)) or (inputs(23)));
    layer0_outputs(3018) <= '0';
    layer0_outputs(3019) <= '1';
    layer0_outputs(3020) <= (inputs(200)) and not (inputs(85));
    layer0_outputs(3021) <= not(inputs(253)) or (inputs(129));
    layer0_outputs(3022) <= not(inputs(200));
    layer0_outputs(3023) <= inputs(107);
    layer0_outputs(3024) <= not((inputs(198)) or (inputs(213)));
    layer0_outputs(3025) <= not(inputs(180)) or (inputs(226));
    layer0_outputs(3026) <= (inputs(50)) xor (inputs(64));
    layer0_outputs(3027) <= (inputs(184)) xor (inputs(50));
    layer0_outputs(3028) <= (inputs(228)) or (inputs(226));
    layer0_outputs(3029) <= (inputs(199)) or (inputs(21));
    layer0_outputs(3030) <= inputs(124);
    layer0_outputs(3031) <= (inputs(208)) xor (inputs(4));
    layer0_outputs(3032) <= '0';
    layer0_outputs(3033) <= (inputs(132)) and not (inputs(126));
    layer0_outputs(3034) <= not((inputs(146)) or (inputs(106)));
    layer0_outputs(3035) <= '1';
    layer0_outputs(3036) <= not((inputs(7)) xor (inputs(73)));
    layer0_outputs(3037) <= not(inputs(69)) or (inputs(241));
    layer0_outputs(3038) <= not((inputs(213)) or (inputs(49)));
    layer0_outputs(3039) <= (inputs(112)) or (inputs(151));
    layer0_outputs(3040) <= not(inputs(105));
    layer0_outputs(3041) <= not((inputs(8)) xor (inputs(119)));
    layer0_outputs(3042) <= not((inputs(46)) xor (inputs(70)));
    layer0_outputs(3043) <= (inputs(9)) xor (inputs(182));
    layer0_outputs(3044) <= not(inputs(90));
    layer0_outputs(3045) <= not((inputs(106)) or (inputs(94)));
    layer0_outputs(3046) <= inputs(167);
    layer0_outputs(3047) <= (inputs(130)) or (inputs(147));
    layer0_outputs(3048) <= inputs(210);
    layer0_outputs(3049) <= '0';
    layer0_outputs(3050) <= (inputs(72)) xor (inputs(255));
    layer0_outputs(3051) <= not(inputs(137)) or (inputs(62));
    layer0_outputs(3052) <= not((inputs(179)) xor (inputs(34)));
    layer0_outputs(3053) <= not((inputs(131)) or (inputs(228)));
    layer0_outputs(3054) <= not(inputs(236));
    layer0_outputs(3055) <= (inputs(106)) xor (inputs(226));
    layer0_outputs(3056) <= (inputs(233)) and not (inputs(211));
    layer0_outputs(3057) <= not((inputs(160)) or (inputs(110)));
    layer0_outputs(3058) <= not((inputs(225)) xor (inputs(37)));
    layer0_outputs(3059) <= not((inputs(181)) or (inputs(220)));
    layer0_outputs(3060) <= not(inputs(164));
    layer0_outputs(3061) <= not((inputs(224)) or (inputs(18)));
    layer0_outputs(3062) <= (inputs(41)) or (inputs(197));
    layer0_outputs(3063) <= not((inputs(173)) or (inputs(68)));
    layer0_outputs(3064) <= (inputs(15)) xor (inputs(1));
    layer0_outputs(3065) <= not(inputs(86));
    layer0_outputs(3066) <= not((inputs(65)) or (inputs(99)));
    layer0_outputs(3067) <= (inputs(174)) xor (inputs(191));
    layer0_outputs(3068) <= not(inputs(166));
    layer0_outputs(3069) <= (inputs(66)) or (inputs(55));
    layer0_outputs(3070) <= not(inputs(230));
    layer0_outputs(3071) <= not(inputs(119));
    layer0_outputs(3072) <= not(inputs(217)) or (inputs(192));
    layer0_outputs(3073) <= not(inputs(136));
    layer0_outputs(3074) <= not((inputs(226)) and (inputs(99)));
    layer0_outputs(3075) <= not(inputs(185)) or (inputs(25));
    layer0_outputs(3076) <= '1';
    layer0_outputs(3077) <= inputs(4);
    layer0_outputs(3078) <= inputs(151);
    layer0_outputs(3079) <= (inputs(90)) and not (inputs(177));
    layer0_outputs(3080) <= not((inputs(230)) or (inputs(172)));
    layer0_outputs(3081) <= not(inputs(38));
    layer0_outputs(3082) <= (inputs(204)) and (inputs(164));
    layer0_outputs(3083) <= not((inputs(221)) and (inputs(109)));
    layer0_outputs(3084) <= not(inputs(90)) or (inputs(254));
    layer0_outputs(3085) <= inputs(181);
    layer0_outputs(3086) <= not(inputs(21)) or (inputs(8));
    layer0_outputs(3087) <= not(inputs(52)) or (inputs(19));
    layer0_outputs(3088) <= (inputs(5)) or (inputs(233));
    layer0_outputs(3089) <= (inputs(61)) or (inputs(232));
    layer0_outputs(3090) <= not(inputs(125));
    layer0_outputs(3091) <= (inputs(195)) or (inputs(156));
    layer0_outputs(3092) <= '1';
    layer0_outputs(3093) <= not(inputs(93)) or (inputs(219));
    layer0_outputs(3094) <= (inputs(57)) or (inputs(178));
    layer0_outputs(3095) <= inputs(120);
    layer0_outputs(3096) <= not(inputs(25)) or (inputs(49));
    layer0_outputs(3097) <= not(inputs(150)) or (inputs(174));
    layer0_outputs(3098) <= inputs(139);
    layer0_outputs(3099) <= not(inputs(79));
    layer0_outputs(3100) <= not((inputs(123)) or (inputs(183)));
    layer0_outputs(3101) <= inputs(201);
    layer0_outputs(3102) <= (inputs(3)) or (inputs(41));
    layer0_outputs(3103) <= (inputs(150)) and not (inputs(214));
    layer0_outputs(3104) <= not((inputs(1)) or (inputs(198)));
    layer0_outputs(3105) <= inputs(117);
    layer0_outputs(3106) <= '0';
    layer0_outputs(3107) <= '1';
    layer0_outputs(3108) <= (inputs(249)) xor (inputs(68));
    layer0_outputs(3109) <= inputs(255);
    layer0_outputs(3110) <= (inputs(194)) xor (inputs(207));
    layer0_outputs(3111) <= not((inputs(206)) and (inputs(67)));
    layer0_outputs(3112) <= not((inputs(177)) or (inputs(228)));
    layer0_outputs(3113) <= (inputs(62)) xor (inputs(82));
    layer0_outputs(3114) <= (inputs(212)) xor (inputs(250));
    layer0_outputs(3115) <= not((inputs(174)) or (inputs(6)));
    layer0_outputs(3116) <= not(inputs(250));
    layer0_outputs(3117) <= not(inputs(171)) or (inputs(255));
    layer0_outputs(3118) <= inputs(197);
    layer0_outputs(3119) <= (inputs(211)) xor (inputs(156));
    layer0_outputs(3120) <= (inputs(232)) and not (inputs(209));
    layer0_outputs(3121) <= '1';
    layer0_outputs(3122) <= (inputs(52)) xor (inputs(81));
    layer0_outputs(3123) <= (inputs(118)) xor (inputs(38));
    layer0_outputs(3124) <= (inputs(168)) xor (inputs(105));
    layer0_outputs(3125) <= not(inputs(212));
    layer0_outputs(3126) <= (inputs(196)) xor (inputs(54));
    layer0_outputs(3127) <= (inputs(68)) and not (inputs(37));
    layer0_outputs(3128) <= (inputs(104)) and not (inputs(77));
    layer0_outputs(3129) <= (inputs(86)) and not (inputs(20));
    layer0_outputs(3130) <= not((inputs(169)) or (inputs(26)));
    layer0_outputs(3131) <= (inputs(19)) or (inputs(190));
    layer0_outputs(3132) <= not(inputs(152));
    layer0_outputs(3133) <= not(inputs(134)) or (inputs(28));
    layer0_outputs(3134) <= not((inputs(248)) or (inputs(174)));
    layer0_outputs(3135) <= not(inputs(5));
    layer0_outputs(3136) <= (inputs(162)) and not (inputs(28));
    layer0_outputs(3137) <= not(inputs(78)) or (inputs(36));
    layer0_outputs(3138) <= not((inputs(83)) and (inputs(184)));
    layer0_outputs(3139) <= (inputs(76)) or (inputs(190));
    layer0_outputs(3140) <= (inputs(199)) or (inputs(113));
    layer0_outputs(3141) <= not(inputs(104)) or (inputs(29));
    layer0_outputs(3142) <= (inputs(242)) xor (inputs(41));
    layer0_outputs(3143) <= not(inputs(186)) or (inputs(27));
    layer0_outputs(3144) <= (inputs(118)) and (inputs(135));
    layer0_outputs(3145) <= (inputs(125)) and not (inputs(253));
    layer0_outputs(3146) <= inputs(210);
    layer0_outputs(3147) <= not((inputs(144)) xor (inputs(121)));
    layer0_outputs(3148) <= (inputs(215)) and not (inputs(45));
    layer0_outputs(3149) <= not((inputs(110)) or (inputs(97)));
    layer0_outputs(3150) <= not(inputs(51));
    layer0_outputs(3151) <= not((inputs(14)) and (inputs(179)));
    layer0_outputs(3152) <= not(inputs(214)) or (inputs(69));
    layer0_outputs(3153) <= (inputs(172)) or (inputs(17));
    layer0_outputs(3154) <= '0';
    layer0_outputs(3155) <= not(inputs(208)) or (inputs(85));
    layer0_outputs(3156) <= not(inputs(31));
    layer0_outputs(3157) <= inputs(151);
    layer0_outputs(3158) <= (inputs(33)) and not (inputs(94));
    layer0_outputs(3159) <= (inputs(223)) or (inputs(23));
    layer0_outputs(3160) <= (inputs(96)) xor (inputs(180));
    layer0_outputs(3161) <= not(inputs(27));
    layer0_outputs(3162) <= not(inputs(193));
    layer0_outputs(3163) <= inputs(197);
    layer0_outputs(3164) <= not(inputs(114)) or (inputs(27));
    layer0_outputs(3165) <= inputs(149);
    layer0_outputs(3166) <= not(inputs(18)) or (inputs(127));
    layer0_outputs(3167) <= '0';
    layer0_outputs(3168) <= (inputs(24)) and not (inputs(95));
    layer0_outputs(3169) <= inputs(102);
    layer0_outputs(3170) <= inputs(245);
    layer0_outputs(3171) <= (inputs(13)) and not (inputs(146));
    layer0_outputs(3172) <= not(inputs(226)) or (inputs(16));
    layer0_outputs(3173) <= not(inputs(19));
    layer0_outputs(3174) <= (inputs(252)) xor (inputs(229));
    layer0_outputs(3175) <= not((inputs(133)) xor (inputs(96)));
    layer0_outputs(3176) <= not(inputs(178));
    layer0_outputs(3177) <= inputs(78);
    layer0_outputs(3178) <= (inputs(174)) or (inputs(140));
    layer0_outputs(3179) <= inputs(36);
    layer0_outputs(3180) <= (inputs(185)) and not (inputs(238));
    layer0_outputs(3181) <= not((inputs(199)) or (inputs(187)));
    layer0_outputs(3182) <= inputs(216);
    layer0_outputs(3183) <= not((inputs(58)) xor (inputs(55)));
    layer0_outputs(3184) <= (inputs(77)) and not (inputs(247));
    layer0_outputs(3185) <= inputs(149);
    layer0_outputs(3186) <= '0';
    layer0_outputs(3187) <= (inputs(71)) xor (inputs(173));
    layer0_outputs(3188) <= not((inputs(223)) and (inputs(0)));
    layer0_outputs(3189) <= not((inputs(141)) or (inputs(147)));
    layer0_outputs(3190) <= '1';
    layer0_outputs(3191) <= (inputs(224)) and not (inputs(63));
    layer0_outputs(3192) <= (inputs(183)) and not (inputs(211));
    layer0_outputs(3193) <= not(inputs(202));
    layer0_outputs(3194) <= not(inputs(178));
    layer0_outputs(3195) <= '1';
    layer0_outputs(3196) <= (inputs(202)) xor (inputs(185));
    layer0_outputs(3197) <= not(inputs(36)) or (inputs(24));
    layer0_outputs(3198) <= (inputs(76)) and not (inputs(244));
    layer0_outputs(3199) <= not(inputs(57));
    layer0_outputs(3200) <= not(inputs(165));
    layer0_outputs(3201) <= not(inputs(217));
    layer0_outputs(3202) <= not(inputs(66)) or (inputs(204));
    layer0_outputs(3203) <= not((inputs(3)) xor (inputs(76)));
    layer0_outputs(3204) <= (inputs(105)) or (inputs(142));
    layer0_outputs(3205) <= not(inputs(242)) or (inputs(254));
    layer0_outputs(3206) <= (inputs(178)) or (inputs(159));
    layer0_outputs(3207) <= (inputs(255)) and not (inputs(226));
    layer0_outputs(3208) <= (inputs(163)) and not (inputs(67));
    layer0_outputs(3209) <= (inputs(207)) and not (inputs(2));
    layer0_outputs(3210) <= inputs(212);
    layer0_outputs(3211) <= inputs(151);
    layer0_outputs(3212) <= (inputs(185)) or (inputs(190));
    layer0_outputs(3213) <= (inputs(21)) and not (inputs(40));
    layer0_outputs(3214) <= inputs(142);
    layer0_outputs(3215) <= '0';
    layer0_outputs(3216) <= (inputs(86)) or (inputs(247));
    layer0_outputs(3217) <= (inputs(154)) xor (inputs(69));
    layer0_outputs(3218) <= not((inputs(93)) or (inputs(189)));
    layer0_outputs(3219) <= (inputs(200)) and not (inputs(36));
    layer0_outputs(3220) <= (inputs(59)) xor (inputs(71));
    layer0_outputs(3221) <= '0';
    layer0_outputs(3222) <= (inputs(213)) and not (inputs(188));
    layer0_outputs(3223) <= not((inputs(117)) or (inputs(17)));
    layer0_outputs(3224) <= not((inputs(140)) or (inputs(184)));
    layer0_outputs(3225) <= not(inputs(136));
    layer0_outputs(3226) <= not(inputs(143));
    layer0_outputs(3227) <= inputs(197);
    layer0_outputs(3228) <= inputs(47);
    layer0_outputs(3229) <= inputs(43);
    layer0_outputs(3230) <= not((inputs(128)) or (inputs(125)));
    layer0_outputs(3231) <= '0';
    layer0_outputs(3232) <= not((inputs(160)) or (inputs(23)));
    layer0_outputs(3233) <= inputs(74);
    layer0_outputs(3234) <= not((inputs(43)) and (inputs(254)));
    layer0_outputs(3235) <= not(inputs(196));
    layer0_outputs(3236) <= (inputs(187)) and not (inputs(229));
    layer0_outputs(3237) <= (inputs(214)) and not (inputs(51));
    layer0_outputs(3238) <= (inputs(30)) or (inputs(231));
    layer0_outputs(3239) <= not((inputs(85)) xor (inputs(249)));
    layer0_outputs(3240) <= (inputs(92)) and not (inputs(1));
    layer0_outputs(3241) <= not(inputs(139)) or (inputs(97));
    layer0_outputs(3242) <= (inputs(195)) or (inputs(209));
    layer0_outputs(3243) <= not((inputs(233)) or (inputs(221)));
    layer0_outputs(3244) <= inputs(191);
    layer0_outputs(3245) <= not((inputs(8)) xor (inputs(128)));
    layer0_outputs(3246) <= not((inputs(128)) xor (inputs(123)));
    layer0_outputs(3247) <= not((inputs(222)) xor (inputs(51)));
    layer0_outputs(3248) <= not(inputs(93));
    layer0_outputs(3249) <= not(inputs(155));
    layer0_outputs(3250) <= not((inputs(107)) xor (inputs(105)));
    layer0_outputs(3251) <= not((inputs(199)) xor (inputs(50)));
    layer0_outputs(3252) <= not((inputs(10)) or (inputs(28)));
    layer0_outputs(3253) <= not(inputs(177));
    layer0_outputs(3254) <= inputs(144);
    layer0_outputs(3255) <= not(inputs(183));
    layer0_outputs(3256) <= inputs(149);
    layer0_outputs(3257) <= not((inputs(187)) xor (inputs(71)));
    layer0_outputs(3258) <= not(inputs(199)) or (inputs(161));
    layer0_outputs(3259) <= (inputs(142)) and (inputs(49));
    layer0_outputs(3260) <= (inputs(255)) or (inputs(202));
    layer0_outputs(3261) <= (inputs(125)) or (inputs(108));
    layer0_outputs(3262) <= (inputs(82)) and not (inputs(209));
    layer0_outputs(3263) <= not(inputs(25));
    layer0_outputs(3264) <= not((inputs(150)) or (inputs(21)));
    layer0_outputs(3265) <= (inputs(37)) or (inputs(57));
    layer0_outputs(3266) <= inputs(22);
    layer0_outputs(3267) <= (inputs(168)) and not (inputs(48));
    layer0_outputs(3268) <= not(inputs(86)) or (inputs(173));
    layer0_outputs(3269) <= inputs(105);
    layer0_outputs(3270) <= (inputs(216)) and not (inputs(9));
    layer0_outputs(3271) <= not((inputs(13)) and (inputs(240)));
    layer0_outputs(3272) <= not(inputs(38)) or (inputs(241));
    layer0_outputs(3273) <= (inputs(14)) and not (inputs(26));
    layer0_outputs(3274) <= inputs(87);
    layer0_outputs(3275) <= inputs(208);
    layer0_outputs(3276) <= (inputs(129)) or (inputs(186));
    layer0_outputs(3277) <= (inputs(20)) or (inputs(88));
    layer0_outputs(3278) <= (inputs(235)) or (inputs(115));
    layer0_outputs(3279) <= (inputs(138)) xor (inputs(108));
    layer0_outputs(3280) <= (inputs(37)) xor (inputs(234));
    layer0_outputs(3281) <= (inputs(215)) and not (inputs(20));
    layer0_outputs(3282) <= not(inputs(63));
    layer0_outputs(3283) <= (inputs(140)) xor (inputs(10));
    layer0_outputs(3284) <= '1';
    layer0_outputs(3285) <= not((inputs(28)) xor (inputs(239)));
    layer0_outputs(3286) <= not(inputs(103));
    layer0_outputs(3287) <= not(inputs(134));
    layer0_outputs(3288) <= not((inputs(178)) or (inputs(174)));
    layer0_outputs(3289) <= inputs(108);
    layer0_outputs(3290) <= inputs(29);
    layer0_outputs(3291) <= (inputs(156)) or (inputs(97));
    layer0_outputs(3292) <= (inputs(196)) or (inputs(197));
    layer0_outputs(3293) <= inputs(164);
    layer0_outputs(3294) <= not(inputs(160));
    layer0_outputs(3295) <= not(inputs(44)) or (inputs(176));
    layer0_outputs(3296) <= not((inputs(110)) xor (inputs(11)));
    layer0_outputs(3297) <= not((inputs(242)) xor (inputs(72)));
    layer0_outputs(3298) <= not((inputs(152)) and (inputs(141)));
    layer0_outputs(3299) <= not((inputs(100)) xor (inputs(70)));
    layer0_outputs(3300) <= not((inputs(33)) xor (inputs(30)));
    layer0_outputs(3301) <= not(inputs(59)) or (inputs(29));
    layer0_outputs(3302) <= not((inputs(147)) xor (inputs(24)));
    layer0_outputs(3303) <= not(inputs(12));
    layer0_outputs(3304) <= (inputs(86)) and not (inputs(57));
    layer0_outputs(3305) <= '1';
    layer0_outputs(3306) <= inputs(102);
    layer0_outputs(3307) <= inputs(20);
    layer0_outputs(3308) <= (inputs(86)) xor (inputs(117));
    layer0_outputs(3309) <= not(inputs(27));
    layer0_outputs(3310) <= not(inputs(137));
    layer0_outputs(3311) <= inputs(73);
    layer0_outputs(3312) <= not(inputs(85));
    layer0_outputs(3313) <= '1';
    layer0_outputs(3314) <= (inputs(191)) and not (inputs(33));
    layer0_outputs(3315) <= not((inputs(130)) and (inputs(162)));
    layer0_outputs(3316) <= inputs(53);
    layer0_outputs(3317) <= (inputs(98)) and (inputs(226));
    layer0_outputs(3318) <= (inputs(40)) xor (inputs(30));
    layer0_outputs(3319) <= (inputs(95)) or (inputs(83));
    layer0_outputs(3320) <= (inputs(65)) and not (inputs(78));
    layer0_outputs(3321) <= (inputs(45)) xor (inputs(36));
    layer0_outputs(3322) <= (inputs(49)) xor (inputs(61));
    layer0_outputs(3323) <= (inputs(177)) and not (inputs(239));
    layer0_outputs(3324) <= not(inputs(118)) or (inputs(2));
    layer0_outputs(3325) <= (inputs(17)) and (inputs(31));
    layer0_outputs(3326) <= inputs(158);
    layer0_outputs(3327) <= not((inputs(250)) or (inputs(25)));
    layer0_outputs(3328) <= inputs(186);
    layer0_outputs(3329) <= (inputs(83)) or (inputs(192));
    layer0_outputs(3330) <= not((inputs(118)) or (inputs(110)));
    layer0_outputs(3331) <= not((inputs(139)) or (inputs(10)));
    layer0_outputs(3332) <= inputs(41);
    layer0_outputs(3333) <= (inputs(143)) and (inputs(20));
    layer0_outputs(3334) <= not((inputs(52)) xor (inputs(65)));
    layer0_outputs(3335) <= (inputs(253)) or (inputs(85));
    layer0_outputs(3336) <= (inputs(117)) and not (inputs(247));
    layer0_outputs(3337) <= not(inputs(169));
    layer0_outputs(3338) <= (inputs(108)) and not (inputs(64));
    layer0_outputs(3339) <= not((inputs(209)) xor (inputs(151)));
    layer0_outputs(3340) <= not(inputs(210)) or (inputs(68));
    layer0_outputs(3341) <= not(inputs(74));
    layer0_outputs(3342) <= inputs(125);
    layer0_outputs(3343) <= not((inputs(159)) xor (inputs(142)));
    layer0_outputs(3344) <= (inputs(101)) xor (inputs(223));
    layer0_outputs(3345) <= (inputs(175)) xor (inputs(116));
    layer0_outputs(3346) <= not(inputs(77));
    layer0_outputs(3347) <= not((inputs(171)) xor (inputs(71)));
    layer0_outputs(3348) <= not(inputs(236)) or (inputs(33));
    layer0_outputs(3349) <= (inputs(209)) xor (inputs(238));
    layer0_outputs(3350) <= (inputs(217)) xor (inputs(78));
    layer0_outputs(3351) <= '1';
    layer0_outputs(3352) <= (inputs(14)) xor (inputs(235));
    layer0_outputs(3353) <= (inputs(230)) or (inputs(113));
    layer0_outputs(3354) <= (inputs(1)) and (inputs(28));
    layer0_outputs(3355) <= not(inputs(239)) or (inputs(39));
    layer0_outputs(3356) <= inputs(63);
    layer0_outputs(3357) <= not(inputs(230));
    layer0_outputs(3358) <= (inputs(67)) or (inputs(149));
    layer0_outputs(3359) <= not((inputs(122)) or (inputs(35)));
    layer0_outputs(3360) <= not(inputs(228));
    layer0_outputs(3361) <= (inputs(156)) or (inputs(141));
    layer0_outputs(3362) <= (inputs(145)) or (inputs(250));
    layer0_outputs(3363) <= not((inputs(191)) and (inputs(108)));
    layer0_outputs(3364) <= (inputs(188)) xor (inputs(79));
    layer0_outputs(3365) <= not((inputs(194)) or (inputs(119)));
    layer0_outputs(3366) <= not((inputs(111)) or (inputs(50)));
    layer0_outputs(3367) <= (inputs(65)) or (inputs(158));
    layer0_outputs(3368) <= not((inputs(226)) xor (inputs(87)));
    layer0_outputs(3369) <= inputs(58);
    layer0_outputs(3370) <= (inputs(229)) xor (inputs(139));
    layer0_outputs(3371) <= inputs(166);
    layer0_outputs(3372) <= not((inputs(78)) xor (inputs(3)));
    layer0_outputs(3373) <= '1';
    layer0_outputs(3374) <= not(inputs(192)) or (inputs(240));
    layer0_outputs(3375) <= (inputs(55)) and not (inputs(235));
    layer0_outputs(3376) <= not((inputs(215)) or (inputs(246)));
    layer0_outputs(3377) <= inputs(250);
    layer0_outputs(3378) <= not(inputs(135));
    layer0_outputs(3379) <= not(inputs(110));
    layer0_outputs(3380) <= not(inputs(187)) or (inputs(215));
    layer0_outputs(3381) <= not((inputs(93)) or (inputs(248)));
    layer0_outputs(3382) <= not(inputs(194));
    layer0_outputs(3383) <= not((inputs(162)) or (inputs(51)));
    layer0_outputs(3384) <= inputs(148);
    layer0_outputs(3385) <= inputs(16);
    layer0_outputs(3386) <= (inputs(176)) and (inputs(52));
    layer0_outputs(3387) <= not(inputs(248));
    layer0_outputs(3388) <= not((inputs(215)) or (inputs(99)));
    layer0_outputs(3389) <= not((inputs(101)) or (inputs(60)));
    layer0_outputs(3390) <= not((inputs(169)) or (inputs(51)));
    layer0_outputs(3391) <= not(inputs(24)) or (inputs(189));
    layer0_outputs(3392) <= (inputs(107)) and not (inputs(243));
    layer0_outputs(3393) <= inputs(3);
    layer0_outputs(3394) <= (inputs(223)) xor (inputs(102));
    layer0_outputs(3395) <= not(inputs(58)) or (inputs(24));
    layer0_outputs(3396) <= (inputs(117)) or (inputs(224));
    layer0_outputs(3397) <= '1';
    layer0_outputs(3398) <= not(inputs(89));
    layer0_outputs(3399) <= inputs(231);
    layer0_outputs(3400) <= not(inputs(182)) or (inputs(108));
    layer0_outputs(3401) <= '1';
    layer0_outputs(3402) <= not((inputs(121)) xor (inputs(225)));
    layer0_outputs(3403) <= not((inputs(45)) or (inputs(46)));
    layer0_outputs(3404) <= not((inputs(128)) or (inputs(173)));
    layer0_outputs(3405) <= '1';
    layer0_outputs(3406) <= not(inputs(99)) or (inputs(127));
    layer0_outputs(3407) <= (inputs(59)) or (inputs(88));
    layer0_outputs(3408) <= '1';
    layer0_outputs(3409) <= not((inputs(12)) or (inputs(123)));
    layer0_outputs(3410) <= not((inputs(210)) xor (inputs(75)));
    layer0_outputs(3411) <= inputs(107);
    layer0_outputs(3412) <= not((inputs(186)) xor (inputs(46)));
    layer0_outputs(3413) <= (inputs(98)) or (inputs(184));
    layer0_outputs(3414) <= '0';
    layer0_outputs(3415) <= inputs(218);
    layer0_outputs(3416) <= not(inputs(172)) or (inputs(238));
    layer0_outputs(3417) <= '1';
    layer0_outputs(3418) <= '0';
    layer0_outputs(3419) <= (inputs(49)) or (inputs(192));
    layer0_outputs(3420) <= (inputs(68)) xor (inputs(123));
    layer0_outputs(3421) <= (inputs(97)) or (inputs(75));
    layer0_outputs(3422) <= (inputs(89)) and (inputs(139));
    layer0_outputs(3423) <= not((inputs(115)) or (inputs(83)));
    layer0_outputs(3424) <= inputs(38);
    layer0_outputs(3425) <= (inputs(185)) or (inputs(12));
    layer0_outputs(3426) <= inputs(95);
    layer0_outputs(3427) <= not((inputs(99)) xor (inputs(16)));
    layer0_outputs(3428) <= (inputs(177)) and (inputs(138));
    layer0_outputs(3429) <= not(inputs(185));
    layer0_outputs(3430) <= (inputs(50)) xor (inputs(230));
    layer0_outputs(3431) <= inputs(137);
    layer0_outputs(3432) <= (inputs(138)) xor (inputs(32));
    layer0_outputs(3433) <= inputs(85);
    layer0_outputs(3434) <= (inputs(165)) xor (inputs(85));
    layer0_outputs(3435) <= not(inputs(201));
    layer0_outputs(3436) <= (inputs(7)) and not (inputs(209));
    layer0_outputs(3437) <= not(inputs(213));
    layer0_outputs(3438) <= not(inputs(61)) or (inputs(82));
    layer0_outputs(3439) <= '0';
    layer0_outputs(3440) <= inputs(54);
    layer0_outputs(3441) <= not((inputs(168)) xor (inputs(206)));
    layer0_outputs(3442) <= not(inputs(105));
    layer0_outputs(3443) <= '1';
    layer0_outputs(3444) <= not(inputs(158));
    layer0_outputs(3445) <= '0';
    layer0_outputs(3446) <= not(inputs(81));
    layer0_outputs(3447) <= (inputs(97)) and not (inputs(7));
    layer0_outputs(3448) <= not((inputs(170)) xor (inputs(91)));
    layer0_outputs(3449) <= inputs(86);
    layer0_outputs(3450) <= (inputs(29)) and not (inputs(218));
    layer0_outputs(3451) <= (inputs(37)) or (inputs(23));
    layer0_outputs(3452) <= (inputs(84)) and not (inputs(174));
    layer0_outputs(3453) <= not(inputs(226));
    layer0_outputs(3454) <= not(inputs(94)) or (inputs(173));
    layer0_outputs(3455) <= not(inputs(132));
    layer0_outputs(3456) <= not(inputs(123));
    layer0_outputs(3457) <= inputs(106);
    layer0_outputs(3458) <= not((inputs(97)) and (inputs(11)));
    layer0_outputs(3459) <= (inputs(183)) and not (inputs(213));
    layer0_outputs(3460) <= (inputs(180)) and not (inputs(222));
    layer0_outputs(3461) <= not(inputs(162));
    layer0_outputs(3462) <= (inputs(140)) or (inputs(222));
    layer0_outputs(3463) <= not(inputs(106)) or (inputs(141));
    layer0_outputs(3464) <= (inputs(198)) or (inputs(172));
    layer0_outputs(3465) <= (inputs(27)) and not (inputs(240));
    layer0_outputs(3466) <= not(inputs(121));
    layer0_outputs(3467) <= not((inputs(2)) and (inputs(14)));
    layer0_outputs(3468) <= (inputs(29)) and not (inputs(111));
    layer0_outputs(3469) <= inputs(120);
    layer0_outputs(3470) <= not((inputs(82)) or (inputs(167)));
    layer0_outputs(3471) <= inputs(60);
    layer0_outputs(3472) <= not(inputs(213)) or (inputs(37));
    layer0_outputs(3473) <= not(inputs(172));
    layer0_outputs(3474) <= inputs(163);
    layer0_outputs(3475) <= (inputs(204)) xor (inputs(192));
    layer0_outputs(3476) <= not(inputs(27));
    layer0_outputs(3477) <= inputs(124);
    layer0_outputs(3478) <= not((inputs(98)) xor (inputs(26)));
    layer0_outputs(3479) <= not((inputs(227)) or (inputs(72)));
    layer0_outputs(3480) <= '0';
    layer0_outputs(3481) <= inputs(131);
    layer0_outputs(3482) <= (inputs(152)) or (inputs(135));
    layer0_outputs(3483) <= inputs(137);
    layer0_outputs(3484) <= '1';
    layer0_outputs(3485) <= (inputs(197)) and not (inputs(113));
    layer0_outputs(3486) <= inputs(110);
    layer0_outputs(3487) <= not(inputs(191));
    layer0_outputs(3488) <= (inputs(172)) or (inputs(109));
    layer0_outputs(3489) <= inputs(3);
    layer0_outputs(3490) <= not(inputs(63)) or (inputs(191));
    layer0_outputs(3491) <= '1';
    layer0_outputs(3492) <= not(inputs(218)) or (inputs(95));
    layer0_outputs(3493) <= (inputs(32)) and not (inputs(206));
    layer0_outputs(3494) <= (inputs(103)) and not (inputs(193));
    layer0_outputs(3495) <= (inputs(95)) and not (inputs(64));
    layer0_outputs(3496) <= '0';
    layer0_outputs(3497) <= not((inputs(233)) xor (inputs(177)));
    layer0_outputs(3498) <= not((inputs(203)) or (inputs(174)));
    layer0_outputs(3499) <= (inputs(22)) and not (inputs(2));
    layer0_outputs(3500) <= not(inputs(141)) or (inputs(94));
    layer0_outputs(3501) <= not(inputs(136));
    layer0_outputs(3502) <= not((inputs(114)) and (inputs(127)));
    layer0_outputs(3503) <= not((inputs(148)) or (inputs(51)));
    layer0_outputs(3504) <= not(inputs(38)) or (inputs(29));
    layer0_outputs(3505) <= (inputs(208)) and not (inputs(244));
    layer0_outputs(3506) <= not((inputs(212)) or (inputs(231)));
    layer0_outputs(3507) <= (inputs(74)) and not (inputs(96));
    layer0_outputs(3508) <= not(inputs(186));
    layer0_outputs(3509) <= (inputs(67)) and not (inputs(246));
    layer0_outputs(3510) <= not(inputs(152)) or (inputs(212));
    layer0_outputs(3511) <= not((inputs(27)) xor (inputs(178)));
    layer0_outputs(3512) <= (inputs(69)) and not (inputs(7));
    layer0_outputs(3513) <= (inputs(154)) xor (inputs(245));
    layer0_outputs(3514) <= not(inputs(225));
    layer0_outputs(3515) <= (inputs(152)) and not (inputs(162));
    layer0_outputs(3516) <= (inputs(180)) and not (inputs(98));
    layer0_outputs(3517) <= inputs(117);
    layer0_outputs(3518) <= inputs(253);
    layer0_outputs(3519) <= (inputs(6)) xor (inputs(201));
    layer0_outputs(3520) <= not((inputs(221)) xor (inputs(224)));
    layer0_outputs(3521) <= not((inputs(139)) or (inputs(124)));
    layer0_outputs(3522) <= (inputs(72)) or (inputs(48));
    layer0_outputs(3523) <= not(inputs(12)) or (inputs(168));
    layer0_outputs(3524) <= not(inputs(143)) or (inputs(2));
    layer0_outputs(3525) <= not(inputs(101));
    layer0_outputs(3526) <= not(inputs(200));
    layer0_outputs(3527) <= inputs(61);
    layer0_outputs(3528) <= (inputs(20)) and not (inputs(2));
    layer0_outputs(3529) <= inputs(200);
    layer0_outputs(3530) <= (inputs(30)) xor (inputs(23));
    layer0_outputs(3531) <= inputs(42);
    layer0_outputs(3532) <= (inputs(159)) and (inputs(255));
    layer0_outputs(3533) <= (inputs(62)) and not (inputs(6));
    layer0_outputs(3534) <= not(inputs(91));
    layer0_outputs(3535) <= (inputs(92)) or (inputs(74));
    layer0_outputs(3536) <= not((inputs(166)) xor (inputs(243)));
    layer0_outputs(3537) <= (inputs(26)) and not (inputs(159));
    layer0_outputs(3538) <= (inputs(193)) or (inputs(232));
    layer0_outputs(3539) <= (inputs(92)) and not (inputs(47));
    layer0_outputs(3540) <= (inputs(154)) or (inputs(202));
    layer0_outputs(3541) <= not((inputs(141)) xor (inputs(112)));
    layer0_outputs(3542) <= (inputs(97)) xor (inputs(147));
    layer0_outputs(3543) <= (inputs(125)) or (inputs(227));
    layer0_outputs(3544) <= (inputs(237)) xor (inputs(56));
    layer0_outputs(3545) <= not((inputs(227)) or (inputs(85)));
    layer0_outputs(3546) <= not((inputs(180)) and (inputs(42)));
    layer0_outputs(3547) <= (inputs(118)) or (inputs(157));
    layer0_outputs(3548) <= (inputs(182)) and not (inputs(30));
    layer0_outputs(3549) <= (inputs(228)) or (inputs(20));
    layer0_outputs(3550) <= (inputs(74)) or (inputs(219));
    layer0_outputs(3551) <= not(inputs(233)) or (inputs(1));
    layer0_outputs(3552) <= not((inputs(225)) xor (inputs(71)));
    layer0_outputs(3553) <= (inputs(152)) or (inputs(28));
    layer0_outputs(3554) <= not((inputs(130)) xor (inputs(249)));
    layer0_outputs(3555) <= not((inputs(117)) xor (inputs(130)));
    layer0_outputs(3556) <= (inputs(145)) or (inputs(38));
    layer0_outputs(3557) <= not(inputs(90)) or (inputs(195));
    layer0_outputs(3558) <= not(inputs(202)) or (inputs(115));
    layer0_outputs(3559) <= (inputs(188)) xor (inputs(238));
    layer0_outputs(3560) <= not(inputs(108));
    layer0_outputs(3561) <= not((inputs(50)) xor (inputs(48)));
    layer0_outputs(3562) <= not((inputs(95)) or (inputs(75)));
    layer0_outputs(3563) <= '1';
    layer0_outputs(3564) <= (inputs(114)) and (inputs(190));
    layer0_outputs(3565) <= inputs(66);
    layer0_outputs(3566) <= not(inputs(132)) or (inputs(24));
    layer0_outputs(3567) <= inputs(215);
    layer0_outputs(3568) <= (inputs(223)) and (inputs(43));
    layer0_outputs(3569) <= not((inputs(148)) or (inputs(83)));
    layer0_outputs(3570) <= not(inputs(53)) or (inputs(115));
    layer0_outputs(3571) <= '1';
    layer0_outputs(3572) <= (inputs(217)) xor (inputs(28));
    layer0_outputs(3573) <= (inputs(156)) or (inputs(102));
    layer0_outputs(3574) <= not(inputs(223));
    layer0_outputs(3575) <= not((inputs(82)) or (inputs(80)));
    layer0_outputs(3576) <= inputs(75);
    layer0_outputs(3577) <= not(inputs(239));
    layer0_outputs(3578) <= not((inputs(85)) or (inputs(212)));
    layer0_outputs(3579) <= not(inputs(138)) or (inputs(220));
    layer0_outputs(3580) <= not(inputs(119));
    layer0_outputs(3581) <= not(inputs(102)) or (inputs(248));
    layer0_outputs(3582) <= not((inputs(199)) and (inputs(185)));
    layer0_outputs(3583) <= inputs(82);
    layer0_outputs(3584) <= (inputs(138)) and not (inputs(175));
    layer0_outputs(3585) <= not(inputs(50)) or (inputs(19));
    layer0_outputs(3586) <= (inputs(27)) xor (inputs(175));
    layer0_outputs(3587) <= not((inputs(103)) or (inputs(222)));
    layer0_outputs(3588) <= inputs(111);
    layer0_outputs(3589) <= (inputs(52)) xor (inputs(140));
    layer0_outputs(3590) <= not(inputs(162)) or (inputs(64));
    layer0_outputs(3591) <= (inputs(20)) and not (inputs(128));
    layer0_outputs(3592) <= not(inputs(55)) or (inputs(132));
    layer0_outputs(3593) <= (inputs(153)) and not (inputs(6));
    layer0_outputs(3594) <= not((inputs(104)) or (inputs(130)));
    layer0_outputs(3595) <= (inputs(221)) or (inputs(249));
    layer0_outputs(3596) <= '0';
    layer0_outputs(3597) <= (inputs(58)) xor (inputs(238));
    layer0_outputs(3598) <= not(inputs(72)) or (inputs(183));
    layer0_outputs(3599) <= inputs(54);
    layer0_outputs(3600) <= not((inputs(98)) xor (inputs(35)));
    layer0_outputs(3601) <= (inputs(197)) and not (inputs(160));
    layer0_outputs(3602) <= not(inputs(170)) or (inputs(211));
    layer0_outputs(3603) <= (inputs(87)) or (inputs(7));
    layer0_outputs(3604) <= inputs(142);
    layer0_outputs(3605) <= (inputs(181)) or (inputs(83));
    layer0_outputs(3606) <= (inputs(65)) and (inputs(3));
    layer0_outputs(3607) <= (inputs(176)) and (inputs(21));
    layer0_outputs(3608) <= inputs(74);
    layer0_outputs(3609) <= not((inputs(14)) or (inputs(37)));
    layer0_outputs(3610) <= not(inputs(166));
    layer0_outputs(3611) <= inputs(88);
    layer0_outputs(3612) <= not((inputs(141)) or (inputs(77)));
    layer0_outputs(3613) <= inputs(120);
    layer0_outputs(3614) <= (inputs(177)) xor (inputs(171));
    layer0_outputs(3615) <= (inputs(43)) or (inputs(4));
    layer0_outputs(3616) <= (inputs(152)) or (inputs(23));
    layer0_outputs(3617) <= (inputs(206)) xor (inputs(176));
    layer0_outputs(3618) <= not((inputs(60)) or (inputs(188)));
    layer0_outputs(3619) <= (inputs(12)) xor (inputs(36));
    layer0_outputs(3620) <= not(inputs(203));
    layer0_outputs(3621) <= (inputs(107)) xor (inputs(49));
    layer0_outputs(3622) <= not(inputs(203)) or (inputs(161));
    layer0_outputs(3623) <= '0';
    layer0_outputs(3624) <= not(inputs(249)) or (inputs(20));
    layer0_outputs(3625) <= not((inputs(208)) xor (inputs(86)));
    layer0_outputs(3626) <= (inputs(62)) and not (inputs(33));
    layer0_outputs(3627) <= (inputs(175)) and not (inputs(12));
    layer0_outputs(3628) <= (inputs(241)) xor (inputs(60));
    layer0_outputs(3629) <= (inputs(160)) and not (inputs(22));
    layer0_outputs(3630) <= not(inputs(52));
    layer0_outputs(3631) <= not((inputs(169)) and (inputs(232)));
    layer0_outputs(3632) <= (inputs(122)) and not (inputs(49));
    layer0_outputs(3633) <= inputs(120);
    layer0_outputs(3634) <= not(inputs(205));
    layer0_outputs(3635) <= inputs(126);
    layer0_outputs(3636) <= inputs(241);
    layer0_outputs(3637) <= (inputs(50)) and not (inputs(219));
    layer0_outputs(3638) <= (inputs(228)) or (inputs(251));
    layer0_outputs(3639) <= not(inputs(136));
    layer0_outputs(3640) <= (inputs(20)) and (inputs(173));
    layer0_outputs(3641) <= not((inputs(74)) xor (inputs(114)));
    layer0_outputs(3642) <= not(inputs(233));
    layer0_outputs(3643) <= not((inputs(222)) xor (inputs(236)));
    layer0_outputs(3644) <= not(inputs(229));
    layer0_outputs(3645) <= inputs(214);
    layer0_outputs(3646) <= not((inputs(26)) or (inputs(185)));
    layer0_outputs(3647) <= (inputs(58)) or (inputs(33));
    layer0_outputs(3648) <= (inputs(58)) and not (inputs(154));
    layer0_outputs(3649) <= not((inputs(125)) xor (inputs(97)));
    layer0_outputs(3650) <= (inputs(175)) xor (inputs(175));
    layer0_outputs(3651) <= (inputs(226)) xor (inputs(31));
    layer0_outputs(3652) <= (inputs(209)) xor (inputs(107));
    layer0_outputs(3653) <= not((inputs(201)) or (inputs(253)));
    layer0_outputs(3654) <= (inputs(186)) or (inputs(91));
    layer0_outputs(3655) <= inputs(120);
    layer0_outputs(3656) <= (inputs(10)) or (inputs(84));
    layer0_outputs(3657) <= inputs(9);
    layer0_outputs(3658) <= inputs(139);
    layer0_outputs(3659) <= inputs(137);
    layer0_outputs(3660) <= (inputs(120)) and (inputs(105));
    layer0_outputs(3661) <= '1';
    layer0_outputs(3662) <= (inputs(106)) and not (inputs(73));
    layer0_outputs(3663) <= inputs(84);
    layer0_outputs(3664) <= (inputs(219)) and not (inputs(51));
    layer0_outputs(3665) <= not((inputs(149)) or (inputs(205)));
    layer0_outputs(3666) <= (inputs(255)) or (inputs(205));
    layer0_outputs(3667) <= (inputs(207)) or (inputs(198));
    layer0_outputs(3668) <= not((inputs(208)) or (inputs(73)));
    layer0_outputs(3669) <= (inputs(133)) and not (inputs(191));
    layer0_outputs(3670) <= (inputs(198)) and not (inputs(15));
    layer0_outputs(3671) <= inputs(237);
    layer0_outputs(3672) <= not((inputs(19)) xor (inputs(205)));
    layer0_outputs(3673) <= not((inputs(16)) or (inputs(235)));
    layer0_outputs(3674) <= (inputs(246)) or (inputs(233));
    layer0_outputs(3675) <= not((inputs(204)) or (inputs(181)));
    layer0_outputs(3676) <= not((inputs(223)) and (inputs(65)));
    layer0_outputs(3677) <= not(inputs(71)) or (inputs(68));
    layer0_outputs(3678) <= not((inputs(2)) or (inputs(83)));
    layer0_outputs(3679) <= (inputs(131)) and not (inputs(6));
    layer0_outputs(3680) <= not(inputs(102));
    layer0_outputs(3681) <= inputs(161);
    layer0_outputs(3682) <= (inputs(187)) and not (inputs(157));
    layer0_outputs(3683) <= (inputs(133)) and not (inputs(240));
    layer0_outputs(3684) <= (inputs(121)) and not (inputs(119));
    layer0_outputs(3685) <= (inputs(172)) or (inputs(22));
    layer0_outputs(3686) <= not(inputs(203));
    layer0_outputs(3687) <= '1';
    layer0_outputs(3688) <= not(inputs(100)) or (inputs(156));
    layer0_outputs(3689) <= not((inputs(211)) or (inputs(26)));
    layer0_outputs(3690) <= (inputs(51)) or (inputs(168));
    layer0_outputs(3691) <= (inputs(37)) or (inputs(70));
    layer0_outputs(3692) <= (inputs(11)) and (inputs(144));
    layer0_outputs(3693) <= not(inputs(116)) or (inputs(246));
    layer0_outputs(3694) <= not((inputs(161)) or (inputs(195)));
    layer0_outputs(3695) <= (inputs(45)) or (inputs(133));
    layer0_outputs(3696) <= not(inputs(204)) or (inputs(66));
    layer0_outputs(3697) <= not(inputs(254));
    layer0_outputs(3698) <= inputs(56);
    layer0_outputs(3699) <= (inputs(169)) or (inputs(205));
    layer0_outputs(3700) <= not(inputs(167)) or (inputs(81));
    layer0_outputs(3701) <= (inputs(151)) and not (inputs(173));
    layer0_outputs(3702) <= (inputs(82)) or (inputs(114));
    layer0_outputs(3703) <= inputs(183);
    layer0_outputs(3704) <= (inputs(242)) or (inputs(56));
    layer0_outputs(3705) <= inputs(187);
    layer0_outputs(3706) <= (inputs(137)) xor (inputs(33));
    layer0_outputs(3707) <= (inputs(59)) and not (inputs(2));
    layer0_outputs(3708) <= '1';
    layer0_outputs(3709) <= not((inputs(221)) or (inputs(133)));
    layer0_outputs(3710) <= not(inputs(134));
    layer0_outputs(3711) <= inputs(21);
    layer0_outputs(3712) <= (inputs(209)) xor (inputs(201));
    layer0_outputs(3713) <= not((inputs(15)) and (inputs(242)));
    layer0_outputs(3714) <= not(inputs(156)) or (inputs(13));
    layer0_outputs(3715) <= inputs(72);
    layer0_outputs(3716) <= not((inputs(4)) and (inputs(95)));
    layer0_outputs(3717) <= (inputs(55)) and (inputs(119));
    layer0_outputs(3718) <= '1';
    layer0_outputs(3719) <= not(inputs(68)) or (inputs(149));
    layer0_outputs(3720) <= (inputs(200)) and (inputs(76));
    layer0_outputs(3721) <= (inputs(79)) or (inputs(252));
    layer0_outputs(3722) <= not(inputs(32));
    layer0_outputs(3723) <= not((inputs(203)) or (inputs(36)));
    layer0_outputs(3724) <= not((inputs(80)) or (inputs(26)));
    layer0_outputs(3725) <= not((inputs(204)) and (inputs(11)));
    layer0_outputs(3726) <= not((inputs(28)) xor (inputs(82)));
    layer0_outputs(3727) <= (inputs(236)) xor (inputs(232));
    layer0_outputs(3728) <= (inputs(220)) or (inputs(175));
    layer0_outputs(3729) <= not((inputs(212)) or (inputs(196)));
    layer0_outputs(3730) <= inputs(150);
    layer0_outputs(3731) <= '0';
    layer0_outputs(3732) <= (inputs(77)) or (inputs(197));
    layer0_outputs(3733) <= (inputs(214)) xor (inputs(77));
    layer0_outputs(3734) <= (inputs(0)) and not (inputs(107));
    layer0_outputs(3735) <= (inputs(249)) and not (inputs(207));
    layer0_outputs(3736) <= inputs(104);
    layer0_outputs(3737) <= (inputs(219)) or (inputs(75));
    layer0_outputs(3738) <= (inputs(167)) and not (inputs(163));
    layer0_outputs(3739) <= (inputs(16)) xor (inputs(230));
    layer0_outputs(3740) <= not(inputs(164)) or (inputs(211));
    layer0_outputs(3741) <= not(inputs(125));
    layer0_outputs(3742) <= (inputs(217)) and not (inputs(113));
    layer0_outputs(3743) <= not(inputs(231));
    layer0_outputs(3744) <= (inputs(205)) and not (inputs(1));
    layer0_outputs(3745) <= (inputs(233)) xor (inputs(111));
    layer0_outputs(3746) <= (inputs(27)) xor (inputs(1));
    layer0_outputs(3747) <= (inputs(165)) xor (inputs(15));
    layer0_outputs(3748) <= (inputs(84)) xor (inputs(214));
    layer0_outputs(3749) <= inputs(28);
    layer0_outputs(3750) <= (inputs(62)) and not (inputs(64));
    layer0_outputs(3751) <= not(inputs(180));
    layer0_outputs(3752) <= not(inputs(99));
    layer0_outputs(3753) <= inputs(233);
    layer0_outputs(3754) <= (inputs(199)) and (inputs(196));
    layer0_outputs(3755) <= (inputs(159)) or (inputs(127));
    layer0_outputs(3756) <= (inputs(61)) and not (inputs(24));
    layer0_outputs(3757) <= (inputs(126)) and not (inputs(137));
    layer0_outputs(3758) <= not(inputs(57)) or (inputs(18));
    layer0_outputs(3759) <= not((inputs(92)) xor (inputs(14)));
    layer0_outputs(3760) <= not((inputs(0)) or (inputs(7)));
    layer0_outputs(3761) <= inputs(109);
    layer0_outputs(3762) <= (inputs(212)) or (inputs(79));
    layer0_outputs(3763) <= not((inputs(4)) xor (inputs(77)));
    layer0_outputs(3764) <= not((inputs(142)) xor (inputs(188)));
    layer0_outputs(3765) <= not((inputs(130)) and (inputs(49)));
    layer0_outputs(3766) <= not(inputs(172));
    layer0_outputs(3767) <= not((inputs(99)) and (inputs(95)));
    layer0_outputs(3768) <= inputs(248);
    layer0_outputs(3769) <= not((inputs(153)) or (inputs(154)));
    layer0_outputs(3770) <= not(inputs(116)) or (inputs(21));
    layer0_outputs(3771) <= not((inputs(25)) or (inputs(52)));
    layer0_outputs(3772) <= not((inputs(17)) or (inputs(238)));
    layer0_outputs(3773) <= (inputs(27)) or (inputs(87));
    layer0_outputs(3774) <= not(inputs(71)) or (inputs(223));
    layer0_outputs(3775) <= inputs(120);
    layer0_outputs(3776) <= (inputs(246)) and not (inputs(12));
    layer0_outputs(3777) <= (inputs(149)) or (inputs(123));
    layer0_outputs(3778) <= (inputs(97)) or (inputs(73));
    layer0_outputs(3779) <= (inputs(184)) and (inputs(154));
    layer0_outputs(3780) <= not(inputs(156));
    layer0_outputs(3781) <= (inputs(248)) xor (inputs(27));
    layer0_outputs(3782) <= inputs(81);
    layer0_outputs(3783) <= not((inputs(138)) or (inputs(66)));
    layer0_outputs(3784) <= inputs(168);
    layer0_outputs(3785) <= inputs(130);
    layer0_outputs(3786) <= not((inputs(189)) xor (inputs(149)));
    layer0_outputs(3787) <= not(inputs(79));
    layer0_outputs(3788) <= '1';
    layer0_outputs(3789) <= inputs(2);
    layer0_outputs(3790) <= not((inputs(84)) xor (inputs(43)));
    layer0_outputs(3791) <= (inputs(25)) or (inputs(114));
    layer0_outputs(3792) <= not((inputs(157)) or (inputs(166)));
    layer0_outputs(3793) <= not(inputs(60));
    layer0_outputs(3794) <= '0';
    layer0_outputs(3795) <= (inputs(166)) or (inputs(129));
    layer0_outputs(3796) <= (inputs(138)) and not (inputs(132));
    layer0_outputs(3797) <= not(inputs(124));
    layer0_outputs(3798) <= (inputs(73)) or (inputs(48));
    layer0_outputs(3799) <= (inputs(47)) xor (inputs(227));
    layer0_outputs(3800) <= (inputs(126)) or (inputs(156));
    layer0_outputs(3801) <= (inputs(26)) and not (inputs(145));
    layer0_outputs(3802) <= (inputs(202)) and not (inputs(46));
    layer0_outputs(3803) <= (inputs(91)) and not (inputs(156));
    layer0_outputs(3804) <= not(inputs(162)) or (inputs(184));
    layer0_outputs(3805) <= not((inputs(196)) xor (inputs(92)));
    layer0_outputs(3806) <= not(inputs(201)) or (inputs(68));
    layer0_outputs(3807) <= not(inputs(173)) or (inputs(250));
    layer0_outputs(3808) <= not((inputs(192)) xor (inputs(105)));
    layer0_outputs(3809) <= (inputs(12)) and not (inputs(79));
    layer0_outputs(3810) <= not((inputs(37)) xor (inputs(20)));
    layer0_outputs(3811) <= not((inputs(132)) or (inputs(205)));
    layer0_outputs(3812) <= not(inputs(88));
    layer0_outputs(3813) <= not(inputs(202)) or (inputs(24));
    layer0_outputs(3814) <= (inputs(240)) and (inputs(252));
    layer0_outputs(3815) <= not(inputs(202)) or (inputs(88));
    layer0_outputs(3816) <= (inputs(97)) xor (inputs(29));
    layer0_outputs(3817) <= inputs(186);
    layer0_outputs(3818) <= (inputs(157)) or (inputs(153));
    layer0_outputs(3819) <= '0';
    layer0_outputs(3820) <= not(inputs(39)) or (inputs(63));
    layer0_outputs(3821) <= inputs(45);
    layer0_outputs(3822) <= (inputs(218)) and (inputs(135));
    layer0_outputs(3823) <= not((inputs(95)) xor (inputs(166)));
    layer0_outputs(3824) <= (inputs(116)) and not (inputs(230));
    layer0_outputs(3825) <= inputs(195);
    layer0_outputs(3826) <= inputs(185);
    layer0_outputs(3827) <= not((inputs(241)) and (inputs(146)));
    layer0_outputs(3828) <= not(inputs(204));
    layer0_outputs(3829) <= '0';
    layer0_outputs(3830) <= inputs(56);
    layer0_outputs(3831) <= not((inputs(192)) or (inputs(147)));
    layer0_outputs(3832) <= inputs(119);
    layer0_outputs(3833) <= not((inputs(186)) or (inputs(35)));
    layer0_outputs(3834) <= not(inputs(213)) or (inputs(81));
    layer0_outputs(3835) <= (inputs(122)) and not (inputs(151));
    layer0_outputs(3836) <= not((inputs(92)) or (inputs(77)));
    layer0_outputs(3837) <= not(inputs(210)) or (inputs(208));
    layer0_outputs(3838) <= (inputs(66)) or (inputs(90));
    layer0_outputs(3839) <= inputs(133);
    layer0_outputs(3840) <= not((inputs(134)) or (inputs(202)));
    layer0_outputs(3841) <= (inputs(55)) xor (inputs(63));
    layer0_outputs(3842) <= not((inputs(176)) xor (inputs(167)));
    layer0_outputs(3843) <= (inputs(216)) or (inputs(28));
    layer0_outputs(3844) <= inputs(66);
    layer0_outputs(3845) <= not(inputs(100)) or (inputs(240));
    layer0_outputs(3846) <= not(inputs(109)) or (inputs(205));
    layer0_outputs(3847) <= inputs(94);
    layer0_outputs(3848) <= not(inputs(61)) or (inputs(113));
    layer0_outputs(3849) <= (inputs(157)) and not (inputs(46));
    layer0_outputs(3850) <= not((inputs(246)) xor (inputs(88)));
    layer0_outputs(3851) <= '1';
    layer0_outputs(3852) <= (inputs(186)) and not (inputs(99));
    layer0_outputs(3853) <= inputs(58);
    layer0_outputs(3854) <= (inputs(218)) and (inputs(206));
    layer0_outputs(3855) <= (inputs(93)) xor (inputs(192));
    layer0_outputs(3856) <= '1';
    layer0_outputs(3857) <= not((inputs(174)) or (inputs(152)));
    layer0_outputs(3858) <= not(inputs(55));
    layer0_outputs(3859) <= not((inputs(233)) or (inputs(178)));
    layer0_outputs(3860) <= not(inputs(83)) or (inputs(245));
    layer0_outputs(3861) <= not(inputs(155)) or (inputs(251));
    layer0_outputs(3862) <= (inputs(179)) or (inputs(254));
    layer0_outputs(3863) <= not(inputs(225));
    layer0_outputs(3864) <= (inputs(28)) xor (inputs(81));
    layer0_outputs(3865) <= not((inputs(6)) or (inputs(251)));
    layer0_outputs(3866) <= not((inputs(104)) or (inputs(235)));
    layer0_outputs(3867) <= (inputs(78)) or (inputs(77));
    layer0_outputs(3868) <= not(inputs(135));
    layer0_outputs(3869) <= not(inputs(133));
    layer0_outputs(3870) <= (inputs(49)) xor (inputs(105));
    layer0_outputs(3871) <= inputs(166);
    layer0_outputs(3872) <= (inputs(243)) and not (inputs(250));
    layer0_outputs(3873) <= not((inputs(147)) or (inputs(37)));
    layer0_outputs(3874) <= not((inputs(147)) xor (inputs(36)));
    layer0_outputs(3875) <= inputs(198);
    layer0_outputs(3876) <= (inputs(95)) and (inputs(210));
    layer0_outputs(3877) <= (inputs(130)) or (inputs(138));
    layer0_outputs(3878) <= not((inputs(81)) or (inputs(124)));
    layer0_outputs(3879) <= '1';
    layer0_outputs(3880) <= not((inputs(112)) or (inputs(184)));
    layer0_outputs(3881) <= (inputs(70)) and not (inputs(235));
    layer0_outputs(3882) <= not(inputs(197)) or (inputs(158));
    layer0_outputs(3883) <= not((inputs(197)) xor (inputs(228)));
    layer0_outputs(3884) <= not((inputs(22)) xor (inputs(108)));
    layer0_outputs(3885) <= inputs(78);
    layer0_outputs(3886) <= not((inputs(246)) and (inputs(20)));
    layer0_outputs(3887) <= not(inputs(47));
    layer0_outputs(3888) <= (inputs(126)) or (inputs(55));
    layer0_outputs(3889) <= not(inputs(104));
    layer0_outputs(3890) <= '0';
    layer0_outputs(3891) <= inputs(120);
    layer0_outputs(3892) <= not(inputs(125));
    layer0_outputs(3893) <= not(inputs(116));
    layer0_outputs(3894) <= not((inputs(21)) xor (inputs(64)));
    layer0_outputs(3895) <= inputs(85);
    layer0_outputs(3896) <= not(inputs(12)) or (inputs(176));
    layer0_outputs(3897) <= (inputs(87)) and not (inputs(82));
    layer0_outputs(3898) <= (inputs(109)) xor (inputs(215));
    layer0_outputs(3899) <= not((inputs(203)) xor (inputs(222)));
    layer0_outputs(3900) <= not((inputs(116)) or (inputs(236)));
    layer0_outputs(3901) <= (inputs(240)) or (inputs(184));
    layer0_outputs(3902) <= (inputs(80)) xor (inputs(172));
    layer0_outputs(3903) <= inputs(253);
    layer0_outputs(3904) <= (inputs(206)) or (inputs(194));
    layer0_outputs(3905) <= (inputs(250)) and not (inputs(243));
    layer0_outputs(3906) <= (inputs(83)) or (inputs(114));
    layer0_outputs(3907) <= (inputs(76)) or (inputs(180));
    layer0_outputs(3908) <= not(inputs(140));
    layer0_outputs(3909) <= not((inputs(233)) xor (inputs(232)));
    layer0_outputs(3910) <= inputs(5);
    layer0_outputs(3911) <= (inputs(67)) or (inputs(182));
    layer0_outputs(3912) <= not((inputs(129)) xor (inputs(145)));
    layer0_outputs(3913) <= (inputs(17)) xor (inputs(201));
    layer0_outputs(3914) <= not((inputs(37)) or (inputs(171)));
    layer0_outputs(3915) <= inputs(122);
    layer0_outputs(3916) <= (inputs(48)) or (inputs(188));
    layer0_outputs(3917) <= (inputs(183)) and not (inputs(211));
    layer0_outputs(3918) <= not((inputs(110)) or (inputs(255)));
    layer0_outputs(3919) <= not((inputs(15)) or (inputs(144)));
    layer0_outputs(3920) <= not((inputs(62)) xor (inputs(47)));
    layer0_outputs(3921) <= not(inputs(24)) or (inputs(128));
    layer0_outputs(3922) <= inputs(219);
    layer0_outputs(3923) <= not(inputs(138));
    layer0_outputs(3924) <= inputs(234);
    layer0_outputs(3925) <= not((inputs(125)) xor (inputs(235)));
    layer0_outputs(3926) <= (inputs(125)) and not (inputs(33));
    layer0_outputs(3927) <= (inputs(72)) or (inputs(38));
    layer0_outputs(3928) <= not(inputs(144)) or (inputs(19));
    layer0_outputs(3929) <= (inputs(94)) xor (inputs(59));
    layer0_outputs(3930) <= '0';
    layer0_outputs(3931) <= (inputs(190)) and not (inputs(2));
    layer0_outputs(3932) <= not(inputs(159));
    layer0_outputs(3933) <= not((inputs(129)) xor (inputs(2)));
    layer0_outputs(3934) <= not((inputs(143)) and (inputs(111)));
    layer0_outputs(3935) <= not(inputs(219));
    layer0_outputs(3936) <= (inputs(243)) and not (inputs(224));
    layer0_outputs(3937) <= not(inputs(17));
    layer0_outputs(3938) <= not((inputs(213)) and (inputs(249)));
    layer0_outputs(3939) <= (inputs(255)) xor (inputs(160));
    layer0_outputs(3940) <= not((inputs(41)) or (inputs(228)));
    layer0_outputs(3941) <= inputs(211);
    layer0_outputs(3942) <= (inputs(71)) xor (inputs(64));
    layer0_outputs(3943) <= not(inputs(93));
    layer0_outputs(3944) <= (inputs(179)) or (inputs(195));
    layer0_outputs(3945) <= inputs(133);
    layer0_outputs(3946) <= not(inputs(116)) or (inputs(33));
    layer0_outputs(3947) <= not(inputs(203));
    layer0_outputs(3948) <= (inputs(121)) and not (inputs(93));
    layer0_outputs(3949) <= (inputs(169)) and not (inputs(247));
    layer0_outputs(3950) <= inputs(132);
    layer0_outputs(3951) <= not((inputs(43)) or (inputs(61)));
    layer0_outputs(3952) <= not((inputs(131)) xor (inputs(8)));
    layer0_outputs(3953) <= not(inputs(165));
    layer0_outputs(3954) <= not(inputs(71)) or (inputs(246));
    layer0_outputs(3955) <= not((inputs(195)) and (inputs(114)));
    layer0_outputs(3956) <= not(inputs(116)) or (inputs(226));
    layer0_outputs(3957) <= not(inputs(135)) or (inputs(24));
    layer0_outputs(3958) <= not(inputs(149)) or (inputs(234));
    layer0_outputs(3959) <= (inputs(195)) or (inputs(44));
    layer0_outputs(3960) <= (inputs(6)) or (inputs(199));
    layer0_outputs(3961) <= not(inputs(5));
    layer0_outputs(3962) <= '0';
    layer0_outputs(3963) <= not(inputs(163));
    layer0_outputs(3964) <= not(inputs(167)) or (inputs(5));
    layer0_outputs(3965) <= not(inputs(71)) or (inputs(8));
    layer0_outputs(3966) <= inputs(165);
    layer0_outputs(3967) <= not(inputs(141)) or (inputs(14));
    layer0_outputs(3968) <= not((inputs(9)) and (inputs(242)));
    layer0_outputs(3969) <= not(inputs(73));
    layer0_outputs(3970) <= inputs(30);
    layer0_outputs(3971) <= (inputs(175)) xor (inputs(25));
    layer0_outputs(3972) <= (inputs(69)) or (inputs(85));
    layer0_outputs(3973) <= not(inputs(23));
    layer0_outputs(3974) <= not(inputs(66));
    layer0_outputs(3975) <= inputs(101);
    layer0_outputs(3976) <= not(inputs(58)) or (inputs(175));
    layer0_outputs(3977) <= not(inputs(90));
    layer0_outputs(3978) <= not(inputs(74));
    layer0_outputs(3979) <= (inputs(84)) and not (inputs(94));
    layer0_outputs(3980) <= (inputs(37)) or (inputs(51));
    layer0_outputs(3981) <= not(inputs(138));
    layer0_outputs(3982) <= not((inputs(111)) or (inputs(181)));
    layer0_outputs(3983) <= not(inputs(166));
    layer0_outputs(3984) <= not(inputs(144));
    layer0_outputs(3985) <= not(inputs(116)) or (inputs(96));
    layer0_outputs(3986) <= not((inputs(36)) and (inputs(145)));
    layer0_outputs(3987) <= (inputs(38)) or (inputs(19));
    layer0_outputs(3988) <= (inputs(179)) or (inputs(60));
    layer0_outputs(3989) <= not((inputs(76)) or (inputs(155)));
    layer0_outputs(3990) <= not(inputs(76)) or (inputs(224));
    layer0_outputs(3991) <= (inputs(212)) xor (inputs(19));
    layer0_outputs(3992) <= (inputs(176)) and (inputs(193));
    layer0_outputs(3993) <= '0';
    layer0_outputs(3994) <= not(inputs(81)) or (inputs(105));
    layer0_outputs(3995) <= not((inputs(249)) and (inputs(130)));
    layer0_outputs(3996) <= (inputs(229)) and not (inputs(223));
    layer0_outputs(3997) <= inputs(227);
    layer0_outputs(3998) <= not(inputs(21)) or (inputs(79));
    layer0_outputs(3999) <= not((inputs(126)) and (inputs(50)));
    layer0_outputs(4000) <= inputs(100);
    layer0_outputs(4001) <= (inputs(80)) and not (inputs(12));
    layer0_outputs(4002) <= not((inputs(43)) or (inputs(173)));
    layer0_outputs(4003) <= not((inputs(83)) or (inputs(248)));
    layer0_outputs(4004) <= not(inputs(106)) or (inputs(240));
    layer0_outputs(4005) <= (inputs(13)) and (inputs(113));
    layer0_outputs(4006) <= not(inputs(48));
    layer0_outputs(4007) <= not((inputs(233)) xor (inputs(61)));
    layer0_outputs(4008) <= (inputs(247)) or (inputs(183));
    layer0_outputs(4009) <= not((inputs(192)) or (inputs(33)));
    layer0_outputs(4010) <= (inputs(37)) or (inputs(63));
    layer0_outputs(4011) <= not(inputs(22));
    layer0_outputs(4012) <= not(inputs(80));
    layer0_outputs(4013) <= not(inputs(72));
    layer0_outputs(4014) <= (inputs(111)) xor (inputs(240));
    layer0_outputs(4015) <= inputs(195);
    layer0_outputs(4016) <= (inputs(55)) xor (inputs(230));
    layer0_outputs(4017) <= (inputs(36)) xor (inputs(89));
    layer0_outputs(4018) <= not((inputs(78)) or (inputs(106)));
    layer0_outputs(4019) <= '0';
    layer0_outputs(4020) <= not(inputs(65));
    layer0_outputs(4021) <= (inputs(155)) and not (inputs(36));
    layer0_outputs(4022) <= inputs(101);
    layer0_outputs(4023) <= (inputs(111)) and not (inputs(227));
    layer0_outputs(4024) <= not((inputs(101)) or (inputs(77)));
    layer0_outputs(4025) <= not((inputs(40)) or (inputs(26)));
    layer0_outputs(4026) <= inputs(86);
    layer0_outputs(4027) <= not(inputs(88));
    layer0_outputs(4028) <= (inputs(176)) and not (inputs(35));
    layer0_outputs(4029) <= (inputs(120)) and not (inputs(16));
    layer0_outputs(4030) <= (inputs(216)) and not (inputs(248));
    layer0_outputs(4031) <= inputs(3);
    layer0_outputs(4032) <= not(inputs(114));
    layer0_outputs(4033) <= (inputs(134)) and not (inputs(108));
    layer0_outputs(4034) <= not(inputs(213));
    layer0_outputs(4035) <= not(inputs(137));
    layer0_outputs(4036) <= (inputs(73)) or (inputs(97));
    layer0_outputs(4037) <= not(inputs(18)) or (inputs(161));
    layer0_outputs(4038) <= inputs(190);
    layer0_outputs(4039) <= (inputs(104)) and not (inputs(167));
    layer0_outputs(4040) <= (inputs(32)) and (inputs(60));
    layer0_outputs(4041) <= (inputs(58)) and not (inputs(38));
    layer0_outputs(4042) <= '0';
    layer0_outputs(4043) <= inputs(139);
    layer0_outputs(4044) <= (inputs(69)) or (inputs(196));
    layer0_outputs(4045) <= not((inputs(34)) or (inputs(164)));
    layer0_outputs(4046) <= (inputs(124)) or (inputs(87));
    layer0_outputs(4047) <= not(inputs(75)) or (inputs(162));
    layer0_outputs(4048) <= not(inputs(105));
    layer0_outputs(4049) <= inputs(140);
    layer0_outputs(4050) <= not(inputs(230));
    layer0_outputs(4051) <= not(inputs(196));
    layer0_outputs(4052) <= (inputs(199)) and not (inputs(249));
    layer0_outputs(4053) <= (inputs(252)) xor (inputs(148));
    layer0_outputs(4054) <= (inputs(172)) or (inputs(176));
    layer0_outputs(4055) <= not((inputs(8)) and (inputs(10)));
    layer0_outputs(4056) <= not(inputs(245)) or (inputs(191));
    layer0_outputs(4057) <= not(inputs(11)) or (inputs(18));
    layer0_outputs(4058) <= not(inputs(85)) or (inputs(163));
    layer0_outputs(4059) <= not(inputs(100)) or (inputs(5));
    layer0_outputs(4060) <= not(inputs(71)) or (inputs(111));
    layer0_outputs(4061) <= not((inputs(114)) and (inputs(228)));
    layer0_outputs(4062) <= (inputs(242)) and not (inputs(176));
    layer0_outputs(4063) <= not(inputs(75)) or (inputs(66));
    layer0_outputs(4064) <= (inputs(107)) or (inputs(176));
    layer0_outputs(4065) <= not((inputs(135)) or (inputs(120)));
    layer0_outputs(4066) <= not(inputs(221));
    layer0_outputs(4067) <= '1';
    layer0_outputs(4068) <= not(inputs(193));
    layer0_outputs(4069) <= inputs(170);
    layer0_outputs(4070) <= inputs(249);
    layer0_outputs(4071) <= (inputs(224)) and not (inputs(140));
    layer0_outputs(4072) <= not((inputs(95)) or (inputs(155)));
    layer0_outputs(4073) <= not(inputs(152));
    layer0_outputs(4074) <= not(inputs(196));
    layer0_outputs(4075) <= not((inputs(26)) xor (inputs(225)));
    layer0_outputs(4076) <= (inputs(204)) or (inputs(177));
    layer0_outputs(4077) <= not((inputs(230)) xor (inputs(67)));
    layer0_outputs(4078) <= not((inputs(48)) xor (inputs(153)));
    layer0_outputs(4079) <= not((inputs(199)) or (inputs(156)));
    layer0_outputs(4080) <= inputs(88);
    layer0_outputs(4081) <= '1';
    layer0_outputs(4082) <= not(inputs(46));
    layer0_outputs(4083) <= (inputs(1)) and not (inputs(250));
    layer0_outputs(4084) <= (inputs(193)) xor (inputs(57));
    layer0_outputs(4085) <= (inputs(79)) xor (inputs(135));
    layer0_outputs(4086) <= (inputs(84)) xor (inputs(133));
    layer0_outputs(4087) <= not(inputs(198)) or (inputs(35));
    layer0_outputs(4088) <= not(inputs(159)) or (inputs(33));
    layer0_outputs(4089) <= not(inputs(162));
    layer0_outputs(4090) <= not(inputs(221));
    layer0_outputs(4091) <= (inputs(13)) and (inputs(204));
    layer0_outputs(4092) <= not(inputs(198)) or (inputs(105));
    layer0_outputs(4093) <= not((inputs(68)) or (inputs(181)));
    layer0_outputs(4094) <= (inputs(137)) and not (inputs(204));
    layer0_outputs(4095) <= (inputs(209)) and not (inputs(63));
    layer0_outputs(4096) <= not((inputs(123)) or (inputs(109)));
    layer0_outputs(4097) <= not(inputs(43)) or (inputs(92));
    layer0_outputs(4098) <= not((inputs(35)) and (inputs(241)));
    layer0_outputs(4099) <= (inputs(231)) and not (inputs(155));
    layer0_outputs(4100) <= inputs(60);
    layer0_outputs(4101) <= (inputs(98)) or (inputs(253));
    layer0_outputs(4102) <= inputs(204);
    layer0_outputs(4103) <= not((inputs(134)) or (inputs(10)));
    layer0_outputs(4104) <= (inputs(36)) xor (inputs(36));
    layer0_outputs(4105) <= not(inputs(235));
    layer0_outputs(4106) <= not((inputs(134)) or (inputs(116)));
    layer0_outputs(4107) <= not(inputs(117)) or (inputs(109));
    layer0_outputs(4108) <= not(inputs(129)) or (inputs(99));
    layer0_outputs(4109) <= not((inputs(56)) or (inputs(114)));
    layer0_outputs(4110) <= '0';
    layer0_outputs(4111) <= not((inputs(180)) or (inputs(204)));
    layer0_outputs(4112) <= (inputs(81)) xor (inputs(240));
    layer0_outputs(4113) <= inputs(59);
    layer0_outputs(4114) <= (inputs(112)) xor (inputs(254));
    layer0_outputs(4115) <= not(inputs(119)) or (inputs(148));
    layer0_outputs(4116) <= not((inputs(149)) or (inputs(164)));
    layer0_outputs(4117) <= not((inputs(119)) or (inputs(63)));
    layer0_outputs(4118) <= not(inputs(84)) or (inputs(227));
    layer0_outputs(4119) <= not(inputs(5)) or (inputs(207));
    layer0_outputs(4120) <= not(inputs(163)) or (inputs(109));
    layer0_outputs(4121) <= not((inputs(43)) xor (inputs(218)));
    layer0_outputs(4122) <= not(inputs(106));
    layer0_outputs(4123) <= inputs(196);
    layer0_outputs(4124) <= inputs(187);
    layer0_outputs(4125) <= not((inputs(113)) xor (inputs(132)));
    layer0_outputs(4126) <= (inputs(192)) and (inputs(127));
    layer0_outputs(4127) <= not((inputs(217)) or (inputs(177)));
    layer0_outputs(4128) <= inputs(83);
    layer0_outputs(4129) <= not((inputs(226)) and (inputs(211)));
    layer0_outputs(4130) <= not(inputs(62));
    layer0_outputs(4131) <= not((inputs(173)) or (inputs(43)));
    layer0_outputs(4132) <= not(inputs(180));
    layer0_outputs(4133) <= not(inputs(81));
    layer0_outputs(4134) <= not(inputs(83));
    layer0_outputs(4135) <= (inputs(171)) and not (inputs(82));
    layer0_outputs(4136) <= inputs(183);
    layer0_outputs(4137) <= (inputs(174)) xor (inputs(14));
    layer0_outputs(4138) <= inputs(145);
    layer0_outputs(4139) <= (inputs(168)) and not (inputs(19));
    layer0_outputs(4140) <= not(inputs(187)) or (inputs(51));
    layer0_outputs(4141) <= not((inputs(200)) or (inputs(207)));
    layer0_outputs(4142) <= not(inputs(69)) or (inputs(122));
    layer0_outputs(4143) <= not(inputs(122)) or (inputs(57));
    layer0_outputs(4144) <= inputs(52);
    layer0_outputs(4145) <= not((inputs(87)) xor (inputs(125)));
    layer0_outputs(4146) <= not((inputs(2)) or (inputs(151)));
    layer0_outputs(4147) <= not((inputs(26)) and (inputs(130)));
    layer0_outputs(4148) <= not(inputs(141));
    layer0_outputs(4149) <= not((inputs(23)) or (inputs(75)));
    layer0_outputs(4150) <= not((inputs(170)) or (inputs(231)));
    layer0_outputs(4151) <= (inputs(161)) xor (inputs(81));
    layer0_outputs(4152) <= not(inputs(181));
    layer0_outputs(4153) <= not((inputs(87)) or (inputs(192)));
    layer0_outputs(4154) <= not((inputs(225)) and (inputs(81)));
    layer0_outputs(4155) <= not((inputs(242)) xor (inputs(246)));
    layer0_outputs(4156) <= not(inputs(133)) or (inputs(39));
    layer0_outputs(4157) <= inputs(209);
    layer0_outputs(4158) <= (inputs(172)) xor (inputs(6));
    layer0_outputs(4159) <= not(inputs(48));
    layer0_outputs(4160) <= not((inputs(174)) and (inputs(26)));
    layer0_outputs(4161) <= not((inputs(123)) xor (inputs(115)));
    layer0_outputs(4162) <= not(inputs(46)) or (inputs(66));
    layer0_outputs(4163) <= not((inputs(4)) or (inputs(107)));
    layer0_outputs(4164) <= not(inputs(136)) or (inputs(106));
    layer0_outputs(4165) <= not(inputs(40));
    layer0_outputs(4166) <= not((inputs(211)) or (inputs(15)));
    layer0_outputs(4167) <= not((inputs(47)) or (inputs(89)));
    layer0_outputs(4168) <= (inputs(117)) and not (inputs(129));
    layer0_outputs(4169) <= (inputs(1)) and not (inputs(27));
    layer0_outputs(4170) <= (inputs(89)) xor (inputs(33));
    layer0_outputs(4171) <= (inputs(48)) or (inputs(102));
    layer0_outputs(4172) <= not((inputs(177)) or (inputs(202)));
    layer0_outputs(4173) <= (inputs(56)) and not (inputs(202));
    layer0_outputs(4174) <= not(inputs(90)) or (inputs(7));
    layer0_outputs(4175) <= (inputs(196)) and not (inputs(115));
    layer0_outputs(4176) <= not((inputs(149)) or (inputs(92)));
    layer0_outputs(4177) <= not(inputs(116)) or (inputs(5));
    layer0_outputs(4178) <= (inputs(134)) xor (inputs(44));
    layer0_outputs(4179) <= not((inputs(90)) xor (inputs(145)));
    layer0_outputs(4180) <= not(inputs(88)) or (inputs(63));
    layer0_outputs(4181) <= not(inputs(121)) or (inputs(113));
    layer0_outputs(4182) <= (inputs(29)) and not (inputs(226));
    layer0_outputs(4183) <= not((inputs(58)) xor (inputs(243)));
    layer0_outputs(4184) <= not(inputs(133));
    layer0_outputs(4185) <= (inputs(21)) or (inputs(223));
    layer0_outputs(4186) <= not(inputs(135));
    layer0_outputs(4187) <= not(inputs(168)) or (inputs(108));
    layer0_outputs(4188) <= (inputs(75)) or (inputs(190));
    layer0_outputs(4189) <= (inputs(121)) and not (inputs(53));
    layer0_outputs(4190) <= not(inputs(137)) or (inputs(109));
    layer0_outputs(4191) <= (inputs(21)) and (inputs(248));
    layer0_outputs(4192) <= (inputs(234)) xor (inputs(146));
    layer0_outputs(4193) <= (inputs(206)) or (inputs(196));
    layer0_outputs(4194) <= '0';
    layer0_outputs(4195) <= not(inputs(198));
    layer0_outputs(4196) <= (inputs(133)) or (inputs(101));
    layer0_outputs(4197) <= (inputs(162)) and not (inputs(65));
    layer0_outputs(4198) <= inputs(198);
    layer0_outputs(4199) <= (inputs(34)) and (inputs(47));
    layer0_outputs(4200) <= not((inputs(232)) xor (inputs(40)));
    layer0_outputs(4201) <= (inputs(244)) and not (inputs(26));
    layer0_outputs(4202) <= (inputs(188)) and not (inputs(48));
    layer0_outputs(4203) <= not(inputs(201));
    layer0_outputs(4204) <= not(inputs(123)) or (inputs(94));
    layer0_outputs(4205) <= '0';
    layer0_outputs(4206) <= not((inputs(108)) xor (inputs(106)));
    layer0_outputs(4207) <= (inputs(32)) and (inputs(226));
    layer0_outputs(4208) <= not(inputs(93));
    layer0_outputs(4209) <= (inputs(117)) xor (inputs(65));
    layer0_outputs(4210) <= (inputs(209)) xor (inputs(40));
    layer0_outputs(4211) <= not((inputs(213)) or (inputs(70)));
    layer0_outputs(4212) <= not(inputs(49));
    layer0_outputs(4213) <= (inputs(141)) or (inputs(41));
    layer0_outputs(4214) <= not(inputs(72));
    layer0_outputs(4215) <= not(inputs(88)) or (inputs(10));
    layer0_outputs(4216) <= not((inputs(135)) xor (inputs(141)));
    layer0_outputs(4217) <= not((inputs(243)) or (inputs(126)));
    layer0_outputs(4218) <= not(inputs(56)) or (inputs(255));
    layer0_outputs(4219) <= inputs(232);
    layer0_outputs(4220) <= not(inputs(92));
    layer0_outputs(4221) <= (inputs(67)) and not (inputs(126));
    layer0_outputs(4222) <= not(inputs(117));
    layer0_outputs(4223) <= (inputs(183)) or (inputs(205));
    layer0_outputs(4224) <= (inputs(199)) or (inputs(111));
    layer0_outputs(4225) <= inputs(120);
    layer0_outputs(4226) <= not(inputs(220)) or (inputs(97));
    layer0_outputs(4227) <= inputs(164);
    layer0_outputs(4228) <= (inputs(116)) and not (inputs(231));
    layer0_outputs(4229) <= not((inputs(149)) or (inputs(117)));
    layer0_outputs(4230) <= (inputs(19)) or (inputs(142));
    layer0_outputs(4231) <= (inputs(71)) or (inputs(204));
    layer0_outputs(4232) <= not(inputs(39)) or (inputs(113));
    layer0_outputs(4233) <= '0';
    layer0_outputs(4234) <= not(inputs(86));
    layer0_outputs(4235) <= not(inputs(133));
    layer0_outputs(4236) <= inputs(182);
    layer0_outputs(4237) <= not(inputs(89));
    layer0_outputs(4238) <= (inputs(89)) or (inputs(253));
    layer0_outputs(4239) <= not((inputs(12)) and (inputs(180)));
    layer0_outputs(4240) <= (inputs(231)) xor (inputs(46));
    layer0_outputs(4241) <= (inputs(176)) xor (inputs(131));
    layer0_outputs(4242) <= not((inputs(52)) or (inputs(134)));
    layer0_outputs(4243) <= inputs(25);
    layer0_outputs(4244) <= (inputs(185)) and not (inputs(94));
    layer0_outputs(4245) <= (inputs(99)) and not (inputs(60));
    layer0_outputs(4246) <= (inputs(37)) or (inputs(242));
    layer0_outputs(4247) <= not((inputs(76)) or (inputs(216)));
    layer0_outputs(4248) <= (inputs(253)) and not (inputs(34));
    layer0_outputs(4249) <= (inputs(48)) xor (inputs(151));
    layer0_outputs(4250) <= (inputs(213)) and not (inputs(52));
    layer0_outputs(4251) <= not((inputs(77)) or (inputs(1)));
    layer0_outputs(4252) <= not((inputs(73)) xor (inputs(121)));
    layer0_outputs(4253) <= inputs(135);
    layer0_outputs(4254) <= (inputs(25)) or (inputs(186));
    layer0_outputs(4255) <= (inputs(150)) and not (inputs(31));
    layer0_outputs(4256) <= not(inputs(214)) or (inputs(249));
    layer0_outputs(4257) <= (inputs(1)) and not (inputs(35));
    layer0_outputs(4258) <= not((inputs(162)) or (inputs(215)));
    layer0_outputs(4259) <= inputs(239);
    layer0_outputs(4260) <= inputs(91);
    layer0_outputs(4261) <= '1';
    layer0_outputs(4262) <= (inputs(225)) xor (inputs(157));
    layer0_outputs(4263) <= inputs(200);
    layer0_outputs(4264) <= (inputs(250)) or (inputs(189));
    layer0_outputs(4265) <= not(inputs(24));
    layer0_outputs(4266) <= (inputs(150)) and not (inputs(213));
    layer0_outputs(4267) <= (inputs(157)) or (inputs(47));
    layer0_outputs(4268) <= not(inputs(69)) or (inputs(209));
    layer0_outputs(4269) <= (inputs(0)) or (inputs(150));
    layer0_outputs(4270) <= (inputs(58)) xor (inputs(179));
    layer0_outputs(4271) <= not(inputs(135)) or (inputs(27));
    layer0_outputs(4272) <= not((inputs(232)) xor (inputs(45)));
    layer0_outputs(4273) <= not(inputs(61)) or (inputs(175));
    layer0_outputs(4274) <= not((inputs(215)) xor (inputs(80)));
    layer0_outputs(4275) <= not(inputs(58)) or (inputs(39));
    layer0_outputs(4276) <= not(inputs(39));
    layer0_outputs(4277) <= (inputs(157)) xor (inputs(184));
    layer0_outputs(4278) <= (inputs(171)) or (inputs(154));
    layer0_outputs(4279) <= (inputs(122)) and not (inputs(45));
    layer0_outputs(4280) <= (inputs(19)) or (inputs(87));
    layer0_outputs(4281) <= not((inputs(104)) xor (inputs(20)));
    layer0_outputs(4282) <= not(inputs(219)) or (inputs(35));
    layer0_outputs(4283) <= not(inputs(213)) or (inputs(252));
    layer0_outputs(4284) <= not(inputs(38));
    layer0_outputs(4285) <= not((inputs(168)) xor (inputs(112)));
    layer0_outputs(4286) <= not(inputs(107));
    layer0_outputs(4287) <= not(inputs(4)) or (inputs(63));
    layer0_outputs(4288) <= (inputs(37)) or (inputs(193));
    layer0_outputs(4289) <= '1';
    layer0_outputs(4290) <= not(inputs(56)) or (inputs(235));
    layer0_outputs(4291) <= inputs(218);
    layer0_outputs(4292) <= (inputs(196)) and not (inputs(225));
    layer0_outputs(4293) <= not(inputs(153)) or (inputs(255));
    layer0_outputs(4294) <= not((inputs(51)) or (inputs(192)));
    layer0_outputs(4295) <= (inputs(51)) or (inputs(149));
    layer0_outputs(4296) <= (inputs(151)) or (inputs(230));
    layer0_outputs(4297) <= (inputs(243)) or (inputs(215));
    layer0_outputs(4298) <= (inputs(72)) and not (inputs(161));
    layer0_outputs(4299) <= '0';
    layer0_outputs(4300) <= (inputs(79)) or (inputs(230));
    layer0_outputs(4301) <= not(inputs(49));
    layer0_outputs(4302) <= '0';
    layer0_outputs(4303) <= not((inputs(14)) xor (inputs(169)));
    layer0_outputs(4304) <= (inputs(113)) xor (inputs(67));
    layer0_outputs(4305) <= not(inputs(12));
    layer0_outputs(4306) <= (inputs(121)) xor (inputs(254));
    layer0_outputs(4307) <= (inputs(71)) and not (inputs(187));
    layer0_outputs(4308) <= (inputs(78)) or (inputs(107));
    layer0_outputs(4309) <= not(inputs(10)) or (inputs(33));
    layer0_outputs(4310) <= (inputs(233)) or (inputs(10));
    layer0_outputs(4311) <= (inputs(187)) and not (inputs(160));
    layer0_outputs(4312) <= (inputs(117)) or (inputs(86));
    layer0_outputs(4313) <= inputs(92);
    layer0_outputs(4314) <= not((inputs(192)) or (inputs(182)));
    layer0_outputs(4315) <= not((inputs(104)) xor (inputs(201)));
    layer0_outputs(4316) <= inputs(160);
    layer0_outputs(4317) <= not(inputs(23));
    layer0_outputs(4318) <= not(inputs(50));
    layer0_outputs(4319) <= (inputs(173)) xor (inputs(152));
    layer0_outputs(4320) <= not((inputs(124)) xor (inputs(62)));
    layer0_outputs(4321) <= not((inputs(157)) or (inputs(212)));
    layer0_outputs(4322) <= (inputs(168)) and not (inputs(195));
    layer0_outputs(4323) <= inputs(229);
    layer0_outputs(4324) <= not(inputs(153));
    layer0_outputs(4325) <= not(inputs(160));
    layer0_outputs(4326) <= not((inputs(59)) or (inputs(205)));
    layer0_outputs(4327) <= (inputs(123)) and not (inputs(2));
    layer0_outputs(4328) <= not(inputs(229)) or (inputs(157));
    layer0_outputs(4329) <= not(inputs(187));
    layer0_outputs(4330) <= inputs(101);
    layer0_outputs(4331) <= (inputs(103)) and not (inputs(130));
    layer0_outputs(4332) <= inputs(222);
    layer0_outputs(4333) <= (inputs(99)) and not (inputs(69));
    layer0_outputs(4334) <= (inputs(109)) and not (inputs(51));
    layer0_outputs(4335) <= (inputs(53)) or (inputs(55));
    layer0_outputs(4336) <= inputs(102);
    layer0_outputs(4337) <= not((inputs(130)) or (inputs(18)));
    layer0_outputs(4338) <= not(inputs(8));
    layer0_outputs(4339) <= not((inputs(151)) xor (inputs(49)));
    layer0_outputs(4340) <= '1';
    layer0_outputs(4341) <= (inputs(31)) xor (inputs(112));
    layer0_outputs(4342) <= (inputs(74)) and (inputs(33));
    layer0_outputs(4343) <= not(inputs(179)) or (inputs(38));
    layer0_outputs(4344) <= (inputs(20)) and not (inputs(104));
    layer0_outputs(4345) <= not((inputs(172)) xor (inputs(255)));
    layer0_outputs(4346) <= not(inputs(122)) or (inputs(205));
    layer0_outputs(4347) <= (inputs(106)) and not (inputs(115));
    layer0_outputs(4348) <= (inputs(79)) and (inputs(174));
    layer0_outputs(4349) <= (inputs(15)) and not (inputs(17));
    layer0_outputs(4350) <= (inputs(254)) and not (inputs(176));
    layer0_outputs(4351) <= not(inputs(65));
    layer0_outputs(4352) <= inputs(67);
    layer0_outputs(4353) <= (inputs(151)) and not (inputs(45));
    layer0_outputs(4354) <= not((inputs(169)) xor (inputs(183)));
    layer0_outputs(4355) <= (inputs(244)) xor (inputs(122));
    layer0_outputs(4356) <= (inputs(90)) and not (inputs(68));
    layer0_outputs(4357) <= not((inputs(141)) or (inputs(200)));
    layer0_outputs(4358) <= not((inputs(142)) xor (inputs(0)));
    layer0_outputs(4359) <= (inputs(187)) or (inputs(80));
    layer0_outputs(4360) <= not((inputs(121)) xor (inputs(242)));
    layer0_outputs(4361) <= not(inputs(107)) or (inputs(149));
    layer0_outputs(4362) <= not(inputs(56)) or (inputs(100));
    layer0_outputs(4363) <= not(inputs(194)) or (inputs(25));
    layer0_outputs(4364) <= not((inputs(10)) or (inputs(90)));
    layer0_outputs(4365) <= not((inputs(234)) xor (inputs(252)));
    layer0_outputs(4366) <= not(inputs(42));
    layer0_outputs(4367) <= not((inputs(55)) xor (inputs(195)));
    layer0_outputs(4368) <= (inputs(246)) or (inputs(103));
    layer0_outputs(4369) <= not((inputs(153)) xor (inputs(13)));
    layer0_outputs(4370) <= not(inputs(92)) or (inputs(22));
    layer0_outputs(4371) <= (inputs(95)) or (inputs(182));
    layer0_outputs(4372) <= inputs(178);
    layer0_outputs(4373) <= not(inputs(36)) or (inputs(109));
    layer0_outputs(4374) <= not(inputs(57));
    layer0_outputs(4375) <= (inputs(145)) or (inputs(85));
    layer0_outputs(4376) <= (inputs(83)) or (inputs(91));
    layer0_outputs(4377) <= not((inputs(125)) or (inputs(180)));
    layer0_outputs(4378) <= (inputs(137)) and not (inputs(225));
    layer0_outputs(4379) <= not(inputs(120));
    layer0_outputs(4380) <= not((inputs(91)) or (inputs(98)));
    layer0_outputs(4381) <= not((inputs(186)) or (inputs(181)));
    layer0_outputs(4382) <= '0';
    layer0_outputs(4383) <= (inputs(117)) or (inputs(62));
    layer0_outputs(4384) <= not(inputs(146));
    layer0_outputs(4385) <= (inputs(200)) xor (inputs(169));
    layer0_outputs(4386) <= (inputs(17)) and not (inputs(228));
    layer0_outputs(4387) <= (inputs(117)) or (inputs(13));
    layer0_outputs(4388) <= (inputs(59)) and not (inputs(247));
    layer0_outputs(4389) <= not((inputs(180)) xor (inputs(34)));
    layer0_outputs(4390) <= (inputs(37)) or (inputs(25));
    layer0_outputs(4391) <= (inputs(32)) and (inputs(35));
    layer0_outputs(4392) <= (inputs(67)) and not (inputs(0));
    layer0_outputs(4393) <= (inputs(24)) and not (inputs(44));
    layer0_outputs(4394) <= (inputs(186)) xor (inputs(33));
    layer0_outputs(4395) <= not(inputs(54));
    layer0_outputs(4396) <= not(inputs(198));
    layer0_outputs(4397) <= not(inputs(106));
    layer0_outputs(4398) <= not(inputs(186)) or (inputs(183));
    layer0_outputs(4399) <= not((inputs(51)) or (inputs(217)));
    layer0_outputs(4400) <= not(inputs(80));
    layer0_outputs(4401) <= not(inputs(3));
    layer0_outputs(4402) <= not(inputs(67));
    layer0_outputs(4403) <= not((inputs(113)) and (inputs(224)));
    layer0_outputs(4404) <= not(inputs(163)) or (inputs(3));
    layer0_outputs(4405) <= inputs(45);
    layer0_outputs(4406) <= not((inputs(248)) and (inputs(57)));
    layer0_outputs(4407) <= inputs(189);
    layer0_outputs(4408) <= (inputs(118)) and not (inputs(17));
    layer0_outputs(4409) <= not(inputs(181));
    layer0_outputs(4410) <= not((inputs(131)) xor (inputs(244)));
    layer0_outputs(4411) <= not((inputs(167)) xor (inputs(147)));
    layer0_outputs(4412) <= not((inputs(29)) or (inputs(60)));
    layer0_outputs(4413) <= (inputs(121)) and not (inputs(62));
    layer0_outputs(4414) <= not(inputs(181)) or (inputs(103));
    layer0_outputs(4415) <= not((inputs(149)) or (inputs(247)));
    layer0_outputs(4416) <= not((inputs(90)) xor (inputs(213)));
    layer0_outputs(4417) <= not(inputs(84)) or (inputs(4));
    layer0_outputs(4418) <= (inputs(170)) and not (inputs(42));
    layer0_outputs(4419) <= inputs(245);
    layer0_outputs(4420) <= not(inputs(162)) or (inputs(125));
    layer0_outputs(4421) <= not((inputs(195)) or (inputs(158)));
    layer0_outputs(4422) <= not(inputs(113));
    layer0_outputs(4423) <= (inputs(239)) xor (inputs(101));
    layer0_outputs(4424) <= inputs(55);
    layer0_outputs(4425) <= inputs(35);
    layer0_outputs(4426) <= not((inputs(83)) or (inputs(36)));
    layer0_outputs(4427) <= not((inputs(106)) or (inputs(215)));
    layer0_outputs(4428) <= not(inputs(23)) or (inputs(222));
    layer0_outputs(4429) <= not((inputs(163)) or (inputs(189)));
    layer0_outputs(4430) <= inputs(56);
    layer0_outputs(4431) <= inputs(131);
    layer0_outputs(4432) <= not(inputs(112)) or (inputs(142));
    layer0_outputs(4433) <= not(inputs(90));
    layer0_outputs(4434) <= inputs(172);
    layer0_outputs(4435) <= not((inputs(102)) xor (inputs(209)));
    layer0_outputs(4436) <= not(inputs(135));
    layer0_outputs(4437) <= not(inputs(244));
    layer0_outputs(4438) <= inputs(73);
    layer0_outputs(4439) <= not((inputs(194)) xor (inputs(32)));
    layer0_outputs(4440) <= not((inputs(210)) or (inputs(205)));
    layer0_outputs(4441) <= not(inputs(225));
    layer0_outputs(4442) <= not(inputs(113));
    layer0_outputs(4443) <= inputs(165);
    layer0_outputs(4444) <= not(inputs(135)) or (inputs(52));
    layer0_outputs(4445) <= (inputs(32)) and (inputs(51));
    layer0_outputs(4446) <= inputs(245);
    layer0_outputs(4447) <= not(inputs(220)) or (inputs(21));
    layer0_outputs(4448) <= not((inputs(61)) or (inputs(32)));
    layer0_outputs(4449) <= not(inputs(181));
    layer0_outputs(4450) <= (inputs(238)) or (inputs(134));
    layer0_outputs(4451) <= not((inputs(94)) xor (inputs(233)));
    layer0_outputs(4452) <= not(inputs(216));
    layer0_outputs(4453) <= not((inputs(99)) xor (inputs(1)));
    layer0_outputs(4454) <= '0';
    layer0_outputs(4455) <= not((inputs(158)) or (inputs(22)));
    layer0_outputs(4456) <= inputs(166);
    layer0_outputs(4457) <= (inputs(127)) or (inputs(251));
    layer0_outputs(4458) <= (inputs(238)) and (inputs(89));
    layer0_outputs(4459) <= inputs(119);
    layer0_outputs(4460) <= (inputs(210)) xor (inputs(231));
    layer0_outputs(4461) <= (inputs(93)) or (inputs(198));
    layer0_outputs(4462) <= not(inputs(68)) or (inputs(235));
    layer0_outputs(4463) <= (inputs(21)) and (inputs(51));
    layer0_outputs(4464) <= inputs(105);
    layer0_outputs(4465) <= not(inputs(155)) or (inputs(109));
    layer0_outputs(4466) <= (inputs(15)) or (inputs(217));
    layer0_outputs(4467) <= (inputs(153)) and not (inputs(177));
    layer0_outputs(4468) <= not(inputs(160));
    layer0_outputs(4469) <= (inputs(94)) and not (inputs(10));
    layer0_outputs(4470) <= not((inputs(253)) xor (inputs(3)));
    layer0_outputs(4471) <= not((inputs(78)) and (inputs(254)));
    layer0_outputs(4472) <= inputs(190);
    layer0_outputs(4473) <= not((inputs(154)) and (inputs(27)));
    layer0_outputs(4474) <= not(inputs(81));
    layer0_outputs(4475) <= inputs(182);
    layer0_outputs(4476) <= (inputs(36)) or (inputs(122));
    layer0_outputs(4477) <= not((inputs(28)) or (inputs(170)));
    layer0_outputs(4478) <= (inputs(3)) or (inputs(134));
    layer0_outputs(4479) <= inputs(57);
    layer0_outputs(4480) <= not(inputs(111));
    layer0_outputs(4481) <= (inputs(78)) xor (inputs(195));
    layer0_outputs(4482) <= not(inputs(59));
    layer0_outputs(4483) <= inputs(95);
    layer0_outputs(4484) <= (inputs(58)) and not (inputs(231));
    layer0_outputs(4485) <= not(inputs(205));
    layer0_outputs(4486) <= (inputs(89)) xor (inputs(159));
    layer0_outputs(4487) <= not(inputs(19));
    layer0_outputs(4488) <= '1';
    layer0_outputs(4489) <= not(inputs(93)) or (inputs(46));
    layer0_outputs(4490) <= (inputs(122)) xor (inputs(49));
    layer0_outputs(4491) <= not(inputs(121));
    layer0_outputs(4492) <= not((inputs(102)) or (inputs(87)));
    layer0_outputs(4493) <= not(inputs(168)) or (inputs(220));
    layer0_outputs(4494) <= (inputs(166)) xor (inputs(103));
    layer0_outputs(4495) <= (inputs(34)) xor (inputs(217));
    layer0_outputs(4496) <= not(inputs(213)) or (inputs(189));
    layer0_outputs(4497) <= not(inputs(39));
    layer0_outputs(4498) <= (inputs(163)) or (inputs(52));
    layer0_outputs(4499) <= not(inputs(255)) or (inputs(29));
    layer0_outputs(4500) <= not(inputs(87)) or (inputs(147));
    layer0_outputs(4501) <= not((inputs(237)) xor (inputs(232)));
    layer0_outputs(4502) <= (inputs(154)) or (inputs(211));
    layer0_outputs(4503) <= (inputs(67)) and not (inputs(124));
    layer0_outputs(4504) <= not((inputs(203)) xor (inputs(34)));
    layer0_outputs(4505) <= not((inputs(41)) or (inputs(119)));
    layer0_outputs(4506) <= inputs(114);
    layer0_outputs(4507) <= inputs(198);
    layer0_outputs(4508) <= not(inputs(170));
    layer0_outputs(4509) <= not((inputs(118)) xor (inputs(222)));
    layer0_outputs(4510) <= (inputs(226)) xor (inputs(157));
    layer0_outputs(4511) <= not(inputs(57));
    layer0_outputs(4512) <= inputs(239);
    layer0_outputs(4513) <= not(inputs(102)) or (inputs(213));
    layer0_outputs(4514) <= not(inputs(133));
    layer0_outputs(4515) <= (inputs(214)) and not (inputs(25));
    layer0_outputs(4516) <= not((inputs(176)) xor (inputs(23)));
    layer0_outputs(4517) <= not(inputs(122)) or (inputs(61));
    layer0_outputs(4518) <= '1';
    layer0_outputs(4519) <= '0';
    layer0_outputs(4520) <= (inputs(167)) xor (inputs(0));
    layer0_outputs(4521) <= not(inputs(183)) or (inputs(227));
    layer0_outputs(4522) <= not((inputs(132)) and (inputs(73)));
    layer0_outputs(4523) <= not((inputs(39)) or (inputs(53)));
    layer0_outputs(4524) <= not((inputs(133)) and (inputs(139)));
    layer0_outputs(4525) <= (inputs(222)) and (inputs(4));
    layer0_outputs(4526) <= not((inputs(53)) or (inputs(39)));
    layer0_outputs(4527) <= not((inputs(193)) xor (inputs(75)));
    layer0_outputs(4528) <= (inputs(181)) and not (inputs(145));
    layer0_outputs(4529) <= (inputs(190)) or (inputs(186));
    layer0_outputs(4530) <= not(inputs(121));
    layer0_outputs(4531) <= not((inputs(41)) or (inputs(210)));
    layer0_outputs(4532) <= not(inputs(122));
    layer0_outputs(4533) <= inputs(197);
    layer0_outputs(4534) <= inputs(116);
    layer0_outputs(4535) <= not(inputs(207));
    layer0_outputs(4536) <= not((inputs(30)) xor (inputs(151)));
    layer0_outputs(4537) <= '0';
    layer0_outputs(4538) <= (inputs(210)) or (inputs(76));
    layer0_outputs(4539) <= not((inputs(64)) and (inputs(48)));
    layer0_outputs(4540) <= not(inputs(218)) or (inputs(238));
    layer0_outputs(4541) <= not((inputs(63)) xor (inputs(199)));
    layer0_outputs(4542) <= inputs(165);
    layer0_outputs(4543) <= not(inputs(57)) or (inputs(192));
    layer0_outputs(4544) <= (inputs(70)) or (inputs(66));
    layer0_outputs(4545) <= (inputs(150)) and not (inputs(50));
    layer0_outputs(4546) <= not(inputs(151)) or (inputs(231));
    layer0_outputs(4547) <= (inputs(146)) and not (inputs(61));
    layer0_outputs(4548) <= (inputs(216)) xor (inputs(140));
    layer0_outputs(4549) <= (inputs(184)) and not (inputs(133));
    layer0_outputs(4550) <= not(inputs(54));
    layer0_outputs(4551) <= (inputs(58)) and not (inputs(35));
    layer0_outputs(4552) <= inputs(207);
    layer0_outputs(4553) <= not((inputs(2)) or (inputs(206)));
    layer0_outputs(4554) <= inputs(120);
    layer0_outputs(4555) <= not((inputs(177)) xor (inputs(53)));
    layer0_outputs(4556) <= (inputs(201)) xor (inputs(237));
    layer0_outputs(4557) <= not((inputs(187)) xor (inputs(154)));
    layer0_outputs(4558) <= (inputs(255)) or (inputs(60));
    layer0_outputs(4559) <= not((inputs(20)) xor (inputs(179)));
    layer0_outputs(4560) <= not(inputs(119)) or (inputs(232));
    layer0_outputs(4561) <= (inputs(57)) xor (inputs(194));
    layer0_outputs(4562) <= '0';
    layer0_outputs(4563) <= inputs(148);
    layer0_outputs(4564) <= not((inputs(248)) xor (inputs(242)));
    layer0_outputs(4565) <= not(inputs(59));
    layer0_outputs(4566) <= (inputs(142)) xor (inputs(94));
    layer0_outputs(4567) <= not(inputs(249)) or (inputs(250));
    layer0_outputs(4568) <= '1';
    layer0_outputs(4569) <= not((inputs(84)) or (inputs(238)));
    layer0_outputs(4570) <= (inputs(90)) and not (inputs(178));
    layer0_outputs(4571) <= (inputs(108)) or (inputs(184));
    layer0_outputs(4572) <= not((inputs(230)) xor (inputs(206)));
    layer0_outputs(4573) <= not((inputs(60)) xor (inputs(69)));
    layer0_outputs(4574) <= not(inputs(148));
    layer0_outputs(4575) <= not((inputs(76)) xor (inputs(247)));
    layer0_outputs(4576) <= not(inputs(16)) or (inputs(80));
    layer0_outputs(4577) <= not(inputs(82));
    layer0_outputs(4578) <= (inputs(13)) and (inputs(251));
    layer0_outputs(4579) <= not(inputs(162)) or (inputs(233));
    layer0_outputs(4580) <= (inputs(116)) or (inputs(214));
    layer0_outputs(4581) <= not((inputs(47)) xor (inputs(100)));
    layer0_outputs(4582) <= (inputs(67)) or (inputs(237));
    layer0_outputs(4583) <= inputs(117);
    layer0_outputs(4584) <= '0';
    layer0_outputs(4585) <= inputs(233);
    layer0_outputs(4586) <= not((inputs(45)) xor (inputs(249)));
    layer0_outputs(4587) <= not((inputs(69)) and (inputs(136)));
    layer0_outputs(4588) <= inputs(48);
    layer0_outputs(4589) <= not(inputs(138));
    layer0_outputs(4590) <= not((inputs(146)) or (inputs(160)));
    layer0_outputs(4591) <= not(inputs(121));
    layer0_outputs(4592) <= inputs(197);
    layer0_outputs(4593) <= not((inputs(201)) and (inputs(215)));
    layer0_outputs(4594) <= (inputs(219)) or (inputs(59));
    layer0_outputs(4595) <= (inputs(134)) or (inputs(230));
    layer0_outputs(4596) <= (inputs(232)) or (inputs(52));
    layer0_outputs(4597) <= (inputs(138)) xor (inputs(145));
    layer0_outputs(4598) <= (inputs(89)) and not (inputs(8));
    layer0_outputs(4599) <= (inputs(134)) and not (inputs(3));
    layer0_outputs(4600) <= (inputs(77)) and not (inputs(22));
    layer0_outputs(4601) <= not((inputs(198)) xor (inputs(77)));
    layer0_outputs(4602) <= (inputs(112)) and not (inputs(158));
    layer0_outputs(4603) <= inputs(147);
    layer0_outputs(4604) <= not(inputs(222)) or (inputs(194));
    layer0_outputs(4605) <= (inputs(232)) and not (inputs(175));
    layer0_outputs(4606) <= inputs(216);
    layer0_outputs(4607) <= not((inputs(171)) xor (inputs(18)));
    layer0_outputs(4608) <= (inputs(219)) or (inputs(124));
    layer0_outputs(4609) <= (inputs(199)) and not (inputs(9));
    layer0_outputs(4610) <= not(inputs(54));
    layer0_outputs(4611) <= (inputs(241)) or (inputs(179));
    layer0_outputs(4612) <= not((inputs(187)) or (inputs(189)));
    layer0_outputs(4613) <= inputs(56);
    layer0_outputs(4614) <= inputs(170);
    layer0_outputs(4615) <= inputs(100);
    layer0_outputs(4616) <= inputs(18);
    layer0_outputs(4617) <= not(inputs(207)) or (inputs(248));
    layer0_outputs(4618) <= (inputs(11)) and not (inputs(2));
    layer0_outputs(4619) <= not(inputs(165));
    layer0_outputs(4620) <= not((inputs(69)) xor (inputs(141)));
    layer0_outputs(4621) <= (inputs(90)) and not (inputs(204));
    layer0_outputs(4622) <= inputs(92);
    layer0_outputs(4623) <= '0';
    layer0_outputs(4624) <= not((inputs(11)) or (inputs(67)));
    layer0_outputs(4625) <= not(inputs(78));
    layer0_outputs(4626) <= inputs(212);
    layer0_outputs(4627) <= not(inputs(107));
    layer0_outputs(4628) <= not((inputs(53)) or (inputs(67)));
    layer0_outputs(4629) <= (inputs(159)) or (inputs(127));
    layer0_outputs(4630) <= (inputs(12)) xor (inputs(15));
    layer0_outputs(4631) <= not((inputs(41)) or (inputs(157)));
    layer0_outputs(4632) <= (inputs(4)) and not (inputs(193));
    layer0_outputs(4633) <= not(inputs(213));
    layer0_outputs(4634) <= (inputs(132)) and not (inputs(55));
    layer0_outputs(4635) <= (inputs(185)) or (inputs(23));
    layer0_outputs(4636) <= (inputs(52)) and not (inputs(33));
    layer0_outputs(4637) <= inputs(133);
    layer0_outputs(4638) <= (inputs(136)) or (inputs(79));
    layer0_outputs(4639) <= not(inputs(80)) or (inputs(206));
    layer0_outputs(4640) <= not(inputs(216));
    layer0_outputs(4641) <= (inputs(54)) and not (inputs(254));
    layer0_outputs(4642) <= (inputs(49)) or (inputs(170));
    layer0_outputs(4643) <= not(inputs(238));
    layer0_outputs(4644) <= inputs(116);
    layer0_outputs(4645) <= inputs(116);
    layer0_outputs(4646) <= not(inputs(107)) or (inputs(175));
    layer0_outputs(4647) <= not(inputs(51));
    layer0_outputs(4648) <= (inputs(194)) or (inputs(177));
    layer0_outputs(4649) <= not(inputs(25));
    layer0_outputs(4650) <= (inputs(150)) and not (inputs(188));
    layer0_outputs(4651) <= (inputs(91)) and not (inputs(226));
    layer0_outputs(4652) <= not((inputs(88)) or (inputs(162)));
    layer0_outputs(4653) <= not(inputs(164)) or (inputs(18));
    layer0_outputs(4654) <= inputs(57);
    layer0_outputs(4655) <= inputs(4);
    layer0_outputs(4656) <= (inputs(179)) and not (inputs(93));
    layer0_outputs(4657) <= inputs(117);
    layer0_outputs(4658) <= not(inputs(125));
    layer0_outputs(4659) <= not(inputs(77)) or (inputs(253));
    layer0_outputs(4660) <= (inputs(225)) and (inputs(83));
    layer0_outputs(4661) <= not(inputs(245));
    layer0_outputs(4662) <= not(inputs(244)) or (inputs(224));
    layer0_outputs(4663) <= inputs(39);
    layer0_outputs(4664) <= (inputs(67)) xor (inputs(243));
    layer0_outputs(4665) <= inputs(117);
    layer0_outputs(4666) <= (inputs(107)) and not (inputs(136));
    layer0_outputs(4667) <= (inputs(246)) and not (inputs(246));
    layer0_outputs(4668) <= (inputs(109)) xor (inputs(172));
    layer0_outputs(4669) <= not(inputs(189));
    layer0_outputs(4670) <= not(inputs(165)) or (inputs(25));
    layer0_outputs(4671) <= not(inputs(162)) or (inputs(159));
    layer0_outputs(4672) <= not(inputs(169)) or (inputs(215));
    layer0_outputs(4673) <= (inputs(243)) and not (inputs(220));
    layer0_outputs(4674) <= inputs(207);
    layer0_outputs(4675) <= (inputs(244)) and not (inputs(176));
    layer0_outputs(4676) <= (inputs(31)) or (inputs(66));
    layer0_outputs(4677) <= not(inputs(57)) or (inputs(88));
    layer0_outputs(4678) <= '0';
    layer0_outputs(4679) <= (inputs(66)) or (inputs(37));
    layer0_outputs(4680) <= (inputs(105)) and not (inputs(162));
    layer0_outputs(4681) <= (inputs(187)) or (inputs(80));
    layer0_outputs(4682) <= not((inputs(1)) or (inputs(226)));
    layer0_outputs(4683) <= not(inputs(146));
    layer0_outputs(4684) <= '0';
    layer0_outputs(4685) <= not((inputs(225)) xor (inputs(68)));
    layer0_outputs(4686) <= (inputs(67)) and not (inputs(19));
    layer0_outputs(4687) <= not((inputs(203)) and (inputs(108)));
    layer0_outputs(4688) <= not((inputs(211)) or (inputs(228)));
    layer0_outputs(4689) <= '1';
    layer0_outputs(4690) <= inputs(219);
    layer0_outputs(4691) <= not((inputs(65)) and (inputs(78)));
    layer0_outputs(4692) <= not(inputs(186));
    layer0_outputs(4693) <= (inputs(72)) xor (inputs(40));
    layer0_outputs(4694) <= (inputs(118)) and not (inputs(236));
    layer0_outputs(4695) <= (inputs(105)) or (inputs(177));
    layer0_outputs(4696) <= inputs(55);
    layer0_outputs(4697) <= inputs(89);
    layer0_outputs(4698) <= not(inputs(121));
    layer0_outputs(4699) <= inputs(99);
    layer0_outputs(4700) <= not((inputs(136)) or (inputs(204)));
    layer0_outputs(4701) <= (inputs(251)) or (inputs(156));
    layer0_outputs(4702) <= (inputs(70)) xor (inputs(49));
    layer0_outputs(4703) <= not((inputs(162)) or (inputs(217)));
    layer0_outputs(4704) <= inputs(227);
    layer0_outputs(4705) <= not(inputs(36)) or (inputs(18));
    layer0_outputs(4706) <= inputs(211);
    layer0_outputs(4707) <= (inputs(236)) and not (inputs(107));
    layer0_outputs(4708) <= not(inputs(63)) or (inputs(161));
    layer0_outputs(4709) <= not(inputs(45)) or (inputs(225));
    layer0_outputs(4710) <= not((inputs(98)) xor (inputs(211)));
    layer0_outputs(4711) <= not(inputs(7)) or (inputs(17));
    layer0_outputs(4712) <= inputs(138);
    layer0_outputs(4713) <= not((inputs(54)) or (inputs(221)));
    layer0_outputs(4714) <= not((inputs(198)) or (inputs(206)));
    layer0_outputs(4715) <= (inputs(168)) and not (inputs(85));
    layer0_outputs(4716) <= inputs(231);
    layer0_outputs(4717) <= not(inputs(152)) or (inputs(156));
    layer0_outputs(4718) <= not((inputs(86)) and (inputs(83)));
    layer0_outputs(4719) <= (inputs(180)) or (inputs(11));
    layer0_outputs(4720) <= (inputs(213)) or (inputs(38));
    layer0_outputs(4721) <= (inputs(235)) and not (inputs(66));
    layer0_outputs(4722) <= (inputs(107)) or (inputs(236));
    layer0_outputs(4723) <= inputs(147);
    layer0_outputs(4724) <= inputs(220);
    layer0_outputs(4725) <= (inputs(63)) and (inputs(29));
    layer0_outputs(4726) <= (inputs(197)) xor (inputs(11));
    layer0_outputs(4727) <= inputs(102);
    layer0_outputs(4728) <= (inputs(234)) and not (inputs(30));
    layer0_outputs(4729) <= inputs(139);
    layer0_outputs(4730) <= inputs(225);
    layer0_outputs(4731) <= (inputs(48)) xor (inputs(60));
    layer0_outputs(4732) <= (inputs(117)) and not (inputs(40));
    layer0_outputs(4733) <= (inputs(89)) or (inputs(40));
    layer0_outputs(4734) <= not((inputs(101)) or (inputs(5)));
    layer0_outputs(4735) <= not((inputs(165)) xor (inputs(192)));
    layer0_outputs(4736) <= not(inputs(147));
    layer0_outputs(4737) <= not(inputs(228));
    layer0_outputs(4738) <= not(inputs(34));
    layer0_outputs(4739) <= (inputs(44)) or (inputs(41));
    layer0_outputs(4740) <= not((inputs(115)) or (inputs(42)));
    layer0_outputs(4741) <= (inputs(111)) and (inputs(51));
    layer0_outputs(4742) <= not(inputs(186)) or (inputs(204));
    layer0_outputs(4743) <= inputs(122);
    layer0_outputs(4744) <= not((inputs(139)) xor (inputs(140)));
    layer0_outputs(4745) <= not(inputs(134));
    layer0_outputs(4746) <= (inputs(215)) and not (inputs(127));
    layer0_outputs(4747) <= not(inputs(197));
    layer0_outputs(4748) <= not((inputs(93)) xor (inputs(90)));
    layer0_outputs(4749) <= inputs(25);
    layer0_outputs(4750) <= not(inputs(148)) or (inputs(193));
    layer0_outputs(4751) <= inputs(104);
    layer0_outputs(4752) <= not((inputs(179)) or (inputs(174)));
    layer0_outputs(4753) <= not(inputs(107)) or (inputs(227));
    layer0_outputs(4754) <= not((inputs(43)) or (inputs(228)));
    layer0_outputs(4755) <= inputs(199);
    layer0_outputs(4756) <= not(inputs(166)) or (inputs(11));
    layer0_outputs(4757) <= not((inputs(164)) xor (inputs(191)));
    layer0_outputs(4758) <= not((inputs(18)) xor (inputs(183)));
    layer0_outputs(4759) <= (inputs(46)) and not (inputs(209));
    layer0_outputs(4760) <= (inputs(173)) and not (inputs(29));
    layer0_outputs(4761) <= not(inputs(242));
    layer0_outputs(4762) <= not(inputs(29)) or (inputs(91));
    layer0_outputs(4763) <= (inputs(44)) xor (inputs(135));
    layer0_outputs(4764) <= (inputs(219)) and not (inputs(238));
    layer0_outputs(4765) <= (inputs(138)) or (inputs(179));
    layer0_outputs(4766) <= (inputs(121)) xor (inputs(24));
    layer0_outputs(4767) <= inputs(222);
    layer0_outputs(4768) <= not((inputs(68)) or (inputs(193)));
    layer0_outputs(4769) <= (inputs(105)) or (inputs(45));
    layer0_outputs(4770) <= (inputs(133)) or (inputs(204));
    layer0_outputs(4771) <= inputs(217);
    layer0_outputs(4772) <= inputs(242);
    layer0_outputs(4773) <= not(inputs(170));
    layer0_outputs(4774) <= not(inputs(86)) or (inputs(50));
    layer0_outputs(4775) <= not(inputs(217)) or (inputs(222));
    layer0_outputs(4776) <= not(inputs(208));
    layer0_outputs(4777) <= not((inputs(61)) or (inputs(160)));
    layer0_outputs(4778) <= inputs(147);
    layer0_outputs(4779) <= not(inputs(185)) or (inputs(145));
    layer0_outputs(4780) <= '1';
    layer0_outputs(4781) <= (inputs(144)) xor (inputs(211));
    layer0_outputs(4782) <= not((inputs(21)) and (inputs(236)));
    layer0_outputs(4783) <= not((inputs(185)) and (inputs(252)));
    layer0_outputs(4784) <= '0';
    layer0_outputs(4785) <= not(inputs(40));
    layer0_outputs(4786) <= inputs(198);
    layer0_outputs(4787) <= not(inputs(226)) or (inputs(178));
    layer0_outputs(4788) <= not((inputs(235)) or (inputs(36)));
    layer0_outputs(4789) <= inputs(73);
    layer0_outputs(4790) <= '1';
    layer0_outputs(4791) <= (inputs(225)) or (inputs(91));
    layer0_outputs(4792) <= inputs(213);
    layer0_outputs(4793) <= not(inputs(49)) or (inputs(254));
    layer0_outputs(4794) <= (inputs(27)) and not (inputs(189));
    layer0_outputs(4795) <= inputs(37);
    layer0_outputs(4796) <= not(inputs(214)) or (inputs(174));
    layer0_outputs(4797) <= (inputs(41)) or (inputs(165));
    layer0_outputs(4798) <= inputs(69);
    layer0_outputs(4799) <= (inputs(68)) and not (inputs(12));
    layer0_outputs(4800) <= inputs(22);
    layer0_outputs(4801) <= not((inputs(137)) xor (inputs(20)));
    layer0_outputs(4802) <= not((inputs(42)) or (inputs(62)));
    layer0_outputs(4803) <= not((inputs(183)) or (inputs(171)));
    layer0_outputs(4804) <= inputs(196);
    layer0_outputs(4805) <= (inputs(85)) and not (inputs(12));
    layer0_outputs(4806) <= inputs(155);
    layer0_outputs(4807) <= (inputs(5)) xor (inputs(15));
    layer0_outputs(4808) <= (inputs(120)) and not (inputs(97));
    layer0_outputs(4809) <= inputs(164);
    layer0_outputs(4810) <= inputs(89);
    layer0_outputs(4811) <= not((inputs(30)) or (inputs(86)));
    layer0_outputs(4812) <= not(inputs(84));
    layer0_outputs(4813) <= not(inputs(252));
    layer0_outputs(4814) <= inputs(41);
    layer0_outputs(4815) <= not(inputs(85)) or (inputs(223));
    layer0_outputs(4816) <= (inputs(176)) xor (inputs(151));
    layer0_outputs(4817) <= inputs(200);
    layer0_outputs(4818) <= (inputs(68)) xor (inputs(140));
    layer0_outputs(4819) <= (inputs(108)) and not (inputs(61));
    layer0_outputs(4820) <= (inputs(187)) xor (inputs(91));
    layer0_outputs(4821) <= not(inputs(16)) or (inputs(241));
    layer0_outputs(4822) <= (inputs(168)) and not (inputs(81));
    layer0_outputs(4823) <= not((inputs(31)) or (inputs(146)));
    layer0_outputs(4824) <= (inputs(213)) or (inputs(215));
    layer0_outputs(4825) <= not(inputs(119));
    layer0_outputs(4826) <= (inputs(224)) xor (inputs(186));
    layer0_outputs(4827) <= (inputs(164)) xor (inputs(71));
    layer0_outputs(4828) <= (inputs(167)) and not (inputs(192));
    layer0_outputs(4829) <= (inputs(199)) and not (inputs(250));
    layer0_outputs(4830) <= (inputs(96)) or (inputs(200));
    layer0_outputs(4831) <= (inputs(121)) and not (inputs(220));
    layer0_outputs(4832) <= not(inputs(109)) or (inputs(62));
    layer0_outputs(4833) <= (inputs(3)) or (inputs(103));
    layer0_outputs(4834) <= (inputs(64)) xor (inputs(233));
    layer0_outputs(4835) <= (inputs(39)) or (inputs(95));
    layer0_outputs(4836) <= not((inputs(46)) xor (inputs(200)));
    layer0_outputs(4837) <= (inputs(111)) xor (inputs(86));
    layer0_outputs(4838) <= (inputs(254)) xor (inputs(75));
    layer0_outputs(4839) <= not((inputs(104)) or (inputs(246)));
    layer0_outputs(4840) <= (inputs(155)) or (inputs(252));
    layer0_outputs(4841) <= not((inputs(182)) or (inputs(188)));
    layer0_outputs(4842) <= not(inputs(55)) or (inputs(102));
    layer0_outputs(4843) <= not((inputs(147)) xor (inputs(249)));
    layer0_outputs(4844) <= not((inputs(6)) xor (inputs(8)));
    layer0_outputs(4845) <= (inputs(203)) and not (inputs(234));
    layer0_outputs(4846) <= not((inputs(54)) or (inputs(31)));
    layer0_outputs(4847) <= not((inputs(61)) xor (inputs(28)));
    layer0_outputs(4848) <= not(inputs(255));
    layer0_outputs(4849) <= not(inputs(59)) or (inputs(96));
    layer0_outputs(4850) <= not((inputs(115)) or (inputs(221)));
    layer0_outputs(4851) <= '1';
    layer0_outputs(4852) <= not((inputs(65)) or (inputs(93)));
    layer0_outputs(4853) <= (inputs(17)) xor (inputs(18));
    layer0_outputs(4854) <= not(inputs(77)) or (inputs(15));
    layer0_outputs(4855) <= not((inputs(230)) xor (inputs(173)));
    layer0_outputs(4856) <= (inputs(185)) xor (inputs(18));
    layer0_outputs(4857) <= inputs(24);
    layer0_outputs(4858) <= (inputs(100)) or (inputs(4));
    layer0_outputs(4859) <= inputs(220);
    layer0_outputs(4860) <= not(inputs(237)) or (inputs(76));
    layer0_outputs(4861) <= (inputs(195)) and not (inputs(223));
    layer0_outputs(4862) <= inputs(226);
    layer0_outputs(4863) <= inputs(91);
    layer0_outputs(4864) <= (inputs(137)) or (inputs(113));
    layer0_outputs(4865) <= not((inputs(123)) xor (inputs(95)));
    layer0_outputs(4866) <= not(inputs(188));
    layer0_outputs(4867) <= not(inputs(166)) or (inputs(195));
    layer0_outputs(4868) <= '0';
    layer0_outputs(4869) <= not(inputs(151));
    layer0_outputs(4870) <= (inputs(16)) and not (inputs(18));
    layer0_outputs(4871) <= inputs(144);
    layer0_outputs(4872) <= (inputs(136)) and not (inputs(124));
    layer0_outputs(4873) <= (inputs(39)) and not (inputs(252));
    layer0_outputs(4874) <= not((inputs(2)) or (inputs(14)));
    layer0_outputs(4875) <= '1';
    layer0_outputs(4876) <= (inputs(71)) and not (inputs(235));
    layer0_outputs(4877) <= (inputs(108)) and not (inputs(146));
    layer0_outputs(4878) <= not((inputs(55)) or (inputs(172)));
    layer0_outputs(4879) <= (inputs(166)) and not (inputs(195));
    layer0_outputs(4880) <= (inputs(120)) and not (inputs(70));
    layer0_outputs(4881) <= (inputs(159)) and not (inputs(248));
    layer0_outputs(4882) <= (inputs(153)) or (inputs(207));
    layer0_outputs(4883) <= (inputs(138)) and not (inputs(171));
    layer0_outputs(4884) <= (inputs(169)) or (inputs(145));
    layer0_outputs(4885) <= not(inputs(174));
    layer0_outputs(4886) <= (inputs(252)) xor (inputs(214));
    layer0_outputs(4887) <= not(inputs(133));
    layer0_outputs(4888) <= (inputs(142)) and not (inputs(237));
    layer0_outputs(4889) <= (inputs(45)) and not (inputs(6));
    layer0_outputs(4890) <= (inputs(40)) or (inputs(150));
    layer0_outputs(4891) <= not(inputs(115));
    layer0_outputs(4892) <= inputs(140);
    layer0_outputs(4893) <= (inputs(1)) and (inputs(1));
    layer0_outputs(4894) <= (inputs(136)) or (inputs(145));
    layer0_outputs(4895) <= (inputs(93)) or (inputs(244));
    layer0_outputs(4896) <= not(inputs(179));
    layer0_outputs(4897) <= not((inputs(129)) and (inputs(210)));
    layer0_outputs(4898) <= (inputs(204)) xor (inputs(158));
    layer0_outputs(4899) <= (inputs(108)) or (inputs(83));
    layer0_outputs(4900) <= not((inputs(73)) xor (inputs(251)));
    layer0_outputs(4901) <= inputs(35);
    layer0_outputs(4902) <= not(inputs(108)) or (inputs(112));
    layer0_outputs(4903) <= not(inputs(88)) or (inputs(92));
    layer0_outputs(4904) <= not((inputs(61)) or (inputs(120)));
    layer0_outputs(4905) <= not(inputs(157));
    layer0_outputs(4906) <= inputs(211);
    layer0_outputs(4907) <= not((inputs(130)) xor (inputs(132)));
    layer0_outputs(4908) <= inputs(83);
    layer0_outputs(4909) <= (inputs(151)) and not (inputs(45));
    layer0_outputs(4910) <= inputs(196);
    layer0_outputs(4911) <= inputs(105);
    layer0_outputs(4912) <= not(inputs(239));
    layer0_outputs(4913) <= not((inputs(104)) or (inputs(177)));
    layer0_outputs(4914) <= '0';
    layer0_outputs(4915) <= not(inputs(215));
    layer0_outputs(4916) <= not((inputs(232)) or (inputs(131)));
    layer0_outputs(4917) <= not(inputs(134)) or (inputs(70));
    layer0_outputs(4918) <= not(inputs(198));
    layer0_outputs(4919) <= (inputs(101)) or (inputs(176));
    layer0_outputs(4920) <= (inputs(191)) and (inputs(236));
    layer0_outputs(4921) <= (inputs(186)) and not (inputs(46));
    layer0_outputs(4922) <= inputs(163);
    layer0_outputs(4923) <= not((inputs(201)) and (inputs(133)));
    layer0_outputs(4924) <= (inputs(18)) and (inputs(49));
    layer0_outputs(4925) <= not((inputs(204)) or (inputs(164)));
    layer0_outputs(4926) <= not(inputs(172)) or (inputs(189));
    layer0_outputs(4927) <= not(inputs(121)) or (inputs(157));
    layer0_outputs(4928) <= not((inputs(243)) and (inputs(37)));
    layer0_outputs(4929) <= not(inputs(219));
    layer0_outputs(4930) <= not(inputs(125)) or (inputs(63));
    layer0_outputs(4931) <= not((inputs(64)) or (inputs(240)));
    layer0_outputs(4932) <= (inputs(70)) and not (inputs(64));
    layer0_outputs(4933) <= not(inputs(165)) or (inputs(146));
    layer0_outputs(4934) <= not((inputs(237)) xor (inputs(229)));
    layer0_outputs(4935) <= inputs(185);
    layer0_outputs(4936) <= '0';
    layer0_outputs(4937) <= (inputs(16)) and not (inputs(241));
    layer0_outputs(4938) <= (inputs(210)) xor (inputs(217));
    layer0_outputs(4939) <= (inputs(79)) or (inputs(153));
    layer0_outputs(4940) <= not(inputs(216));
    layer0_outputs(4941) <= inputs(40);
    layer0_outputs(4942) <= not(inputs(98));
    layer0_outputs(4943) <= not((inputs(109)) xor (inputs(225)));
    layer0_outputs(4944) <= (inputs(51)) or (inputs(96));
    layer0_outputs(4945) <= not((inputs(143)) xor (inputs(191)));
    layer0_outputs(4946) <= not(inputs(16)) or (inputs(190));
    layer0_outputs(4947) <= not(inputs(53));
    layer0_outputs(4948) <= not(inputs(171)) or (inputs(30));
    layer0_outputs(4949) <= not(inputs(26));
    layer0_outputs(4950) <= not(inputs(0));
    layer0_outputs(4951) <= '0';
    layer0_outputs(4952) <= not(inputs(136)) or (inputs(230));
    layer0_outputs(4953) <= not(inputs(42));
    layer0_outputs(4954) <= inputs(49);
    layer0_outputs(4955) <= (inputs(158)) or (inputs(9));
    layer0_outputs(4956) <= not((inputs(129)) and (inputs(185)));
    layer0_outputs(4957) <= inputs(178);
    layer0_outputs(4958) <= not(inputs(40)) or (inputs(160));
    layer0_outputs(4959) <= not((inputs(167)) or (inputs(58)));
    layer0_outputs(4960) <= not(inputs(186));
    layer0_outputs(4961) <= not(inputs(118)) or (inputs(230));
    layer0_outputs(4962) <= (inputs(66)) and not (inputs(14));
    layer0_outputs(4963) <= not(inputs(41));
    layer0_outputs(4964) <= not((inputs(23)) or (inputs(103)));
    layer0_outputs(4965) <= inputs(164);
    layer0_outputs(4966) <= not(inputs(69)) or (inputs(24));
    layer0_outputs(4967) <= (inputs(69)) and not (inputs(116));
    layer0_outputs(4968) <= not((inputs(78)) xor (inputs(46)));
    layer0_outputs(4969) <= inputs(163);
    layer0_outputs(4970) <= inputs(138);
    layer0_outputs(4971) <= not(inputs(54));
    layer0_outputs(4972) <= not(inputs(242));
    layer0_outputs(4973) <= not(inputs(84)) or (inputs(205));
    layer0_outputs(4974) <= not((inputs(252)) or (inputs(8)));
    layer0_outputs(4975) <= not((inputs(112)) xor (inputs(145)));
    layer0_outputs(4976) <= (inputs(54)) and not (inputs(6));
    layer0_outputs(4977) <= not(inputs(133)) or (inputs(62));
    layer0_outputs(4978) <= not(inputs(156));
    layer0_outputs(4979) <= not(inputs(197));
    layer0_outputs(4980) <= not(inputs(10));
    layer0_outputs(4981) <= (inputs(93)) xor (inputs(221));
    layer0_outputs(4982) <= inputs(18);
    layer0_outputs(4983) <= inputs(166);
    layer0_outputs(4984) <= not(inputs(184));
    layer0_outputs(4985) <= not(inputs(141)) or (inputs(65));
    layer0_outputs(4986) <= (inputs(11)) or (inputs(231));
    layer0_outputs(4987) <= (inputs(35)) xor (inputs(169));
    layer0_outputs(4988) <= '0';
    layer0_outputs(4989) <= not((inputs(246)) xor (inputs(131)));
    layer0_outputs(4990) <= not((inputs(26)) or (inputs(191)));
    layer0_outputs(4991) <= not((inputs(109)) or (inputs(61)));
    layer0_outputs(4992) <= not(inputs(105));
    layer0_outputs(4993) <= (inputs(182)) and not (inputs(44));
    layer0_outputs(4994) <= (inputs(178)) xor (inputs(248));
    layer0_outputs(4995) <= not(inputs(207));
    layer0_outputs(4996) <= (inputs(140)) xor (inputs(20));
    layer0_outputs(4997) <= not((inputs(61)) xor (inputs(80)));
    layer0_outputs(4998) <= not(inputs(60)) or (inputs(28));
    layer0_outputs(4999) <= (inputs(70)) and not (inputs(22));
    layer0_outputs(5000) <= not(inputs(125));
    layer0_outputs(5001) <= (inputs(22)) and not (inputs(146));
    layer0_outputs(5002) <= inputs(202);
    layer0_outputs(5003) <= (inputs(27)) or (inputs(185));
    layer0_outputs(5004) <= (inputs(170)) and not (inputs(175));
    layer0_outputs(5005) <= not(inputs(209));
    layer0_outputs(5006) <= (inputs(191)) and not (inputs(144));
    layer0_outputs(5007) <= inputs(131);
    layer0_outputs(5008) <= not((inputs(135)) and (inputs(57)));
    layer0_outputs(5009) <= (inputs(84)) and not (inputs(54));
    layer0_outputs(5010) <= not((inputs(28)) xor (inputs(12)));
    layer0_outputs(5011) <= inputs(69);
    layer0_outputs(5012) <= (inputs(98)) or (inputs(183));
    layer0_outputs(5013) <= (inputs(220)) xor (inputs(251));
    layer0_outputs(5014) <= (inputs(157)) or (inputs(255));
    layer0_outputs(5015) <= not((inputs(78)) xor (inputs(49)));
    layer0_outputs(5016) <= (inputs(50)) and (inputs(241));
    layer0_outputs(5017) <= not(inputs(173)) or (inputs(21));
    layer0_outputs(5018) <= not((inputs(107)) xor (inputs(115)));
    layer0_outputs(5019) <= (inputs(225)) and not (inputs(148));
    layer0_outputs(5020) <= not(inputs(120)) or (inputs(17));
    layer0_outputs(5021) <= '0';
    layer0_outputs(5022) <= (inputs(127)) or (inputs(181));
    layer0_outputs(5023) <= not((inputs(174)) or (inputs(20)));
    layer0_outputs(5024) <= (inputs(77)) and not (inputs(69));
    layer0_outputs(5025) <= '1';
    layer0_outputs(5026) <= '0';
    layer0_outputs(5027) <= (inputs(83)) xor (inputs(179));
    layer0_outputs(5028) <= '0';
    layer0_outputs(5029) <= not(inputs(114)) or (inputs(70));
    layer0_outputs(5030) <= not(inputs(55));
    layer0_outputs(5031) <= not(inputs(164));
    layer0_outputs(5032) <= (inputs(44)) or (inputs(196));
    layer0_outputs(5033) <= inputs(197);
    layer0_outputs(5034) <= not((inputs(245)) xor (inputs(155)));
    layer0_outputs(5035) <= '0';
    layer0_outputs(5036) <= (inputs(154)) or (inputs(15));
    layer0_outputs(5037) <= inputs(167);
    layer0_outputs(5038) <= not((inputs(124)) or (inputs(89)));
    layer0_outputs(5039) <= (inputs(61)) xor (inputs(150));
    layer0_outputs(5040) <= not((inputs(169)) or (inputs(16)));
    layer0_outputs(5041) <= not(inputs(25));
    layer0_outputs(5042) <= not(inputs(90)) or (inputs(141));
    layer0_outputs(5043) <= not((inputs(0)) xor (inputs(111)));
    layer0_outputs(5044) <= not(inputs(244));
    layer0_outputs(5045) <= not(inputs(55)) or (inputs(64));
    layer0_outputs(5046) <= not(inputs(166));
    layer0_outputs(5047) <= inputs(117);
    layer0_outputs(5048) <= not(inputs(89));
    layer0_outputs(5049) <= (inputs(93)) xor (inputs(17));
    layer0_outputs(5050) <= (inputs(112)) or (inputs(60));
    layer0_outputs(5051) <= (inputs(56)) or (inputs(247));
    layer0_outputs(5052) <= '1';
    layer0_outputs(5053) <= not(inputs(134)) or (inputs(220));
    layer0_outputs(5054) <= inputs(39);
    layer0_outputs(5055) <= not(inputs(10)) or (inputs(60));
    layer0_outputs(5056) <= not(inputs(22)) or (inputs(80));
    layer0_outputs(5057) <= not((inputs(208)) or (inputs(97)));
    layer0_outputs(5058) <= (inputs(89)) and not (inputs(171));
    layer0_outputs(5059) <= not(inputs(227)) or (inputs(192));
    layer0_outputs(5060) <= inputs(156);
    layer0_outputs(5061) <= (inputs(161)) and not (inputs(223));
    layer0_outputs(5062) <= '1';
    layer0_outputs(5063) <= not((inputs(10)) xor (inputs(149)));
    layer0_outputs(5064) <= not(inputs(157)) or (inputs(2));
    layer0_outputs(5065) <= not(inputs(231)) or (inputs(190));
    layer0_outputs(5066) <= not((inputs(223)) xor (inputs(41)));
    layer0_outputs(5067) <= (inputs(97)) xor (inputs(188));
    layer0_outputs(5068) <= '0';
    layer0_outputs(5069) <= not(inputs(187)) or (inputs(82));
    layer0_outputs(5070) <= (inputs(136)) and (inputs(136));
    layer0_outputs(5071) <= inputs(43);
    layer0_outputs(5072) <= (inputs(110)) and not (inputs(243));
    layer0_outputs(5073) <= not(inputs(176));
    layer0_outputs(5074) <= '0';
    layer0_outputs(5075) <= not((inputs(172)) or (inputs(96)));
    layer0_outputs(5076) <= (inputs(215)) or (inputs(40));
    layer0_outputs(5077) <= inputs(54);
    layer0_outputs(5078) <= not(inputs(22));
    layer0_outputs(5079) <= (inputs(1)) and not (inputs(62));
    layer0_outputs(5080) <= not((inputs(97)) or (inputs(187)));
    layer0_outputs(5081) <= '0';
    layer0_outputs(5082) <= (inputs(137)) and not (inputs(68));
    layer0_outputs(5083) <= (inputs(167)) and not (inputs(224));
    layer0_outputs(5084) <= (inputs(224)) or (inputs(205));
    layer0_outputs(5085) <= not((inputs(138)) or (inputs(146)));
    layer0_outputs(5086) <= not(inputs(23));
    layer0_outputs(5087) <= (inputs(112)) xor (inputs(105));
    layer0_outputs(5088) <= (inputs(124)) and not (inputs(234));
    layer0_outputs(5089) <= not(inputs(170));
    layer0_outputs(5090) <= not((inputs(90)) xor (inputs(189)));
    layer0_outputs(5091) <= (inputs(177)) or (inputs(211));
    layer0_outputs(5092) <= inputs(22);
    layer0_outputs(5093) <= not((inputs(195)) xor (inputs(5)));
    layer0_outputs(5094) <= not(inputs(119));
    layer0_outputs(5095) <= (inputs(247)) xor (inputs(224));
    layer0_outputs(5096) <= (inputs(2)) or (inputs(76));
    layer0_outputs(5097) <= not((inputs(161)) xor (inputs(57)));
    layer0_outputs(5098) <= (inputs(40)) or (inputs(163));
    layer0_outputs(5099) <= inputs(165);
    layer0_outputs(5100) <= inputs(181);
    layer0_outputs(5101) <= not(inputs(5)) or (inputs(147));
    layer0_outputs(5102) <= not(inputs(193)) or (inputs(238));
    layer0_outputs(5103) <= (inputs(254)) or (inputs(90));
    layer0_outputs(5104) <= not(inputs(200)) or (inputs(11));
    layer0_outputs(5105) <= not((inputs(235)) or (inputs(237)));
    layer0_outputs(5106) <= not((inputs(156)) or (inputs(139)));
    layer0_outputs(5107) <= not(inputs(140));
    layer0_outputs(5108) <= inputs(55);
    layer0_outputs(5109) <= not((inputs(101)) xor (inputs(114)));
    layer0_outputs(5110) <= not(inputs(32));
    layer0_outputs(5111) <= inputs(164);
    layer0_outputs(5112) <= (inputs(122)) xor (inputs(142));
    layer0_outputs(5113) <= not(inputs(150));
    layer0_outputs(5114) <= (inputs(171)) and not (inputs(114));
    layer0_outputs(5115) <= (inputs(131)) and not (inputs(247));
    layer0_outputs(5116) <= (inputs(22)) xor (inputs(143));
    layer0_outputs(5117) <= not(inputs(174));
    layer0_outputs(5118) <= not(inputs(139)) or (inputs(32));
    layer0_outputs(5119) <= (inputs(3)) and not (inputs(144));
    outputs(0) <= (layer0_outputs(4090)) xor (layer0_outputs(4751));
    outputs(1) <= (layer0_outputs(2188)) xor (layer0_outputs(3085));
    outputs(2) <= not(layer0_outputs(1224));
    outputs(3) <= (layer0_outputs(3792)) xor (layer0_outputs(4442));
    outputs(4) <= (layer0_outputs(801)) xor (layer0_outputs(1110));
    outputs(5) <= (layer0_outputs(2215)) and (layer0_outputs(5059));
    outputs(6) <= layer0_outputs(2519);
    outputs(7) <= (layer0_outputs(2540)) xor (layer0_outputs(4021));
    outputs(8) <= not(layer0_outputs(4223));
    outputs(9) <= (layer0_outputs(1615)) xor (layer0_outputs(3363));
    outputs(10) <= not((layer0_outputs(3077)) or (layer0_outputs(1829)));
    outputs(11) <= not(layer0_outputs(2953));
    outputs(12) <= not((layer0_outputs(4386)) xor (layer0_outputs(2901)));
    outputs(13) <= layer0_outputs(3311);
    outputs(14) <= not((layer0_outputs(4459)) or (layer0_outputs(3662)));
    outputs(15) <= layer0_outputs(2241);
    outputs(16) <= layer0_outputs(4526);
    outputs(17) <= (layer0_outputs(4228)) and (layer0_outputs(3554));
    outputs(18) <= (layer0_outputs(3989)) xor (layer0_outputs(4590));
    outputs(19) <= layer0_outputs(2187);
    outputs(20) <= not((layer0_outputs(3928)) and (layer0_outputs(4995)));
    outputs(21) <= layer0_outputs(4146);
    outputs(22) <= not(layer0_outputs(4832));
    outputs(23) <= not((layer0_outputs(5079)) xor (layer0_outputs(5018)));
    outputs(24) <= not(layer0_outputs(206)) or (layer0_outputs(489));
    outputs(25) <= not(layer0_outputs(1980)) or (layer0_outputs(712));
    outputs(26) <= not(layer0_outputs(748)) or (layer0_outputs(526));
    outputs(27) <= (layer0_outputs(2853)) or (layer0_outputs(950));
    outputs(28) <= not(layer0_outputs(1329)) or (layer0_outputs(927));
    outputs(29) <= not((layer0_outputs(2739)) xor (layer0_outputs(999)));
    outputs(30) <= not((layer0_outputs(1720)) xor (layer0_outputs(2535)));
    outputs(31) <= not(layer0_outputs(3203)) or (layer0_outputs(886));
    outputs(32) <= not((layer0_outputs(4155)) and (layer0_outputs(2271)));
    outputs(33) <= (layer0_outputs(5019)) or (layer0_outputs(2744));
    outputs(34) <= (layer0_outputs(2404)) xor (layer0_outputs(3532));
    outputs(35) <= not(layer0_outputs(1162));
    outputs(36) <= not((layer0_outputs(4648)) xor (layer0_outputs(3109)));
    outputs(37) <= (layer0_outputs(2218)) xor (layer0_outputs(3727));
    outputs(38) <= not(layer0_outputs(4322));
    outputs(39) <= not(layer0_outputs(1197));
    outputs(40) <= (layer0_outputs(453)) xor (layer0_outputs(3061));
    outputs(41) <= (layer0_outputs(1917)) and (layer0_outputs(4025));
    outputs(42) <= (layer0_outputs(4868)) or (layer0_outputs(4755));
    outputs(43) <= not((layer0_outputs(1736)) or (layer0_outputs(3528)));
    outputs(44) <= (layer0_outputs(1469)) xor (layer0_outputs(3460));
    outputs(45) <= layer0_outputs(4997);
    outputs(46) <= not(layer0_outputs(1626)) or (layer0_outputs(364));
    outputs(47) <= layer0_outputs(67);
    outputs(48) <= not(layer0_outputs(3258));
    outputs(49) <= not(layer0_outputs(1206));
    outputs(50) <= not(layer0_outputs(4977));
    outputs(51) <= not(layer0_outputs(5087)) or (layer0_outputs(407));
    outputs(52) <= not((layer0_outputs(5093)) xor (layer0_outputs(2858)));
    outputs(53) <= not(layer0_outputs(256));
    outputs(54) <= (layer0_outputs(1067)) and (layer0_outputs(4455));
    outputs(55) <= not((layer0_outputs(3453)) and (layer0_outputs(4100)));
    outputs(56) <= not(layer0_outputs(1066));
    outputs(57) <= not((layer0_outputs(3437)) xor (layer0_outputs(103)));
    outputs(58) <= layer0_outputs(531);
    outputs(59) <= not(layer0_outputs(1258));
    outputs(60) <= not(layer0_outputs(3482));
    outputs(61) <= layer0_outputs(3610);
    outputs(62) <= layer0_outputs(624);
    outputs(63) <= not(layer0_outputs(4522));
    outputs(64) <= not((layer0_outputs(4670)) and (layer0_outputs(2348)));
    outputs(65) <= layer0_outputs(176);
    outputs(66) <= (layer0_outputs(3130)) xor (layer0_outputs(2773));
    outputs(67) <= not((layer0_outputs(2227)) xor (layer0_outputs(3699)));
    outputs(68) <= not((layer0_outputs(3307)) or (layer0_outputs(2882)));
    outputs(69) <= layer0_outputs(416);
    outputs(70) <= (layer0_outputs(1712)) xor (layer0_outputs(3924));
    outputs(71) <= layer0_outputs(1079);
    outputs(72) <= not(layer0_outputs(2940)) or (layer0_outputs(342));
    outputs(73) <= not(layer0_outputs(2220));
    outputs(74) <= not(layer0_outputs(798));
    outputs(75) <= layer0_outputs(3592);
    outputs(76) <= (layer0_outputs(4818)) and not (layer0_outputs(4636));
    outputs(77) <= layer0_outputs(3501);
    outputs(78) <= not(layer0_outputs(1896)) or (layer0_outputs(993));
    outputs(79) <= layer0_outputs(3830);
    outputs(80) <= not((layer0_outputs(3585)) xor (layer0_outputs(1450)));
    outputs(81) <= not(layer0_outputs(820));
    outputs(82) <= (layer0_outputs(4135)) and not (layer0_outputs(3430));
    outputs(83) <= '1';
    outputs(84) <= not(layer0_outputs(386));
    outputs(85) <= layer0_outputs(4892);
    outputs(86) <= not(layer0_outputs(833)) or (layer0_outputs(726));
    outputs(87) <= layer0_outputs(4561);
    outputs(88) <= not((layer0_outputs(3123)) xor (layer0_outputs(1187)));
    outputs(89) <= not((layer0_outputs(1805)) xor (layer0_outputs(759)));
    outputs(90) <= not(layer0_outputs(2111));
    outputs(91) <= not(layer0_outputs(3759));
    outputs(92) <= layer0_outputs(4563);
    outputs(93) <= not(layer0_outputs(5034));
    outputs(94) <= layer0_outputs(836);
    outputs(95) <= (layer0_outputs(3310)) or (layer0_outputs(4042));
    outputs(96) <= not(layer0_outputs(1303)) or (layer0_outputs(2084));
    outputs(97) <= not(layer0_outputs(3249));
    outputs(98) <= not((layer0_outputs(1161)) and (layer0_outputs(3910)));
    outputs(99) <= not((layer0_outputs(2367)) and (layer0_outputs(4736)));
    outputs(100) <= not(layer0_outputs(2889)) or (layer0_outputs(1253));
    outputs(101) <= not((layer0_outputs(4092)) xor (layer0_outputs(4472)));
    outputs(102) <= layer0_outputs(1314);
    outputs(103) <= not(layer0_outputs(1138));
    outputs(104) <= not((layer0_outputs(1610)) xor (layer0_outputs(4232)));
    outputs(105) <= not(layer0_outputs(2547)) or (layer0_outputs(4018));
    outputs(106) <= not(layer0_outputs(2719));
    outputs(107) <= not(layer0_outputs(4793)) or (layer0_outputs(2144));
    outputs(108) <= not(layer0_outputs(960));
    outputs(109) <= not(layer0_outputs(1580));
    outputs(110) <= (layer0_outputs(957)) or (layer0_outputs(1834));
    outputs(111) <= not(layer0_outputs(1538)) or (layer0_outputs(4172));
    outputs(112) <= not((layer0_outputs(3920)) xor (layer0_outputs(4713)));
    outputs(113) <= not((layer0_outputs(2825)) xor (layer0_outputs(3126)));
    outputs(114) <= not((layer0_outputs(5109)) xor (layer0_outputs(1536)));
    outputs(115) <= not(layer0_outputs(4898));
    outputs(116) <= not(layer0_outputs(4392));
    outputs(117) <= layer0_outputs(3700);
    outputs(118) <= '1';
    outputs(119) <= layer0_outputs(1137);
    outputs(120) <= not(layer0_outputs(3976));
    outputs(121) <= (layer0_outputs(3292)) xor (layer0_outputs(4951));
    outputs(122) <= layer0_outputs(3667);
    outputs(123) <= (layer0_outputs(2389)) and (layer0_outputs(4394));
    outputs(124) <= layer0_outputs(1961);
    outputs(125) <= (layer0_outputs(2900)) or (layer0_outputs(3916));
    outputs(126) <= layer0_outputs(3178);
    outputs(127) <= not((layer0_outputs(312)) or (layer0_outputs(905)));
    outputs(128) <= not(layer0_outputs(4176));
    outputs(129) <= (layer0_outputs(766)) and not (layer0_outputs(4799));
    outputs(130) <= not((layer0_outputs(676)) xor (layer0_outputs(511)));
    outputs(131) <= not(layer0_outputs(3483)) or (layer0_outputs(2640));
    outputs(132) <= layer0_outputs(4510);
    outputs(133) <= layer0_outputs(2398);
    outputs(134) <= not(layer0_outputs(1642)) or (layer0_outputs(1526));
    outputs(135) <= not((layer0_outputs(3367)) xor (layer0_outputs(3016)));
    outputs(136) <= layer0_outputs(400);
    outputs(137) <= (layer0_outputs(4425)) xor (layer0_outputs(3403));
    outputs(138) <= not((layer0_outputs(3680)) xor (layer0_outputs(2632)));
    outputs(139) <= layer0_outputs(606);
    outputs(140) <= layer0_outputs(2525);
    outputs(141) <= (layer0_outputs(1239)) xor (layer0_outputs(3533));
    outputs(142) <= (layer0_outputs(3335)) and (layer0_outputs(516));
    outputs(143) <= not(layer0_outputs(453));
    outputs(144) <= layer0_outputs(685);
    outputs(145) <= not(layer0_outputs(977));
    outputs(146) <= not((layer0_outputs(1654)) xor (layer0_outputs(2447)));
    outputs(147) <= layer0_outputs(4733);
    outputs(148) <= (layer0_outputs(4838)) and not (layer0_outputs(1));
    outputs(149) <= (layer0_outputs(3194)) and not (layer0_outputs(2954));
    outputs(150) <= (layer0_outputs(2730)) and not (layer0_outputs(2860));
    outputs(151) <= (layer0_outputs(2457)) xor (layer0_outputs(3795));
    outputs(152) <= (layer0_outputs(2169)) xor (layer0_outputs(1518));
    outputs(153) <= not(layer0_outputs(2740));
    outputs(154) <= not(layer0_outputs(1550));
    outputs(155) <= not(layer0_outputs(1881)) or (layer0_outputs(1679));
    outputs(156) <= not(layer0_outputs(5031));
    outputs(157) <= not(layer0_outputs(120));
    outputs(158) <= (layer0_outputs(4936)) xor (layer0_outputs(4052));
    outputs(159) <= not((layer0_outputs(3259)) xor (layer0_outputs(2694)));
    outputs(160) <= not(layer0_outputs(2403));
    outputs(161) <= not(layer0_outputs(3590)) or (layer0_outputs(1161));
    outputs(162) <= layer0_outputs(702);
    outputs(163) <= not((layer0_outputs(673)) or (layer0_outputs(1291)));
    outputs(164) <= (layer0_outputs(221)) and not (layer0_outputs(2399));
    outputs(165) <= not((layer0_outputs(3112)) xor (layer0_outputs(3149)));
    outputs(166) <= not(layer0_outputs(4496));
    outputs(167) <= not(layer0_outputs(3456)) or (layer0_outputs(1666));
    outputs(168) <= not(layer0_outputs(4967));
    outputs(169) <= (layer0_outputs(2603)) or (layer0_outputs(1503));
    outputs(170) <= (layer0_outputs(3310)) and not (layer0_outputs(4101));
    outputs(171) <= not((layer0_outputs(4605)) xor (layer0_outputs(3549)));
    outputs(172) <= not((layer0_outputs(4931)) and (layer0_outputs(2295)));
    outputs(173) <= not((layer0_outputs(687)) xor (layer0_outputs(4777)));
    outputs(174) <= (layer0_outputs(2860)) xor (layer0_outputs(708));
    outputs(175) <= not(layer0_outputs(747));
    outputs(176) <= not((layer0_outputs(2218)) xor (layer0_outputs(2856)));
    outputs(177) <= layer0_outputs(2769);
    outputs(178) <= layer0_outputs(652);
    outputs(179) <= layer0_outputs(1638);
    outputs(180) <= not(layer0_outputs(1877));
    outputs(181) <= not(layer0_outputs(4137)) or (layer0_outputs(3762));
    outputs(182) <= not((layer0_outputs(645)) and (layer0_outputs(3521)));
    outputs(183) <= (layer0_outputs(5105)) and (layer0_outputs(1132));
    outputs(184) <= not((layer0_outputs(3617)) and (layer0_outputs(4233)));
    outputs(185) <= not(layer0_outputs(1987));
    outputs(186) <= not((layer0_outputs(5017)) and (layer0_outputs(1715)));
    outputs(187) <= not(layer0_outputs(984));
    outputs(188) <= not(layer0_outputs(4255));
    outputs(189) <= (layer0_outputs(569)) and not (layer0_outputs(2335));
    outputs(190) <= (layer0_outputs(4627)) xor (layer0_outputs(1078));
    outputs(191) <= not((layer0_outputs(127)) and (layer0_outputs(1546)));
    outputs(192) <= not(layer0_outputs(966)) or (layer0_outputs(2974));
    outputs(193) <= not(layer0_outputs(1731)) or (layer0_outputs(988));
    outputs(194) <= layer0_outputs(2429);
    outputs(195) <= (layer0_outputs(2338)) and not (layer0_outputs(3591));
    outputs(196) <= layer0_outputs(5088);
    outputs(197) <= not(layer0_outputs(4907));
    outputs(198) <= (layer0_outputs(1598)) and not (layer0_outputs(2501));
    outputs(199) <= (layer0_outputs(498)) and not (layer0_outputs(1923));
    outputs(200) <= not((layer0_outputs(3273)) xor (layer0_outputs(394)));
    outputs(201) <= layer0_outputs(778);
    outputs(202) <= (layer0_outputs(4950)) and not (layer0_outputs(3211));
    outputs(203) <= not(layer0_outputs(1002));
    outputs(204) <= layer0_outputs(639);
    outputs(205) <= not((layer0_outputs(4988)) xor (layer0_outputs(2708)));
    outputs(206) <= layer0_outputs(2752);
    outputs(207) <= not(layer0_outputs(1700));
    outputs(208) <= not((layer0_outputs(4667)) xor (layer0_outputs(1384)));
    outputs(209) <= (layer0_outputs(3219)) or (layer0_outputs(5060));
    outputs(210) <= not((layer0_outputs(1123)) and (layer0_outputs(3189)));
    outputs(211) <= not((layer0_outputs(4902)) xor (layer0_outputs(81)));
    outputs(212) <= not(layer0_outputs(1612));
    outputs(213) <= (layer0_outputs(1400)) and (layer0_outputs(869));
    outputs(214) <= not((layer0_outputs(4055)) xor (layer0_outputs(3464)));
    outputs(215) <= layer0_outputs(2507);
    outputs(216) <= not(layer0_outputs(5075)) or (layer0_outputs(4083));
    outputs(217) <= layer0_outputs(3748);
    outputs(218) <= layer0_outputs(4048);
    outputs(219) <= (layer0_outputs(2189)) xor (layer0_outputs(3110));
    outputs(220) <= layer0_outputs(311);
    outputs(221) <= layer0_outputs(516);
    outputs(222) <= layer0_outputs(968);
    outputs(223) <= not(layer0_outputs(872));
    outputs(224) <= not(layer0_outputs(1888));
    outputs(225) <= not(layer0_outputs(1063)) or (layer0_outputs(75));
    outputs(226) <= layer0_outputs(808);
    outputs(227) <= layer0_outputs(750);
    outputs(228) <= not(layer0_outputs(1085)) or (layer0_outputs(705));
    outputs(229) <= layer0_outputs(295);
    outputs(230) <= (layer0_outputs(3966)) and not (layer0_outputs(0));
    outputs(231) <= not(layer0_outputs(4923)) or (layer0_outputs(3273));
    outputs(232) <= not((layer0_outputs(3692)) xor (layer0_outputs(3200)));
    outputs(233) <= not(layer0_outputs(189));
    outputs(234) <= layer0_outputs(3140);
    outputs(235) <= (layer0_outputs(1801)) xor (layer0_outputs(1535));
    outputs(236) <= not((layer0_outputs(1073)) and (layer0_outputs(3892)));
    outputs(237) <= not((layer0_outputs(2268)) xor (layer0_outputs(2341)));
    outputs(238) <= not((layer0_outputs(1546)) and (layer0_outputs(1847)));
    outputs(239) <= layer0_outputs(4965);
    outputs(240) <= (layer0_outputs(4604)) and (layer0_outputs(2752));
    outputs(241) <= '1';
    outputs(242) <= layer0_outputs(4532);
    outputs(243) <= (layer0_outputs(779)) and not (layer0_outputs(688));
    outputs(244) <= layer0_outputs(4969);
    outputs(245) <= (layer0_outputs(492)) or (layer0_outputs(3514));
    outputs(246) <= (layer0_outputs(2365)) and (layer0_outputs(4090));
    outputs(247) <= layer0_outputs(4651);
    outputs(248) <= not(layer0_outputs(4907));
    outputs(249) <= not((layer0_outputs(3730)) xor (layer0_outputs(1635)));
    outputs(250) <= not((layer0_outputs(614)) xor (layer0_outputs(2731)));
    outputs(251) <= not(layer0_outputs(1816));
    outputs(252) <= (layer0_outputs(1340)) xor (layer0_outputs(295));
    outputs(253) <= not((layer0_outputs(2724)) and (layer0_outputs(914)));
    outputs(254) <= (layer0_outputs(665)) and not (layer0_outputs(4392));
    outputs(255) <= (layer0_outputs(4196)) and (layer0_outputs(2162));
    outputs(256) <= not(layer0_outputs(4129)) or (layer0_outputs(1634));
    outputs(257) <= layer0_outputs(1513);
    outputs(258) <= (layer0_outputs(3390)) xor (layer0_outputs(2179));
    outputs(259) <= not((layer0_outputs(2931)) xor (layer0_outputs(2682)));
    outputs(260) <= (layer0_outputs(1458)) and (layer0_outputs(2279));
    outputs(261) <= (layer0_outputs(1608)) xor (layer0_outputs(3984));
    outputs(262) <= layer0_outputs(2558);
    outputs(263) <= not((layer0_outputs(4128)) or (layer0_outputs(2388)));
    outputs(264) <= (layer0_outputs(1186)) and not (layer0_outputs(297));
    outputs(265) <= layer0_outputs(4080);
    outputs(266) <= layer0_outputs(4628);
    outputs(267) <= layer0_outputs(4295);
    outputs(268) <= (layer0_outputs(4838)) and (layer0_outputs(240));
    outputs(269) <= not(layer0_outputs(4374));
    outputs(270) <= not(layer0_outputs(3811));
    outputs(271) <= (layer0_outputs(4201)) or (layer0_outputs(1472));
    outputs(272) <= not(layer0_outputs(2893));
    outputs(273) <= (layer0_outputs(4789)) and (layer0_outputs(3160));
    outputs(274) <= not(layer0_outputs(2988));
    outputs(275) <= '1';
    outputs(276) <= (layer0_outputs(735)) xor (layer0_outputs(3173));
    outputs(277) <= layer0_outputs(2566);
    outputs(278) <= (layer0_outputs(1156)) xor (layer0_outputs(3698));
    outputs(279) <= layer0_outputs(401);
    outputs(280) <= not(layer0_outputs(737));
    outputs(281) <= not((layer0_outputs(64)) xor (layer0_outputs(3329)));
    outputs(282) <= not(layer0_outputs(1380));
    outputs(283) <= layer0_outputs(4847);
    outputs(284) <= not(layer0_outputs(1720)) or (layer0_outputs(746));
    outputs(285) <= layer0_outputs(311);
    outputs(286) <= not((layer0_outputs(1296)) xor (layer0_outputs(4277)));
    outputs(287) <= not((layer0_outputs(1884)) xor (layer0_outputs(3845)));
    outputs(288) <= (layer0_outputs(2222)) or (layer0_outputs(3185));
    outputs(289) <= (layer0_outputs(4551)) and not (layer0_outputs(3755));
    outputs(290) <= not((layer0_outputs(2516)) or (layer0_outputs(3786)));
    outputs(291) <= not(layer0_outputs(2716));
    outputs(292) <= (layer0_outputs(3888)) and not (layer0_outputs(4288));
    outputs(293) <= (layer0_outputs(505)) and not (layer0_outputs(4585));
    outputs(294) <= (layer0_outputs(4474)) and not (layer0_outputs(3775));
    outputs(295) <= not(layer0_outputs(118));
    outputs(296) <= not((layer0_outputs(774)) or (layer0_outputs(636)));
    outputs(297) <= not((layer0_outputs(3742)) and (layer0_outputs(4470)));
    outputs(298) <= not(layer0_outputs(3834)) or (layer0_outputs(4054));
    outputs(299) <= layer0_outputs(838);
    outputs(300) <= (layer0_outputs(122)) xor (layer0_outputs(1025));
    outputs(301) <= layer0_outputs(3923);
    outputs(302) <= not((layer0_outputs(5097)) and (layer0_outputs(1779)));
    outputs(303) <= (layer0_outputs(3380)) and not (layer0_outputs(1642));
    outputs(304) <= not(layer0_outputs(2260));
    outputs(305) <= (layer0_outputs(3045)) or (layer0_outputs(3256));
    outputs(306) <= layer0_outputs(3384);
    outputs(307) <= not(layer0_outputs(59));
    outputs(308) <= not(layer0_outputs(3967));
    outputs(309) <= layer0_outputs(4904);
    outputs(310) <= layer0_outputs(3783);
    outputs(311) <= (layer0_outputs(196)) xor (layer0_outputs(1288));
    outputs(312) <= layer0_outputs(1311);
    outputs(313) <= not(layer0_outputs(704));
    outputs(314) <= layer0_outputs(1106);
    outputs(315) <= not(layer0_outputs(4859));
    outputs(316) <= not((layer0_outputs(4206)) or (layer0_outputs(62)));
    outputs(317) <= (layer0_outputs(2362)) or (layer0_outputs(1264));
    outputs(318) <= not(layer0_outputs(4766));
    outputs(319) <= layer0_outputs(4356);
    outputs(320) <= not((layer0_outputs(3075)) and (layer0_outputs(833)));
    outputs(321) <= not(layer0_outputs(2692)) or (layer0_outputs(3007));
    outputs(322) <= not(layer0_outputs(5070));
    outputs(323) <= not(layer0_outputs(2301));
    outputs(324) <= not(layer0_outputs(2181));
    outputs(325) <= not(layer0_outputs(4983));
    outputs(326) <= not((layer0_outputs(4360)) xor (layer0_outputs(1966)));
    outputs(327) <= (layer0_outputs(702)) or (layer0_outputs(2138));
    outputs(328) <= not((layer0_outputs(692)) or (layer0_outputs(1479)));
    outputs(329) <= layer0_outputs(4696);
    outputs(330) <= not((layer0_outputs(1428)) xor (layer0_outputs(2227)));
    outputs(331) <= not(layer0_outputs(1273));
    outputs(332) <= layer0_outputs(3147);
    outputs(333) <= (layer0_outputs(4388)) xor (layer0_outputs(2201));
    outputs(334) <= (layer0_outputs(2662)) or (layer0_outputs(2959));
    outputs(335) <= (layer0_outputs(1232)) xor (layer0_outputs(876));
    outputs(336) <= layer0_outputs(3481);
    outputs(337) <= (layer0_outputs(3277)) or (layer0_outputs(18));
    outputs(338) <= layer0_outputs(4651);
    outputs(339) <= not(layer0_outputs(678)) or (layer0_outputs(1532));
    outputs(340) <= layer0_outputs(5111);
    outputs(341) <= not((layer0_outputs(1469)) xor (layer0_outputs(4060)));
    outputs(342) <= not(layer0_outputs(1391)) or (layer0_outputs(4327));
    outputs(343) <= not(layer0_outputs(2161));
    outputs(344) <= not(layer0_outputs(2877));
    outputs(345) <= (layer0_outputs(3507)) and not (layer0_outputs(803));
    outputs(346) <= not(layer0_outputs(1710)) or (layer0_outputs(1186));
    outputs(347) <= not((layer0_outputs(4834)) or (layer0_outputs(4900)));
    outputs(348) <= (layer0_outputs(2283)) and (layer0_outputs(1569));
    outputs(349) <= (layer0_outputs(2757)) and (layer0_outputs(2645));
    outputs(350) <= (layer0_outputs(1749)) or (layer0_outputs(2261));
    outputs(351) <= not((layer0_outputs(2657)) and (layer0_outputs(3248)));
    outputs(352) <= not((layer0_outputs(4161)) or (layer0_outputs(820)));
    outputs(353) <= not(layer0_outputs(180)) or (layer0_outputs(3707));
    outputs(354) <= not((layer0_outputs(2046)) or (layer0_outputs(765)));
    outputs(355) <= not(layer0_outputs(811)) or (layer0_outputs(959));
    outputs(356) <= not((layer0_outputs(3690)) or (layer0_outputs(733)));
    outputs(357) <= not((layer0_outputs(4001)) xor (layer0_outputs(1594)));
    outputs(358) <= (layer0_outputs(4369)) and (layer0_outputs(711));
    outputs(359) <= not((layer0_outputs(2276)) or (layer0_outputs(1920)));
    outputs(360) <= not((layer0_outputs(3128)) or (layer0_outputs(2472)));
    outputs(361) <= not((layer0_outputs(1860)) xor (layer0_outputs(1014)));
    outputs(362) <= (layer0_outputs(1701)) and (layer0_outputs(4608));
    outputs(363) <= (layer0_outputs(2585)) xor (layer0_outputs(652));
    outputs(364) <= not((layer0_outputs(3637)) or (layer0_outputs(1476)));
    outputs(365) <= layer0_outputs(4726);
    outputs(366) <= not(layer0_outputs(4290));
    outputs(367) <= layer0_outputs(3094);
    outputs(368) <= layer0_outputs(4387);
    outputs(369) <= not(layer0_outputs(4541));
    outputs(370) <= layer0_outputs(4913);
    outputs(371) <= layer0_outputs(2230);
    outputs(372) <= (layer0_outputs(2260)) xor (layer0_outputs(1301));
    outputs(373) <= (layer0_outputs(1232)) xor (layer0_outputs(2527));
    outputs(374) <= not(layer0_outputs(178));
    outputs(375) <= layer0_outputs(2679);
    outputs(376) <= (layer0_outputs(2786)) xor (layer0_outputs(4318));
    outputs(377) <= not(layer0_outputs(1028));
    outputs(378) <= not(layer0_outputs(795));
    outputs(379) <= not(layer0_outputs(3473)) or (layer0_outputs(4817));
    outputs(380) <= layer0_outputs(4914);
    outputs(381) <= (layer0_outputs(2355)) xor (layer0_outputs(3321));
    outputs(382) <= not(layer0_outputs(210));
    outputs(383) <= (layer0_outputs(3535)) and (layer0_outputs(3732));
    outputs(384) <= not(layer0_outputs(4735)) or (layer0_outputs(823));
    outputs(385) <= not(layer0_outputs(187));
    outputs(386) <= layer0_outputs(1565);
    outputs(387) <= not((layer0_outputs(1158)) and (layer0_outputs(1558)));
    outputs(388) <= not(layer0_outputs(4520));
    outputs(389) <= not((layer0_outputs(37)) and (layer0_outputs(1818)));
    outputs(390) <= layer0_outputs(4797);
    outputs(391) <= not(layer0_outputs(456)) or (layer0_outputs(2475));
    outputs(392) <= not((layer0_outputs(496)) and (layer0_outputs(3500)));
    outputs(393) <= layer0_outputs(4443);
    outputs(394) <= layer0_outputs(3808);
    outputs(395) <= layer0_outputs(2121);
    outputs(396) <= layer0_outputs(3935);
    outputs(397) <= not((layer0_outputs(445)) and (layer0_outputs(1501)));
    outputs(398) <= not(layer0_outputs(2552)) or (layer0_outputs(548));
    outputs(399) <= not(layer0_outputs(264)) or (layer0_outputs(3418));
    outputs(400) <= (layer0_outputs(7)) xor (layer0_outputs(2173));
    outputs(401) <= not(layer0_outputs(806));
    outputs(402) <= layer0_outputs(4501);
    outputs(403) <= not((layer0_outputs(3527)) or (layer0_outputs(1480)));
    outputs(404) <= (layer0_outputs(4507)) and (layer0_outputs(2177));
    outputs(405) <= (layer0_outputs(2059)) and not (layer0_outputs(4185));
    outputs(406) <= (layer0_outputs(371)) and not (layer0_outputs(3882));
    outputs(407) <= not(layer0_outputs(1637));
    outputs(408) <= layer0_outputs(2019);
    outputs(409) <= not(layer0_outputs(5000));
    outputs(410) <= (layer0_outputs(4661)) and not (layer0_outputs(307));
    outputs(411) <= not(layer0_outputs(3075));
    outputs(412) <= layer0_outputs(344);
    outputs(413) <= not(layer0_outputs(1774)) or (layer0_outputs(4394));
    outputs(414) <= not(layer0_outputs(3192));
    outputs(415) <= layer0_outputs(4354);
    outputs(416) <= not(layer0_outputs(2049));
    outputs(417) <= not((layer0_outputs(4923)) and (layer0_outputs(3976)));
    outputs(418) <= not(layer0_outputs(610));
    outputs(419) <= layer0_outputs(296);
    outputs(420) <= (layer0_outputs(2105)) xor (layer0_outputs(953));
    outputs(421) <= not(layer0_outputs(4248)) or (layer0_outputs(2480));
    outputs(422) <= layer0_outputs(4560);
    outputs(423) <= not((layer0_outputs(206)) or (layer0_outputs(2406)));
    outputs(424) <= layer0_outputs(1420);
    outputs(425) <= not(layer0_outputs(2132)) or (layer0_outputs(4491));
    outputs(426) <= (layer0_outputs(3290)) xor (layer0_outputs(4046));
    outputs(427) <= (layer0_outputs(3222)) and not (layer0_outputs(228));
    outputs(428) <= (layer0_outputs(4425)) or (layer0_outputs(1005));
    outputs(429) <= (layer0_outputs(2920)) and not (layer0_outputs(4179));
    outputs(430) <= not((layer0_outputs(3846)) and (layer0_outputs(2987)));
    outputs(431) <= not((layer0_outputs(3509)) or (layer0_outputs(4757)));
    outputs(432) <= layer0_outputs(4166);
    outputs(433) <= layer0_outputs(2213);
    outputs(434) <= not(layer0_outputs(3395)) or (layer0_outputs(4205));
    outputs(435) <= layer0_outputs(42);
    outputs(436) <= (layer0_outputs(4050)) and not (layer0_outputs(3152));
    outputs(437) <= layer0_outputs(906);
    outputs(438) <= layer0_outputs(4424);
    outputs(439) <= layer0_outputs(1304);
    outputs(440) <= (layer0_outputs(2997)) and (layer0_outputs(591));
    outputs(441) <= layer0_outputs(353);
    outputs(442) <= not(layer0_outputs(1140));
    outputs(443) <= not(layer0_outputs(44));
    outputs(444) <= not((layer0_outputs(3846)) and (layer0_outputs(4496)));
    outputs(445) <= not(layer0_outputs(3908));
    outputs(446) <= not(layer0_outputs(764)) or (layer0_outputs(4754));
    outputs(447) <= not(layer0_outputs(4943)) or (layer0_outputs(3289));
    outputs(448) <= not(layer0_outputs(2300));
    outputs(449) <= '0';
    outputs(450) <= not((layer0_outputs(2865)) and (layer0_outputs(1279)));
    outputs(451) <= (layer0_outputs(684)) or (layer0_outputs(588));
    outputs(452) <= (layer0_outputs(4017)) xor (layer0_outputs(3003));
    outputs(453) <= not((layer0_outputs(2886)) xor (layer0_outputs(3253)));
    outputs(454) <= not((layer0_outputs(4553)) xor (layer0_outputs(4723)));
    outputs(455) <= (layer0_outputs(763)) xor (layer0_outputs(5005));
    outputs(456) <= not(layer0_outputs(2228));
    outputs(457) <= not(layer0_outputs(3591)) or (layer0_outputs(723));
    outputs(458) <= (layer0_outputs(3676)) xor (layer0_outputs(3917));
    outputs(459) <= (layer0_outputs(2688)) or (layer0_outputs(5040));
    outputs(460) <= layer0_outputs(858);
    outputs(461) <= (layer0_outputs(3442)) xor (layer0_outputs(1086));
    outputs(462) <= not(layer0_outputs(4882));
    outputs(463) <= layer0_outputs(4628);
    outputs(464) <= layer0_outputs(4103);
    outputs(465) <= not(layer0_outputs(2600));
    outputs(466) <= layer0_outputs(5100);
    outputs(467) <= not((layer0_outputs(1837)) and (layer0_outputs(2898)));
    outputs(468) <= layer0_outputs(2802);
    outputs(469) <= layer0_outputs(3091);
    outputs(470) <= not(layer0_outputs(3850));
    outputs(471) <= (layer0_outputs(4306)) xor (layer0_outputs(4709));
    outputs(472) <= layer0_outputs(3225);
    outputs(473) <= not((layer0_outputs(14)) or (layer0_outputs(4970)));
    outputs(474) <= not(layer0_outputs(661)) or (layer0_outputs(3172));
    outputs(475) <= not(layer0_outputs(2693));
    outputs(476) <= not(layer0_outputs(683)) or (layer0_outputs(4227));
    outputs(477) <= not((layer0_outputs(4460)) xor (layer0_outputs(3468)));
    outputs(478) <= not(layer0_outputs(1786));
    outputs(479) <= not(layer0_outputs(3467)) or (layer0_outputs(2717));
    outputs(480) <= layer0_outputs(2789);
    outputs(481) <= not(layer0_outputs(2805));
    outputs(482) <= not((layer0_outputs(2328)) xor (layer0_outputs(4800)));
    outputs(483) <= not(layer0_outputs(3483));
    outputs(484) <= not((layer0_outputs(2193)) and (layer0_outputs(1614)));
    outputs(485) <= not(layer0_outputs(1332));
    outputs(486) <= (layer0_outputs(2577)) or (layer0_outputs(1471));
    outputs(487) <= layer0_outputs(3492);
    outputs(488) <= layer0_outputs(477);
    outputs(489) <= layer0_outputs(4121);
    outputs(490) <= layer0_outputs(4922);
    outputs(491) <= not((layer0_outputs(1422)) xor (layer0_outputs(3072)));
    outputs(492) <= (layer0_outputs(4855)) and (layer0_outputs(1414));
    outputs(493) <= (layer0_outputs(4665)) and not (layer0_outputs(3224));
    outputs(494) <= not(layer0_outputs(519));
    outputs(495) <= not(layer0_outputs(815)) or (layer0_outputs(1390));
    outputs(496) <= not(layer0_outputs(1760));
    outputs(497) <= layer0_outputs(804);
    outputs(498) <= not(layer0_outputs(3325));
    outputs(499) <= (layer0_outputs(418)) or (layer0_outputs(2460));
    outputs(500) <= (layer0_outputs(4019)) or (layer0_outputs(3354));
    outputs(501) <= not((layer0_outputs(2487)) or (layer0_outputs(4692)));
    outputs(502) <= not(layer0_outputs(1955));
    outputs(503) <= (layer0_outputs(32)) and not (layer0_outputs(3452));
    outputs(504) <= layer0_outputs(319);
    outputs(505) <= not(layer0_outputs(2552));
    outputs(506) <= not((layer0_outputs(3331)) xor (layer0_outputs(3671)));
    outputs(507) <= layer0_outputs(230);
    outputs(508) <= not(layer0_outputs(1520));
    outputs(509) <= not(layer0_outputs(3152));
    outputs(510) <= not(layer0_outputs(4541));
    outputs(511) <= not((layer0_outputs(2340)) and (layer0_outputs(2452)));
    outputs(512) <= layer0_outputs(2060);
    outputs(513) <= (layer0_outputs(4677)) and (layer0_outputs(253));
    outputs(514) <= layer0_outputs(1998);
    outputs(515) <= layer0_outputs(2764);
    outputs(516) <= (layer0_outputs(850)) xor (layer0_outputs(368));
    outputs(517) <= (layer0_outputs(961)) xor (layer0_outputs(1566));
    outputs(518) <= (layer0_outputs(2108)) and not (layer0_outputs(2892));
    outputs(519) <= not((layer0_outputs(3400)) or (layer0_outputs(363)));
    outputs(520) <= (layer0_outputs(3245)) and (layer0_outputs(3287));
    outputs(521) <= (layer0_outputs(3884)) and (layer0_outputs(2470));
    outputs(522) <= not(layer0_outputs(4383));
    outputs(523) <= (layer0_outputs(241)) and (layer0_outputs(4211));
    outputs(524) <= (layer0_outputs(3287)) and not (layer0_outputs(908));
    outputs(525) <= not(layer0_outputs(127));
    outputs(526) <= not((layer0_outputs(4827)) or (layer0_outputs(2044)));
    outputs(527) <= not(layer0_outputs(1421));
    outputs(528) <= (layer0_outputs(4190)) and (layer0_outputs(3766));
    outputs(529) <= (layer0_outputs(4555)) and not (layer0_outputs(3706));
    outputs(530) <= (layer0_outputs(3381)) and (layer0_outputs(1019));
    outputs(531) <= (layer0_outputs(3740)) and (layer0_outputs(405));
    outputs(532) <= (layer0_outputs(3086)) xor (layer0_outputs(4312));
    outputs(533) <= not((layer0_outputs(3099)) or (layer0_outputs(4447)));
    outputs(534) <= not((layer0_outputs(475)) xor (layer0_outputs(393)));
    outputs(535) <= (layer0_outputs(3498)) and not (layer0_outputs(4359));
    outputs(536) <= not(layer0_outputs(4467)) or (layer0_outputs(4001));
    outputs(537) <= '0';
    outputs(538) <= (layer0_outputs(2264)) and not (layer0_outputs(1455));
    outputs(539) <= layer0_outputs(1189);
    outputs(540) <= (layer0_outputs(397)) and not (layer0_outputs(3184));
    outputs(541) <= (layer0_outputs(4072)) and not (layer0_outputs(4884));
    outputs(542) <= (layer0_outputs(4235)) and not (layer0_outputs(2166));
    outputs(543) <= not((layer0_outputs(4036)) xor (layer0_outputs(1552)));
    outputs(544) <= layer0_outputs(981);
    outputs(545) <= '0';
    outputs(546) <= (layer0_outputs(4935)) xor (layer0_outputs(1379));
    outputs(547) <= not((layer0_outputs(3289)) or (layer0_outputs(1087)));
    outputs(548) <= not((layer0_outputs(898)) xor (layer0_outputs(163)));
    outputs(549) <= (layer0_outputs(425)) and (layer0_outputs(2450));
    outputs(550) <= (layer0_outputs(1786)) and (layer0_outputs(1592));
    outputs(551) <= (layer0_outputs(2920)) and (layer0_outputs(1014));
    outputs(552) <= (layer0_outputs(309)) and (layer0_outputs(367));
    outputs(553) <= (layer0_outputs(2140)) xor (layer0_outputs(1770));
    outputs(554) <= not(layer0_outputs(3304)) or (layer0_outputs(2962));
    outputs(555) <= (layer0_outputs(112)) and not (layer0_outputs(3430));
    outputs(556) <= not((layer0_outputs(2993)) xor (layer0_outputs(2737)));
    outputs(557) <= not(layer0_outputs(459));
    outputs(558) <= not(layer0_outputs(2787));
    outputs(559) <= not((layer0_outputs(2702)) or (layer0_outputs(2753)));
    outputs(560) <= (layer0_outputs(1814)) xor (layer0_outputs(3629));
    outputs(561) <= not(layer0_outputs(2672));
    outputs(562) <= '0';
    outputs(563) <= not((layer0_outputs(135)) xor (layer0_outputs(1182)));
    outputs(564) <= not(layer0_outputs(4044));
    outputs(565) <= layer0_outputs(4815);
    outputs(566) <= (layer0_outputs(1058)) xor (layer0_outputs(2424));
    outputs(567) <= not((layer0_outputs(2520)) or (layer0_outputs(3292)));
    outputs(568) <= not((layer0_outputs(3614)) and (layer0_outputs(3351)));
    outputs(569) <= not((layer0_outputs(1831)) or (layer0_outputs(269)));
    outputs(570) <= layer0_outputs(5071);
    outputs(571) <= (layer0_outputs(243)) and (layer0_outputs(1381));
    outputs(572) <= (layer0_outputs(3020)) and not (layer0_outputs(4731));
    outputs(573) <= layer0_outputs(3910);
    outputs(574) <= not((layer0_outputs(3750)) or (layer0_outputs(508)));
    outputs(575) <= (layer0_outputs(1963)) and not (layer0_outputs(1300));
    outputs(576) <= (layer0_outputs(3079)) xor (layer0_outputs(4133));
    outputs(577) <= (layer0_outputs(2417)) and not (layer0_outputs(1473));
    outputs(578) <= layer0_outputs(1784);
    outputs(579) <= (layer0_outputs(1710)) and not (layer0_outputs(4636));
    outputs(580) <= (layer0_outputs(5078)) and not (layer0_outputs(1474));
    outputs(581) <= (layer0_outputs(2143)) and (layer0_outputs(577));
    outputs(582) <= (layer0_outputs(821)) and (layer0_outputs(818));
    outputs(583) <= (layer0_outputs(4772)) and not (layer0_outputs(2982));
    outputs(584) <= (layer0_outputs(131)) and (layer0_outputs(601));
    outputs(585) <= (layer0_outputs(1579)) and not (layer0_outputs(882));
    outputs(586) <= (layer0_outputs(354)) and not (layer0_outputs(4921));
    outputs(587) <= (layer0_outputs(3423)) and not (layer0_outputs(700));
    outputs(588) <= (layer0_outputs(3709)) and not (layer0_outputs(2263));
    outputs(589) <= not((layer0_outputs(4556)) or (layer0_outputs(2247)));
    outputs(590) <= layer0_outputs(1056);
    outputs(591) <= (layer0_outputs(4444)) xor (layer0_outputs(2797));
    outputs(592) <= not((layer0_outputs(128)) or (layer0_outputs(1432)));
    outputs(593) <= not(layer0_outputs(4877));
    outputs(594) <= not(layer0_outputs(2444));
    outputs(595) <= layer0_outputs(4429);
    outputs(596) <= (layer0_outputs(1489)) and not (layer0_outputs(3419));
    outputs(597) <= (layer0_outputs(4736)) and not (layer0_outputs(3474));
    outputs(598) <= layer0_outputs(2829);
    outputs(599) <= not(layer0_outputs(1492));
    outputs(600) <= (layer0_outputs(1977)) and not (layer0_outputs(2298));
    outputs(601) <= (layer0_outputs(2864)) and not (layer0_outputs(5047));
    outputs(602) <= (layer0_outputs(4462)) and not (layer0_outputs(906));
    outputs(603) <= (layer0_outputs(4380)) and not (layer0_outputs(3659));
    outputs(604) <= not(layer0_outputs(3141));
    outputs(605) <= (layer0_outputs(1261)) xor (layer0_outputs(3408));
    outputs(606) <= layer0_outputs(4091);
    outputs(607) <= not((layer0_outputs(694)) or (layer0_outputs(548)));
    outputs(608) <= '0';
    outputs(609) <= not(layer0_outputs(750));
    outputs(610) <= not((layer0_outputs(2353)) or (layer0_outputs(2378)));
    outputs(611) <= not((layer0_outputs(4972)) and (layer0_outputs(1467)));
    outputs(612) <= not((layer0_outputs(5089)) xor (layer0_outputs(291)));
    outputs(613) <= not((layer0_outputs(3196)) or (layer0_outputs(4436)));
    outputs(614) <= not(layer0_outputs(4536));
    outputs(615) <= layer0_outputs(2621);
    outputs(616) <= layer0_outputs(4324);
    outputs(617) <= (layer0_outputs(2748)) and not (layer0_outputs(4826));
    outputs(618) <= (layer0_outputs(4035)) and (layer0_outputs(302));
    outputs(619) <= layer0_outputs(2309);
    outputs(620) <= (layer0_outputs(4673)) and not (layer0_outputs(3661));
    outputs(621) <= (layer0_outputs(766)) and (layer0_outputs(3080));
    outputs(622) <= (layer0_outputs(970)) and not (layer0_outputs(2571));
    outputs(623) <= (layer0_outputs(2806)) and (layer0_outputs(1198));
    outputs(624) <= (layer0_outputs(3128)) and not (layer0_outputs(834));
    outputs(625) <= (layer0_outputs(2879)) xor (layer0_outputs(2025));
    outputs(626) <= not((layer0_outputs(2020)) or (layer0_outputs(4954)));
    outputs(627) <= '0';
    outputs(628) <= layer0_outputs(4132);
    outputs(629) <= layer0_outputs(4357);
    outputs(630) <= not((layer0_outputs(1125)) or (layer0_outputs(3038)));
    outputs(631) <= (layer0_outputs(3708)) and not (layer0_outputs(2828));
    outputs(632) <= not((layer0_outputs(3107)) or (layer0_outputs(136)));
    outputs(633) <= (layer0_outputs(4919)) xor (layer0_outputs(2880));
    outputs(634) <= not(layer0_outputs(3912));
    outputs(635) <= not((layer0_outputs(1778)) or (layer0_outputs(1173)));
    outputs(636) <= (layer0_outputs(4139)) and not (layer0_outputs(463));
    outputs(637) <= not(layer0_outputs(3639));
    outputs(638) <= not((layer0_outputs(3685)) or (layer0_outputs(693)));
    outputs(639) <= not(layer0_outputs(3335));
    outputs(640) <= (layer0_outputs(4734)) and not (layer0_outputs(4010));
    outputs(641) <= (layer0_outputs(1259)) and (layer0_outputs(3878));
    outputs(642) <= not((layer0_outputs(3745)) or (layer0_outputs(2044)));
    outputs(643) <= not((layer0_outputs(1903)) or (layer0_outputs(279)));
    outputs(644) <= (layer0_outputs(3025)) and not (layer0_outputs(3398));
    outputs(645) <= (layer0_outputs(3553)) and (layer0_outputs(2611));
    outputs(646) <= not((layer0_outputs(952)) xor (layer0_outputs(888)));
    outputs(647) <= not(layer0_outputs(782));
    outputs(648) <= layer0_outputs(339);
    outputs(649) <= layer0_outputs(3429);
    outputs(650) <= layer0_outputs(1120);
    outputs(651) <= layer0_outputs(1181);
    outputs(652) <= not((layer0_outputs(184)) or (layer0_outputs(3984)));
    outputs(653) <= (layer0_outputs(2014)) and not (layer0_outputs(3988));
    outputs(654) <= not(layer0_outputs(4164));
    outputs(655) <= not(layer0_outputs(1467));
    outputs(656) <= (layer0_outputs(3400)) xor (layer0_outputs(2267));
    outputs(657) <= not(layer0_outputs(3522));
    outputs(658) <= layer0_outputs(4248);
    outputs(659) <= not(layer0_outputs(4069));
    outputs(660) <= (layer0_outputs(93)) and not (layer0_outputs(1599));
    outputs(661) <= not(layer0_outputs(1887));
    outputs(662) <= (layer0_outputs(3518)) and (layer0_outputs(4807));
    outputs(663) <= not(layer0_outputs(2508));
    outputs(664) <= (layer0_outputs(1976)) and not (layer0_outputs(720));
    outputs(665) <= layer0_outputs(4751);
    outputs(666) <= (layer0_outputs(4903)) xor (layer0_outputs(4586));
    outputs(667) <= layer0_outputs(2785);
    outputs(668) <= (layer0_outputs(1718)) and not (layer0_outputs(2097));
    outputs(669) <= (layer0_outputs(3815)) and (layer0_outputs(1872));
    outputs(670) <= (layer0_outputs(2483)) and not (layer0_outputs(4158));
    outputs(671) <= (layer0_outputs(3810)) and (layer0_outputs(2152));
    outputs(672) <= (layer0_outputs(354)) and not (layer0_outputs(1285));
    outputs(673) <= (layer0_outputs(4795)) xor (layer0_outputs(2937));
    outputs(674) <= (layer0_outputs(3758)) and not (layer0_outputs(4618));
    outputs(675) <= not(layer0_outputs(3894));
    outputs(676) <= not((layer0_outputs(3415)) or (layer0_outputs(179)));
    outputs(677) <= not(layer0_outputs(2122));
    outputs(678) <= layer0_outputs(4537);
    outputs(679) <= not((layer0_outputs(4899)) or (layer0_outputs(4431)));
    outputs(680) <= (layer0_outputs(2130)) and not (layer0_outputs(175));
    outputs(681) <= not((layer0_outputs(4818)) or (layer0_outputs(48)));
    outputs(682) <= (layer0_outputs(2151)) and not (layer0_outputs(869));
    outputs(683) <= (layer0_outputs(790)) and (layer0_outputs(313));
    outputs(684) <= not(layer0_outputs(1651)) or (layer0_outputs(1135));
    outputs(685) <= (layer0_outputs(3032)) and not (layer0_outputs(3526));
    outputs(686) <= layer0_outputs(1788);
    outputs(687) <= layer0_outputs(4040);
    outputs(688) <= '0';
    outputs(689) <= (layer0_outputs(1085)) or (layer0_outputs(3211));
    outputs(690) <= (layer0_outputs(938)) and (layer0_outputs(197));
    outputs(691) <= not((layer0_outputs(2070)) xor (layer0_outputs(5094)));
    outputs(692) <= not(layer0_outputs(2286));
    outputs(693) <= not(layer0_outputs(1094)) or (layer0_outputs(2219));
    outputs(694) <= not(layer0_outputs(4478));
    outputs(695) <= (layer0_outputs(2464)) and not (layer0_outputs(846));
    outputs(696) <= (layer0_outputs(2863)) and not (layer0_outputs(2570));
    outputs(697) <= layer0_outputs(2211);
    outputs(698) <= not(layer0_outputs(232));
    outputs(699) <= (layer0_outputs(1735)) and (layer0_outputs(1838));
    outputs(700) <= not((layer0_outputs(2095)) or (layer0_outputs(4086)));
    outputs(701) <= (layer0_outputs(4846)) and not (layer0_outputs(2498));
    outputs(702) <= (layer0_outputs(1037)) and not (layer0_outputs(4423));
    outputs(703) <= not(layer0_outputs(4932));
    outputs(704) <= not(layer0_outputs(2529));
    outputs(705) <= (layer0_outputs(3718)) and not (layer0_outputs(4945));
    outputs(706) <= (layer0_outputs(1683)) and not (layer0_outputs(4538));
    outputs(707) <= (layer0_outputs(3633)) xor (layer0_outputs(2163));
    outputs(708) <= (layer0_outputs(3967)) and (layer0_outputs(1963));
    outputs(709) <= (layer0_outputs(1672)) and (layer0_outputs(1374));
    outputs(710) <= (layer0_outputs(2369)) and (layer0_outputs(156));
    outputs(711) <= not(layer0_outputs(1325));
    outputs(712) <= (layer0_outputs(3859)) and not (layer0_outputs(627));
    outputs(713) <= layer0_outputs(3740);
    outputs(714) <= (layer0_outputs(1958)) and not (layer0_outputs(316));
    outputs(715) <= not((layer0_outputs(4771)) or (layer0_outputs(1119)));
    outputs(716) <= (layer0_outputs(415)) and (layer0_outputs(2395));
    outputs(717) <= not(layer0_outputs(635));
    outputs(718) <= (layer0_outputs(1730)) and (layer0_outputs(4808));
    outputs(719) <= (layer0_outputs(292)) and not (layer0_outputs(2659));
    outputs(720) <= not(layer0_outputs(1603));
    outputs(721) <= (layer0_outputs(4138)) and (layer0_outputs(433));
    outputs(722) <= not(layer0_outputs(686)) or (layer0_outputs(4324));
    outputs(723) <= (layer0_outputs(137)) xor (layer0_outputs(1676));
    outputs(724) <= not(layer0_outputs(1195));
    outputs(725) <= (layer0_outputs(1932)) and not (layer0_outputs(3056));
    outputs(726) <= (layer0_outputs(2178)) and (layer0_outputs(1907));
    outputs(727) <= not(layer0_outputs(2741));
    outputs(728) <= not(layer0_outputs(2824));
    outputs(729) <= (layer0_outputs(1029)) and not (layer0_outputs(2009));
    outputs(730) <= (layer0_outputs(1313)) and not (layer0_outputs(2906));
    outputs(731) <= (layer0_outputs(1631)) and (layer0_outputs(2379));
    outputs(732) <= layer0_outputs(774);
    outputs(733) <= (layer0_outputs(2670)) xor (layer0_outputs(1525));
    outputs(734) <= not(layer0_outputs(2223));
    outputs(735) <= not(layer0_outputs(4701));
    outputs(736) <= not(layer0_outputs(2528));
    outputs(737) <= layer0_outputs(149);
    outputs(738) <= layer0_outputs(4286);
    outputs(739) <= (layer0_outputs(2619)) and (layer0_outputs(1695));
    outputs(740) <= (layer0_outputs(3921)) and (layer0_outputs(2782));
    outputs(741) <= (layer0_outputs(1719)) and not (layer0_outputs(4291));
    outputs(742) <= not(layer0_outputs(5108));
    outputs(743) <= not(layer0_outputs(4586));
    outputs(744) <= not((layer0_outputs(4642)) or (layer0_outputs(3543)));
    outputs(745) <= not(layer0_outputs(860));
    outputs(746) <= (layer0_outputs(3598)) and not (layer0_outputs(3033));
    outputs(747) <= '0';
    outputs(748) <= (layer0_outputs(603)) and (layer0_outputs(2817));
    outputs(749) <= (layer0_outputs(3790)) xor (layer0_outputs(1605));
    outputs(750) <= (layer0_outputs(2767)) xor (layer0_outputs(4548));
    outputs(751) <= (layer0_outputs(5057)) xor (layer0_outputs(4693));
    outputs(752) <= layer0_outputs(2174);
    outputs(753) <= not(layer0_outputs(5112));
    outputs(754) <= (layer0_outputs(1789)) and not (layer0_outputs(3432));
    outputs(755) <= (layer0_outputs(1033)) and not (layer0_outputs(1603));
    outputs(756) <= not((layer0_outputs(493)) xor (layer0_outputs(1733)));
    outputs(757) <= (layer0_outputs(4163)) and not (layer0_outputs(293));
    outputs(758) <= layer0_outputs(2790);
    outputs(759) <= (layer0_outputs(1411)) and (layer0_outputs(4682));
    outputs(760) <= (layer0_outputs(3878)) and not (layer0_outputs(1919));
    outputs(761) <= layer0_outputs(3114);
    outputs(762) <= layer0_outputs(690);
    outputs(763) <= (layer0_outputs(666)) and (layer0_outputs(1926));
    outputs(764) <= not(layer0_outputs(2058));
    outputs(765) <= (layer0_outputs(3302)) and not (layer0_outputs(3031));
    outputs(766) <= not((layer0_outputs(356)) or (layer0_outputs(2883)));
    outputs(767) <= (layer0_outputs(759)) and not (layer0_outputs(198));
    outputs(768) <= (layer0_outputs(379)) and (layer0_outputs(3642));
    outputs(769) <= (layer0_outputs(2393)) and (layer0_outputs(2798));
    outputs(770) <= (layer0_outputs(5090)) and not (layer0_outputs(1895));
    outputs(771) <= (layer0_outputs(1422)) and (layer0_outputs(1164));
    outputs(772) <= not((layer0_outputs(1780)) or (layer0_outputs(2648)));
    outputs(773) <= (layer0_outputs(3381)) and (layer0_outputs(1527));
    outputs(774) <= (layer0_outputs(2074)) and not (layer0_outputs(4542));
    outputs(775) <= (layer0_outputs(3736)) xor (layer0_outputs(2827));
    outputs(776) <= (layer0_outputs(435)) and (layer0_outputs(3406));
    outputs(777) <= layer0_outputs(1286);
    outputs(778) <= layer0_outputs(1596);
    outputs(779) <= not((layer0_outputs(2069)) or (layer0_outputs(4198)));
    outputs(780) <= '0';
    outputs(781) <= (layer0_outputs(4872)) and not (layer0_outputs(1530));
    outputs(782) <= layer0_outputs(2831);
    outputs(783) <= layer0_outputs(4660);
    outputs(784) <= (layer0_outputs(1081)) and (layer0_outputs(398));
    outputs(785) <= not((layer0_outputs(4837)) or (layer0_outputs(1221)));
    outputs(786) <= (layer0_outputs(1554)) and not (layer0_outputs(4255));
    outputs(787) <= (layer0_outputs(2468)) and (layer0_outputs(3845));
    outputs(788) <= not((layer0_outputs(3968)) or (layer0_outputs(3904)));
    outputs(789) <= (layer0_outputs(578)) and not (layer0_outputs(3547));
    outputs(790) <= not((layer0_outputs(3820)) and (layer0_outputs(4488)));
    outputs(791) <= not((layer0_outputs(521)) or (layer0_outputs(4264)));
    outputs(792) <= (layer0_outputs(1055)) and not (layer0_outputs(1775));
    outputs(793) <= (layer0_outputs(4364)) and not (layer0_outputs(5072));
    outputs(794) <= (layer0_outputs(3039)) and not (layer0_outputs(3488));
    outputs(795) <= layer0_outputs(1452);
    outputs(796) <= (layer0_outputs(1039)) and not (layer0_outputs(3800));
    outputs(797) <= not((layer0_outputs(1032)) or (layer0_outputs(1479)));
    outputs(798) <= layer0_outputs(1061);
    outputs(799) <= layer0_outputs(5085);
    outputs(800) <= layer0_outputs(1016);
    outputs(801) <= layer0_outputs(2885);
    outputs(802) <= not(layer0_outputs(3877));
    outputs(803) <= (layer0_outputs(2536)) and not (layer0_outputs(2718));
    outputs(804) <= not((layer0_outputs(1270)) or (layer0_outputs(1316)));
    outputs(805) <= (layer0_outputs(1436)) and not (layer0_outputs(2113));
    outputs(806) <= layer0_outputs(1251);
    outputs(807) <= not(layer0_outputs(830));
    outputs(808) <= not((layer0_outputs(1559)) or (layer0_outputs(653)));
    outputs(809) <= (layer0_outputs(3162)) and not (layer0_outputs(714));
    outputs(810) <= not((layer0_outputs(3942)) xor (layer0_outputs(4183)));
    outputs(811) <= not((layer0_outputs(4375)) or (layer0_outputs(2026)));
    outputs(812) <= not((layer0_outputs(1093)) or (layer0_outputs(1336)));
    outputs(813) <= (layer0_outputs(29)) and not (layer0_outputs(3997));
    outputs(814) <= (layer0_outputs(4773)) and not (layer0_outputs(3361));
    outputs(815) <= (layer0_outputs(2019)) and not (layer0_outputs(3294));
    outputs(816) <= not((layer0_outputs(5022)) or (layer0_outputs(2685)));
    outputs(817) <= (layer0_outputs(3300)) and (layer0_outputs(3052));
    outputs(818) <= not((layer0_outputs(1736)) or (layer0_outputs(4595)));
    outputs(819) <= (layer0_outputs(687)) and not (layer0_outputs(1293));
    outputs(820) <= (layer0_outputs(1417)) and not (layer0_outputs(499));
    outputs(821) <= not((layer0_outputs(2655)) xor (layer0_outputs(3013)));
    outputs(822) <= not((layer0_outputs(3139)) or (layer0_outputs(1306)));
    outputs(823) <= (layer0_outputs(2985)) and (layer0_outputs(3359));
    outputs(824) <= (layer0_outputs(2872)) xor (layer0_outputs(3652));
    outputs(825) <= (layer0_outputs(3701)) and not (layer0_outputs(2633));
    outputs(826) <= not(layer0_outputs(2738));
    outputs(827) <= not((layer0_outputs(4988)) or (layer0_outputs(2947)));
    outputs(828) <= (layer0_outputs(949)) and (layer0_outputs(2712));
    outputs(829) <= not(layer0_outputs(4432));
    outputs(830) <= (layer0_outputs(3797)) and not (layer0_outputs(2874));
    outputs(831) <= layer0_outputs(2923);
    outputs(832) <= layer0_outputs(4242);
    outputs(833) <= not((layer0_outputs(4318)) xor (layer0_outputs(3163)));
    outputs(834) <= (layer0_outputs(4142)) and not (layer0_outputs(4285));
    outputs(835) <= not(layer0_outputs(245));
    outputs(836) <= not((layer0_outputs(943)) or (layer0_outputs(4600)));
    outputs(837) <= (layer0_outputs(3620)) and (layer0_outputs(185));
    outputs(838) <= (layer0_outputs(2700)) and (layer0_outputs(2143));
    outputs(839) <= not(layer0_outputs(3392));
    outputs(840) <= not((layer0_outputs(2284)) xor (layer0_outputs(745)));
    outputs(841) <= not((layer0_outputs(4679)) or (layer0_outputs(1129)));
    outputs(842) <= (layer0_outputs(1688)) and not (layer0_outputs(5054));
    outputs(843) <= (layer0_outputs(854)) and (layer0_outputs(1482));
    outputs(844) <= (layer0_outputs(2624)) and not (layer0_outputs(3801));
    outputs(845) <= (layer0_outputs(1628)) and not (layer0_outputs(2706));
    outputs(846) <= not(layer0_outputs(1496));
    outputs(847) <= (layer0_outputs(4106)) and (layer0_outputs(2847));
    outputs(848) <= (layer0_outputs(1294)) and not (layer0_outputs(4725));
    outputs(849) <= layer0_outputs(2412);
    outputs(850) <= not((layer0_outputs(3216)) or (layer0_outputs(4834)));
    outputs(851) <= (layer0_outputs(1986)) xor (layer0_outputs(258));
    outputs(852) <= layer0_outputs(3861);
    outputs(853) <= not(layer0_outputs(4903));
    outputs(854) <= not(layer0_outputs(154)) or (layer0_outputs(3436));
    outputs(855) <= not(layer0_outputs(52));
    outputs(856) <= not((layer0_outputs(3384)) or (layer0_outputs(2154)));
    outputs(857) <= layer0_outputs(3062);
    outputs(858) <= (layer0_outputs(655)) xor (layer0_outputs(4216));
    outputs(859) <= layer0_outputs(2017);
    outputs(860) <= (layer0_outputs(2991)) and not (layer0_outputs(4529));
    outputs(861) <= not((layer0_outputs(327)) or (layer0_outputs(3476)));
    outputs(862) <= (layer0_outputs(194)) and (layer0_outputs(4889));
    outputs(863) <= not(layer0_outputs(4490));
    outputs(864) <= (layer0_outputs(2764)) and not (layer0_outputs(1269));
    outputs(865) <= (layer0_outputs(769)) and not (layer0_outputs(2036));
    outputs(866) <= not((layer0_outputs(2482)) or (layer0_outputs(2015)));
    outputs(867) <= not((layer0_outputs(2171)) or (layer0_outputs(1293)));
    outputs(868) <= layer0_outputs(3655);
    outputs(869) <= not((layer0_outputs(3055)) xor (layer0_outputs(1665)));
    outputs(870) <= not((layer0_outputs(4746)) or (layer0_outputs(950)));
    outputs(871) <= not((layer0_outputs(4595)) or (layer0_outputs(3108)));
    outputs(872) <= (layer0_outputs(3077)) and not (layer0_outputs(2569));
    outputs(873) <= (layer0_outputs(3314)) and not (layer0_outputs(2648));
    outputs(874) <= (layer0_outputs(3473)) and not (layer0_outputs(1776));
    outputs(875) <= (layer0_outputs(3791)) and not (layer0_outputs(777));
    outputs(876) <= not((layer0_outputs(1400)) or (layer0_outputs(2068)));
    outputs(877) <= (layer0_outputs(5058)) and (layer0_outputs(987));
    outputs(878) <= layer0_outputs(2390);
    outputs(879) <= not(layer0_outputs(794));
    outputs(880) <= not((layer0_outputs(1551)) or (layer0_outputs(2363)));
    outputs(881) <= (layer0_outputs(3644)) and not (layer0_outputs(1755));
    outputs(882) <= (layer0_outputs(213)) and (layer0_outputs(4960));
    outputs(883) <= not((layer0_outputs(4635)) or (layer0_outputs(4372)));
    outputs(884) <= (layer0_outputs(212)) and (layer0_outputs(1797));
    outputs(885) <= (layer0_outputs(2812)) and (layer0_outputs(1557));
    outputs(886) <= not((layer0_outputs(2528)) or (layer0_outputs(319)));
    outputs(887) <= (layer0_outputs(111)) and (layer0_outputs(4110));
    outputs(888) <= layer0_outputs(178);
    outputs(889) <= (layer0_outputs(1590)) and not (layer0_outputs(4681));
    outputs(890) <= (layer0_outputs(4343)) and not (layer0_outputs(4198));
    outputs(891) <= not((layer0_outputs(17)) or (layer0_outputs(3972)));
    outputs(892) <= layer0_outputs(3769);
    outputs(893) <= layer0_outputs(2442);
    outputs(894) <= (layer0_outputs(4182)) and (layer0_outputs(1053));
    outputs(895) <= layer0_outputs(4191);
    outputs(896) <= not(layer0_outputs(2607)) or (layer0_outputs(3158));
    outputs(897) <= (layer0_outputs(4050)) and not (layer0_outputs(2368));
    outputs(898) <= not(layer0_outputs(4240));
    outputs(899) <= (layer0_outputs(792)) and (layer0_outputs(3993));
    outputs(900) <= not((layer0_outputs(2191)) or (layer0_outputs(4185)));
    outputs(901) <= layer0_outputs(3636);
    outputs(902) <= (layer0_outputs(5006)) and not (layer0_outputs(3816));
    outputs(903) <= layer0_outputs(3989);
    outputs(904) <= (layer0_outputs(1965)) and not (layer0_outputs(2274));
    outputs(905) <= not((layer0_outputs(4957)) or (layer0_outputs(1841)));
    outputs(906) <= (layer0_outputs(2088)) and not (layer0_outputs(1042));
    outputs(907) <= (layer0_outputs(372)) and not (layer0_outputs(1771));
    outputs(908) <= (layer0_outputs(1338)) and (layer0_outputs(3012));
    outputs(909) <= not(layer0_outputs(2557));
    outputs(910) <= not(layer0_outputs(805));
    outputs(911) <= not(layer0_outputs(3767));
    outputs(912) <= not((layer0_outputs(524)) or (layer0_outputs(2214)));
    outputs(913) <= not(layer0_outputs(4133)) or (layer0_outputs(5037));
    outputs(914) <= '0';
    outputs(915) <= (layer0_outputs(2284)) and not (layer0_outputs(3071));
    outputs(916) <= not((layer0_outputs(4355)) or (layer0_outputs(1105)));
    outputs(917) <= not((layer0_outputs(329)) xor (layer0_outputs(1664)));
    outputs(918) <= layer0_outputs(4416);
    outputs(919) <= (layer0_outputs(2495)) and not (layer0_outputs(2403));
    outputs(920) <= not(layer0_outputs(762));
    outputs(921) <= (layer0_outputs(4774)) and not (layer0_outputs(1925));
    outputs(922) <= not(layer0_outputs(2757));
    outputs(923) <= not((layer0_outputs(3539)) or (layer0_outputs(3842)));
    outputs(924) <= layer0_outputs(1267);
    outputs(925) <= (layer0_outputs(2518)) xor (layer0_outputs(3834));
    outputs(926) <= not((layer0_outputs(4091)) or (layer0_outputs(2148)));
    outputs(927) <= not(layer0_outputs(1213));
    outputs(928) <= layer0_outputs(2057);
    outputs(929) <= (layer0_outputs(4381)) and (layer0_outputs(1752));
    outputs(930) <= layer0_outputs(2884);
    outputs(931) <= (layer0_outputs(3207)) and (layer0_outputs(4908));
    outputs(932) <= (layer0_outputs(3448)) and (layer0_outputs(1765));
    outputs(933) <= (layer0_outputs(3034)) and not (layer0_outputs(4944));
    outputs(934) <= not((layer0_outputs(668)) xor (layer0_outputs(570)));
    outputs(935) <= (layer0_outputs(4500)) and not (layer0_outputs(1648));
    outputs(936) <= not((layer0_outputs(2026)) or (layer0_outputs(1948)));
    outputs(937) <= not(layer0_outputs(2171)) or (layer0_outputs(4126));
    outputs(938) <= layer0_outputs(1796);
    outputs(939) <= layer0_outputs(2237);
    outputs(940) <= layer0_outputs(2054);
    outputs(941) <= layer0_outputs(983);
    outputs(942) <= (layer0_outputs(2051)) and (layer0_outputs(743));
    outputs(943) <= (layer0_outputs(3243)) and not (layer0_outputs(570));
    outputs(944) <= not((layer0_outputs(4645)) or (layer0_outputs(956)));
    outputs(945) <= layer0_outputs(4302);
    outputs(946) <= (layer0_outputs(3241)) and (layer0_outputs(4268));
    outputs(947) <= not((layer0_outputs(434)) xor (layer0_outputs(390)));
    outputs(948) <= (layer0_outputs(2239)) and not (layer0_outputs(4760));
    outputs(949) <= not(layer0_outputs(1079));
    outputs(950) <= (layer0_outputs(299)) and not (layer0_outputs(2154));
    outputs(951) <= (layer0_outputs(4494)) and not (layer0_outputs(1625));
    outputs(952) <= not(layer0_outputs(4851)) or (layer0_outputs(1323));
    outputs(953) <= not(layer0_outputs(2992));
    outputs(954) <= layer0_outputs(4229);
    outputs(955) <= not((layer0_outputs(1737)) xor (layer0_outputs(1421)));
    outputs(956) <= (layer0_outputs(2271)) and not (layer0_outputs(2524));
    outputs(957) <= (layer0_outputs(2505)) and (layer0_outputs(4742));
    outputs(958) <= (layer0_outputs(2493)) xor (layer0_outputs(2526));
    outputs(959) <= (layer0_outputs(2713)) and not (layer0_outputs(5115));
    outputs(960) <= (layer0_outputs(2226)) and (layer0_outputs(4428));
    outputs(961) <= (layer0_outputs(985)) xor (layer0_outputs(164));
    outputs(962) <= not(layer0_outputs(145));
    outputs(963) <= (layer0_outputs(3701)) and not (layer0_outputs(3238));
    outputs(964) <= (layer0_outputs(608)) and not (layer0_outputs(1690));
    outputs(965) <= (layer0_outputs(2598)) and (layer0_outputs(965));
    outputs(966) <= not((layer0_outputs(3240)) or (layer0_outputs(1308)));
    outputs(967) <= not(layer0_outputs(4746));
    outputs(968) <= not((layer0_outputs(2996)) or (layer0_outputs(2588)));
    outputs(969) <= (layer0_outputs(1211)) and not (layer0_outputs(3345));
    outputs(970) <= not(layer0_outputs(3174));
    outputs(971) <= (layer0_outputs(2856)) and (layer0_outputs(3977));
    outputs(972) <= (layer0_outputs(507)) and (layer0_outputs(3859));
    outputs(973) <= not((layer0_outputs(2958)) xor (layer0_outputs(907)));
    outputs(974) <= layer0_outputs(2047);
    outputs(975) <= not(layer0_outputs(3654));
    outputs(976) <= layer0_outputs(1946);
    outputs(977) <= not((layer0_outputs(4594)) xor (layer0_outputs(4703)));
    outputs(978) <= not(layer0_outputs(4498));
    outputs(979) <= (layer0_outputs(2426)) and not (layer0_outputs(3632));
    outputs(980) <= (layer0_outputs(1950)) and not (layer0_outputs(4292));
    outputs(981) <= not(layer0_outputs(2375));
    outputs(982) <= (layer0_outputs(3810)) and (layer0_outputs(2027));
    outputs(983) <= not((layer0_outputs(3295)) or (layer0_outputs(3715)));
    outputs(984) <= not((layer0_outputs(2090)) xor (layer0_outputs(2080)));
    outputs(985) <= (layer0_outputs(3002)) and (layer0_outputs(277));
    outputs(986) <= (layer0_outputs(698)) and not (layer0_outputs(411));
    outputs(987) <= layer0_outputs(2372);
    outputs(988) <= not((layer0_outputs(2322)) or (layer0_outputs(35)));
    outputs(989) <= (layer0_outputs(1585)) and not (layer0_outputs(3333));
    outputs(990) <= not(layer0_outputs(552));
    outputs(991) <= (layer0_outputs(1210)) and not (layer0_outputs(4196));
    outputs(992) <= not((layer0_outputs(664)) or (layer0_outputs(2053)));
    outputs(993) <= (layer0_outputs(44)) and not (layer0_outputs(4798));
    outputs(994) <= not((layer0_outputs(266)) or (layer0_outputs(4662)));
    outputs(995) <= not(layer0_outputs(2134));
    outputs(996) <= not(layer0_outputs(1806));
    outputs(997) <= (layer0_outputs(1215)) and not (layer0_outputs(3852));
    outputs(998) <= not(layer0_outputs(2481));
    outputs(999) <= (layer0_outputs(2436)) and (layer0_outputs(3359));
    outputs(1000) <= (layer0_outputs(1918)) xor (layer0_outputs(1385));
    outputs(1001) <= (layer0_outputs(2314)) and (layer0_outputs(4880));
    outputs(1002) <= layer0_outputs(358);
    outputs(1003) <= (layer0_outputs(1352)) and (layer0_outputs(862));
    outputs(1004) <= not(layer0_outputs(151));
    outputs(1005) <= (layer0_outputs(406)) and not (layer0_outputs(5011));
    outputs(1006) <= layer0_outputs(4176);
    outputs(1007) <= (layer0_outputs(2616)) and not (layer0_outputs(4308));
    outputs(1008) <= (layer0_outputs(1240)) and not (layer0_outputs(1847));
    outputs(1009) <= (layer0_outputs(5040)) xor (layer0_outputs(2201));
    outputs(1010) <= not((layer0_outputs(4870)) xor (layer0_outputs(1657)));
    outputs(1011) <= not(layer0_outputs(1031));
    outputs(1012) <= not((layer0_outputs(2421)) or (layer0_outputs(585)));
    outputs(1013) <= '0';
    outputs(1014) <= (layer0_outputs(4150)) and (layer0_outputs(4891));
    outputs(1015) <= (layer0_outputs(2161)) and not (layer0_outputs(63));
    outputs(1016) <= layer0_outputs(4116);
    outputs(1017) <= layer0_outputs(1272);
    outputs(1018) <= (layer0_outputs(1202)) or (layer0_outputs(275));
    outputs(1019) <= (layer0_outputs(4619)) and (layer0_outputs(539));
    outputs(1020) <= not(layer0_outputs(3960));
    outputs(1021) <= not((layer0_outputs(1369)) or (layer0_outputs(190)));
    outputs(1022) <= (layer0_outputs(3053)) and not (layer0_outputs(1050));
    outputs(1023) <= not(layer0_outputs(2247));
    outputs(1024) <= not(layer0_outputs(2522)) or (layer0_outputs(1783));
    outputs(1025) <= not((layer0_outputs(1853)) xor (layer0_outputs(4259)));
    outputs(1026) <= not(layer0_outputs(258));
    outputs(1027) <= not((layer0_outputs(2120)) or (layer0_outputs(3832)));
    outputs(1028) <= layer0_outputs(1175);
    outputs(1029) <= not(layer0_outputs(4363)) or (layer0_outputs(3065));
    outputs(1030) <= not(layer0_outputs(3433));
    outputs(1031) <= not(layer0_outputs(324));
    outputs(1032) <= not(layer0_outputs(510));
    outputs(1033) <= layer0_outputs(1118);
    outputs(1034) <= layer0_outputs(4115);
    outputs(1035) <= not(layer0_outputs(1117)) or (layer0_outputs(4888));
    outputs(1036) <= not(layer0_outputs(1171)) or (layer0_outputs(2654));
    outputs(1037) <= not(layer0_outputs(4250)) or (layer0_outputs(1486));
    outputs(1038) <= not(layer0_outputs(2203)) or (layer0_outputs(2245));
    outputs(1039) <= (layer0_outputs(3223)) or (layer0_outputs(345));
    outputs(1040) <= not((layer0_outputs(2680)) and (layer0_outputs(878)));
    outputs(1041) <= (layer0_outputs(2568)) xor (layer0_outputs(2491));
    outputs(1042) <= (layer0_outputs(2740)) and not (layer0_outputs(4959));
    outputs(1043) <= not((layer0_outputs(54)) and (layer0_outputs(1030)));
    outputs(1044) <= not((layer0_outputs(1622)) xor (layer0_outputs(2832)));
    outputs(1045) <= not(layer0_outputs(4637));
    outputs(1046) <= not(layer0_outputs(3748));
    outputs(1047) <= layer0_outputs(3485);
    outputs(1048) <= not((layer0_outputs(3168)) xor (layer0_outputs(989)));
    outputs(1049) <= layer0_outputs(2356);
    outputs(1050) <= (layer0_outputs(1571)) xor (layer0_outputs(1179));
    outputs(1051) <= (layer0_outputs(3568)) xor (layer0_outputs(4));
    outputs(1052) <= not((layer0_outputs(2542)) xor (layer0_outputs(2099)));
    outputs(1053) <= not(layer0_outputs(1000));
    outputs(1054) <= not(layer0_outputs(3150));
    outputs(1055) <= not((layer0_outputs(3177)) xor (layer0_outputs(1627)));
    outputs(1056) <= (layer0_outputs(777)) and not (layer0_outputs(564));
    outputs(1057) <= layer0_outputs(2228);
    outputs(1058) <= (layer0_outputs(3027)) or (layer0_outputs(823));
    outputs(1059) <= not(layer0_outputs(1445));
    outputs(1060) <= (layer0_outputs(4314)) xor (layer0_outputs(2690));
    outputs(1061) <= layer0_outputs(1373);
    outputs(1062) <= layer0_outputs(4222);
    outputs(1063) <= not(layer0_outputs(2681)) or (layer0_outputs(3784));
    outputs(1064) <= layer0_outputs(2698);
    outputs(1065) <= layer0_outputs(5099);
    outputs(1066) <= (layer0_outputs(3949)) and not (layer0_outputs(2541));
    outputs(1067) <= layer0_outputs(4451);
    outputs(1068) <= (layer0_outputs(1824)) or (layer0_outputs(4514));
    outputs(1069) <= not(layer0_outputs(2094));
    outputs(1070) <= (layer0_outputs(593)) xor (layer0_outputs(2957));
    outputs(1071) <= not((layer0_outputs(4632)) or (layer0_outputs(1178)));
    outputs(1072) <= (layer0_outputs(2880)) and (layer0_outputs(3605));
    outputs(1073) <= not(layer0_outputs(730)) or (layer0_outputs(2625));
    outputs(1074) <= not(layer0_outputs(4408));
    outputs(1075) <= layer0_outputs(2758);
    outputs(1076) <= not(layer0_outputs(213));
    outputs(1077) <= not(layer0_outputs(2211));
    outputs(1078) <= not(layer0_outputs(3182));
    outputs(1079) <= not(layer0_outputs(1843));
    outputs(1080) <= not((layer0_outputs(1248)) xor (layer0_outputs(4303)));
    outputs(1081) <= (layer0_outputs(5059)) and not (layer0_outputs(133));
    outputs(1082) <= not(layer0_outputs(1978)) or (layer0_outputs(636));
    outputs(1083) <= layer0_outputs(187);
    outputs(1084) <= (layer0_outputs(1661)) and not (layer0_outputs(3729));
    outputs(1085) <= not(layer0_outputs(30));
    outputs(1086) <= layer0_outputs(4993);
    outputs(1087) <= not(layer0_outputs(3843));
    outputs(1088) <= not((layer0_outputs(2919)) xor (layer0_outputs(4702)));
    outputs(1089) <= not(layer0_outputs(3609));
    outputs(1090) <= layer0_outputs(1924);
    outputs(1091) <= not(layer0_outputs(4653)) or (layer0_outputs(409));
    outputs(1092) <= layer0_outputs(3649);
    outputs(1093) <= not(layer0_outputs(3144));
    outputs(1094) <= (layer0_outputs(5109)) and not (layer0_outputs(1003));
    outputs(1095) <= not(layer0_outputs(3095)) or (layer0_outputs(117));
    outputs(1096) <= layer0_outputs(935);
    outputs(1097) <= not(layer0_outputs(4307));
    outputs(1098) <= (layer0_outputs(574)) xor (layer0_outputs(505));
    outputs(1099) <= not((layer0_outputs(359)) xor (layer0_outputs(3978)));
    outputs(1100) <= not(layer0_outputs(4131)) or (layer0_outputs(4229));
    outputs(1101) <= not(layer0_outputs(3344));
    outputs(1102) <= not((layer0_outputs(1168)) or (layer0_outputs(2165)));
    outputs(1103) <= (layer0_outputs(3993)) or (layer0_outputs(4539));
    outputs(1104) <= layer0_outputs(1148);
    outputs(1105) <= not((layer0_outputs(1937)) and (layer0_outputs(2938)));
    outputs(1106) <= layer0_outputs(1348);
    outputs(1107) <= layer0_outputs(1545);
    outputs(1108) <= not(layer0_outputs(4669));
    outputs(1109) <= (layer0_outputs(507)) xor (layer0_outputs(4301));
    outputs(1110) <= not(layer0_outputs(2861)) or (layer0_outputs(437));
    outputs(1111) <= not(layer0_outputs(3197)) or (layer0_outputs(975));
    outputs(1112) <= layer0_outputs(3559);
    outputs(1113) <= not((layer0_outputs(2112)) and (layer0_outputs(2144)));
    outputs(1114) <= (layer0_outputs(272)) and not (layer0_outputs(1662));
    outputs(1115) <= not(layer0_outputs(4971));
    outputs(1116) <= not(layer0_outputs(4550));
    outputs(1117) <= not(layer0_outputs(1641));
    outputs(1118) <= not(layer0_outputs(654));
    outputs(1119) <= not(layer0_outputs(4218));
    outputs(1120) <= (layer0_outputs(2574)) and not (layer0_outputs(742));
    outputs(1121) <= not(layer0_outputs(3350));
    outputs(1122) <= not(layer0_outputs(840));
    outputs(1123) <= (layer0_outputs(2232)) or (layer0_outputs(5092));
    outputs(1124) <= not(layer0_outputs(931));
    outputs(1125) <= not((layer0_outputs(381)) or (layer0_outputs(2246)));
    outputs(1126) <= not(layer0_outputs(2985)) or (layer0_outputs(1761));
    outputs(1127) <= layer0_outputs(4592);
    outputs(1128) <= not(layer0_outputs(1835)) or (layer0_outputs(3110));
    outputs(1129) <= layer0_outputs(1636);
    outputs(1130) <= (layer0_outputs(696)) or (layer0_outputs(3424));
    outputs(1131) <= not(layer0_outputs(3679));
    outputs(1132) <= not(layer0_outputs(2802)) or (layer0_outputs(4598));
    outputs(1133) <= (layer0_outputs(2544)) and not (layer0_outputs(200));
    outputs(1134) <= not((layer0_outputs(1168)) and (layer0_outputs(3562)));
    outputs(1135) <= not((layer0_outputs(4885)) xor (layer0_outputs(1509)));
    outputs(1136) <= layer0_outputs(5067);
    outputs(1137) <= layer0_outputs(3802);
    outputs(1138) <= (layer0_outputs(4569)) and not (layer0_outputs(4925));
    outputs(1139) <= not((layer0_outputs(4699)) xor (layer0_outputs(1164)));
    outputs(1140) <= layer0_outputs(4180);
    outputs(1141) <= not((layer0_outputs(1170)) xor (layer0_outputs(1219)));
    outputs(1142) <= not(layer0_outputs(1781)) or (layer0_outputs(4236));
    outputs(1143) <= not((layer0_outputs(1910)) xor (layer0_outputs(3074)));
    outputs(1144) <= not(layer0_outputs(1098));
    outputs(1145) <= (layer0_outputs(3577)) and not (layer0_outputs(2541));
    outputs(1146) <= not(layer0_outputs(19)) or (layer0_outputs(4807));
    outputs(1147) <= (layer0_outputs(4734)) and (layer0_outputs(4581));
    outputs(1148) <= not(layer0_outputs(2619)) or (layer0_outputs(1628));
    outputs(1149) <= not(layer0_outputs(1892));
    outputs(1150) <= not(layer0_outputs(1687));
    outputs(1151) <= not(layer0_outputs(94)) or (layer0_outputs(275));
    outputs(1152) <= (layer0_outputs(3153)) or (layer0_outputs(2385));
    outputs(1153) <= layer0_outputs(1885);
    outputs(1154) <= not(layer0_outputs(1208));
    outputs(1155) <= layer0_outputs(2427);
    outputs(1156) <= layer0_outputs(5037);
    outputs(1157) <= layer0_outputs(4549);
    outputs(1158) <= (layer0_outputs(1714)) xor (layer0_outputs(1233));
    outputs(1159) <= (layer0_outputs(4999)) or (layer0_outputs(919));
    outputs(1160) <= not((layer0_outputs(1484)) or (layer0_outputs(2840)));
    outputs(1161) <= not(layer0_outputs(4415));
    outputs(1162) <= (layer0_outputs(3204)) xor (layer0_outputs(4597));
    outputs(1163) <= not(layer0_outputs(204)) or (layer0_outputs(4246));
    outputs(1164) <= not((layer0_outputs(4003)) and (layer0_outputs(1742)));
    outputs(1165) <= layer0_outputs(2944);
    outputs(1166) <= not((layer0_outputs(842)) xor (layer0_outputs(847)));
    outputs(1167) <= not(layer0_outputs(2989));
    outputs(1168) <= not(layer0_outputs(984)) or (layer0_outputs(1452));
    outputs(1169) <= layer0_outputs(3046);
    outputs(1170) <= not(layer0_outputs(230)) or (layer0_outputs(4457));
    outputs(1171) <= not(layer0_outputs(1284));
    outputs(1172) <= (layer0_outputs(4568)) and not (layer0_outputs(3609));
    outputs(1173) <= not(layer0_outputs(4219));
    outputs(1174) <= (layer0_outputs(788)) or (layer0_outputs(5077));
    outputs(1175) <= not(layer0_outputs(5117)) or (layer0_outputs(1103));
    outputs(1176) <= (layer0_outputs(3671)) xor (layer0_outputs(3103));
    outputs(1177) <= not(layer0_outputs(2828));
    outputs(1178) <= not(layer0_outputs(2186));
    outputs(1179) <= (layer0_outputs(1237)) and not (layer0_outputs(2183));
    outputs(1180) <= (layer0_outputs(1783)) or (layer0_outputs(4991));
    outputs(1181) <= (layer0_outputs(2819)) xor (layer0_outputs(3481));
    outputs(1182) <= (layer0_outputs(3680)) and (layer0_outputs(922));
    outputs(1183) <= (layer0_outputs(3421)) xor (layer0_outputs(3720));
    outputs(1184) <= (layer0_outputs(4701)) xor (layer0_outputs(3101));
    outputs(1185) <= (layer0_outputs(4641)) or (layer0_outputs(989));
    outputs(1186) <= layer0_outputs(4498);
    outputs(1187) <= layer0_outputs(4679);
    outputs(1188) <= not(layer0_outputs(3958)) or (layer0_outputs(4359));
    outputs(1189) <= not(layer0_outputs(3341));
    outputs(1190) <= not(layer0_outputs(2627));
    outputs(1191) <= layer0_outputs(4873);
    outputs(1192) <= (layer0_outputs(4238)) or (layer0_outputs(2525));
    outputs(1193) <= not((layer0_outputs(3537)) or (layer0_outputs(3068)));
    outputs(1194) <= layer0_outputs(1078);
    outputs(1195) <= layer0_outputs(250);
    outputs(1196) <= (layer0_outputs(4400)) and not (layer0_outputs(4323));
    outputs(1197) <= not(layer0_outputs(414)) or (layer0_outputs(4292));
    outputs(1198) <= layer0_outputs(958);
    outputs(1199) <= not(layer0_outputs(4420));
    outputs(1200) <= layer0_outputs(4715);
    outputs(1201) <= not(layer0_outputs(698));
    outputs(1202) <= not((layer0_outputs(2842)) xor (layer0_outputs(4946)));
    outputs(1203) <= (layer0_outputs(2313)) xor (layer0_outputs(2035));
    outputs(1204) <= not(layer0_outputs(4276));
    outputs(1205) <= not(layer0_outputs(3669));
    outputs(1206) <= not((layer0_outputs(4574)) and (layer0_outputs(4093)));
    outputs(1207) <= layer0_outputs(3286);
    outputs(1208) <= layer0_outputs(571);
    outputs(1209) <= not((layer0_outputs(255)) and (layer0_outputs(1382)));
    outputs(1210) <= not(layer0_outputs(2762)) or (layer0_outputs(2169));
    outputs(1211) <= not((layer0_outputs(978)) xor (layer0_outputs(1936)));
    outputs(1212) <= layer0_outputs(848);
    outputs(1213) <= not((layer0_outputs(4262)) xor (layer0_outputs(1817)));
    outputs(1214) <= (layer0_outputs(1768)) and (layer0_outputs(1308));
    outputs(1215) <= not(layer0_outputs(1283));
    outputs(1216) <= not(layer0_outputs(980));
    outputs(1217) <= (layer0_outputs(5102)) or (layer0_outputs(278));
    outputs(1218) <= not(layer0_outputs(3571)) or (layer0_outputs(4158));
    outputs(1219) <= not(layer0_outputs(3932)) or (layer0_outputs(2598));
    outputs(1220) <= (layer0_outputs(73)) xor (layer0_outputs(515));
    outputs(1221) <= not(layer0_outputs(3487)) or (layer0_outputs(5002));
    outputs(1222) <= layer0_outputs(2423);
    outputs(1223) <= (layer0_outputs(2618)) and not (layer0_outputs(2360));
    outputs(1224) <= not(layer0_outputs(4704));
    outputs(1225) <= (layer0_outputs(280)) and (layer0_outputs(4032));
    outputs(1226) <= (layer0_outputs(1848)) or (layer0_outputs(1402));
    outputs(1227) <= not(layer0_outputs(1755)) or (layer0_outputs(3691));
    outputs(1228) <= not((layer0_outputs(878)) and (layer0_outputs(2319)));
    outputs(1229) <= layer0_outputs(1430);
    outputs(1230) <= not(layer0_outputs(2207));
    outputs(1231) <= (layer0_outputs(902)) or (layer0_outputs(5110));
    outputs(1232) <= (layer0_outputs(2189)) and (layer0_outputs(2903));
    outputs(1233) <= not(layer0_outputs(3734)) or (layer0_outputs(3596));
    outputs(1234) <= layer0_outputs(3236);
    outputs(1235) <= layer0_outputs(4193);
    outputs(1236) <= not(layer0_outputs(3504));
    outputs(1237) <= (layer0_outputs(2455)) xor (layer0_outputs(4302));
    outputs(1238) <= layer0_outputs(1345);
    outputs(1239) <= not(layer0_outputs(3974)) or (layer0_outputs(3293));
    outputs(1240) <= layer0_outputs(1065);
    outputs(1241) <= not(layer0_outputs(1507));
    outputs(1242) <= not(layer0_outputs(1843));
    outputs(1243) <= not(layer0_outputs(1170)) or (layer0_outputs(2149));
    outputs(1244) <= not((layer0_outputs(3320)) xor (layer0_outputs(1595)));
    outputs(1245) <= (layer0_outputs(1672)) and not (layer0_outputs(4868));
    outputs(1246) <= (layer0_outputs(1353)) xor (layer0_outputs(502));
    outputs(1247) <= not(layer0_outputs(4049));
    outputs(1248) <= (layer0_outputs(4456)) or (layer0_outputs(3482));
    outputs(1249) <= layer0_outputs(42);
    outputs(1250) <= not((layer0_outputs(3753)) or (layer0_outputs(995)));
    outputs(1251) <= (layer0_outputs(1105)) or (layer0_outputs(3841));
    outputs(1252) <= layer0_outputs(3869);
    outputs(1253) <= not(layer0_outputs(3831)) or (layer0_outputs(602));
    outputs(1254) <= (layer0_outputs(3555)) and not (layer0_outputs(404));
    outputs(1255) <= (layer0_outputs(912)) xor (layer0_outputs(2756));
    outputs(1256) <= (layer0_outputs(1548)) xor (layer0_outputs(4167));
    outputs(1257) <= (layer0_outputs(4277)) or (layer0_outputs(694));
    outputs(1258) <= layer0_outputs(2845);
    outputs(1259) <= '1';
    outputs(1260) <= layer0_outputs(3316);
    outputs(1261) <= not(layer0_outputs(2200));
    outputs(1262) <= layer0_outputs(2679);
    outputs(1263) <= layer0_outputs(2004);
    outputs(1264) <= (layer0_outputs(2651)) xor (layer0_outputs(2926));
    outputs(1265) <= not((layer0_outputs(4979)) or (layer0_outputs(4300)));
    outputs(1266) <= layer0_outputs(1294);
    outputs(1267) <= not(layer0_outputs(3098));
    outputs(1268) <= not(layer0_outputs(2253));
    outputs(1269) <= layer0_outputs(3046);
    outputs(1270) <= not(layer0_outputs(1361));
    outputs(1271) <= layer0_outputs(2128);
    outputs(1272) <= not(layer0_outputs(736)) or (layer0_outputs(1858));
    outputs(1273) <= not(layer0_outputs(2226)) or (layer0_outputs(1173));
    outputs(1274) <= (layer0_outputs(3251)) or (layer0_outputs(1062));
    outputs(1275) <= not(layer0_outputs(488));
    outputs(1276) <= not(layer0_outputs(3914)) or (layer0_outputs(5065));
    outputs(1277) <= not(layer0_outputs(3342));
    outputs(1278) <= (layer0_outputs(3014)) xor (layer0_outputs(4305));
    outputs(1279) <= not((layer0_outputs(3665)) and (layer0_outputs(3382)));
    outputs(1280) <= not(layer0_outputs(3463)) or (layer0_outputs(1157));
    outputs(1281) <= (layer0_outputs(2608)) or (layer0_outputs(2514));
    outputs(1282) <= (layer0_outputs(3217)) or (layer0_outputs(3604));
    outputs(1283) <= not(layer0_outputs(3821)) or (layer0_outputs(705));
    outputs(1284) <= (layer0_outputs(1036)) and (layer0_outputs(3525));
    outputs(1285) <= layer0_outputs(2564);
    outputs(1286) <= layer0_outputs(696);
    outputs(1287) <= not((layer0_outputs(2001)) or (layer0_outputs(793)));
    outputs(1288) <= layer0_outputs(1930);
    outputs(1289) <= layer0_outputs(4084);
    outputs(1290) <= layer0_outputs(2758);
    outputs(1291) <= layer0_outputs(2327);
    outputs(1292) <= not(layer0_outputs(1622)) or (layer0_outputs(2064));
    outputs(1293) <= (layer0_outputs(4317)) xor (layer0_outputs(4382));
    outputs(1294) <= not(layer0_outputs(1241)) or (layer0_outputs(4856));
    outputs(1295) <= (layer0_outputs(1233)) and not (layer0_outputs(4209));
    outputs(1296) <= not((layer0_outputs(4358)) xor (layer0_outputs(2901)));
    outputs(1297) <= layer0_outputs(4443);
    outputs(1298) <= not(layer0_outputs(2005));
    outputs(1299) <= (layer0_outputs(2009)) or (layer0_outputs(3420));
    outputs(1300) <= layer0_outputs(1541);
    outputs(1301) <= layer0_outputs(3371);
    outputs(1302) <= (layer0_outputs(328)) xor (layer0_outputs(637));
    outputs(1303) <= (layer0_outputs(1365)) or (layer0_outputs(2309));
    outputs(1304) <= not(layer0_outputs(2490));
    outputs(1305) <= layer0_outputs(3580);
    outputs(1306) <= (layer0_outputs(4104)) xor (layer0_outputs(286));
    outputs(1307) <= (layer0_outputs(1379)) and (layer0_outputs(659));
    outputs(1308) <= (layer0_outputs(1281)) xor (layer0_outputs(629));
    outputs(1309) <= (layer0_outputs(4682)) and not (layer0_outputs(1305));
    outputs(1310) <= layer0_outputs(4296);
    outputs(1311) <= (layer0_outputs(3206)) or (layer0_outputs(4969));
    outputs(1312) <= (layer0_outputs(675)) and (layer0_outputs(4910));
    outputs(1313) <= layer0_outputs(4865);
    outputs(1314) <= not(layer0_outputs(3237));
    outputs(1315) <= layer0_outputs(2073);
    outputs(1316) <= layer0_outputs(1639);
    outputs(1317) <= not((layer0_outputs(2024)) and (layer0_outputs(2641)));
    outputs(1318) <= (layer0_outputs(4106)) and not (layer0_outputs(2508));
    outputs(1319) <= (layer0_outputs(4317)) xor (layer0_outputs(2778));
    outputs(1320) <= layer0_outputs(1002);
    outputs(1321) <= (layer0_outputs(3067)) xor (layer0_outputs(751));
    outputs(1322) <= layer0_outputs(3455);
    outputs(1323) <= not(layer0_outputs(1483));
    outputs(1324) <= layer0_outputs(4398);
    outputs(1325) <= layer0_outputs(4059);
    outputs(1326) <= layer0_outputs(3102);
    outputs(1327) <= (layer0_outputs(2614)) and not (layer0_outputs(2363));
    outputs(1328) <= (layer0_outputs(4825)) and not (layer0_outputs(1741));
    outputs(1329) <= layer0_outputs(3944);
    outputs(1330) <= not(layer0_outputs(1106));
    outputs(1331) <= not(layer0_outputs(436));
    outputs(1332) <= not(layer0_outputs(4823)) or (layer0_outputs(3424));
    outputs(1333) <= not(layer0_outputs(3695));
    outputs(1334) <= not(layer0_outputs(2785));
    outputs(1335) <= not(layer0_outputs(1850)) or (layer0_outputs(596));
    outputs(1336) <= (layer0_outputs(3348)) and (layer0_outputs(2051));
    outputs(1337) <= (layer0_outputs(3157)) and not (layer0_outputs(4986));
    outputs(1338) <= (layer0_outputs(4783)) and not (layer0_outputs(1488));
    outputs(1339) <= layer0_outputs(4269);
    outputs(1340) <= not(layer0_outputs(4414));
    outputs(1341) <= not(layer0_outputs(450)) or (layer0_outputs(2650));
    outputs(1342) <= (layer0_outputs(3348)) and not (layer0_outputs(2986));
    outputs(1343) <= (layer0_outputs(3434)) and (layer0_outputs(3908));
    outputs(1344) <= not(layer0_outputs(4268));
    outputs(1345) <= not(layer0_outputs(3030));
    outputs(1346) <= layer0_outputs(173);
    outputs(1347) <= (layer0_outputs(972)) xor (layer0_outputs(4207));
    outputs(1348) <= not(layer0_outputs(4329));
    outputs(1349) <= not(layer0_outputs(205));
    outputs(1350) <= not((layer0_outputs(3024)) xor (layer0_outputs(4426)));
    outputs(1351) <= not(layer0_outputs(2192));
    outputs(1352) <= not(layer0_outputs(1474));
    outputs(1353) <= layer0_outputs(157);
    outputs(1354) <= not((layer0_outputs(2185)) or (layer0_outputs(3120)));
    outputs(1355) <= (layer0_outputs(4475)) and not (layer0_outputs(1299));
    outputs(1356) <= not(layer0_outputs(1309)) or (layer0_outputs(4456));
    outputs(1357) <= not((layer0_outputs(757)) xor (layer0_outputs(36)));
    outputs(1358) <= not((layer0_outputs(4043)) or (layer0_outputs(417)));
    outputs(1359) <= not(layer0_outputs(284)) or (layer0_outputs(5053));
    outputs(1360) <= layer0_outputs(300);
    outputs(1361) <= layer0_outputs(4890);
    outputs(1362) <= layer0_outputs(2070);
    outputs(1363) <= not(layer0_outputs(2115));
    outputs(1364) <= not(layer0_outputs(2778));
    outputs(1365) <= layer0_outputs(326);
    outputs(1366) <= not(layer0_outputs(2866)) or (layer0_outputs(3744));
    outputs(1367) <= not(layer0_outputs(2939));
    outputs(1368) <= not(layer0_outputs(1177)) or (layer0_outputs(1897));
    outputs(1369) <= not((layer0_outputs(4775)) xor (layer0_outputs(3125)));
    outputs(1370) <= not((layer0_outputs(3484)) and (layer0_outputs(4714)));
    outputs(1371) <= (layer0_outputs(4693)) and not (layer0_outputs(1112));
    outputs(1372) <= not(layer0_outputs(4179));
    outputs(1373) <= not(layer0_outputs(2613));
    outputs(1374) <= not(layer0_outputs(1049)) or (layer0_outputs(2454));
    outputs(1375) <= not((layer0_outputs(346)) xor (layer0_outputs(2749)));
    outputs(1376) <= not((layer0_outputs(4336)) and (layer0_outputs(5025)));
    outputs(1377) <= not(layer0_outputs(4880));
    outputs(1378) <= not(layer0_outputs(2916));
    outputs(1379) <= not(layer0_outputs(5097));
    outputs(1380) <= not(layer0_outputs(4030));
    outputs(1381) <= layer0_outputs(2610);
    outputs(1382) <= not(layer0_outputs(3926));
    outputs(1383) <= (layer0_outputs(1629)) and (layer0_outputs(853));
    outputs(1384) <= (layer0_outputs(4489)) and not (layer0_outputs(2800));
    outputs(1385) <= (layer0_outputs(3008)) and not (layer0_outputs(3733));
    outputs(1386) <= layer0_outputs(2846);
    outputs(1387) <= layer0_outputs(2944);
    outputs(1388) <= not(layer0_outputs(2190));
    outputs(1389) <= not(layer0_outputs(472));
    outputs(1390) <= layer0_outputs(2462);
    outputs(1391) <= (layer0_outputs(3460)) or (layer0_outputs(2065));
    outputs(1392) <= not(layer0_outputs(3675));
    outputs(1393) <= not(layer0_outputs(175));
    outputs(1394) <= not(layer0_outputs(819));
    outputs(1395) <= layer0_outputs(1442);
    outputs(1396) <= not(layer0_outputs(632));
    outputs(1397) <= not(layer0_outputs(753));
    outputs(1398) <= not(layer0_outputs(1162)) or (layer0_outputs(5006));
    outputs(1399) <= layer0_outputs(4760);
    outputs(1400) <= layer0_outputs(3065);
    outputs(1401) <= '1';
    outputs(1402) <= (layer0_outputs(369)) xor (layer0_outputs(1495));
    outputs(1403) <= not(layer0_outputs(1310));
    outputs(1404) <= not((layer0_outputs(2830)) or (layer0_outputs(4316)));
    outputs(1405) <= not(layer0_outputs(4508));
    outputs(1406) <= not(layer0_outputs(1152));
    outputs(1407) <= (layer0_outputs(222)) xor (layer0_outputs(1481));
    outputs(1408) <= (layer0_outputs(1103)) and not (layer0_outputs(2414));
    outputs(1409) <= not((layer0_outputs(3063)) and (layer0_outputs(4497)));
    outputs(1410) <= not((layer0_outputs(212)) and (layer0_outputs(1718)));
    outputs(1411) <= layer0_outputs(3078);
    outputs(1412) <= (layer0_outputs(11)) and not (layer0_outputs(2212));
    outputs(1413) <= layer0_outputs(5118);
    outputs(1414) <= layer0_outputs(1365);
    outputs(1415) <= (layer0_outputs(3924)) xor (layer0_outputs(4946));
    outputs(1416) <= not(layer0_outputs(3111)) or (layer0_outputs(3451));
    outputs(1417) <= (layer0_outputs(3485)) and not (layer0_outputs(3450));
    outputs(1418) <= (layer0_outputs(798)) and not (layer0_outputs(2360));
    outputs(1419) <= layer0_outputs(107);
    outputs(1420) <= not(layer0_outputs(3169));
    outputs(1421) <= layer0_outputs(2129);
    outputs(1422) <= not((layer0_outputs(3266)) xor (layer0_outputs(1341)));
    outputs(1423) <= not(layer0_outputs(4824));
    outputs(1424) <= not(layer0_outputs(2973)) or (layer0_outputs(4870));
    outputs(1425) <= not((layer0_outputs(4698)) xor (layer0_outputs(760)));
    outputs(1426) <= not(layer0_outputs(2059)) or (layer0_outputs(441));
    outputs(1427) <= not(layer0_outputs(758));
    outputs(1428) <= layer0_outputs(4295);
    outputs(1429) <= not((layer0_outputs(2312)) and (layer0_outputs(1882)));
    outputs(1430) <= (layer0_outputs(1402)) or (layer0_outputs(2473));
    outputs(1431) <= (layer0_outputs(3599)) and (layer0_outputs(1967));
    outputs(1432) <= layer0_outputs(4127);
    outputs(1433) <= (layer0_outputs(3286)) or (layer0_outputs(3916));
    outputs(1434) <= not(layer0_outputs(2313));
    outputs(1435) <= layer0_outputs(3927);
    outputs(1436) <= not(layer0_outputs(567));
    outputs(1437) <= (layer0_outputs(2055)) and not (layer0_outputs(728));
    outputs(1438) <= (layer0_outputs(3995)) and not (layer0_outputs(341));
    outputs(1439) <= (layer0_outputs(643)) and not (layer0_outputs(1311));
    outputs(1440) <= layer0_outputs(2364);
    outputs(1441) <= not(layer0_outputs(1912));
    outputs(1442) <= (layer0_outputs(3066)) and not (layer0_outputs(793));
    outputs(1443) <= layer0_outputs(2514);
    outputs(1444) <= not((layer0_outputs(130)) or (layer0_outputs(3983)));
    outputs(1445) <= not(layer0_outputs(2943)) or (layer0_outputs(2066));
    outputs(1446) <= not(layer0_outputs(617)) or (layer0_outputs(4814));
    outputs(1447) <= not(layer0_outputs(4120));
    outputs(1448) <= (layer0_outputs(4758)) xor (layer0_outputs(3714));
    outputs(1449) <= not(layer0_outputs(1904)) or (layer0_outputs(3806));
    outputs(1450) <= (layer0_outputs(1821)) or (layer0_outputs(2270));
    outputs(1451) <= not(layer0_outputs(2921));
    outputs(1452) <= layer0_outputs(2599);
    outputs(1453) <= not(layer0_outputs(3416)) or (layer0_outputs(5020));
    outputs(1454) <= layer0_outputs(914);
    outputs(1455) <= not(layer0_outputs(1490)) or (layer0_outputs(157));
    outputs(1456) <= not(layer0_outputs(2299)) or (layer0_outputs(2278));
    outputs(1457) <= (layer0_outputs(4659)) xor (layer0_outputs(1505));
    outputs(1458) <= not(layer0_outputs(1663));
    outputs(1459) <= not(layer0_outputs(2483)) or (layer0_outputs(3598));
    outputs(1460) <= layer0_outputs(1625);
    outputs(1461) <= '1';
    outputs(1462) <= not(layer0_outputs(3955)) or (layer0_outputs(2770));
    outputs(1463) <= not(layer0_outputs(1470));
    outputs(1464) <= layer0_outputs(1673);
    outputs(1465) <= not((layer0_outputs(2685)) xor (layer0_outputs(3114)));
    outputs(1466) <= not(layer0_outputs(4841)) or (layer0_outputs(4054));
    outputs(1467) <= layer0_outputs(125);
    outputs(1468) <= layer0_outputs(5107);
    outputs(1469) <= (layer0_outputs(760)) and (layer0_outputs(3752));
    outputs(1470) <= not((layer0_outputs(4304)) xor (layer0_outputs(4422)));
    outputs(1471) <= layer0_outputs(1435);
    outputs(1472) <= layer0_outputs(1200);
    outputs(1473) <= layer0_outputs(2769);
    outputs(1474) <= (layer0_outputs(4305)) xor (layer0_outputs(4749));
    outputs(1475) <= (layer0_outputs(2485)) and not (layer0_outputs(3756));
    outputs(1476) <= not((layer0_outputs(23)) and (layer0_outputs(1839)));
    outputs(1477) <= not(layer0_outputs(3573));
    outputs(1478) <= not((layer0_outputs(4615)) or (layer0_outputs(2765)));
    outputs(1479) <= (layer0_outputs(214)) and not (layer0_outputs(976));
    outputs(1480) <= (layer0_outputs(589)) or (layer0_outputs(3136));
    outputs(1481) <= (layer0_outputs(2405)) or (layer0_outputs(4264));
    outputs(1482) <= not((layer0_outputs(2630)) and (layer0_outputs(3068)));
    outputs(1483) <= not((layer0_outputs(2351)) and (layer0_outputs(4757)));
    outputs(1484) <= not(layer0_outputs(1133));
    outputs(1485) <= not(layer0_outputs(3084));
    outputs(1486) <= not((layer0_outputs(3858)) or (layer0_outputs(4580)));
    outputs(1487) <= layer0_outputs(4710);
    outputs(1488) <= not(layer0_outputs(3350));
    outputs(1489) <= not((layer0_outputs(1959)) and (layer0_outputs(489)));
    outputs(1490) <= layer0_outputs(814);
    outputs(1491) <= layer0_outputs(4252);
    outputs(1492) <= (layer0_outputs(4280)) xor (layer0_outputs(1891));
    outputs(1493) <= not(layer0_outputs(1587));
    outputs(1494) <= not(layer0_outputs(3773));
    outputs(1495) <= (layer0_outputs(3636)) xor (layer0_outputs(152));
    outputs(1496) <= not(layer0_outputs(305)) or (layer0_outputs(1650));
    outputs(1497) <= not(layer0_outputs(2434));
    outputs(1498) <= (layer0_outputs(1121)) xor (layer0_outputs(3607));
    outputs(1499) <= not(layer0_outputs(3572));
    outputs(1500) <= not(layer0_outputs(2873)) or (layer0_outputs(4839));
    outputs(1501) <= (layer0_outputs(2834)) and (layer0_outputs(3889));
    outputs(1502) <= not(layer0_outputs(2176));
    outputs(1503) <= layer0_outputs(4492);
    outputs(1504) <= not(layer0_outputs(1832)) or (layer0_outputs(827));
    outputs(1505) <= not((layer0_outputs(3611)) or (layer0_outputs(1466)));
    outputs(1506) <= not(layer0_outputs(1263));
    outputs(1507) <= not(layer0_outputs(21)) or (layer0_outputs(1113));
    outputs(1508) <= not(layer0_outputs(395));
    outputs(1509) <= (layer0_outputs(4968)) xor (layer0_outputs(1287));
    outputs(1510) <= not(layer0_outputs(1604));
    outputs(1511) <= not(layer0_outputs(3081));
    outputs(1512) <= not((layer0_outputs(2823)) xor (layer0_outputs(2372)));
    outputs(1513) <= not((layer0_outputs(2001)) or (layer0_outputs(2840)));
    outputs(1514) <= not((layer0_outputs(4956)) and (layer0_outputs(378)));
    outputs(1515) <= not(layer0_outputs(873)) or (layer0_outputs(5021));
    outputs(1516) <= not(layer0_outputs(3344)) or (layer0_outputs(4781));
    outputs(1517) <= (layer0_outputs(3227)) or (layer0_outputs(3179));
    outputs(1518) <= not((layer0_outputs(767)) or (layer0_outputs(4449)));
    outputs(1519) <= (layer0_outputs(3697)) xor (layer0_outputs(2804));
    outputs(1520) <= layer0_outputs(170);
    outputs(1521) <= (layer0_outputs(2321)) and not (layer0_outputs(85));
    outputs(1522) <= layer0_outputs(1759);
    outputs(1523) <= (layer0_outputs(69)) xor (layer0_outputs(2214));
    outputs(1524) <= (layer0_outputs(2263)) and (layer0_outputs(2337));
    outputs(1525) <= (layer0_outputs(4234)) and not (layer0_outputs(3407));
    outputs(1526) <= not((layer0_outputs(3964)) or (layer0_outputs(4099)));
    outputs(1527) <= layer0_outputs(3647);
    outputs(1528) <= not(layer0_outputs(3394));
    outputs(1529) <= layer0_outputs(565);
    outputs(1530) <= layer0_outputs(4208);
    outputs(1531) <= (layer0_outputs(3644)) and not (layer0_outputs(898));
    outputs(1532) <= layer0_outputs(554);
    outputs(1533) <= layer0_outputs(2912);
    outputs(1534) <= not(layer0_outputs(1522));
    outputs(1535) <= (layer0_outputs(720)) and not (layer0_outputs(2800));
    outputs(1536) <= not(layer0_outputs(3435));
    outputs(1537) <= not(layer0_outputs(4232));
    outputs(1538) <= layer0_outputs(2731);
    outputs(1539) <= not(layer0_outputs(3784));
    outputs(1540) <= (layer0_outputs(2755)) xor (layer0_outputs(969));
    outputs(1541) <= (layer0_outputs(3672)) or (layer0_outputs(4192));
    outputs(1542) <= (layer0_outputs(867)) and not (layer0_outputs(285));
    outputs(1543) <= not(layer0_outputs(429)) or (layer0_outputs(1939));
    outputs(1544) <= not(layer0_outputs(2748));
    outputs(1545) <= layer0_outputs(3893);
    outputs(1546) <= layer0_outputs(3704);
    outputs(1547) <= layer0_outputs(4378);
    outputs(1548) <= not(layer0_outputs(2855)) or (layer0_outputs(4503));
    outputs(1549) <= (layer0_outputs(3583)) xor (layer0_outputs(317));
    outputs(1550) <= (layer0_outputs(4584)) or (layer0_outputs(3633));
    outputs(1551) <= (layer0_outputs(3897)) xor (layer0_outputs(4066));
    outputs(1552) <= not(layer0_outputs(3561)) or (layer0_outputs(1771));
    outputs(1553) <= not(layer0_outputs(1319));
    outputs(1554) <= not(layer0_outputs(543)) or (layer0_outputs(4874));
    outputs(1555) <= (layer0_outputs(74)) xor (layer0_outputs(2254));
    outputs(1556) <= not(layer0_outputs(4398));
    outputs(1557) <= (layer0_outputs(39)) and not (layer0_outputs(3666));
    outputs(1558) <= (layer0_outputs(249)) and not (layer0_outputs(2869));
    outputs(1559) <= not(layer0_outputs(524));
    outputs(1560) <= layer0_outputs(3100);
    outputs(1561) <= (layer0_outputs(4854)) and not (layer0_outputs(4038));
    outputs(1562) <= not(layer0_outputs(1167));
    outputs(1563) <= not(layer0_outputs(2834));
    outputs(1564) <= (layer0_outputs(4502)) and not (layer0_outputs(463));
    outputs(1565) <= not(layer0_outputs(3365));
    outputs(1566) <= not(layer0_outputs(1751));
    outputs(1567) <= layer0_outputs(4039);
    outputs(1568) <= (layer0_outputs(3628)) xor (layer0_outputs(1331));
    outputs(1569) <= not(layer0_outputs(4689)) or (layer0_outputs(525));
    outputs(1570) <= not(layer0_outputs(4666));
    outputs(1571) <= layer0_outputs(2721);
    outputs(1572) <= (layer0_outputs(889)) xor (layer0_outputs(2282));
    outputs(1573) <= not(layer0_outputs(2028));
    outputs(1574) <= not(layer0_outputs(2575));
    outputs(1575) <= (layer0_outputs(2919)) and (layer0_outputs(4670));
    outputs(1576) <= not(layer0_outputs(4506));
    outputs(1577) <= (layer0_outputs(2195)) and (layer0_outputs(2198));
    outputs(1578) <= not(layer0_outputs(3458)) or (layer0_outputs(2623));
    outputs(1579) <= (layer0_outputs(5048)) xor (layer0_outputs(3643));
    outputs(1580) <= not(layer0_outputs(80));
    outputs(1581) <= (layer0_outputs(1926)) xor (layer0_outputs(336));
    outputs(1582) <= not((layer0_outputs(392)) or (layer0_outputs(2318)));
    outputs(1583) <= layer0_outputs(4740);
    outputs(1584) <= (layer0_outputs(81)) xor (layer0_outputs(390));
    outputs(1585) <= not(layer0_outputs(2445));
    outputs(1586) <= not((layer0_outputs(3871)) or (layer0_outputs(412)));
    outputs(1587) <= not(layer0_outputs(3906)) or (layer0_outputs(751));
    outputs(1588) <= not(layer0_outputs(405));
    outputs(1589) <= (layer0_outputs(885)) and not (layer0_outputs(4822));
    outputs(1590) <= layer0_outputs(3951);
    outputs(1591) <= (layer0_outputs(3094)) and not (layer0_outputs(2852));
    outputs(1592) <= layer0_outputs(1038);
    outputs(1593) <= (layer0_outputs(3514)) and not (layer0_outputs(4637));
    outputs(1594) <= not(layer0_outputs(2437));
    outputs(1595) <= not(layer0_outputs(2446));
    outputs(1596) <= layer0_outputs(3132);
    outputs(1597) <= not((layer0_outputs(388)) xor (layer0_outputs(60)));
    outputs(1598) <= layer0_outputs(3009);
    outputs(1599) <= not(layer0_outputs(5080));
    outputs(1600) <= (layer0_outputs(3423)) and not (layer0_outputs(706));
    outputs(1601) <= not(layer0_outputs(4089)) or (layer0_outputs(2577));
    outputs(1602) <= not(layer0_outputs(4671)) or (layer0_outputs(4932));
    outputs(1603) <= layer0_outputs(3705);
    outputs(1604) <= not((layer0_outputs(868)) or (layer0_outputs(4809)));
    outputs(1605) <= not(layer0_outputs(3895)) or (layer0_outputs(4906));
    outputs(1606) <= not(layer0_outputs(1584));
    outputs(1607) <= not((layer0_outputs(2563)) xor (layer0_outputs(259)));
    outputs(1608) <= not(layer0_outputs(1721));
    outputs(1609) <= not(layer0_outputs(2202)) or (layer0_outputs(4499));
    outputs(1610) <= not((layer0_outputs(4300)) xor (layer0_outputs(2167)));
    outputs(1611) <= (layer0_outputs(4347)) xor (layer0_outputs(4454));
    outputs(1612) <= layer0_outputs(2660);
    outputs(1613) <= not((layer0_outputs(4022)) xor (layer0_outputs(2927)));
    outputs(1614) <= not((layer0_outputs(1852)) xor (layer0_outputs(2381)));
    outputs(1615) <= (layer0_outputs(4676)) or (layer0_outputs(4917));
    outputs(1616) <= (layer0_outputs(4073)) and not (layer0_outputs(144));
    outputs(1617) <= not(layer0_outputs(2325));
    outputs(1618) <= (layer0_outputs(4366)) xor (layer0_outputs(963));
    outputs(1619) <= layer0_outputs(1328);
    outputs(1620) <= layer0_outputs(2090);
    outputs(1621) <= layer0_outputs(3242);
    outputs(1622) <= not(layer0_outputs(2998)) or (layer0_outputs(2656));
    outputs(1623) <= layer0_outputs(2425);
    outputs(1624) <= (layer0_outputs(5023)) xor (layer0_outputs(4243));
    outputs(1625) <= not(layer0_outputs(440));
    outputs(1626) <= not(layer0_outputs(1740));
    outputs(1627) <= layer0_outputs(4776);
    outputs(1628) <= not(layer0_outputs(3147));
    outputs(1629) <= not(layer0_outputs(1953));
    outputs(1630) <= not(layer0_outputs(2279));
    outputs(1631) <= not(layer0_outputs(3306));
    outputs(1632) <= (layer0_outputs(1132)) and (layer0_outputs(1201));
    outputs(1633) <= not(layer0_outputs(2152));
    outputs(1634) <= not(layer0_outputs(1138));
    outputs(1635) <= not((layer0_outputs(2890)) and (layer0_outputs(2183)));
    outputs(1636) <= not(layer0_outputs(2549)) or (layer0_outputs(541));
    outputs(1637) <= (layer0_outputs(960)) and (layer0_outputs(1957));
    outputs(1638) <= (layer0_outputs(322)) and (layer0_outputs(50));
    outputs(1639) <= not(layer0_outputs(1165));
    outputs(1640) <= not(layer0_outputs(4432)) or (layer0_outputs(3601));
    outputs(1641) <= layer0_outputs(3754);
    outputs(1642) <= not((layer0_outputs(1041)) or (layer0_outputs(4423)));
    outputs(1643) <= (layer0_outputs(2122)) and not (layer0_outputs(2420));
    outputs(1644) <= not(layer0_outputs(2862)) or (layer0_outputs(2386));
    outputs(1645) <= not(layer0_outputs(3129)) or (layer0_outputs(3822));
    outputs(1646) <= not(layer0_outputs(164));
    outputs(1647) <= not((layer0_outputs(2437)) or (layer0_outputs(5014)));
    outputs(1648) <= (layer0_outputs(332)) and (layer0_outputs(3551));
    outputs(1649) <= (layer0_outputs(3140)) or (layer0_outputs(2810));
    outputs(1650) <= not(layer0_outputs(3466));
    outputs(1651) <= not(layer0_outputs(3085));
    outputs(1652) <= layer0_outputs(1465);
    outputs(1653) <= (layer0_outputs(1520)) and not (layer0_outputs(3728));
    outputs(1654) <= layer0_outputs(4499);
    outputs(1655) <= layer0_outputs(1649);
    outputs(1656) <= (layer0_outputs(1109)) xor (layer0_outputs(3301));
    outputs(1657) <= not((layer0_outputs(3558)) or (layer0_outputs(1131)));
    outputs(1658) <= not((layer0_outputs(3106)) and (layer0_outputs(4672)));
    outputs(1659) <= layer0_outputs(5087);
    outputs(1660) <= not(layer0_outputs(2575));
    outputs(1661) <= not((layer0_outputs(2327)) and (layer0_outputs(2186)));
    outputs(1662) <= (layer0_outputs(246)) and not (layer0_outputs(1772));
    outputs(1663) <= layer0_outputs(1320);
    outputs(1664) <= not((layer0_outputs(3912)) and (layer0_outputs(1275)));
    outputs(1665) <= not((layer0_outputs(1176)) xor (layer0_outputs(447)));
    outputs(1666) <= not(layer0_outputs(321));
    outputs(1667) <= (layer0_outputs(2430)) or (layer0_outputs(3677));
    outputs(1668) <= layer0_outputs(235);
    outputs(1669) <= layer0_outputs(120);
    outputs(1670) <= layer0_outputs(853);
    outputs(1671) <= not((layer0_outputs(1277)) and (layer0_outputs(4762)));
    outputs(1672) <= not(layer0_outputs(501)) or (layer0_outputs(3776));
    outputs(1673) <= not(layer0_outputs(891));
    outputs(1674) <= not(layer0_outputs(4947));
    outputs(1675) <= not(layer0_outputs(1676));
    outputs(1676) <= (layer0_outputs(1679)) or (layer0_outputs(3220));
    outputs(1677) <= not((layer0_outputs(1350)) and (layer0_outputs(2867)));
    outputs(1678) <= (layer0_outputs(849)) and (layer0_outputs(4891));
    outputs(1679) <= '1';
    outputs(1680) <= (layer0_outputs(3947)) and not (layer0_outputs(65));
    outputs(1681) <= (layer0_outputs(1230)) and (layer0_outputs(1968));
    outputs(1682) <= (layer0_outputs(3471)) xor (layer0_outputs(4886));
    outputs(1683) <= (layer0_outputs(3180)) and not (layer0_outputs(812));
    outputs(1684) <= not(layer0_outputs(769));
    outputs(1685) <= (layer0_outputs(2727)) and (layer0_outputs(1959));
    outputs(1686) <= not(layer0_outputs(297));
    outputs(1687) <= not(layer0_outputs(2273));
    outputs(1688) <= not((layer0_outputs(679)) xor (layer0_outputs(4006)));
    outputs(1689) <= not((layer0_outputs(3178)) or (layer0_outputs(117)));
    outputs(1690) <= not(layer0_outputs(6));
    outputs(1691) <= (layer0_outputs(1459)) xor (layer0_outputs(3145));
    outputs(1692) <= not((layer0_outputs(2370)) xor (layer0_outputs(2910)));
    outputs(1693) <= (layer0_outputs(167)) and (layer0_outputs(4804));
    outputs(1694) <= not(layer0_outputs(4610));
    outputs(1695) <= layer0_outputs(184);
    outputs(1696) <= not((layer0_outputs(5070)) xor (layer0_outputs(3137)));
    outputs(1697) <= (layer0_outputs(83)) xor (layer0_outputs(49));
    outputs(1698) <= (layer0_outputs(406)) and not (layer0_outputs(293));
    outputs(1699) <= layer0_outputs(1295);
    outputs(1700) <= not(layer0_outputs(1549));
    outputs(1701) <= not((layer0_outputs(259)) or (layer0_outputs(3947)));
    outputs(1702) <= not(layer0_outputs(3272));
    outputs(1703) <= (layer0_outputs(1971)) and (layer0_outputs(2573));
    outputs(1704) <= not(layer0_outputs(674));
    outputs(1705) <= not((layer0_outputs(3663)) or (layer0_outputs(1927)));
    outputs(1706) <= not(layer0_outputs(1893));
    outputs(1707) <= not(layer0_outputs(831));
    outputs(1708) <= (layer0_outputs(2853)) and (layer0_outputs(4815));
    outputs(1709) <= layer0_outputs(3964);
    outputs(1710) <= not((layer0_outputs(2918)) or (layer0_outputs(5050)));
    outputs(1711) <= layer0_outputs(3069);
    outputs(1712) <= not((layer0_outputs(4665)) or (layer0_outputs(3477)));
    outputs(1713) <= layer0_outputs(4906);
    outputs(1714) <= (layer0_outputs(619)) xor (layer0_outputs(784));
    outputs(1715) <= not(layer0_outputs(4141));
    outputs(1716) <= (layer0_outputs(3269)) and (layer0_outputs(2024));
    outputs(1717) <= (layer0_outputs(1948)) or (layer0_outputs(2744));
    outputs(1718) <= (layer0_outputs(95)) and not (layer0_outputs(2822));
    outputs(1719) <= (layer0_outputs(1851)) and not (layer0_outputs(2336));
    outputs(1720) <= layer0_outputs(4831);
    outputs(1721) <= not((layer0_outputs(4620)) and (layer0_outputs(3977)));
    outputs(1722) <= layer0_outputs(3825);
    outputs(1723) <= not((layer0_outputs(1436)) xor (layer0_outputs(2329)));
    outputs(1724) <= (layer0_outputs(1188)) and (layer0_outputs(2977));
    outputs(1725) <= layer0_outputs(3985);
    outputs(1726) <= not(layer0_outputs(3030));
    outputs(1727) <= (layer0_outputs(4744)) and (layer0_outputs(3438));
    outputs(1728) <= not(layer0_outputs(4034)) or (layer0_outputs(404));
    outputs(1729) <= layer0_outputs(3709);
    outputs(1730) <= not(layer0_outputs(1790)) or (layer0_outputs(455));
    outputs(1731) <= layer0_outputs(689);
    outputs(1732) <= not(layer0_outputs(802));
    outputs(1733) <= layer0_outputs(3717);
    outputs(1734) <= not((layer0_outputs(3005)) or (layer0_outputs(2200)));
    outputs(1735) <= layer0_outputs(3239);
    outputs(1736) <= not(layer0_outputs(1531));
    outputs(1737) <= not((layer0_outputs(333)) xor (layer0_outputs(4186)));
    outputs(1738) <= not(layer0_outputs(1020));
    outputs(1739) <= not(layer0_outputs(3998)) or (layer0_outputs(2238));
    outputs(1740) <= layer0_outputs(2971);
    outputs(1741) <= (layer0_outputs(1927)) xor (layer0_outputs(2538));
    outputs(1742) <= not(layer0_outputs(4276));
    outputs(1743) <= (layer0_outputs(761)) and not (layer0_outputs(2460));
    outputs(1744) <= layer0_outputs(35);
    outputs(1745) <= layer0_outputs(3327);
    outputs(1746) <= (layer0_outputs(3900)) and not (layer0_outputs(4530));
    outputs(1747) <= not(layer0_outputs(1482));
    outputs(1748) <= (layer0_outputs(2042)) and not (layer0_outputs(673));
    outputs(1749) <= (layer0_outputs(3300)) xor (layer0_outputs(1597));
    outputs(1750) <= layer0_outputs(4339);
    outputs(1751) <= layer0_outputs(3948);
    outputs(1752) <= (layer0_outputs(4753)) xor (layer0_outputs(2801));
    outputs(1753) <= layer0_outputs(1338);
    outputs(1754) <= layer0_outputs(1420);
    outputs(1755) <= not((layer0_outputs(161)) xor (layer0_outputs(2155)));
    outputs(1756) <= not(layer0_outputs(2167));
    outputs(1757) <= not(layer0_outputs(4685));
    outputs(1758) <= not(layer0_outputs(4258));
    outputs(1759) <= layer0_outputs(176);
    outputs(1760) <= layer0_outputs(455);
    outputs(1761) <= not(layer0_outputs(4000));
    outputs(1762) <= layer0_outputs(4521);
    outputs(1763) <= not(layer0_outputs(1345));
    outputs(1764) <= not((layer0_outputs(4763)) xor (layer0_outputs(101)));
    outputs(1765) <= layer0_outputs(2779);
    outputs(1766) <= not((layer0_outputs(4291)) xor (layer0_outputs(3530)));
    outputs(1767) <= (layer0_outputs(2307)) and not (layer0_outputs(2839));
    outputs(1768) <= layer0_outputs(4795);
    outputs(1769) <= not((layer0_outputs(2836)) xor (layer0_outputs(3588)));
    outputs(1770) <= (layer0_outputs(4726)) and not (layer0_outputs(4601));
    outputs(1771) <= layer0_outputs(4503);
    outputs(1772) <= not((layer0_outputs(3648)) xor (layer0_outputs(3352)));
    outputs(1773) <= not((layer0_outputs(4567)) xor (layer0_outputs(691)));
    outputs(1774) <= not(layer0_outputs(4796)) or (layer0_outputs(1354));
    outputs(1775) <= layer0_outputs(3469);
    outputs(1776) <= layer0_outputs(4335);
    outputs(1777) <= not(layer0_outputs(1408));
    outputs(1778) <= '1';
    outputs(1779) <= (layer0_outputs(1692)) xor (layer0_outputs(826));
    outputs(1780) <= not(layer0_outputs(3383));
    outputs(1781) <= (layer0_outputs(1723)) xor (layer0_outputs(1974));
    outputs(1782) <= not(layer0_outputs(4692));
    outputs(1783) <= not((layer0_outputs(1633)) and (layer0_outputs(5038)));
    outputs(1784) <= (layer0_outputs(135)) and not (layer0_outputs(4136));
    outputs(1785) <= not(layer0_outputs(4433));
    outputs(1786) <= not(layer0_outputs(493)) or (layer0_outputs(2053));
    outputs(1787) <= not(layer0_outputs(323));
    outputs(1788) <= not((layer0_outputs(2076)) and (layer0_outputs(619)));
    outputs(1789) <= not(layer0_outputs(2683));
    outputs(1790) <= not((layer0_outputs(1833)) xor (layer0_outputs(2886)));
    outputs(1791) <= (layer0_outputs(4125)) and not (layer0_outputs(709));
    outputs(1792) <= not(layer0_outputs(4927));
    outputs(1793) <= not((layer0_outputs(2714)) xor (layer0_outputs(3297)));
    outputs(1794) <= not((layer0_outputs(3818)) and (layer0_outputs(4373)));
    outputs(1795) <= not(layer0_outputs(752)) or (layer0_outputs(541));
    outputs(1796) <= (layer0_outputs(1505)) xor (layer0_outputs(3973));
    outputs(1797) <= not(layer0_outputs(864)) or (layer0_outputs(1416));
    outputs(1798) <= not(layer0_outputs(2343));
    outputs(1799) <= (layer0_outputs(1512)) or (layer0_outputs(4720));
    outputs(1800) <= (layer0_outputs(1254)) and (layer0_outputs(330));
    outputs(1801) <= (layer0_outputs(4202)) xor (layer0_outputs(3247));
    outputs(1802) <= (layer0_outputs(1276)) and not (layer0_outputs(5039));
    outputs(1803) <= not(layer0_outputs(968));
    outputs(1804) <= not((layer0_outputs(2732)) xor (layer0_outputs(2173)));
    outputs(1805) <= not((layer0_outputs(2401)) xor (layer0_outputs(4754)));
    outputs(1806) <= layer0_outputs(3122);
    outputs(1807) <= not(layer0_outputs(2855));
    outputs(1808) <= (layer0_outputs(3612)) and not (layer0_outputs(4256));
    outputs(1809) <= not((layer0_outputs(239)) or (layer0_outputs(1488)));
    outputs(1810) <= not(layer0_outputs(2028));
    outputs(1811) <= not(layer0_outputs(2903)) or (layer0_outputs(1401));
    outputs(1812) <= layer0_outputs(360);
    outputs(1813) <= (layer0_outputs(2530)) and not (layer0_outputs(3727));
    outputs(1814) <= (layer0_outputs(2915)) xor (layer0_outputs(667));
    outputs(1815) <= not((layer0_outputs(857)) xor (layer0_outputs(358)));
    outputs(1816) <= (layer0_outputs(3884)) and (layer0_outputs(3148));
    outputs(1817) <= not((layer0_outputs(3047)) or (layer0_outputs(1107)));
    outputs(1818) <= (layer0_outputs(2939)) or (layer0_outputs(3153));
    outputs(1819) <= not((layer0_outputs(1169)) xor (layer0_outputs(3139)));
    outputs(1820) <= not((layer0_outputs(2489)) xor (layer0_outputs(5091)));
    outputs(1821) <= not(layer0_outputs(2109)) or (layer0_outputs(844));
    outputs(1822) <= (layer0_outputs(2324)) and (layer0_outputs(4451));
    outputs(1823) <= not(layer0_outputs(1933)) or (layer0_outputs(697));
    outputs(1824) <= not(layer0_outputs(4936));
    outputs(1825) <= not(layer0_outputs(470)) or (layer0_outputs(431));
    outputs(1826) <= not((layer0_outputs(5049)) or (layer0_outputs(775)));
    outputs(1827) <= layer0_outputs(3000);
    outputs(1828) <= (layer0_outputs(4224)) xor (layer0_outputs(2678));
    outputs(1829) <= not(layer0_outputs(1377));
    outputs(1830) <= (layer0_outputs(3894)) xor (layer0_outputs(1900));
    outputs(1831) <= not((layer0_outputs(1068)) xor (layer0_outputs(4616)));
    outputs(1832) <= not((layer0_outputs(4866)) xor (layer0_outputs(3698)));
    outputs(1833) <= not((layer0_outputs(2075)) or (layer0_outputs(4109)));
    outputs(1834) <= (layer0_outputs(1333)) xor (layer0_outputs(4871));
    outputs(1835) <= not(layer0_outputs(177)) or (layer0_outputs(107));
    outputs(1836) <= not((layer0_outputs(4885)) xor (layer0_outputs(5066)));
    outputs(1837) <= not(layer0_outputs(2672));
    outputs(1838) <= not(layer0_outputs(437)) or (layer0_outputs(2447));
    outputs(1839) <= not(layer0_outputs(1808)) or (layer0_outputs(1895));
    outputs(1840) <= layer0_outputs(3733);
    outputs(1841) <= not(layer0_outputs(1059)) or (layer0_outputs(2142));
    outputs(1842) <= (layer0_outputs(703)) xor (layer0_outputs(1902));
    outputs(1843) <= (layer0_outputs(3345)) xor (layer0_outputs(2861));
    outputs(1844) <= not((layer0_outputs(2071)) xor (layer0_outputs(2378)));
    outputs(1845) <= layer0_outputs(2005);
    outputs(1846) <= (layer0_outputs(4571)) xor (layer0_outputs(708));
    outputs(1847) <= not(layer0_outputs(2102)) or (layer0_outputs(3122));
    outputs(1848) <= not(layer0_outputs(4274));
    outputs(1849) <= not(layer0_outputs(1924));
    outputs(1850) <= layer0_outputs(1401);
    outputs(1851) <= not(layer0_outputs(432));
    outputs(1852) <= not((layer0_outputs(313)) and (layer0_outputs(1746)));
    outputs(1853) <= not((layer0_outputs(514)) xor (layer0_outputs(3998)));
    outputs(1854) <= (layer0_outputs(5113)) and (layer0_outputs(3625));
    outputs(1855) <= (layer0_outputs(3266)) xor (layer0_outputs(1539));
    outputs(1856) <= layer0_outputs(1328);
    outputs(1857) <= layer0_outputs(3257);
    outputs(1858) <= (layer0_outputs(2788)) and (layer0_outputs(3613));
    outputs(1859) <= not((layer0_outputs(223)) xor (layer0_outputs(4695)));
    outputs(1860) <= '1';
    outputs(1861) <= not(layer0_outputs(2125));
    outputs(1862) <= layer0_outputs(4930);
    outputs(1863) <= not(layer0_outputs(2002));
    outputs(1864) <= not(layer0_outputs(3216));
    outputs(1865) <= (layer0_outputs(2007)) or (layer0_outputs(1082));
    outputs(1866) <= layer0_outputs(2936);
    outputs(1867) <= layer0_outputs(1497);
    outputs(1868) <= '1';
    outputs(1869) <= not(layer0_outputs(3813));
    outputs(1870) <= not((layer0_outputs(2433)) and (layer0_outputs(836)));
    outputs(1871) <= (layer0_outputs(2380)) and not (layer0_outputs(736));
    outputs(1872) <= not(layer0_outputs(2132));
    outputs(1873) <= not((layer0_outputs(130)) xor (layer0_outputs(3864)));
    outputs(1874) <= (layer0_outputs(1207)) and not (layer0_outputs(4724));
    outputs(1875) <= not((layer0_outputs(503)) or (layer0_outputs(4858)));
    outputs(1876) <= layer0_outputs(1678);
    outputs(1877) <= not(layer0_outputs(1508));
    outputs(1878) <= (layer0_outputs(2889)) and (layer0_outputs(2806));
    outputs(1879) <= (layer0_outputs(2307)) and not (layer0_outputs(1425));
    outputs(1880) <= (layer0_outputs(356)) or (layer0_outputs(910));
    outputs(1881) <= not(layer0_outputs(4274));
    outputs(1882) <= not((layer0_outputs(1381)) xor (layer0_outputs(1441)));
    outputs(1883) <= not((layer0_outputs(2017)) and (layer0_outputs(4395)));
    outputs(1884) <= not((layer0_outputs(586)) xor (layer0_outputs(3164)));
    outputs(1885) <= (layer0_outputs(3991)) or (layer0_outputs(5011));
    outputs(1886) <= not((layer0_outputs(813)) xor (layer0_outputs(4244)));
    outputs(1887) <= not((layer0_outputs(3719)) and (layer0_outputs(4022)));
    outputs(1888) <= not(layer0_outputs(940));
    outputs(1889) <= (layer0_outputs(4638)) and (layer0_outputs(388));
    outputs(1890) <= not(layer0_outputs(2109));
    outputs(1891) <= layer0_outputs(587);
    outputs(1892) <= layer0_outputs(2373);
    outputs(1893) <= not(layer0_outputs(1273));
    outputs(1894) <= not(layer0_outputs(1604));
    outputs(1895) <= layer0_outputs(4989);
    outputs(1896) <= layer0_outputs(746);
    outputs(1897) <= layer0_outputs(4515);
    outputs(1898) <= layer0_outputs(901);
    outputs(1899) <= not(layer0_outputs(5066)) or (layer0_outputs(1159));
    outputs(1900) <= (layer0_outputs(3224)) and (layer0_outputs(4148));
    outputs(1901) <= (layer0_outputs(4851)) and (layer0_outputs(1217));
    outputs(1902) <= not(layer0_outputs(980));
    outputs(1903) <= layer0_outputs(3660);
    outputs(1904) <= layer0_outputs(3312);
    outputs(1905) <= not(layer0_outputs(4209)) or (layer0_outputs(4648));
    outputs(1906) <= layer0_outputs(1615);
    outputs(1907) <= layer0_outputs(4949);
    outputs(1908) <= not((layer0_outputs(876)) or (layer0_outputs(748)));
    outputs(1909) <= not(layer0_outputs(4249));
    outputs(1910) <= not(layer0_outputs(4079)) or (layer0_outputs(5119));
    outputs(1911) <= layer0_outputs(3175);
    outputs(1912) <= not(layer0_outputs(2674)) or (layer0_outputs(4767));
    outputs(1913) <= not(layer0_outputs(5084));
    outputs(1914) <= (layer0_outputs(4649)) and (layer0_outputs(3952));
    outputs(1915) <= layer0_outputs(2439);
    outputs(1916) <= layer0_outputs(3566);
    outputs(1917) <= (layer0_outputs(2506)) and not (layer0_outputs(4283));
    outputs(1918) <= not(layer0_outputs(3371));
    outputs(1919) <= (layer0_outputs(1734)) xor (layer0_outputs(3814));
    outputs(1920) <= (layer0_outputs(3682)) or (layer0_outputs(2270));
    outputs(1921) <= not(layer0_outputs(4402));
    outputs(1922) <= (layer0_outputs(3031)) or (layer0_outputs(1089));
    outputs(1923) <= layer0_outputs(3700);
    outputs(1924) <= layer0_outputs(896);
    outputs(1925) <= layer0_outputs(5114);
    outputs(1926) <= not(layer0_outputs(592));
    outputs(1927) <= not((layer0_outputs(1070)) and (layer0_outputs(1332)));
    outputs(1928) <= not(layer0_outputs(3526));
    outputs(1929) <= layer0_outputs(791);
    outputs(1930) <= (layer0_outputs(2136)) and not (layer0_outputs(3003));
    outputs(1931) <= layer0_outputs(1744);
    outputs(1932) <= (layer0_outputs(4118)) and not (layer0_outputs(4350));
    outputs(1933) <= layer0_outputs(5046);
    outputs(1934) <= not((layer0_outputs(4028)) or (layer0_outputs(276)));
    outputs(1935) <= layer0_outputs(1027);
    outputs(1936) <= not((layer0_outputs(1749)) xor (layer0_outputs(432)));
    outputs(1937) <= not(layer0_outputs(3226)) or (layer0_outputs(4830));
    outputs(1938) <= layer0_outputs(1507);
    outputs(1939) <= not(layer0_outputs(4996)) or (layer0_outputs(3019));
    outputs(1940) <= layer0_outputs(1814);
    outputs(1941) <= not(layer0_outputs(3267));
    outputs(1942) <= not(layer0_outputs(2652));
    outputs(1943) <= not(layer0_outputs(4013));
    outputs(1944) <= (layer0_outputs(1888)) xor (layer0_outputs(2457));
    outputs(1945) <= layer0_outputs(3741);
    outputs(1946) <= layer0_outputs(4107);
    outputs(1947) <= not(layer0_outputs(4526));
    outputs(1948) <= layer0_outputs(1762);
    outputs(1949) <= layer0_outputs(3148);
    outputs(1950) <= (layer0_outputs(1005)) xor (layer0_outputs(4349));
    outputs(1951) <= (layer0_outputs(4654)) and (layer0_outputs(2530));
    outputs(1952) <= (layer0_outputs(2168)) xor (layer0_outputs(703));
    outputs(1953) <= not(layer0_outputs(2844));
    outputs(1954) <= not((layer0_outputs(3360)) and (layer0_outputs(2453)));
    outputs(1955) <= not(layer0_outputs(1034));
    outputs(1956) <= not((layer0_outputs(1272)) or (layer0_outputs(428)));
    outputs(1957) <= layer0_outputs(4911);
    outputs(1958) <= not(layer0_outputs(362)) or (layer0_outputs(278));
    outputs(1959) <= not(layer0_outputs(4023));
    outputs(1960) <= (layer0_outputs(2238)) or (layer0_outputs(301));
    outputs(1961) <= (layer0_outputs(3268)) and not (layer0_outputs(780));
    outputs(1962) <= layer0_outputs(2910);
    outputs(1963) <= not(layer0_outputs(2418));
    outputs(1964) <= not((layer0_outputs(4571)) xor (layer0_outputs(3615)));
    outputs(1965) <= not(layer0_outputs(5090));
    outputs(1966) <= not((layer0_outputs(1955)) and (layer0_outputs(918)));
    outputs(1967) <= not(layer0_outputs(108));
    outputs(1968) <= layer0_outputs(2458);
    outputs(1969) <= (layer0_outputs(2567)) or (layer0_outputs(2693));
    outputs(1970) <= layer0_outputs(2254);
    outputs(1971) <= not(layer0_outputs(3687)) or (layer0_outputs(2308));
    outputs(1972) <= not((layer0_outputs(102)) xor (layer0_outputs(977)));
    outputs(1973) <= not((layer0_outputs(1389)) xor (layer0_outputs(2714)));
    outputs(1974) <= '1';
    outputs(1975) <= (layer0_outputs(1398)) xor (layer0_outputs(2825));
    outputs(1976) <= not((layer0_outputs(2527)) and (layer0_outputs(3694)));
    outputs(1977) <= (layer0_outputs(2576)) and not (layer0_outputs(338));
    outputs(1978) <= not(layer0_outputs(4166)) or (layer0_outputs(2765));
    outputs(1979) <= '1';
    outputs(1980) <= not((layer0_outputs(2999)) or (layer0_outputs(1342)));
    outputs(1981) <= not((layer0_outputs(4707)) or (layer0_outputs(1211)));
    outputs(1982) <= (layer0_outputs(970)) and not (layer0_outputs(2892));
    outputs(1983) <= not(layer0_outputs(556));
    outputs(1984) <= layer0_outputs(3811);
    outputs(1985) <= not(layer0_outputs(491));
    outputs(1986) <= not(layer0_outputs(483));
    outputs(1987) <= not(layer0_outputs(704));
    outputs(1988) <= not((layer0_outputs(1938)) xor (layer0_outputs(2229)));
    outputs(1989) <= (layer0_outputs(4468)) and not (layer0_outputs(4801));
    outputs(1990) <= (layer0_outputs(4427)) xor (layer0_outputs(4488));
    outputs(1991) <= (layer0_outputs(3095)) and not (layer0_outputs(3442));
    outputs(1992) <= not((layer0_outputs(3595)) xor (layer0_outputs(4249)));
    outputs(1993) <= not((layer0_outputs(1119)) and (layer0_outputs(1911)));
    outputs(1994) <= not(layer0_outputs(2868)) or (layer0_outputs(2763));
    outputs(1995) <= not((layer0_outputs(3563)) and (layer0_outputs(2994)));
    outputs(1996) <= layer0_outputs(4750);
    outputs(1997) <= not(layer0_outputs(2596));
    outputs(1998) <= not((layer0_outputs(4244)) xor (layer0_outputs(3282)));
    outputs(1999) <= (layer0_outputs(40)) and not (layer0_outputs(215));
    outputs(2000) <= (layer0_outputs(2352)) and not (layer0_outputs(1650));
    outputs(2001) <= not((layer0_outputs(835)) and (layer0_outputs(2948)));
    outputs(2002) <= (layer0_outputs(738)) xor (layer0_outputs(4422));
    outputs(2003) <= (layer0_outputs(4314)) and not (layer0_outputs(3595));
    outputs(2004) <= (layer0_outputs(3520)) xor (layer0_outputs(4150));
    outputs(2005) <= layer0_outputs(1480);
    outputs(2006) <= layer0_outputs(4272);
    outputs(2007) <= not((layer0_outputs(2377)) xor (layer0_outputs(1125)));
    outputs(2008) <= (layer0_outputs(3303)) and not (layer0_outputs(2952));
    outputs(2009) <= not((layer0_outputs(281)) and (layer0_outputs(1275)));
    outputs(2010) <= (layer0_outputs(3454)) and (layer0_outputs(1390));
    outputs(2011) <= (layer0_outputs(2427)) or (layer0_outputs(1496));
    outputs(2012) <= not(layer0_outputs(3477));
    outputs(2013) <= not((layer0_outputs(3396)) xor (layer0_outputs(1454)));
    outputs(2014) <= not(layer0_outputs(4362)) or (layer0_outputs(5072));
    outputs(2015) <= layer0_outputs(1478);
    outputs(2016) <= not(layer0_outputs(4117));
    outputs(2017) <= not((layer0_outputs(3829)) xor (layer0_outputs(385)));
    outputs(2018) <= (layer0_outputs(1685)) and not (layer0_outputs(1915));
    outputs(2019) <= layer0_outputs(3898);
    outputs(2020) <= (layer0_outputs(268)) or (layer0_outputs(3843));
    outputs(2021) <= not((layer0_outputs(1602)) xor (layer0_outputs(918)));
    outputs(2022) <= (layer0_outputs(1011)) and not (layer0_outputs(3051));
    outputs(2023) <= layer0_outputs(1708);
    outputs(2024) <= layer0_outputs(153);
    outputs(2025) <= layer0_outputs(4789);
    outputs(2026) <= layer0_outputs(1940);
    outputs(2027) <= layer0_outputs(2316);
    outputs(2028) <= not(layer0_outputs(1900));
    outputs(2029) <= not((layer0_outputs(340)) or (layer0_outputs(555)));
    outputs(2030) <= not(layer0_outputs(1515));
    outputs(2031) <= not((layer0_outputs(2699)) and (layer0_outputs(2578)));
    outputs(2032) <= not(layer0_outputs(4465));
    outputs(2033) <= not(layer0_outputs(1491));
    outputs(2034) <= not((layer0_outputs(728)) xor (layer0_outputs(4346)));
    outputs(2035) <= (layer0_outputs(4029)) and (layer0_outputs(5051));
    outputs(2036) <= (layer0_outputs(1954)) and (layer0_outputs(5003));
    outputs(2037) <= not(layer0_outputs(3504)) or (layer0_outputs(3608));
    outputs(2038) <= not(layer0_outputs(2240));
    outputs(2039) <= not(layer0_outputs(4203));
    outputs(2040) <= not((layer0_outputs(3006)) or (layer0_outputs(3868)));
    outputs(2041) <= not(layer0_outputs(2250));
    outputs(2042) <= layer0_outputs(3010);
    outputs(2043) <= '1';
    outputs(2044) <= (layer0_outputs(2955)) or (layer0_outputs(3464));
    outputs(2045) <= layer0_outputs(3440);
    outputs(2046) <= not(layer0_outputs(4199)) or (layer0_outputs(474));
    outputs(2047) <= (layer0_outputs(3281)) or (layer0_outputs(2188));
    outputs(2048) <= layer0_outputs(2013);
    outputs(2049) <= not(layer0_outputs(3891)) or (layer0_outputs(4157));
    outputs(2050) <= layer0_outputs(4178);
    outputs(2051) <= (layer0_outputs(1654)) and not (layer0_outputs(3337));
    outputs(2052) <= layer0_outputs(3662);
    outputs(2053) <= not((layer0_outputs(1978)) or (layer0_outputs(995)));
    outputs(2054) <= not(layer0_outputs(1524)) or (layer0_outputs(1864));
    outputs(2055) <= not((layer0_outputs(2794)) xor (layer0_outputs(2796)));
    outputs(2056) <= layer0_outputs(4816);
    outputs(2057) <= (layer0_outputs(436)) and not (layer0_outputs(3354));
    outputs(2058) <= layer0_outputs(2736);
    outputs(2059) <= not(layer0_outputs(791));
    outputs(2060) <= not((layer0_outputs(271)) or (layer0_outputs(4722)));
    outputs(2061) <= (layer0_outputs(4168)) and not (layer0_outputs(633));
    outputs(2062) <= not((layer0_outputs(1822)) xor (layer0_outputs(3090)));
    outputs(2063) <= (layer0_outputs(476)) and (layer0_outputs(449));
    outputs(2064) <= not((layer0_outputs(4026)) or (layer0_outputs(1242)));
    outputs(2065) <= not((layer0_outputs(4647)) xor (layer0_outputs(4737)));
    outputs(2066) <= not((layer0_outputs(4672)) and (layer0_outputs(1298)));
    outputs(2067) <= (layer0_outputs(3365)) and not (layer0_outputs(2383));
    outputs(2068) <= not(layer0_outputs(4231));
    outputs(2069) <= layer0_outputs(2187);
    outputs(2070) <= (layer0_outputs(4694)) and not (layer0_outputs(658));
    outputs(2071) <= (layer0_outputs(1494)) or (layer0_outputs(754));
    outputs(2072) <= not(layer0_outputs(546));
    outputs(2073) <= not(layer0_outputs(613)) or (layer0_outputs(3231));
    outputs(2074) <= (layer0_outputs(2916)) xor (layer0_outputs(500));
    outputs(2075) <= not((layer0_outputs(4782)) xor (layer0_outputs(1327)));
    outputs(2076) <= (layer0_outputs(4949)) and not (layer0_outputs(4069));
    outputs(2077) <= (layer0_outputs(3855)) xor (layer0_outputs(3535));
    outputs(2078) <= (layer0_outputs(1716)) and not (layer0_outputs(3353));
    outputs(2079) <= not(layer0_outputs(1811));
    outputs(2080) <= (layer0_outputs(2499)) xor (layer0_outputs(1351));
    outputs(2081) <= (layer0_outputs(4881)) and not (layer0_outputs(2677));
    outputs(2082) <= not(layer0_outputs(1410)) or (layer0_outputs(3527));
    outputs(2083) <= not(layer0_outputs(866));
    outputs(2084) <= not(layer0_outputs(4411));
    outputs(2085) <= layer0_outputs(671);
    outputs(2086) <= (layer0_outputs(277)) and (layer0_outputs(4718));
    outputs(2087) <= not((layer0_outputs(2406)) or (layer0_outputs(3131)));
    outputs(2088) <= not(layer0_outputs(3175));
    outputs(2089) <= layer0_outputs(2796);
    outputs(2090) <= not((layer0_outputs(3770)) and (layer0_outputs(3389)));
    outputs(2091) <= (layer0_outputs(2961)) and not (layer0_outputs(1378));
    outputs(2092) <= (layer0_outputs(2684)) and not (layer0_outputs(4861));
    outputs(2093) <= not(layer0_outputs(3133));
    outputs(2094) <= (layer0_outputs(635)) xor (layer0_outputs(2704));
    outputs(2095) <= not((layer0_outputs(225)) or (layer0_outputs(3862)));
    outputs(2096) <= (layer0_outputs(882)) and (layer0_outputs(4404));
    outputs(2097) <= (layer0_outputs(3863)) xor (layer0_outputs(4655));
    outputs(2098) <= not((layer0_outputs(2206)) or (layer0_outputs(2231)));
    outputs(2099) <= not(layer0_outputs(4887));
    outputs(2100) <= not(layer0_outputs(810));
    outputs(2101) <= (layer0_outputs(3363)) and not (layer0_outputs(473));
    outputs(2102) <= not(layer0_outputs(4098)) or (layer0_outputs(761));
    outputs(2103) <= layer0_outputs(530);
    outputs(2104) <= not(layer0_outputs(182));
    outputs(2105) <= layer0_outputs(2098);
    outputs(2106) <= layer0_outputs(1128);
    outputs(2107) <= not(layer0_outputs(1498));
    outputs(2108) <= (layer0_outputs(1982)) and not (layer0_outputs(201));
    outputs(2109) <= not(layer0_outputs(431));
    outputs(2110) <= (layer0_outputs(4266)) and not (layer0_outputs(2449));
    outputs(2111) <= not(layer0_outputs(3126));
    outputs(2112) <= (layer0_outputs(1907)) and (layer0_outputs(3443));
    outputs(2113) <= layer0_outputs(794);
    outputs(2114) <= (layer0_outputs(691)) and not (layer0_outputs(4494));
    outputs(2115) <= (layer0_outputs(171)) and (layer0_outputs(4915));
    outputs(2116) <= not((layer0_outputs(2452)) xor (layer0_outputs(4745)));
    outputs(2117) <= layer0_outputs(1121);
    outputs(2118) <= (layer0_outputs(1540)) and not (layer0_outputs(2735));
    outputs(2119) <= (layer0_outputs(1424)) and (layer0_outputs(3161));
    outputs(2120) <= (layer0_outputs(2341)) and not (layer0_outputs(4994));
    outputs(2121) <= layer0_outputs(1844);
    outputs(2122) <= not(layer0_outputs(4384)) or (layer0_outputs(5024));
    outputs(2123) <= layer0_outputs(3641);
    outputs(2124) <= (layer0_outputs(2511)) xor (layer0_outputs(2474));
    outputs(2125) <= layer0_outputs(3679);
    outputs(2126) <= (layer0_outputs(3713)) xor (layer0_outputs(4514));
    outputs(2127) <= not((layer0_outputs(4763)) xor (layer0_outputs(2)));
    outputs(2128) <= not(layer0_outputs(2795));
    outputs(2129) <= not(layer0_outputs(822));
    outputs(2130) <= layer0_outputs(2303);
    outputs(2131) <= (layer0_outputs(2112)) and not (layer0_outputs(3597));
    outputs(2132) <= not((layer0_outputs(459)) xor (layer0_outputs(4769)));
    outputs(2133) <= not((layer0_outputs(2691)) and (layer0_outputs(1813)));
    outputs(2134) <= layer0_outputs(4188);
    outputs(2135) <= layer0_outputs(5115);
    outputs(2136) <= layer0_outputs(4615);
    outputs(2137) <= (layer0_outputs(2232)) xor (layer0_outputs(1606));
    outputs(2138) <= layer0_outputs(1663);
    outputs(2139) <= (layer0_outputs(2088)) xor (layer0_outputs(394));
    outputs(2140) <= not((layer0_outputs(3870)) xor (layer0_outputs(990)));
    outputs(2141) <= layer0_outputs(1511);
    outputs(2142) <= (layer0_outputs(1394)) and not (layer0_outputs(2771));
    outputs(2143) <= not(layer0_outputs(2129));
    outputs(2144) <= not((layer0_outputs(4632)) xor (layer0_outputs(1979)));
    outputs(2145) <= layer0_outputs(4964);
    outputs(2146) <= (layer0_outputs(2591)) or (layer0_outputs(1567));
    outputs(2147) <= (layer0_outputs(1990)) and not (layer0_outputs(3316));
    outputs(2148) <= (layer0_outputs(15)) xor (layer0_outputs(1228));
    outputs(2149) <= (layer0_outputs(4583)) and (layer0_outputs(3017));
    outputs(2150) <= (layer0_outputs(3149)) and (layer0_outputs(3341));
    outputs(2151) <= (layer0_outputs(4895)) xor (layer0_outputs(1965));
    outputs(2152) <= (layer0_outputs(1244)) and (layer0_outputs(3478));
    outputs(2153) <= not((layer0_outputs(3093)) xor (layer0_outputs(3164)));
    outputs(2154) <= (layer0_outputs(4738)) and (layer0_outputs(4492));
    outputs(2155) <= not(layer0_outputs(1322)) or (layer0_outputs(419));
    outputs(2156) <= not((layer0_outputs(1996)) xor (layer0_outputs(5025)));
    outputs(2157) <= not(layer0_outputs(3934)) or (layer0_outputs(4821));
    outputs(2158) <= (layer0_outputs(3158)) xor (layer0_outputs(138));
    outputs(2159) <= (layer0_outputs(90)) and not (layer0_outputs(2639));
    outputs(2160) <= layer0_outputs(2662);
    outputs(2161) <= not((layer0_outputs(5076)) xor (layer0_outputs(1274)));
    outputs(2162) <= not((layer0_outputs(2997)) xor (layer0_outputs(2407)));
    outputs(2163) <= layer0_outputs(1849);
    outputs(2164) <= layer0_outputs(3953);
    outputs(2165) <= layer0_outputs(2857);
    outputs(2166) <= layer0_outputs(1781);
    outputs(2167) <= not((layer0_outputs(2296)) or (layer0_outputs(2041)));
    outputs(2168) <= layer0_outputs(2439);
    outputs(2169) <= not((layer0_outputs(3537)) xor (layer0_outputs(1995)));
    outputs(2170) <= (layer0_outputs(1554)) and not (layer0_outputs(1260));
    outputs(2171) <= not((layer0_outputs(3655)) and (layer0_outputs(3561)));
    outputs(2172) <= not((layer0_outputs(2783)) or (layer0_outputs(499)));
    outputs(2173) <= not(layer0_outputs(4412));
    outputs(2174) <= not(layer0_outputs(4154));
    outputs(2175) <= (layer0_outputs(1740)) and (layer0_outputs(4894));
    outputs(2176) <= not(layer0_outputs(3173)) or (layer0_outputs(3932));
    outputs(2177) <= not(layer0_outputs(1902));
    outputs(2178) <= (layer0_outputs(3563)) and not (layer0_outputs(575));
    outputs(2179) <= (layer0_outputs(266)) and not (layer0_outputs(2503));
    outputs(2180) <= not(layer0_outputs(162)) or (layer0_outputs(1484));
    outputs(2181) <= (layer0_outputs(4519)) or (layer0_outputs(1823));
    outputs(2182) <= not((layer0_outputs(1100)) xor (layer0_outputs(4354)));
    outputs(2183) <= not((layer0_outputs(2249)) and (layer0_outputs(655)));
    outputs(2184) <= layer0_outputs(3432);
    outputs(2185) <= not((layer0_outputs(1651)) xor (layer0_outputs(2963)));
    outputs(2186) <= not((layer0_outputs(2918)) xor (layer0_outputs(2820)));
    outputs(2187) <= (layer0_outputs(4855)) and not (layer0_outputs(2969));
    outputs(2188) <= layer0_outputs(445);
    outputs(2189) <= (layer0_outputs(4284)) and (layer0_outputs(4027));
    outputs(2190) <= not(layer0_outputs(3043));
    outputs(2191) <= layer0_outputs(5104);
    outputs(2192) <= not(layer0_outputs(4334));
    outputs(2193) <= layer0_outputs(3866);
    outputs(2194) <= not((layer0_outputs(1443)) and (layer0_outputs(2178)));
    outputs(2195) <= (layer0_outputs(2703)) and not (layer0_outputs(4942));
    outputs(2196) <= (layer0_outputs(1288)) and not (layer0_outputs(3086));
    outputs(2197) <= layer0_outputs(3431);
    outputs(2198) <= not(layer0_outputs(1685));
    outputs(2199) <= not(layer0_outputs(3494));
    outputs(2200) <= (layer0_outputs(923)) and not (layer0_outputs(4418));
    outputs(2201) <= layer0_outputs(3824);
    outputs(2202) <= (layer0_outputs(1110)) xor (layer0_outputs(4528));
    outputs(2203) <= (layer0_outputs(4725)) xor (layer0_outputs(2582));
    outputs(2204) <= not(layer0_outputs(3451));
    outputs(2205) <= not(layer0_outputs(926));
    outputs(2206) <= not(layer0_outputs(310));
    outputs(2207) <= layer0_outputs(2207);
    outputs(2208) <= (layer0_outputs(1960)) and not (layer0_outputs(1590));
    outputs(2209) <= not(layer0_outputs(5012));
    outputs(2210) <= layer0_outputs(4650);
    outputs(2211) <= not((layer0_outputs(3106)) xor (layer0_outputs(3575)));
    outputs(2212) <= not((layer0_outputs(3187)) or (layer0_outputs(3832)));
    outputs(2213) <= not((layer0_outputs(3125)) xor (layer0_outputs(1009)));
    outputs(2214) <= (layer0_outputs(1277)) and (layer0_outputs(1035));
    outputs(2215) <= not(layer0_outputs(1448));
    outputs(2216) <= (layer0_outputs(2283)) and (layer0_outputs(1825));
    outputs(2217) <= layer0_outputs(3457);
    outputs(2218) <= not((layer0_outputs(1733)) xor (layer0_outputs(4017)));
    outputs(2219) <= layer0_outputs(1174);
    outputs(2220) <= layer0_outputs(1024);
    outputs(2221) <= not((layer0_outputs(2467)) xor (layer0_outputs(3842)));
    outputs(2222) <= layer0_outputs(1611);
    outputs(2223) <= (layer0_outputs(471)) and (layer0_outputs(4978));
    outputs(2224) <= layer0_outputs(979);
    outputs(2225) <= not((layer0_outputs(546)) xor (layer0_outputs(3992)));
    outputs(2226) <= not((layer0_outputs(3515)) xor (layer0_outputs(3994)));
    outputs(2227) <= not(layer0_outputs(1465));
    outputs(2228) <= (layer0_outputs(1892)) and not (layer0_outputs(4544));
    outputs(2229) <= not((layer0_outputs(2204)) xor (layer0_outputs(3635)));
    outputs(2230) <= (layer0_outputs(4680)) and (layer0_outputs(1607));
    outputs(2231) <= layer0_outputs(596);
    outputs(2232) <= layer0_outputs(5064);
    outputs(2233) <= layer0_outputs(4281);
    outputs(2234) <= not((layer0_outputs(341)) xor (layer0_outputs(1397)));
    outputs(2235) <= not(layer0_outputs(479));
    outputs(2236) <= not(layer0_outputs(1347));
    outputs(2237) <= (layer0_outputs(5068)) xor (layer0_outputs(3867));
    outputs(2238) <= (layer0_outputs(2298)) and not (layer0_outputs(5001));
    outputs(2239) <= layer0_outputs(4000);
    outputs(2240) <= not(layer0_outputs(3825));
    outputs(2241) <= (layer0_outputs(1922)) and (layer0_outputs(4572));
    outputs(2242) <= not(layer0_outputs(3566));
    outputs(2243) <= (layer0_outputs(3517)) and (layer0_outputs(979));
    outputs(2244) <= not((layer0_outputs(1220)) xor (layer0_outputs(1160)));
    outputs(2245) <= layer0_outputs(2547);
    outputs(2246) <= not((layer0_outputs(2708)) xor (layer0_outputs(4730)));
    outputs(2247) <= (layer0_outputs(2156)) xor (layer0_outputs(2497));
    outputs(2248) <= (layer0_outputs(1697)) xor (layer0_outputs(2093));
    outputs(2249) <= not(layer0_outputs(3946));
    outputs(2250) <= '0';
    outputs(2251) <= (layer0_outputs(1793)) xor (layer0_outputs(2131));
    outputs(2252) <= (layer0_outputs(4971)) xor (layer0_outputs(2509));
    outputs(2253) <= layer0_outputs(4214);
    outputs(2254) <= not((layer0_outputs(537)) xor (layer0_outputs(161)));
    outputs(2255) <= not((layer0_outputs(1317)) or (layer0_outputs(87)));
    outputs(2256) <= (layer0_outputs(1262)) xor (layer0_outputs(2813));
    outputs(2257) <= (layer0_outputs(4212)) and (layer0_outputs(2550));
    outputs(2258) <= layer0_outputs(1245);
    outputs(2259) <= not(layer0_outputs(4817));
    outputs(2260) <= not((layer0_outputs(3470)) or (layer0_outputs(2312)));
    outputs(2261) <= (layer0_outputs(3317)) xor (layer0_outputs(2601));
    outputs(2262) <= not((layer0_outputs(2854)) xor (layer0_outputs(4104)));
    outputs(2263) <= not(layer0_outputs(1287));
    outputs(2264) <= not(layer0_outputs(3787)) or (layer0_outputs(1953));
    outputs(2265) <= not(layer0_outputs(2110));
    outputs(2266) <= not((layer0_outputs(1815)) xor (layer0_outputs(4393)));
    outputs(2267) <= (layer0_outputs(1573)) and (layer0_outputs(1516));
    outputs(2268) <= not(layer0_outputs(4513));
    outputs(2269) <= not((layer0_outputs(4297)) or (layer0_outputs(1146)));
    outputs(2270) <= not((layer0_outputs(714)) and (layer0_outputs(1753)));
    outputs(2271) <= not(layer0_outputs(1349));
    outputs(2272) <= (layer0_outputs(89)) and not (layer0_outputs(1757));
    outputs(2273) <= not((layer0_outputs(4258)) xor (layer0_outputs(3649)));
    outputs(2274) <= (layer0_outputs(2495)) and (layer0_outputs(874));
    outputs(2275) <= not(layer0_outputs(2959));
    outputs(2276) <= not((layer0_outputs(3221)) or (layer0_outputs(994)));
    outputs(2277) <= not(layer0_outputs(2707));
    outputs(2278) <= (layer0_outputs(129)) xor (layer0_outputs(3867));
    outputs(2279) <= not(layer0_outputs(4961));
    outputs(2280) <= layer0_outputs(3668);
    outputs(2281) <= not(layer0_outputs(3898));
    outputs(2282) <= (layer0_outputs(4813)) and not (layer0_outputs(4099));
    outputs(2283) <= not(layer0_outputs(5033));
    outputs(2284) <= (layer0_outputs(2874)) and not (layer0_outputs(218));
    outputs(2285) <= (layer0_outputs(4743)) and (layer0_outputs(4322));
    outputs(2286) <= (layer0_outputs(4761)) and (layer0_outputs(195));
    outputs(2287) <= not((layer0_outputs(4213)) or (layer0_outputs(1804)));
    outputs(2288) <= layer0_outputs(4100);
    outputs(2289) <= '1';
    outputs(2290) <= (layer0_outputs(3621)) and not (layer0_outputs(991));
    outputs(2291) <= not((layer0_outputs(920)) xor (layer0_outputs(1404)));
    outputs(2292) <= layer0_outputs(4918);
    outputs(2293) <= (layer0_outputs(233)) and not (layer0_outputs(830));
    outputs(2294) <= layer0_outputs(1726);
    outputs(2295) <= layer0_outputs(1700);
    outputs(2296) <= not((layer0_outputs(616)) xor (layer0_outputs(2771)));
    outputs(2297) <= not(layer0_outputs(191));
    outputs(2298) <= layer0_outputs(4770);
    outputs(2299) <= layer0_outputs(1047);
    outputs(2300) <= (layer0_outputs(2574)) xor (layer0_outputs(4848));
    outputs(2301) <= not(layer0_outputs(1497));
    outputs(2302) <= layer0_outputs(4583);
    outputs(2303) <= layer0_outputs(1706);
    outputs(2304) <= not(layer0_outputs(4716)) or (layer0_outputs(3198));
    outputs(2305) <= (layer0_outputs(1527)) and not (layer0_outputs(1255));
    outputs(2306) <= (layer0_outputs(84)) and not (layer0_outputs(1217));
    outputs(2307) <= not((layer0_outputs(859)) xor (layer0_outputs(2742)));
    outputs(2308) <= not(layer0_outputs(1282));
    outputs(2309) <= (layer0_outputs(4500)) and (layer0_outputs(4142));
    outputs(2310) <= not(layer0_outputs(4998)) or (layer0_outputs(2413));
    outputs(2311) <= not((layer0_outputs(849)) xor (layer0_outputs(786)));
    outputs(2312) <= layer0_outputs(1490);
    outputs(2313) <= (layer0_outputs(2726)) and (layer0_outputs(2681));
    outputs(2314) <= (layer0_outputs(3581)) xor (layer0_outputs(4130));
    outputs(2315) <= not(layer0_outputs(3337));
    outputs(2316) <= not(layer0_outputs(3778));
    outputs(2317) <= not(layer0_outputs(3101));
    outputs(2318) <= (layer0_outputs(4883)) and not (layer0_outputs(4611));
    outputs(2319) <= (layer0_outputs(1886)) and not (layer0_outputs(3971));
    outputs(2320) <= (layer0_outputs(2646)) and (layer0_outputs(4034));
    outputs(2321) <= not((layer0_outputs(441)) or (layer0_outputs(3538)));
    outputs(2322) <= layer0_outputs(1399);
    outputs(2323) <= not((layer0_outputs(3369)) xor (layer0_outputs(3026)));
    outputs(2324) <= layer0_outputs(2925);
    outputs(2325) <= not((layer0_outputs(3670)) or (layer0_outputs(537)));
    outputs(2326) <= layer0_outputs(771);
    outputs(2327) <= (layer0_outputs(1031)) xor (layer0_outputs(3112));
    outputs(2328) <= (layer0_outputs(3571)) and not (layer0_outputs(4445));
    outputs(2329) <= not(layer0_outputs(1021));
    outputs(2330) <= not(layer0_outputs(1866));
    outputs(2331) <= (layer0_outputs(2580)) and not (layer0_outputs(1341));
    outputs(2332) <= layer0_outputs(353);
    outputs(2333) <= (layer0_outputs(2991)) and not (layer0_outputs(1962));
    outputs(2334) <= layer0_outputs(1007);
    outputs(2335) <= layer0_outputs(4396);
    outputs(2336) <= layer0_outputs(4200);
    outputs(2337) <= layer0_outputs(839);
    outputs(2338) <= not(layer0_outputs(4481));
    outputs(2339) <= layer0_outputs(1960);
    outputs(2340) <= layer0_outputs(1617);
    outputs(2341) <= not(layer0_outputs(933));
    outputs(2342) <= not((layer0_outputs(2904)) or (layer0_outputs(2342)));
    outputs(2343) <= not(layer0_outputs(2727));
    outputs(2344) <= not((layer0_outputs(4518)) and (layer0_outputs(491)));
    outputs(2345) <= not(layer0_outputs(4804));
    outputs(2346) <= layer0_outputs(1000);
    outputs(2347) <= not((layer0_outputs(2712)) xor (layer0_outputs(826)));
    outputs(2348) <= (layer0_outputs(2395)) xor (layer0_outputs(4138));
    outputs(2349) <= not((layer0_outputs(3234)) xor (layer0_outputs(2900)));
    outputs(2350) <= not((layer0_outputs(49)) xor (layer0_outputs(545)));
    outputs(2351) <= (layer0_outputs(2808)) xor (layer0_outputs(2981));
    outputs(2352) <= (layer0_outputs(855)) or (layer0_outputs(3322));
    outputs(2353) <= layer0_outputs(1846);
    outputs(2354) <= not(layer0_outputs(1030));
    outputs(2355) <= not(layer0_outputs(4507));
    outputs(2356) <= not((layer0_outputs(3753)) xor (layer0_outputs(1157)));
    outputs(2357) <= (layer0_outputs(2032)) and not (layer0_outputs(4368));
    outputs(2358) <= (layer0_outputs(3560)) and not (layer0_outputs(1728));
    outputs(2359) <= layer0_outputs(1575);
    outputs(2360) <= not((layer0_outputs(2223)) xor (layer0_outputs(4680)));
    outputs(2361) <= '0';
    outputs(2362) <= not(layer0_outputs(3174));
    outputs(2363) <= not((layer0_outputs(3506)) xor (layer0_outputs(4844)));
    outputs(2364) <= (layer0_outputs(281)) and not (layer0_outputs(3798));
    outputs(2365) <= (layer0_outputs(609)) and not (layer0_outputs(261));
    outputs(2366) <= not(layer0_outputs(1001));
    outputs(2367) <= not((layer0_outputs(2684)) or (layer0_outputs(809)));
    outputs(2368) <= not(layer0_outputs(3280));
    outputs(2369) <= (layer0_outputs(2699)) and not (layer0_outputs(1471));
    outputs(2370) <= (layer0_outputs(1047)) and not (layer0_outputs(965));
    outputs(2371) <= not((layer0_outputs(5012)) or (layer0_outputs(1748)));
    outputs(2372) <= not((layer0_outputs(3329)) xor (layer0_outputs(2339)));
    outputs(2373) <= layer0_outputs(2056);
    outputs(2374) <= not(layer0_outputs(3979)) or (layer0_outputs(1660));
    outputs(2375) <= not((layer0_outputs(951)) and (layer0_outputs(549)));
    outputs(2376) <= layer0_outputs(1550);
    outputs(2377) <= layer0_outputs(5020);
    outputs(2378) <= not((layer0_outputs(4667)) xor (layer0_outputs(2831)));
    outputs(2379) <= layer0_outputs(239);
    outputs(2380) <= not(layer0_outputs(2162));
    outputs(2381) <= not((layer0_outputs(937)) xor (layer0_outputs(843)));
    outputs(2382) <= layer0_outputs(1646);
    outputs(2383) <= layer0_outputs(1198);
    outputs(2384) <= (layer0_outputs(1678)) and not (layer0_outputs(2321));
    outputs(2385) <= (layer0_outputs(2069)) xor (layer0_outputs(4646));
    outputs(2386) <= not((layer0_outputs(1707)) xor (layer0_outputs(28)));
    outputs(2387) <= not((layer0_outputs(4609)) xor (layer0_outputs(1951)));
    outputs(2388) <= (layer0_outputs(2030)) and not (layer0_outputs(392));
    outputs(2389) <= not((layer0_outputs(4730)) xor (layer0_outputs(1836)));
    outputs(2390) <= not((layer0_outputs(591)) and (layer0_outputs(832)));
    outputs(2391) <= (layer0_outputs(4743)) and (layer0_outputs(3837));
    outputs(2392) <= not(layer0_outputs(1193)) or (layer0_outputs(1156));
    outputs(2393) <= (layer0_outputs(5048)) and not (layer0_outputs(123));
    outputs(2394) <= (layer0_outputs(4558)) and not (layer0_outputs(641));
    outputs(2395) <= layer0_outputs(2409);
    outputs(2396) <= not((layer0_outputs(920)) xor (layer0_outputs(4330)));
    outputs(2397) <= layer0_outputs(1406);
    outputs(2398) <= layer0_outputs(1726);
    outputs(2399) <= not(layer0_outputs(1259));
    outputs(2400) <= not((layer0_outputs(630)) xor (layer0_outputs(48)));
    outputs(2401) <= (layer0_outputs(734)) xor (layer0_outputs(5022));
    outputs(2402) <= not(layer0_outputs(5054));
    outputs(2403) <= not(layer0_outputs(2291));
    outputs(2404) <= (layer0_outputs(1445)) and not (layer0_outputs(2960));
    outputs(2405) <= layer0_outputs(2320);
    outputs(2406) <= layer0_outputs(1398);
    outputs(2407) <= layer0_outputs(4109);
    outputs(2408) <= (layer0_outputs(2040)) xor (layer0_outputs(701));
    outputs(2409) <= '1';
    outputs(2410) <= not((layer0_outputs(3685)) or (layer0_outputs(2561)));
    outputs(2411) <= (layer0_outputs(4014)) xor (layer0_outputs(1935));
    outputs(2412) <= (layer0_outputs(2197)) and not (layer0_outputs(3277));
    outputs(2413) <= (layer0_outputs(355)) and not (layer0_outputs(5081));
    outputs(2414) <= not((layer0_outputs(3441)) or (layer0_outputs(1707)));
    outputs(2415) <= layer0_outputs(1367);
    outputs(2416) <= not((layer0_outputs(5026)) xor (layer0_outputs(3156)));
    outputs(2417) <= (layer0_outputs(4958)) and not (layer0_outputs(1409));
    outputs(2418) <= (layer0_outputs(1017)) and not (layer0_outputs(2127));
    outputs(2419) <= (layer0_outputs(4593)) and (layer0_outputs(710));
    outputs(2420) <= not(layer0_outputs(469));
    outputs(2421) <= (layer0_outputs(4447)) xor (layer0_outputs(3579));
    outputs(2422) <= (layer0_outputs(304)) and not (layer0_outputs(4201));
    outputs(2423) <= not((layer0_outputs(2089)) or (layer0_outputs(1640)));
    outputs(2424) <= layer0_outputs(260);
    outputs(2425) <= (layer0_outputs(3729)) xor (layer0_outputs(1826));
    outputs(2426) <= (layer0_outputs(2083)) xor (layer0_outputs(11));
    outputs(2427) <= layer0_outputs(183);
    outputs(2428) <= not((layer0_outputs(1260)) or (layer0_outputs(3238)));
    outputs(2429) <= not((layer0_outputs(835)) or (layer0_outputs(1334)));
    outputs(2430) <= (layer0_outputs(2389)) and (layer0_outputs(2446));
    outputs(2431) <= layer0_outputs(2012);
    outputs(2432) <= layer0_outputs(2297);
    outputs(2433) <= (layer0_outputs(1313)) or (layer0_outputs(2203));
    outputs(2434) <= (layer0_outputs(3858)) xor (layer0_outputs(5024));
    outputs(2435) <= (layer0_outputs(811)) and not (layer0_outputs(1521));
    outputs(2436) <= not(layer0_outputs(4941));
    outputs(2437) <= (layer0_outputs(4878)) or (layer0_outputs(462));
    outputs(2438) <= (layer0_outputs(3096)) and (layer0_outputs(1393));
    outputs(2439) <= (layer0_outputs(3138)) and (layer0_outputs(3839));
    outputs(2440) <= not((layer0_outputs(267)) and (layer0_outputs(2637)));
    outputs(2441) <= not((layer0_outputs(4729)) xor (layer0_outputs(3021)));
    outputs(2442) <= not((layer0_outputs(4753)) or (layer0_outputs(1702)));
    outputs(2443) <= not(layer0_outputs(3492)) or (layer0_outputs(4420));
    outputs(2444) <= not(layer0_outputs(1820));
    outputs(2445) <= not(layer0_outputs(610));
    outputs(2446) <= not((layer0_outputs(1589)) or (layer0_outputs(747)));
    outputs(2447) <= not(layer0_outputs(2332));
    outputs(2448) <= not(layer0_outputs(1339));
    outputs(2449) <= not(layer0_outputs(2157));
    outputs(2450) <= not(layer0_outputs(2027));
    outputs(2451) <= (layer0_outputs(2315)) and not (layer0_outputs(2488));
    outputs(2452) <= (layer0_outputs(5065)) xor (layer0_outputs(3136));
    outputs(2453) <= (layer0_outputs(5030)) and not (layer0_outputs(3510));
    outputs(2454) <= (layer0_outputs(3357)) and not (layer0_outputs(4385));
    outputs(2455) <= (layer0_outputs(3115)) and not (layer0_outputs(67));
    outputs(2456) <= not(layer0_outputs(1029));
    outputs(2457) <= (layer0_outputs(787)) xor (layer0_outputs(4547));
    outputs(2458) <= (layer0_outputs(39)) and not (layer0_outputs(3332));
    outputs(2459) <= (layer0_outputs(4678)) or (layer0_outputs(2262));
    outputs(2460) <= (layer0_outputs(4882)) and not (layer0_outputs(486));
    outputs(2461) <= layer0_outputs(678);
    outputs(2462) <= not(layer0_outputs(2899));
    outputs(2463) <= (layer0_outputs(1101)) xor (layer0_outputs(1880));
    outputs(2464) <= not((layer0_outputs(1247)) or (layer0_outputs(3702)));
    outputs(2465) <= layer0_outputs(690);
    outputs(2466) <= (layer0_outputs(1512)) xor (layer0_outputs(1203));
    outputs(2467) <= not(layer0_outputs(3118));
    outputs(2468) <= not(layer0_outputs(3693)) or (layer0_outputs(2330));
    outputs(2469) <= not((layer0_outputs(3958)) and (layer0_outputs(4061)));
    outputs(2470) <= not(layer0_outputs(3390));
    outputs(2471) <= layer0_outputs(2521);
    outputs(2472) <= (layer0_outputs(4802)) and not (layer0_outputs(1761));
    outputs(2473) <= not((layer0_outputs(1360)) and (layer0_outputs(2968)));
    outputs(2474) <= layer0_outputs(3593);
    outputs(2475) <= (layer0_outputs(1438)) and (layer0_outputs(928));
    outputs(2476) <= layer0_outputs(5103);
    outputs(2477) <= (layer0_outputs(171)) xor (layer0_outputs(1440));
    outputs(2478) <= not((layer0_outputs(4919)) xor (layer0_outputs(3305)));
    outputs(2479) <= not(layer0_outputs(4143)) or (layer0_outputs(3681));
    outputs(2480) <= not((layer0_outputs(4457)) xor (layer0_outputs(2776)));
    outputs(2481) <= not((layer0_outputs(4124)) or (layer0_outputs(3905)));
    outputs(2482) <= layer0_outputs(2767);
    outputs(2483) <= (layer0_outputs(4896)) and not (layer0_outputs(3674));
    outputs(2484) <= (layer0_outputs(631)) and not (layer0_outputs(160));
    outputs(2485) <= not(layer0_outputs(3981));
    outputs(2486) <= (layer0_outputs(2956)) and not (layer0_outputs(4797));
    outputs(2487) <= layer0_outputs(4060);
    outputs(2488) <= layer0_outputs(2762);
    outputs(2489) <= (layer0_outputs(3134)) and not (layer0_outputs(4156));
    outputs(2490) <= (layer0_outputs(4321)) and not (layer0_outputs(2617));
    outputs(2491) <= (layer0_outputs(1386)) and not (layer0_outputs(2148));
    outputs(2492) <= not(layer0_outputs(2696));
    outputs(2493) <= not((layer0_outputs(69)) or (layer0_outputs(2818)));
    outputs(2494) <= '0';
    outputs(2495) <= (layer0_outputs(2977)) and (layer0_outputs(2097));
    outputs(2496) <= (layer0_outputs(2120)) and (layer0_outputs(3387));
    outputs(2497) <= (layer0_outputs(2030)) and (layer0_outputs(4872));
    outputs(2498) <= not((layer0_outputs(3750)) or (layer0_outputs(5084)));
    outputs(2499) <= layer0_outputs(4234);
    outputs(2500) <= (layer0_outputs(427)) xor (layer0_outputs(2851));
    outputs(2501) <= not(layer0_outputs(2698));
    outputs(2502) <= '0';
    outputs(2503) <= (layer0_outputs(932)) xor (layer0_outputs(2251));
    outputs(2504) <= layer0_outputs(2063);
    outputs(2505) <= layer0_outputs(4836);
    outputs(2506) <= not(layer0_outputs(4528));
    outputs(2507) <= not(layer0_outputs(4952));
    outputs(2508) <= not((layer0_outputs(4935)) xor (layer0_outputs(3131)));
    outputs(2509) <= layer0_outputs(3945);
    outputs(2510) <= not((layer0_outputs(3931)) xor (layer0_outputs(1458)));
    outputs(2511) <= (layer0_outputs(732)) and not (layer0_outputs(22));
    outputs(2512) <= (layer0_outputs(4186)) xor (layer0_outputs(3760));
    outputs(2513) <= layer0_outputs(4211);
    outputs(2514) <= (layer0_outputs(1851)) and not (layer0_outputs(2891));
    outputs(2515) <= not((layer0_outputs(4684)) xor (layer0_outputs(2149)));
    outputs(2516) <= (layer0_outputs(4396)) and not (layer0_outputs(2512));
    outputs(2517) <= layer0_outputs(4237);
    outputs(2518) <= not((layer0_outputs(2632)) xor (layer0_outputs(509)));
    outputs(2519) <= not(layer0_outputs(5042));
    outputs(2520) <= not(layer0_outputs(2768));
    outputs(2521) <= not(layer0_outputs(3770));
    outputs(2522) <= layer0_outputs(3258);
    outputs(2523) <= not((layer0_outputs(4440)) xor (layer0_outputs(727)));
    outputs(2524) <= (layer0_outputs(1226)) xor (layer0_outputs(1144));
    outputs(2525) <= not(layer0_outputs(3638));
    outputs(2526) <= (layer0_outputs(2139)) xor (layer0_outputs(3576));
    outputs(2527) <= not((layer0_outputs(3515)) xor (layer0_outputs(514)));
    outputs(2528) <= not(layer0_outputs(4016));
    outputs(2529) <= not((layer0_outputs(1197)) xor (layer0_outputs(1185)));
    outputs(2530) <= layer0_outputs(3022);
    outputs(2531) <= not((layer0_outputs(2045)) and (layer0_outputs(4786)));
    outputs(2532) <= (layer0_outputs(4108)) and not (layer0_outputs(1448));
    outputs(2533) <= (layer0_outputs(3792)) and (layer0_outputs(2817));
    outputs(2534) <= not(layer0_outputs(3280));
    outputs(2535) <= not(layer0_outputs(1562));
    outputs(2536) <= layer0_outputs(1972);
    outputs(2537) <= (layer0_outputs(1528)) and not (layer0_outputs(2471));
    outputs(2538) <= not(layer0_outputs(3020));
    outputs(2539) <= layer0_outputs(743);
    outputs(2540) <= (layer0_outputs(3288)) and not (layer0_outputs(3927));
    outputs(2541) <= not((layer0_outputs(1899)) xor (layer0_outputs(3505)));
    outputs(2542) <= layer0_outputs(4043);
    outputs(2543) <= layer0_outputs(366);
    outputs(2544) <= (layer0_outputs(3837)) xor (layer0_outputs(1526));
    outputs(2545) <= not(layer0_outputs(1447));
    outputs(2546) <= not(layer0_outputs(4574));
    outputs(2547) <= not((layer0_outputs(3135)) and (layer0_outputs(1218)));
    outputs(2548) <= layer0_outputs(956);
    outputs(2549) <= (layer0_outputs(1747)) and not (layer0_outputs(3265));
    outputs(2550) <= (layer0_outputs(41)) xor (layer0_outputs(3581));
    outputs(2551) <= not((layer0_outputs(3385)) xor (layer0_outputs(579)));
    outputs(2552) <= '0';
    outputs(2553) <= not((layer0_outputs(3167)) xor (layer0_outputs(3057)));
    outputs(2554) <= not((layer0_outputs(126)) or (layer0_outputs(4962)));
    outputs(2555) <= not(layer0_outputs(229));
    outputs(2556) <= not(layer0_outputs(4225));
    outputs(2557) <= (layer0_outputs(4640)) xor (layer0_outputs(3620));
    outputs(2558) <= layer0_outputs(4341);
    outputs(2559) <= (layer0_outputs(3632)) and (layer0_outputs(227));
    outputs(2560) <= (layer0_outputs(3083)) or (layer0_outputs(545));
    outputs(2561) <= (layer0_outputs(3484)) and not (layer0_outputs(1185));
    outputs(2562) <= not((layer0_outputs(4733)) xor (layer0_outputs(1705)));
    outputs(2563) <= layer0_outputs(4627);
    outputs(2564) <= not((layer0_outputs(621)) xor (layer0_outputs(1928)));
    outputs(2565) <= not((layer0_outputs(4177)) and (layer0_outputs(4130)));
    outputs(2566) <= (layer0_outputs(4105)) xor (layer0_outputs(68));
    outputs(2567) <= not((layer0_outputs(940)) xor (layer0_outputs(443)));
    outputs(2568) <= layer0_outputs(208);
    outputs(2569) <= not(layer0_outputs(1004));
    outputs(2570) <= layer0_outputs(4428);
    outputs(2571) <= layer0_outputs(3925);
    outputs(2572) <= not((layer0_outputs(4603)) or (layer0_outputs(3531)));
    outputs(2573) <= layer0_outputs(4005);
    outputs(2574) <= layer0_outputs(3150);
    outputs(2575) <= layer0_outputs(3669);
    outputs(2576) <= not(layer0_outputs(2288));
    outputs(2577) <= layer0_outputs(4178);
    outputs(2578) <= not((layer0_outputs(626)) or (layer0_outputs(2729)));
    outputs(2579) <= (layer0_outputs(4683)) and not (layer0_outputs(5010));
    outputs(2580) <= not((layer0_outputs(1634)) or (layer0_outputs(3358)));
    outputs(2581) <= layer0_outputs(3087);
    outputs(2582) <= not(layer0_outputs(958));
    outputs(2583) <= not((layer0_outputs(2325)) or (layer0_outputs(904)));
    outputs(2584) <= (layer0_outputs(3968)) and not (layer0_outputs(4241));
    outputs(2585) <= not((layer0_outputs(2103)) or (layer0_outputs(508)));
    outputs(2586) <= (layer0_outputs(4165)) and (layer0_outputs(4768));
    outputs(2587) <= layer0_outputs(3260);
    outputs(2588) <= (layer0_outputs(3576)) and (layer0_outputs(583));
    outputs(2589) <= not(layer0_outputs(3653)) or (layer0_outputs(2344));
    outputs(2590) <= not(layer0_outputs(310)) or (layer0_outputs(2134));
    outputs(2591) <= not(layer0_outputs(2242));
    outputs(2592) <= (layer0_outputs(2534)) and (layer0_outputs(2324));
    outputs(2593) <= not(layer0_outputs(349));
    outputs(2594) <= not(layer0_outputs(1532));
    outputs(2595) <= not(layer0_outputs(360));
    outputs(2596) <= layer0_outputs(3503);
    outputs(2597) <= not((layer0_outputs(1609)) xor (layer0_outputs(4342)));
    outputs(2598) <= not((layer0_outputs(1898)) xor (layer0_outputs(233)));
    outputs(2599) <= (layer0_outputs(1025)) and not (layer0_outputs(4127));
    outputs(2600) <= not(layer0_outputs(1378));
    outputs(2601) <= (layer0_outputs(3697)) and not (layer0_outputs(254));
    outputs(2602) <= layer0_outputs(3182);
    outputs(2603) <= layer0_outputs(1904);
    outputs(2604) <= not(layer0_outputs(1088));
    outputs(2605) <= not(layer0_outputs(3990));
    outputs(2606) <= not((layer0_outputs(3293)) xor (layer0_outputs(4092)));
    outputs(2607) <= not(layer0_outputs(926));
    outputs(2608) <= not(layer0_outputs(598));
    outputs(2609) <= not(layer0_outputs(783)) or (layer0_outputs(3568));
    outputs(2610) <= not(layer0_outputs(1600));
    outputs(2611) <= not((layer0_outputs(3189)) xor (layer0_outputs(529)));
    outputs(2612) <= not((layer0_outputs(2838)) or (layer0_outputs(503)));
    outputs(2613) <= not((layer0_outputs(79)) and (layer0_outputs(1447)));
    outputs(2614) <= layer0_outputs(4004);
    outputs(2615) <= not(layer0_outputs(2345));
    outputs(2616) <= (layer0_outputs(4261)) and not (layer0_outputs(4197));
    outputs(2617) <= not(layer0_outputs(2320)) or (layer0_outputs(1756));
    outputs(2618) <= (layer0_outputs(4811)) xor (layer0_outputs(1468));
    outputs(2619) <= (layer0_outputs(620)) or (layer0_outputs(2273));
    outputs(2620) <= not(layer0_outputs(1283)) or (layer0_outputs(4937));
    outputs(2621) <= not(layer0_outputs(3104));
    outputs(2622) <= not((layer0_outputs(1803)) xor (layer0_outputs(3176)));
    outputs(2623) <= (layer0_outputs(2697)) or (layer0_outputs(1587));
    outputs(2624) <= not(layer0_outputs(57)) or (layer0_outputs(2480));
    outputs(2625) <= not(layer0_outputs(1425));
    outputs(2626) <= not((layer0_outputs(385)) xor (layer0_outputs(520)));
    outputs(2627) <= (layer0_outputs(4985)) and not (layer0_outputs(2347));
    outputs(2628) <= not((layer0_outputs(471)) xor (layer0_outputs(4599)));
    outputs(2629) <= (layer0_outputs(1816)) and (layer0_outputs(1906));
    outputs(2630) <= not(layer0_outputs(3457));
    outputs(2631) <= (layer0_outputs(3322)) or (layer0_outputs(1021));
    outputs(2632) <= not((layer0_outputs(3296)) or (layer0_outputs(414)));
    outputs(2633) <= (layer0_outputs(1411)) xor (layer0_outputs(3143));
    outputs(2634) <= not((layer0_outputs(24)) or (layer0_outputs(2738)));
    outputs(2635) <= not((layer0_outputs(3540)) xor (layer0_outputs(4225)));
    outputs(2636) <= not(layer0_outputs(3997)) or (layer0_outputs(1346));
    outputs(2637) <= not((layer0_outputs(737)) xor (layer0_outputs(1879)));
    outputs(2638) <= not((layer0_outputs(4491)) xor (layer0_outputs(1478)));
    outputs(2639) <= not(layer0_outputs(4315));
    outputs(2640) <= not(layer0_outputs(47));
    outputs(2641) <= layer0_outputs(2929);
    outputs(2642) <= not(layer0_outputs(262)) or (layer0_outputs(2322));
    outputs(2643) <= (layer0_outputs(1636)) and (layer0_outputs(2357));
    outputs(2644) <= '0';
    outputs(2645) <= not(layer0_outputs(3745)) or (layer0_outputs(1131));
    outputs(2646) <= not(layer0_outputs(1789)) or (layer0_outputs(4044));
    outputs(2647) <= (layer0_outputs(234)) and not (layer0_outputs(2967));
    outputs(2648) <= (layer0_outputs(401)) xor (layer0_outputs(2780));
    outputs(2649) <= not(layer0_outputs(2435));
    outputs(2650) <= not(layer0_outputs(3502)) or (layer0_outputs(3726));
    outputs(2651) <= layer0_outputs(2781);
    outputs(2652) <= '1';
    outputs(2653) <= layer0_outputs(1208);
    outputs(2654) <= not((layer0_outputs(4684)) xor (layer0_outputs(2114)));
    outputs(2655) <= not((layer0_outputs(139)) or (layer0_outputs(4778)));
    outputs(2656) <= not((layer0_outputs(4125)) xor (layer0_outputs(880)));
    outputs(2657) <= layer0_outputs(442);
    outputs(2658) <= layer0_outputs(1709);
    outputs(2659) <= layer0_outputs(3034);
    outputs(2660) <= (layer0_outputs(4862)) and (layer0_outputs(3973));
    outputs(2661) <= layer0_outputs(1134);
    outputs(2662) <= not(layer0_outputs(3041)) or (layer0_outputs(2408));
    outputs(2663) <= layer0_outputs(4536);
    outputs(2664) <= not(layer0_outputs(4912));
    outputs(2665) <= layer0_outputs(3881);
    outputs(2666) <= not(layer0_outputs(1206));
    outputs(2667) <= not((layer0_outputs(4024)) or (layer0_outputs(563)));
    outputs(2668) <= not((layer0_outputs(4678)) and (layer0_outputs(1111)));
    outputs(2669) <= not(layer0_outputs(1184)) or (layer0_outputs(2668));
    outputs(2670) <= layer0_outputs(4727);
    outputs(2671) <= layer0_outputs(1149);
    outputs(2672) <= not(layer0_outputs(2937));
    outputs(2673) <= layer0_outputs(3682);
    outputs(2674) <= not((layer0_outputs(1567)) or (layer0_outputs(5007)));
    outputs(2675) <= (layer0_outputs(1257)) and not (layer0_outputs(3883));
    outputs(2676) <= (layer0_outputs(2842)) xor (layer0_outputs(4487));
    outputs(2677) <= layer0_outputs(4698);
    outputs(2678) <= (layer0_outputs(4478)) and (layer0_outputs(1568));
    outputs(2679) <= (layer0_outputs(3129)) and (layer0_outputs(4974));
    outputs(2680) <= (layer0_outputs(2617)) xor (layer0_outputs(4990));
    outputs(2681) <= (layer0_outputs(4214)) and not (layer0_outputs(2732));
    outputs(2682) <= (layer0_outputs(2098)) and not (layer0_outputs(5009));
    outputs(2683) <= not(layer0_outputs(101));
    outputs(2684) <= not(layer0_outputs(1312));
    outputs(2685) <= (layer0_outputs(4261)) xor (layer0_outputs(3358));
    outputs(2686) <= not((layer0_outputs(3235)) and (layer0_outputs(4959)));
    outputs(2687) <= not((layer0_outputs(306)) or (layer0_outputs(2586)));
    outputs(2688) <= not(layer0_outputs(1225));
    outputs(2689) <= (layer0_outputs(4756)) and not (layer0_outputs(4563));
    outputs(2690) <= layer0_outputs(3264);
    outputs(2691) <= not(layer0_outputs(1224)) or (layer0_outputs(3756));
    outputs(2692) <= (layer0_outputs(1426)) and (layer0_outputs(3134));
    outputs(2693) <= (layer0_outputs(1235)) or (layer0_outputs(3749));
    outputs(2694) <= not(layer0_outputs(561));
    outputs(2695) <= layer0_outputs(1290);
    outputs(2696) <= (layer0_outputs(608)) xor (layer0_outputs(1637));
    outputs(2697) <= not((layer0_outputs(3541)) xor (layer0_outputs(686)));
    outputs(2698) <= (layer0_outputs(152)) xor (layer0_outputs(2743));
    outputs(2699) <= (layer0_outputs(327)) xor (layer0_outputs(2913));
    outputs(2700) <= layer0_outputs(1671);
    outputs(2701) <= not((layer0_outputs(2494)) xor (layer0_outputs(3377)));
    outputs(2702) <= (layer0_outputs(3549)) xor (layer0_outputs(4303));
    outputs(2703) <= not(layer0_outputs(2297)) or (layer0_outputs(4981));
    outputs(2704) <= not(layer0_outputs(4230));
    outputs(2705) <= layer0_outputs(5063);
    outputs(2706) <= layer0_outputs(3183);
    outputs(2707) <= not(layer0_outputs(4625));
    outputs(2708) <= not((layer0_outputs(3195)) xor (layer0_outputs(3503)));
    outputs(2709) <= not((layer0_outputs(3508)) xor (layer0_outputs(2366)));
    outputs(2710) <= not((layer0_outputs(4550)) and (layer0_outputs(2430)));
    outputs(2711) <= not(layer0_outputs(1729));
    outputs(2712) <= (layer0_outputs(2932)) or (layer0_outputs(3765));
    outputs(2713) <= not(layer0_outputs(2368));
    outputs(2714) <= (layer0_outputs(62)) or (layer0_outputs(226));
    outputs(2715) <= (layer0_outputs(220)) and (layer0_outputs(2371));
    outputs(2716) <= not((layer0_outputs(1684)) xor (layer0_outputs(1292)));
    outputs(2717) <= (layer0_outputs(2392)) xor (layer0_outputs(1020));
    outputs(2718) <= not(layer0_outputs(4714));
    outputs(2719) <= (layer0_outputs(1518)) and not (layer0_outputs(391));
    outputs(2720) <= not((layer0_outputs(3467)) xor (layer0_outputs(2827)));
    outputs(2721) <= (layer0_outputs(660)) xor (layer0_outputs(4675));
    outputs(2722) <= layer0_outputs(4820);
    outputs(2723) <= not(layer0_outputs(3920)) or (layer0_outputs(3569));
    outputs(2724) <= not(layer0_outputs(4527));
    outputs(2725) <= (layer0_outputs(4395)) xor (layer0_outputs(3957));
    outputs(2726) <= (layer0_outputs(374)) and not (layer0_outputs(4344));
    outputs(2727) <= (layer0_outputs(1819)) and not (layer0_outputs(1555));
    outputs(2728) <= not(layer0_outputs(4111));
    outputs(2729) <= not((layer0_outputs(4407)) xor (layer0_outputs(1159)));
    outputs(2730) <= not(layer0_outputs(2686));
    outputs(2731) <= (layer0_outputs(4796)) xor (layer0_outputs(3491));
    outputs(2732) <= layer0_outputs(86);
    outputs(2733) <= not(layer0_outputs(4449));
    outputs(2734) <= not(layer0_outputs(3324));
    outputs(2735) <= (layer0_outputs(2208)) or (layer0_outputs(1147));
    outputs(2736) <= layer0_outputs(4517);
    outputs(2737) <= layer0_outputs(3200);
    outputs(2738) <= not((layer0_outputs(1931)) and (layer0_outputs(3899)));
    outputs(2739) <= not((layer0_outputs(976)) or (layer0_outputs(638)));
    outputs(2740) <= not((layer0_outputs(3137)) and (layer0_outputs(5017)));
    outputs(2741) <= layer0_outputs(8);
    outputs(2742) <= not(layer0_outputs(4847));
    outputs(2743) <= not((layer0_outputs(315)) xor (layer0_outputs(456)));
    outputs(2744) <= (layer0_outputs(2854)) and not (layer0_outputs(3098));
    outputs(2745) <= not(layer0_outputs(91));
    outputs(2746) <= (layer0_outputs(4579)) and not (layer0_outputs(1428));
    outputs(2747) <= not(layer0_outputs(713)) or (layer0_outputs(3449));
    outputs(2748) <= not(layer0_outputs(3686)) or (layer0_outputs(416));
    outputs(2749) <= (layer0_outputs(4718)) and (layer0_outputs(4165));
    outputs(2750) <= layer0_outputs(1172);
    outputs(2751) <= not((layer0_outputs(2722)) or (layer0_outputs(1939)));
    outputs(2752) <= layer0_outputs(4426);
    outputs(2753) <= (layer0_outputs(5045)) xor (layer0_outputs(3960));
    outputs(2754) <= not((layer0_outputs(134)) or (layer0_outputs(4828)));
    outputs(2755) <= layer0_outputs(1143);
    outputs(2756) <= not(layer0_outputs(3660));
    outputs(2757) <= layer0_outputs(1348);
    outputs(2758) <= layer0_outputs(5038);
    outputs(2759) <= (layer0_outputs(4254)) and not (layer0_outputs(1528));
    outputs(2760) <= (layer0_outputs(4649)) and not (layer0_outputs(1375));
    outputs(2761) <= (layer0_outputs(4591)) xor (layer0_outputs(4976));
    outputs(2762) <= (layer0_outputs(4992)) or (layer0_outputs(2399));
    outputs(2763) <= not(layer0_outputs(3893));
    outputs(2764) <= (layer0_outputs(2078)) xor (layer0_outputs(1574));
    outputs(2765) <= layer0_outputs(3754);
    outputs(2766) <= not(layer0_outputs(3793));
    outputs(2767) <= not(layer0_outputs(842));
    outputs(2768) <= not((layer0_outputs(2107)) xor (layer0_outputs(1928)));
    outputs(2769) <= layer0_outputs(2894);
    outputs(2770) <= not((layer0_outputs(3921)) xor (layer0_outputs(4783)));
    outputs(2771) <= layer0_outputs(1003);
    outputs(2772) <= not((layer0_outputs(4351)) xor (layer0_outputs(4231)));
    outputs(2773) <= not(layer0_outputs(2990));
    outputs(2774) <= layer0_outputs(381);
    outputs(2775) <= not(layer0_outputs(3684));
    outputs(2776) <= not((layer0_outputs(3420)) and (layer0_outputs(29)));
    outputs(2777) <= (layer0_outputs(4397)) and (layer0_outputs(2141));
    outputs(2778) <= not(layer0_outputs(4115)) or (layer0_outputs(4741));
    outputs(2779) <= not((layer0_outputs(4582)) and (layer0_outputs(4929)));
    outputs(2780) <= not(layer0_outputs(556));
    outputs(2781) <= not((layer0_outputs(467)) and (layer0_outputs(2798)));
    outputs(2782) <= layer0_outputs(4833);
    outputs(2783) <= not(layer0_outputs(644));
    outputs(2784) <= layer0_outputs(4748);
    outputs(2785) <= layer0_outputs(217);
    outputs(2786) <= not((layer0_outputs(2932)) or (layer0_outputs(3738)));
    outputs(2787) <= layer0_outputs(2615);
    outputs(2788) <= (layer0_outputs(5057)) or (layer0_outputs(1449));
    outputs(2789) <= not(layer0_outputs(2709)) or (layer0_outputs(2902));
    outputs(2790) <= not(layer0_outputs(576));
    outputs(2791) <= not((layer0_outputs(4047)) and (layer0_outputs(1165)));
    outputs(2792) <= (layer0_outputs(50)) and not (layer0_outputs(4849));
    outputs(2793) <= not(layer0_outputs(3431)) or (layer0_outputs(4532));
    outputs(2794) <= (layer0_outputs(4524)) and not (layer0_outputs(1004));
    outputs(2795) <= not(layer0_outputs(2585));
    outputs(2796) <= not((layer0_outputs(3663)) xor (layer0_outputs(2531)));
    outputs(2797) <= not(layer0_outputs(4279));
    outputs(2798) <= not(layer0_outputs(373)) or (layer0_outputs(1392));
    outputs(2799) <= not(layer0_outputs(4915));
    outputs(2800) <= layer0_outputs(4599);
    outputs(2801) <= layer0_outputs(108);
    outputs(2802) <= not((layer0_outputs(2076)) xor (layer0_outputs(2600)));
    outputs(2803) <= not((layer0_outputs(4549)) xor (layer0_outputs(41)));
    outputs(2804) <= (layer0_outputs(3119)) xor (layer0_outputs(867));
    outputs(2805) <= (layer0_outputs(2634)) and (layer0_outputs(5117));
    outputs(2806) <= not((layer0_outputs(4629)) xor (layer0_outputs(3513)));
    outputs(2807) <= not(layer0_outputs(4747));
    outputs(2808) <= not((layer0_outputs(2881)) xor (layer0_outputs(1745)));
    outputs(2809) <= not((layer0_outputs(997)) xor (layer0_outputs(4559)));
    outputs(2810) <= layer0_outputs(3952);
    outputs(2811) <= not(layer0_outputs(82));
    outputs(2812) <= not((layer0_outputs(204)) xor (layer0_outputs(1367)));
    outputs(2813) <= not((layer0_outputs(2382)) or (layer0_outputs(2899)));
    outputs(2814) <= not(layer0_outputs(143)) or (layer0_outputs(4681));
    outputs(2815) <= layer0_outputs(1880);
    outputs(2816) <= not(layer0_outputs(3587));
    outputs(2817) <= layer0_outputs(2943);
    outputs(2818) <= not(layer0_outputs(4266));
    outputs(2819) <= not(layer0_outputs(599)) or (layer0_outputs(3475));
    outputs(2820) <= layer0_outputs(1983);
    outputs(2821) <= not((layer0_outputs(3687)) xor (layer0_outputs(3969)));
    outputs(2822) <= layer0_outputs(3336);
    outputs(2823) <= (layer0_outputs(323)) and (layer0_outputs(2669));
    outputs(2824) <= (layer0_outputs(2934)) and not (layer0_outputs(2022));
    outputs(2825) <= (layer0_outputs(3232)) and (layer0_outputs(1561));
    outputs(2826) <= not((layer0_outputs(2046)) xor (layer0_outputs(4850)));
    outputs(2827) <= layer0_outputs(567);
    outputs(2828) <= (layer0_outputs(4912)) and not (layer0_outputs(51));
    outputs(2829) <= not(layer0_outputs(4810));
    outputs(2830) <= layer0_outputs(2023);
    outputs(2831) <= layer0_outputs(283);
    outputs(2832) <= layer0_outputs(796);
    outputs(2833) <= (layer0_outputs(1730)) and not (layer0_outputs(1442));
    outputs(2834) <= (layer0_outputs(3291)) xor (layer0_outputs(4374));
    outputs(2835) <= (layer0_outputs(1994)) and not (layer0_outputs(128));
    outputs(2836) <= (layer0_outputs(2569)) and (layer0_outputs(1091));
    outputs(2837) <= (layer0_outputs(518)) and (layer0_outputs(150));
    outputs(2838) <= not((layer0_outputs(4944)) or (layer0_outputs(1657)));
    outputs(2839) <= (layer0_outputs(5063)) and not (layer0_outputs(1800));
    outputs(2840) <= layer0_outputs(1453);
    outputs(2841) <= layer0_outputs(216);
    outputs(2842) <= layer0_outputs(4842);
    outputs(2843) <= layer0_outputs(3010);
    outputs(2844) <= (layer0_outputs(739)) xor (layer0_outputs(680));
    outputs(2845) <= not((layer0_outputs(2521)) xor (layer0_outputs(1481)));
    outputs(2846) <= not((layer0_outputs(3718)) xor (layer0_outputs(1577)));
    outputs(2847) <= not(layer0_outputs(955));
    outputs(2848) <= not((layer0_outputs(3542)) or (layer0_outputs(3589)));
    outputs(2849) <= not(layer0_outputs(228));
    outputs(2850) <= not(layer0_outputs(1524));
    outputs(2851) <= (layer0_outputs(1129)) and not (layer0_outputs(3926));
    outputs(2852) <= (layer0_outputs(758)) xor (layer0_outputs(1566));
    outputs(2853) <= not((layer0_outputs(1683)) xor (layer0_outputs(3600)));
    outputs(2854) <= not(layer0_outputs(56)) or (layer0_outputs(2905));
    outputs(2855) <= not((layer0_outputs(185)) xor (layer0_outputs(573)));
    outputs(2856) <= not(layer0_outputs(4939));
    outputs(2857) <= not(layer0_outputs(454));
    outputs(2858) <= not((layer0_outputs(2185)) or (layer0_outputs(1243)));
    outputs(2859) <= layer0_outputs(3892);
    outputs(2860) <= not((layer0_outputs(2579)) xor (layer0_outputs(2837)));
    outputs(2861) <= layer0_outputs(3402);
    outputs(2862) <= (layer0_outputs(890)) xor (layer0_outputs(1104));
    outputs(2863) <= (layer0_outputs(1645)) xor (layer0_outputs(1883));
    outputs(2864) <= not(layer0_outputs(2741)) or (layer0_outputs(3415));
    outputs(2865) <= not((layer0_outputs(1945)) and (layer0_outputs(4713)));
    outputs(2866) <= not(layer0_outputs(3704)) or (layer0_outputs(3529));
    outputs(2867) <= not((layer0_outputs(2644)) or (layer0_outputs(2126)));
    outputs(2868) <= not((layer0_outputs(3820)) xor (layer0_outputs(4468)));
    outputs(2869) <= layer0_outputs(3510);
    outputs(2870) <= layer0_outputs(63);
    outputs(2871) <= layer0_outputs(364);
    outputs(2872) <= not(layer0_outputs(148));
    outputs(2873) <= (layer0_outputs(513)) and not (layer0_outputs(1107));
    outputs(2874) <= '1';
    outputs(2875) <= (layer0_outputs(1671)) and (layer0_outputs(1857));
    outputs(2876) <= not((layer0_outputs(1427)) or (layer0_outputs(3192)));
    outputs(2877) <= (layer0_outputs(3409)) and not (layer0_outputs(125));
    outputs(2878) <= not((layer0_outputs(140)) or (layer0_outputs(1910)));
    outputs(2879) <= not((layer0_outputs(3794)) xor (layer0_outputs(3422)));
    outputs(2880) <= not((layer0_outputs(1583)) and (layer0_outputs(648)));
    outputs(2881) <= not(layer0_outputs(1817));
    outputs(2882) <= (layer0_outputs(1372)) xor (layer0_outputs(481));
    outputs(2883) <= not((layer0_outputs(116)) xor (layer0_outputs(2333)));
    outputs(2884) <= layer0_outputs(89);
    outputs(2885) <= not((layer0_outputs(3804)) xor (layer0_outputs(301)));
    outputs(2886) <= not(layer0_outputs(4140)) or (layer0_outputs(4609));
    outputs(2887) <= (layer0_outputs(156)) and not (layer0_outputs(174));
    outputs(2888) <= not(layer0_outputs(2373));
    outputs(2889) <= layer0_outputs(3089);
    outputs(2890) <= layer0_outputs(584);
    outputs(2891) <= not(layer0_outputs(871));
    outputs(2892) <= layer0_outputs(4180);
    outputs(2893) <= not((layer0_outputs(4383)) xor (layer0_outputs(1416)));
    outputs(2894) <= not(layer0_outputs(3312));
    outputs(2895) <= layer0_outputs(1321);
    outputs(2896) <= (layer0_outputs(1405)) or (layer0_outputs(4853));
    outputs(2897) <= layer0_outputs(2928);
    outputs(2898) <= layer0_outputs(4984);
    outputs(2899) <= not((layer0_outputs(1698)) or (layer0_outputs(3939)));
    outputs(2900) <= layer0_outputs(753);
    outputs(2901) <= not((layer0_outputs(26)) or (layer0_outputs(2276)));
    outputs(2902) <= not((layer0_outputs(3052)) and (layer0_outputs(4343)));
    outputs(2903) <= not(layer0_outputs(1543)) or (layer0_outputs(899));
    outputs(2904) <= not((layer0_outputs(504)) xor (layer0_outputs(2661)));
    outputs(2905) <= not((layer0_outputs(2548)) or (layer0_outputs(2385)));
    outputs(2906) <= not((layer0_outputs(288)) and (layer0_outputs(4617)));
    outputs(2907) <= not(layer0_outputs(2747));
    outputs(2908) <= (layer0_outputs(3940)) and not (layer0_outputs(3278));
    outputs(2909) <= not(layer0_outputs(2429));
    outputs(2910) <= not((layer0_outputs(1855)) and (layer0_outputs(553)));
    outputs(2911) <= not(layer0_outputs(2560));
    outputs(2912) <= layer0_outputs(1510);
    outputs(2913) <= layer0_outputs(4175);
    outputs(2914) <= not((layer0_outputs(4696)) xor (layer0_outputs(4215)));
    outputs(2915) <= not(layer0_outputs(3840));
    outputs(2916) <= not((layer0_outputs(382)) xor (layer0_outputs(2442)));
    outputs(2917) <= (layer0_outputs(528)) xor (layer0_outputs(3971));
    outputs(2918) <= not((layer0_outputs(3472)) and (layer0_outputs(3212)));
    outputs(2919) <= not(layer0_outputs(3012)) or (layer0_outputs(4587));
    outputs(2920) <= layer0_outputs(2881);
    outputs(2921) <= not(layer0_outputs(2219));
    outputs(2922) <= not(layer0_outputs(3652)) or (layer0_outputs(377));
    outputs(2923) <= layer0_outputs(1431);
    outputs(2924) <= layer0_outputs(3945);
    outputs(2925) <= not(layer0_outputs(2826));
    outputs(2926) <= (layer0_outputs(4876)) or (layer0_outputs(3788));
    outputs(2927) <= not(layer0_outputs(1753));
    outputs(2928) <= layer0_outputs(3603);
    outputs(2929) <= (layer0_outputs(710)) xor (layer0_outputs(2441));
    outputs(2930) <= not(layer0_outputs(3915));
    outputs(2931) <= (layer0_outputs(2972)) xor (layer0_outputs(1314));
    outputs(2932) <= (layer0_outputs(1826)) xor (layer0_outputs(3276));
    outputs(2933) <= not((layer0_outputs(2346)) xor (layer0_outputs(2581)));
    outputs(2934) <= (layer0_outputs(1879)) xor (layer0_outputs(4256));
    outputs(2935) <= layer0_outputs(4577);
    outputs(2936) <= not(layer0_outputs(1798));
    outputs(2937) <= not(layer0_outputs(3805)) or (layer0_outputs(4981));
    outputs(2938) <= not((layer0_outputs(2210)) or (layer0_outputs(3499)));
    outputs(2939) <= (layer0_outputs(2911)) and not (layer0_outputs(1530));
    outputs(2940) <= (layer0_outputs(4779)) and not (layer0_outputs(3844));
    outputs(2941) <= (layer0_outputs(1290)) and (layer0_outputs(2628));
    outputs(2942) <= (layer0_outputs(3247)) and (layer0_outputs(4293));
    outputs(2943) <= not((layer0_outputs(682)) xor (layer0_outputs(1419)));
    outputs(2944) <= (layer0_outputs(4827)) xor (layer0_outputs(900));
    outputs(2945) <= not(layer0_outputs(1630));
    outputs(2946) <= not((layer0_outputs(896)) and (layer0_outputs(94)));
    outputs(2947) <= (layer0_outputs(2803)) and not (layer0_outputs(0));
    outputs(2948) <= not(layer0_outputs(3330));
    outputs(2949) <= not(layer0_outputs(4210)) or (layer0_outputs(2867));
    outputs(2950) <= not(layer0_outputs(3552));
    outputs(2951) <= not(layer0_outputs(1218));
    outputs(2952) <= not((layer0_outputs(4630)) xor (layer0_outputs(2349)));
    outputs(2953) <= not(layer0_outputs(4476));
    outputs(2954) <= not(layer0_outputs(4968));
    outputs(2955) <= layer0_outputs(779);
    outputs(2956) <= (layer0_outputs(4582)) xor (layer0_outputs(1070));
    outputs(2957) <= (layer0_outputs(3631)) and not (layer0_outputs(1582));
    outputs(2958) <= layer0_outputs(160);
    outputs(2959) <= not(layer0_outputs(523));
    outputs(2960) <= (layer0_outputs(808)) xor (layer0_outputs(3812));
    outputs(2961) <= layer0_outputs(612);
    outputs(2962) <= not(layer0_outputs(2150));
    outputs(2963) <= not(layer0_outputs(1838));
    outputs(2964) <= not(layer0_outputs(3871));
    outputs(2965) <= (layer0_outputs(287)) or (layer0_outputs(4263));
    outputs(2966) <= not((layer0_outputs(1166)) xor (layer0_outputs(4212)));
    outputs(2967) <= not(layer0_outputs(1081));
    outputs(2968) <= not(layer0_outputs(3261));
    outputs(2969) <= (layer0_outputs(4843)) and (layer0_outputs(283));
    outputs(2970) <= layer0_outputs(4820);
    outputs(2971) <= layer0_outputs(612);
    outputs(2972) <= not(layer0_outputs(1387)) or (layer0_outputs(452));
    outputs(2973) <= not((layer0_outputs(3661)) xor (layer0_outputs(3275)));
    outputs(2974) <= not((layer0_outputs(1215)) and (layer0_outputs(2281)));
    outputs(2975) <= (layer0_outputs(5101)) and not (layer0_outputs(1872));
    outputs(2976) <= not((layer0_outputs(24)) or (layer0_outputs(2180)));
    outputs(2977) <= not(layer0_outputs(4893)) or (layer0_outputs(997));
    outputs(2978) <= not((layer0_outputs(3060)) xor (layer0_outputs(224)));
    outputs(2979) <= (layer0_outputs(4893)) or (layer0_outputs(336));
    outputs(2980) <= layer0_outputs(4122);
    outputs(2981) <= layer0_outputs(119);
    outputs(2982) <= (layer0_outputs(4788)) and not (layer0_outputs(4350));
    outputs(2983) <= not(layer0_outputs(4854));
    outputs(2984) <= (layer0_outputs(2788)) and (layer0_outputs(3554));
    outputs(2985) <= layer0_outputs(4135);
    outputs(2986) <= not((layer0_outputs(1584)) and (layer0_outputs(3372)));
    outputs(2987) <= (layer0_outputs(2863)) and not (layer0_outputs(2180));
    outputs(2988) <= (layer0_outputs(4564)) and (layer0_outputs(1941));
    outputs(2989) <= (layer0_outputs(1983)) xor (layer0_outputs(3903));
    outputs(2990) <= layer0_outputs(3572);
    outputs(2991) <= not((layer0_outputs(3544)) xor (layer0_outputs(4839)));
    outputs(2992) <= layer0_outputs(4805);
    outputs(2993) <= not(layer0_outputs(1667)) or (layer0_outputs(1344));
    outputs(2994) <= (layer0_outputs(656)) and not (layer0_outputs(607));
    outputs(2995) <= (layer0_outputs(2157)) and not (layer0_outputs(4139));
    outputs(2996) <= not((layer0_outputs(3594)) xor (layer0_outputs(3887)));
    outputs(2997) <= not(layer0_outputs(988)) or (layer0_outputs(4205));
    outputs(2998) <= layer0_outputs(2784);
    outputs(2999) <= layer0_outputs(1703);
    outputs(3000) <= not((layer0_outputs(1412)) or (layer0_outputs(1695)));
    outputs(3001) <= (layer0_outputs(1108)) xor (layer0_outputs(3624));
    outputs(3002) <= not(layer0_outputs(3410)) or (layer0_outputs(4515));
    outputs(3003) <= (layer0_outputs(662)) or (layer0_outputs(4466));
    outputs(3004) <= layer0_outputs(3988);
    outputs(3005) <= not(layer0_outputs(3093)) or (layer0_outputs(2018));
    outputs(3006) <= not((layer0_outputs(17)) xor (layer0_outputs(600)));
    outputs(3007) <= not((layer0_outputs(4482)) and (layer0_outputs(3587)));
    outputs(3008) <= not(layer0_outputs(1461));
    outputs(3009) <= layer0_outputs(3610);
    outputs(3010) <= not((layer0_outputs(3854)) xor (layer0_outputs(3826)));
    outputs(3011) <= not((layer0_outputs(883)) or (layer0_outputs(2912)));
    outputs(3012) <= layer0_outputs(1238);
    outputs(3013) <= not(layer0_outputs(2504));
    outputs(3014) <= not(layer0_outputs(3616));
    outputs(3015) <= not(layer0_outputs(2453)) or (layer0_outputs(196));
    outputs(3016) <= layer0_outputs(942);
    outputs(3017) <= (layer0_outputs(2338)) and (layer0_outputs(129));
    outputs(3018) <= (layer0_outputs(4055)) xor (layer0_outputs(724));
    outputs(3019) <= (layer0_outputs(1399)) and not (layer0_outputs(4552));
    outputs(3020) <= (layer0_outputs(3270)) and (layer0_outputs(3343));
    outputs(3021) <= not((layer0_outputs(1711)) or (layer0_outputs(4828)));
    outputs(3022) <= (layer0_outputs(4934)) or (layer0_outputs(2418));
    outputs(3023) <= (layer0_outputs(642)) and not (layer0_outputs(4811));
    outputs(3024) <= (layer0_outputs(4126)) xor (layer0_outputs(924));
    outputs(3025) <= layer0_outputs(1326);
    outputs(3026) <= layer0_outputs(540);
    outputs(3027) <= not(layer0_outputs(3848));
    outputs(3028) <= not(layer0_outputs(3042)) or (layer0_outputs(999));
    outputs(3029) <= (layer0_outputs(3528)) xor (layer0_outputs(4129));
    outputs(3030) <= layer0_outputs(4461);
    outputs(3031) <= not(layer0_outputs(2469));
    outputs(3032) <= not(layer0_outputs(2314)) or (layer0_outputs(2713));
    outputs(3033) <= layer0_outputs(4161);
    outputs(3034) <= (layer0_outputs(2394)) and (layer0_outputs(2946));
    outputs(3035) <= '0';
    outputs(3036) <= not((layer0_outputs(2984)) xor (layer0_outputs(2715)));
    outputs(3037) <= (layer0_outputs(4508)) xor (layer0_outputs(473));
    outputs(3038) <= not(layer0_outputs(2865)) or (layer0_outputs(4858));
    outputs(3039) <= not(layer0_outputs(1995));
    outputs(3040) <= not(layer0_outputs(4894));
    outputs(3041) <= layer0_outputs(944);
    outputs(3042) <= not((layer0_outputs(1583)) xor (layer0_outputs(650)));
    outputs(3043) <= not(layer0_outputs(911));
    outputs(3044) <= layer0_outputs(3922);
    outputs(3045) <= not(layer0_outputs(140)) or (layer0_outputs(3494));
    outputs(3046) <= (layer0_outputs(1449)) or (layer0_outputs(1246));
    outputs(3047) <= layer0_outputs(4171);
    outputs(3048) <= layer0_outputs(5032);
    outputs(3049) <= not(layer0_outputs(4527));
    outputs(3050) <= not((layer0_outputs(1908)) xor (layer0_outputs(1305)));
    outputs(3051) <= layer0_outputs(366);
    outputs(3052) <= not(layer0_outputs(2266));
    outputs(3053) <= layer0_outputs(670);
    outputs(3054) <= layer0_outputs(3929);
    outputs(3055) <= layer0_outputs(4410);
    outputs(3056) <= (layer0_outputs(4768)) xor (layer0_outputs(5116));
    outputs(3057) <= not(layer0_outputs(3948));
    outputs(3058) <= (layer0_outputs(4051)) xor (layer0_outputs(1144));
    outputs(3059) <= not(layer0_outputs(3849));
    outputs(3060) <= not(layer0_outputs(2444));
    outputs(3061) <= not(layer0_outputs(1690)) or (layer0_outputs(3512));
    outputs(3062) <= not(layer0_outputs(4509));
    outputs(3063) <= layer0_outputs(447);
    outputs(3064) <= (layer0_outputs(3154)) xor (layer0_outputs(642));
    outputs(3065) <= not((layer0_outputs(1357)) xor (layer0_outputs(3703)));
    outputs(3066) <= layer0_outputs(3875);
    outputs(3067) <= not((layer0_outputs(4096)) xor (layer0_outputs(4523)));
    outputs(3068) <= not(layer0_outputs(3919)) or (layer0_outputs(3597));
    outputs(3069) <= not(layer0_outputs(1018)) or (layer0_outputs(3263));
    outputs(3070) <= layer0_outputs(538);
    outputs(3071) <= not(layer0_outputs(599));
    outputs(3072) <= not((layer0_outputs(1017)) and (layer0_outputs(1523)));
    outputs(3073) <= (layer0_outputs(253)) and not (layer0_outputs(1122));
    outputs(3074) <= not(layer0_outputs(325));
    outputs(3075) <= not((layer0_outputs(3555)) or (layer0_outputs(2302)));
    outputs(3076) <= (layer0_outputs(4511)) and not (layer0_outputs(38));
    outputs(3077) <= not((layer0_outputs(1321)) or (layer0_outputs(2975)));
    outputs(3078) <= layer0_outputs(2356);
    outputs(3079) <= layer0_outputs(931);
    outputs(3080) <= layer0_outputs(1252);
    outputs(3081) <= (layer0_outputs(242)) xor (layer0_outputs(268));
    outputs(3082) <= not((layer0_outputs(1456)) and (layer0_outputs(1035)));
    outputs(3083) <= layer0_outputs(374);
    outputs(3084) <= not((layer0_outputs(20)) xor (layer0_outputs(526)));
    outputs(3085) <= layer0_outputs(5082);
    outputs(3086) <= not((layer0_outputs(73)) and (layer0_outputs(3263)));
    outputs(3087) <= layer0_outputs(2087);
    outputs(3088) <= not((layer0_outputs(291)) xor (layer0_outputs(1429)));
    outputs(3089) <= not((layer0_outputs(3014)) xor (layer0_outputs(207)));
    outputs(3090) <= (layer0_outputs(3716)) and not (layer0_outputs(3230));
    outputs(3091) <= (layer0_outputs(1992)) xor (layer0_outputs(1015));
    outputs(3092) <= not(layer0_outputs(5010)) or (layer0_outputs(4410));
    outputs(3093) <= (layer0_outputs(4123)) xor (layer0_outputs(2315));
    outputs(3094) <= not(layer0_outputs(238));
    outputs(3095) <= layer0_outputs(3917);
    outputs(3096) <= (layer0_outputs(3121)) and (layer0_outputs(5018));
    outputs(3097) <= (layer0_outputs(3619)) xor (layer0_outputs(1812));
    outputs(3098) <= (layer0_outputs(423)) or (layer0_outputs(2124));
    outputs(3099) <= (layer0_outputs(3301)) xor (layer0_outputs(4588));
    outputs(3100) <= not((layer0_outputs(903)) xor (layer0_outputs(1024)));
    outputs(3101) <= (layer0_outputs(2641)) and not (layer0_outputs(824));
    outputs(3102) <= not(layer0_outputs(873));
    outputs(3103) <= (layer0_outputs(2915)) and not (layer0_outputs(2496));
    outputs(3104) <= not((layer0_outputs(5061)) xor (layer0_outputs(553)));
    outputs(3105) <= (layer0_outputs(1265)) and not (layer0_outputs(1920));
    outputs(3106) <= layer0_outputs(4520);
    outputs(3107) <= (layer0_outputs(1997)) and (layer0_outputs(2104));
    outputs(3108) <= not((layer0_outputs(1919)) and (layer0_outputs(2701)));
    outputs(3109) <= (layer0_outputs(1689)) or (layer0_outputs(3962));
    outputs(3110) <= not((layer0_outputs(2917)) or (layer0_outputs(146)));
    outputs(3111) <= (layer0_outputs(19)) and not (layer0_outputs(1));
    outputs(3112) <= not(layer0_outputs(4613));
    outputs(3113) <= not((layer0_outputs(572)) and (layer0_outputs(2221)));
    outputs(3114) <= not(layer0_outputs(3391));
    outputs(3115) <= not(layer0_outputs(4238));
    outputs(3116) <= not(layer0_outputs(1142));
    outputs(3117) <= (layer0_outputs(1216)) and not (layer0_outputs(1342));
    outputs(3118) <= not((layer0_outputs(4685)) xor (layer0_outputs(2976)));
    outputs(3119) <= layer0_outputs(2216);
    outputs(3120) <= not((layer0_outputs(677)) and (layer0_outputs(2259)));
    outputs(3121) <= not(layer0_outputs(365));
    outputs(3122) <= (layer0_outputs(4012)) and not (layer0_outputs(4123));
    outputs(3123) <= not(layer0_outputs(3638));
    outputs(3124) <= not(layer0_outputs(4953));
    outputs(3125) <= not(layer0_outputs(4611));
    outputs(3126) <= layer0_outputs(4816);
    outputs(3127) <= not(layer0_outputs(4479));
    outputs(3128) <= not((layer0_outputs(4948)) or (layer0_outputs(10)));
    outputs(3129) <= (layer0_outputs(3000)) or (layer0_outputs(1697));
    outputs(3130) <= not(layer0_outputs(32)) or (layer0_outputs(1245));
    outputs(3131) <= not((layer0_outputs(2994)) and (layer0_outputs(1139)));
    outputs(3132) <= not(layer0_outputs(4631));
    outputs(3133) <= not((layer0_outputs(104)) xor (layer0_outputs(5044)));
    outputs(3134) <= not(layer0_outputs(2101));
    outputs(3135) <= (layer0_outputs(4655)) xor (layer0_outputs(254));
    outputs(3136) <= not((layer0_outputs(2728)) xor (layer0_outputs(3360)));
    outputs(3137) <= not((layer0_outputs(2636)) xor (layer0_outputs(945)));
    outputs(3138) <= layer0_outputs(1236);
    outputs(3139) <= not(layer0_outputs(4557));
    outputs(3140) <= (layer0_outputs(1745)) and not (layer0_outputs(457));
    outputs(3141) <= not(layer0_outputs(4146));
    outputs(3142) <= (layer0_outputs(4879)) and not (layer0_outputs(3637));
    outputs(3143) <= not(layer0_outputs(1552));
    outputs(3144) <= not(layer0_outputs(308));
    outputs(3145) <= (layer0_outputs(4659)) and not (layer0_outputs(380));
    outputs(3146) <= not(layer0_outputs(569));
    outputs(3147) <= not(layer0_outputs(1578));
    outputs(3148) <= (layer0_outputs(4614)) and (layer0_outputs(4703));
    outputs(3149) <= (layer0_outputs(3199)) and (layer0_outputs(4852));
    outputs(3150) <= layer0_outputs(399);
    outputs(3151) <= layer0_outputs(2664);
    outputs(3152) <= not(layer0_outputs(986));
    outputs(3153) <= layer0_outputs(1551);
    outputs(3154) <= not(layer0_outputs(476));
    outputs(3155) <= not((layer0_outputs(3716)) and (layer0_outputs(240)));
    outputs(3156) <= not(layer0_outputs(4719));
    outputs(3157) <= (layer0_outputs(3270)) xor (layer0_outputs(4849));
    outputs(3158) <= not(layer0_outputs(3780));
    outputs(3159) <= layer0_outputs(4078);
    outputs(3160) <= not(layer0_outputs(718));
    outputs(3161) <= not(layer0_outputs(2671));
    outputs(3162) <= layer0_outputs(2913);
    outputs(3163) <= not((layer0_outputs(3249)) or (layer0_outputs(4113)));
    outputs(3164) <= (layer0_outputs(2995)) xor (layer0_outputs(1664));
    outputs(3165) <= not((layer0_outputs(4623)) xor (layer0_outputs(1064)));
    outputs(3166) <= not(layer0_outputs(3117));
    outputs(3167) <= layer0_outputs(2925);
    outputs(3168) <= (layer0_outputs(2728)) and not (layer0_outputs(4039));
    outputs(3169) <= not(layer0_outputs(2688));
    outputs(3170) <= not(layer0_outputs(4905));
    outputs(3171) <= layer0_outputs(236);
    outputs(3172) <= not(layer0_outputs(4204)) or (layer0_outputs(3712));
    outputs(3173) <= (layer0_outputs(3388)) and (layer0_outputs(4237));
    outputs(3174) <= not(layer0_outputs(4605));
    outputs(3175) <= layer0_outputs(46);
    outputs(3176) <= layer0_outputs(3459);
    outputs(3177) <= not(layer0_outputs(4742));
    outputs(3178) <= not(layer0_outputs(3847));
    outputs(3179) <= (layer0_outputs(1180)) xor (layer0_outputs(3349));
    outputs(3180) <= not((layer0_outputs(1075)) xor (layer0_outputs(209)));
    outputs(3181) <= not((layer0_outputs(4587)) xor (layer0_outputs(421)));
    outputs(3182) <= layer0_outputs(782);
    outputs(3183) <= not(layer0_outputs(983));
    outputs(3184) <= not(layer0_outputs(492));
    outputs(3185) <= not(layer0_outputs(1203));
    outputs(3186) <= (layer0_outputs(317)) and (layer0_outputs(4290));
    outputs(3187) <= not(layer0_outputs(616));
    outputs(3188) <= layer0_outputs(2816);
    outputs(3189) <= not((layer0_outputs(4785)) and (layer0_outputs(298)));
    outputs(3190) <= (layer0_outputs(4089)) and not (layer0_outputs(1670));
    outputs(3191) <= (layer0_outputs(350)) xor (layer0_outputs(4650));
    outputs(3192) <= not((layer0_outputs(3896)) xor (layer0_outputs(4459)));
    outputs(3193) <= (layer0_outputs(4218)) and not (layer0_outputs(271));
    outputs(3194) <= not(layer0_outputs(3088)) or (layer0_outputs(337));
    outputs(3195) <= (layer0_outputs(542)) xor (layer0_outputs(4512));
    outputs(3196) <= not((layer0_outputs(4602)) xor (layer0_outputs(2717)));
    outputs(3197) <= (layer0_outputs(3382)) and (layer0_outputs(3805));
    outputs(3198) <= not(layer0_outputs(2145)) or (layer0_outputs(3027));
    outputs(3199) <= (layer0_outputs(3138)) xor (layer0_outputs(368));
    outputs(3200) <= not(layer0_outputs(1451));
    outputs(3201) <= not(layer0_outputs(4513));
    outputs(3202) <= (layer0_outputs(4927)) and not (layer0_outputs(700));
    outputs(3203) <= layer0_outputs(1026);
    outputs(3204) <= (layer0_outputs(1012)) and not (layer0_outputs(100));
    outputs(3205) <= (layer0_outputs(224)) and not (layer0_outputs(3146));
    outputs(3206) <= not(layer0_outputs(1214));
    outputs(3207) <= layer0_outputs(4640);
    outputs(3208) <= layer0_outputs(1981);
    outputs(3209) <= layer0_outputs(741);
    outputs(3210) <= not((layer0_outputs(3607)) or (layer0_outputs(4952)));
    outputs(3211) <= (layer0_outputs(3703)) or (layer0_outputs(4224));
    outputs(3212) <= (layer0_outputs(3407)) xor (layer0_outputs(424));
    outputs(3213) <= not(layer0_outputs(773)) or (layer0_outputs(756));
    outputs(3214) <= not((layer0_outputs(2308)) or (layer0_outputs(2791)));
    outputs(3215) <= layer0_outputs(1049);
    outputs(3216) <= (layer0_outputs(1464)) and not (layer0_outputs(83));
    outputs(3217) <= not(layer0_outputs(3936)) or (layer0_outputs(4108));
    outputs(3218) <= not((layer0_outputs(4391)) or (layer0_outputs(2513)));
    outputs(3219) <= (layer0_outputs(582)) and not (layer0_outputs(2753));
    outputs(3220) <= layer0_outputs(1770);
    outputs(3221) <= layer0_outputs(3592);
    outputs(3222) <= layer0_outputs(2084);
    outputs(3223) <= layer0_outputs(818);
    outputs(3224) <= (layer0_outputs(3747)) and not (layer0_outputs(2843));
    outputs(3225) <= layer0_outputs(622);
    outputs(3226) <= not(layer0_outputs(3225));
    outputs(3227) <= not((layer0_outputs(2711)) or (layer0_outputs(4600)));
    outputs(3228) <= not((layer0_outputs(3517)) xor (layer0_outputs(2677)));
    outputs(3229) <= not(layer0_outputs(4580)) or (layer0_outputs(837));
    outputs(3230) <= (layer0_outputs(4082)) and (layer0_outputs(1767));
    outputs(3231) <= not(layer0_outputs(4381));
    outputs(3232) <= (layer0_outputs(2175)) and not (layer0_outputs(4233));
    outputs(3233) <= (layer0_outputs(1961)) or (layer0_outputs(895));
    outputs(3234) <= layer0_outputs(2652);
    outputs(3235) <= layer0_outputs(3250);
    outputs(3236) <= not((layer0_outputs(790)) and (layer0_outputs(3940)));
    outputs(3237) <= not((layer0_outputs(2391)) or (layer0_outputs(523)));
    outputs(3238) <= not(layer0_outputs(2477)) or (layer0_outputs(4293));
    outputs(3239) <= (layer0_outputs(3857)) xor (layer0_outputs(5073));
    outputs(3240) <= (layer0_outputs(2182)) and not (layer0_outputs(2594));
    outputs(3241) <= not(layer0_outputs(173));
    outputs(3242) <= layer0_outputs(3388);
    outputs(3243) <= (layer0_outputs(3808)) and (layer0_outputs(5039));
    outputs(3244) <= not(layer0_outputs(3946)) or (layer0_outputs(72));
    outputs(3245) <= not(layer0_outputs(1500));
    outputs(3246) <= not(layer0_outputs(2468));
    outputs(3247) <= layer0_outputs(174);
    outputs(3248) <= not((layer0_outputs(1337)) or (layer0_outputs(679)));
    outputs(3249) <= not((layer0_outputs(628)) xor (layer0_outputs(4887)));
    outputs(3250) <= (layer0_outputs(167)) and (layer0_outputs(2793));
    outputs(3251) <= (layer0_outputs(5095)) xor (layer0_outputs(5105));
    outputs(3252) <= not(layer0_outputs(3541));
    outputs(3253) <= not(layer0_outputs(446));
    outputs(3254) <= not((layer0_outputs(4375)) xor (layer0_outputs(3794)));
    outputs(3255) <= (layer0_outputs(3961)) xor (layer0_outputs(1118));
    outputs(3256) <= (layer0_outputs(4347)) xor (layer0_outputs(1438));
    outputs(3257) <= not(layer0_outputs(2983));
    outputs(3258) <= not(layer0_outputs(1595));
    outputs(3259) <= not(layer0_outputs(5027));
    outputs(3260) <= not((layer0_outputs(380)) or (layer0_outputs(3198)));
    outputs(3261) <= not(layer0_outputs(1575)) or (layer0_outputs(4173));
    outputs(3262) <= not(layer0_outputs(1785));
    outputs(3263) <= layer0_outputs(2014);
    outputs(3264) <= (layer0_outputs(4370)) and not (layer0_outputs(1455));
    outputs(3265) <= not((layer0_outputs(3523)) and (layer0_outputs(1533)));
    outputs(3266) <= (layer0_outputs(478)) xor (layer0_outputs(2613));
    outputs(3267) <= layer0_outputs(509);
    outputs(3268) <= layer0_outputs(709);
    outputs(3269) <= (layer0_outputs(56)) and not (layer0_outputs(2532));
    outputs(3270) <= not(layer0_outputs(2277)) or (layer0_outputs(26));
    outputs(3271) <= (layer0_outputs(2546)) xor (layer0_outputs(158));
    outputs(3272) <= layer0_outputs(4254);
    outputs(3273) <= layer0_outputs(2330);
    outputs(3274) <= (layer0_outputs(2942)) and not (layer0_outputs(907));
    outputs(3275) <= not((layer0_outputs(418)) or (layer0_outputs(2691)));
    outputs(3276) <= layer0_outputs(1732);
    outputs(3277) <= not((layer0_outputs(4152)) or (layer0_outputs(4895)));
    outputs(3278) <= not((layer0_outputs(2876)) or (layer0_outputs(1160)));
    outputs(3279) <= not((layer0_outputs(2249)) xor (layer0_outputs(3058)));
    outputs(3280) <= (layer0_outputs(2945)) or (layer0_outputs(3493));
    outputs(3281) <= (layer0_outputs(2725)) xor (layer0_outputs(1742));
    outputs(3282) <= (layer0_outputs(2515)) and (layer0_outputs(4983));
    outputs(3283) <= not((layer0_outputs(1947)) or (layer0_outputs(800)));
    outputs(3284) <= (layer0_outputs(2237)) and not (layer0_outputs(1461));
    outputs(3285) <= layer0_outputs(4965);
    outputs(3286) <= not((layer0_outputs(1982)) xor (layer0_outputs(3573)));
    outputs(3287) <= not((layer0_outputs(4791)) xor (layer0_outputs(2318)));
    outputs(3288) <= not((layer0_outputs(2398)) and (layer0_outputs(2720)));
    outputs(3289) <= not((layer0_outputs(2537)) xor (layer0_outputs(88)));
    outputs(3290) <= not((layer0_outputs(4207)) and (layer0_outputs(3553)));
    outputs(3291) <= not(layer0_outputs(2870));
    outputs(3292) <= not((layer0_outputs(5030)) xor (layer0_outputs(236)));
    outputs(3293) <= (layer0_outputs(2522)) and not (layer0_outputs(4464));
    outputs(3294) <= not(layer0_outputs(1172));
    outputs(3295) <= not((layer0_outputs(1591)) and (layer0_outputs(3083)));
    outputs(3296) <= (layer0_outputs(488)) and (layer0_outputs(3562));
    outputs(3297) <= not((layer0_outputs(3181)) and (layer0_outputs(435)));
    outputs(3298) <= (layer0_outputs(60)) xor (layer0_outputs(3412));
    outputs(3299) <= (layer0_outputs(3368)) xor (layer0_outputs(2033));
    outputs(3300) <= (layer0_outputs(3342)) xor (layer0_outputs(626));
    outputs(3301) <= (layer0_outputs(3199)) xor (layer0_outputs(3299));
    outputs(3302) <= not(layer0_outputs(4533));
    outputs(3303) <= not((layer0_outputs(3490)) and (layer0_outputs(3404)));
    outputs(3304) <= not(layer0_outputs(1999));
    outputs(3305) <= layer0_outputs(1369);
    outputs(3306) <= layer0_outputs(1333);
    outputs(3307) <= not((layer0_outputs(715)) and (layer0_outputs(3767)));
    outputs(3308) <= layer0_outputs(3594);
    outputs(3309) <= (layer0_outputs(3667)) or (layer0_outputs(3757));
    outputs(3310) <= not((layer0_outputs(162)) and (layer0_outputs(3161)));
    outputs(3311) <= (layer0_outputs(4555)) and not (layer0_outputs(263));
    outputs(3312) <= (layer0_outputs(3913)) xor (layer0_outputs(3339));
    outputs(3313) <= (layer0_outputs(786)) and not (layer0_outputs(4771));
    outputs(3314) <= (layer0_outputs(1069)) and not (layer0_outputs(1092));
    outputs(3315) <= (layer0_outputs(2072)) xor (layer0_outputs(511));
    outputs(3316) <= (layer0_outputs(4642)) and (layer0_outputs(2003));
    outputs(3317) <= layer0_outputs(879);
    outputs(3318) <= not((layer0_outputs(4015)) or (layer0_outputs(452)));
    outputs(3319) <= not((layer0_outputs(554)) xor (layer0_outputs(3205)));
    outputs(3320) <= not(layer0_outputs(2176));
    outputs(3321) <= layer0_outputs(1096);
    outputs(3322) <= not((layer0_outputs(457)) xor (layer0_outputs(462)));
    outputs(3323) <= not((layer0_outputs(1011)) or (layer0_outputs(2678)));
    outputs(3324) <= layer0_outputs(669);
    outputs(3325) <= not(layer0_outputs(3540)) or (layer0_outputs(3711));
    outputs(3326) <= not((layer0_outputs(3741)) xor (layer0_outputs(602)));
    outputs(3327) <= layer0_outputs(3180);
    outputs(3328) <= (layer0_outputs(810)) and not (layer0_outputs(2972));
    outputs(3329) <= not((layer0_outputs(106)) xor (layer0_outputs(1744)));
    outputs(3330) <= not(layer0_outputs(2929));
    outputs(3331) <= not((layer0_outputs(852)) or (layer0_outputs(3104)));
    outputs(3332) <= (layer0_outputs(3874)) and (layer0_outputs(1018));
    outputs(3333) <= not(layer0_outputs(1797)) or (layer0_outputs(1864));
    outputs(3334) <= not((layer0_outputs(2964)) xor (layer0_outputs(1059)));
    outputs(3335) <= not(layer0_outputs(1576));
    outputs(3336) <= layer0_outputs(2473);
    outputs(3337) <= not(layer0_outputs(5104));
    outputs(3338) <= layer0_outputs(3534);
    outputs(3339) <= (layer0_outputs(4990)) xor (layer0_outputs(3951));
    outputs(3340) <= layer0_outputs(5014);
    outputs(3341) <= (layer0_outputs(4577)) xor (layer0_outputs(4483));
    outputs(3342) <= not(layer0_outputs(3295)) or (layer0_outputs(2950));
    outputs(3343) <= not((layer0_outputs(4962)) xor (layer0_outputs(4466)));
    outputs(3344) <= layer0_outputs(2922);
    outputs(3345) <= (layer0_outputs(4941)) and (layer0_outputs(1151));
    outputs(3346) <= not(layer0_outputs(4750));
    outputs(3347) <= layer0_outputs(5100);
    outputs(3348) <= not(layer0_outputs(917)) or (layer0_outputs(2542));
    outputs(3349) <= not((layer0_outputs(4424)) xor (layer0_outputs(2184)));
    outputs(3350) <= layer0_outputs(4210);
    outputs(3351) <= not(layer0_outputs(2067)) or (layer0_outputs(4657));
    outputs(3352) <= (layer0_outputs(909)) and not (layer0_outputs(2554));
    outputs(3353) <= not((layer0_outputs(2676)) xor (layer0_outputs(1201)));
    outputs(3354) <= layer0_outputs(4729);
    outputs(3355) <= not((layer0_outputs(3861)) or (layer0_outputs(4064)));
    outputs(3356) <= layer0_outputs(618);
    outputs(3357) <= layer0_outputs(2354);
    outputs(3358) <= not(layer0_outputs(159)) or (layer0_outputs(177));
    outputs(3359) <= layer0_outputs(3668);
    outputs(3360) <= (layer0_outputs(5106)) xor (layer0_outputs(2106));
    outputs(3361) <= not(layer0_outputs(467)) or (layer0_outputs(1330));
    outputs(3362) <= layer0_outputs(3376);
    outputs(3363) <= (layer0_outputs(1499)) xor (layer0_outputs(3362));
    outputs(3364) <= not(layer0_outputs(340));
    outputs(3365) <= layer0_outputs(4879);
    outputs(3366) <= layer0_outputs(2963);
    outputs(3367) <= (layer0_outputs(1324)) xor (layer0_outputs(4413));
    outputs(3368) <= not(layer0_outputs(1871));
    outputs(3369) <= layer0_outputs(3201);
    outputs(3370) <= (layer0_outputs(801)) and not (layer0_outputs(296));
    outputs(3371) <= not((layer0_outputs(92)) xor (layer0_outputs(348)));
    outputs(3372) <= (layer0_outputs(2830)) and (layer0_outputs(4590));
    outputs(3373) <= not((layer0_outputs(520)) or (layer0_outputs(4779)));
    outputs(3374) <= layer0_outputs(91);
    outputs(3375) <= layer0_outputs(1073);
    outputs(3376) <= not(layer0_outputs(4874)) or (layer0_outputs(2265));
    outputs(3377) <= layer0_outputs(2205);
    outputs(3378) <= not(layer0_outputs(25)) or (layer0_outputs(3169));
    outputs(3379) <= layer0_outputs(3283);
    outputs(3380) <= layer0_outputs(2610);
    outputs(3381) <= not((layer0_outputs(151)) or (layer0_outputs(865)));
    outputs(3382) <= not(layer0_outputs(2209));
    outputs(3383) <= not(layer0_outputs(1561));
    outputs(3384) <= layer0_outputs(3437);
    outputs(3385) <= layer0_outputs(1633);
    outputs(3386) <= (layer0_outputs(4145)) xor (layer0_outputs(4024));
    outputs(3387) <= layer0_outputs(5004);
    outputs(3388) <= not(layer0_outputs(3233));
    outputs(3389) <= not(layer0_outputs(2657));
    outputs(3390) <= layer0_outputs(3826);
    outputs(3391) <= (layer0_outputs(3883)) and not (layer0_outputs(1659));
    outputs(3392) <= (layer0_outputs(3980)) xor (layer0_outputs(1485));
    outputs(3393) <= layer0_outputs(1508);
    outputs(3394) <= not((layer0_outputs(3468)) xor (layer0_outputs(4148)));
    outputs(3395) <= not((layer0_outputs(3298)) and (layer0_outputs(1246)));
    outputs(3396) <= not(layer0_outputs(4250));
    outputs(3397) <= (layer0_outputs(2415)) and not (layer0_outputs(3929));
    outputs(3398) <= layer0_outputs(3866);
    outputs(3399) <= not(layer0_outputs(5041));
    outputs(3400) <= not((layer0_outputs(4153)) xor (layer0_outputs(205)));
    outputs(3401) <= layer0_outputs(3194);
    outputs(3402) <= not((layer0_outputs(4003)) xor (layer0_outputs(3943)));
    outputs(3403) <= not(layer0_outputs(1716)) or (layer0_outputs(1647));
    outputs(3404) <= not(layer0_outputs(1229));
    outputs(3405) <= not((layer0_outputs(2194)) xor (layer0_outputs(3043)));
    outputs(3406) <= layer0_outputs(4267);
    outputs(3407) <= (layer0_outputs(3317)) xor (layer0_outputs(3889));
    outputs(3408) <= layer0_outputs(723);
    outputs(3409) <= layer0_outputs(1760);
    outputs(3410) <= not((layer0_outputs(2166)) xor (layer0_outputs(2015)));
    outputs(3411) <= layer0_outputs(3949);
    outputs(3412) <= layer0_outputs(4404);
    outputs(3413) <= not(layer0_outputs(31));
    outputs(3414) <= not(layer0_outputs(2726));
    outputs(3415) <= (layer0_outputs(934)) and not (layer0_outputs(1302));
    outputs(3416) <= (layer0_outputs(2539)) xor (layer0_outputs(2472));
    outputs(3417) <= layer0_outputs(3836);
    outputs(3418) <= not(layer0_outputs(4666));
    outputs(3419) <= not((layer0_outputs(4197)) xor (layer0_outputs(4221)));
    outputs(3420) <= layer0_outputs(868);
    outputs(3421) <= not(layer0_outputs(2361));
    outputs(3422) <= not(layer0_outputs(427));
    outputs(3423) <= (layer0_outputs(1315)) or (layer0_outputs(4525));
    outputs(3424) <= not((layer0_outputs(2170)) xor (layer0_outputs(3956)));
    outputs(3425) <= not(layer0_outputs(4917));
    outputs(3426) <= not((layer0_outputs(2513)) xor (layer0_outputs(2955)));
    outputs(3427) <= (layer0_outputs(5003)) and not (layer0_outputs(4102));
    outputs(3428) <= (layer0_outputs(1727)) xor (layer0_outputs(1930));
    outputs(3429) <= (layer0_outputs(1426)) xor (layer0_outputs(2745));
    outputs(3430) <= not(layer0_outputs(4516)) or (layer0_outputs(2198));
    outputs(3431) <= not((layer0_outputs(3245)) xor (layer0_outputs(4826)));
    outputs(3432) <= layer0_outputs(3029);
    outputs(3433) <= layer0_outputs(2258);
    outputs(3434) <= not((layer0_outputs(883)) xor (layer0_outputs(5053)));
    outputs(3435) <= layer0_outputs(1115);
    outputs(3436) <= not((layer0_outputs(3262)) or (layer0_outputs(1602)));
    outputs(3437) <= not((layer0_outputs(3089)) xor (layer0_outputs(3352)));
    outputs(3438) <= not(layer0_outputs(4409)) or (layer0_outputs(4749));
    outputs(3439) <= (layer0_outputs(2052)) and not (layer0_outputs(2121));
    outputs(3440) <= not(layer0_outputs(2622));
    outputs(3441) <= layer0_outputs(2639);
    outputs(3442) <= layer0_outputs(2435);
    outputs(3443) <= (layer0_outputs(948)) and not (layer0_outputs(3448));
    outputs(3444) <= not(layer0_outputs(4926));
    outputs(3445) <= layer0_outputs(2673);
    outputs(3446) <= not((layer0_outputs(4660)) xor (layer0_outputs(3319)));
    outputs(3447) <= not(layer0_outputs(3536)) or (layer0_outputs(961));
    outputs(3448) <= not(layer0_outputs(2909));
    outputs(3449) <= not(layer0_outputs(2983));
    outputs(3450) <= layer0_outputs(4007);
    outputs(3451) <= not((layer0_outputs(351)) or (layer0_outputs(4938)));
    outputs(3452) <= not((layer0_outputs(2592)) or (layer0_outputs(566)));
    outputs(3453) <= (layer0_outputs(2560)) and not (layer0_outputs(4297));
    outputs(3454) <= not(layer0_outputs(2209));
    outputs(3455) <= (layer0_outputs(4495)) xor (layer0_outputs(2820));
    outputs(3456) <= not((layer0_outputs(4406)) xor (layer0_outputs(182)));
    outputs(3457) <= (layer0_outputs(4543)) and not (layer0_outputs(4954));
    outputs(3458) <= (layer0_outputs(3427)) and not (layer0_outputs(1869));
    outputs(3459) <= not(layer0_outputs(2067));
    outputs(3460) <= not(layer0_outputs(487));
    outputs(3461) <= layer0_outputs(3398);
    outputs(3462) <= (layer0_outputs(4101)) xor (layer0_outputs(895));
    outputs(3463) <= (layer0_outputs(4918)) xor (layer0_outputs(1453));
    outputs(3464) <= layer0_outputs(795);
    outputs(3465) <= layer0_outputs(1285);
    outputs(3466) <= not((layer0_outputs(2917)) or (layer0_outputs(3982)));
    outputs(3467) <= not((layer0_outputs(2391)) or (layer0_outputs(1477)));
    outputs(3468) <= not((layer0_outputs(478)) xor (layer0_outputs(1659)));
    outputs(3469) <= not((layer0_outputs(4776)) and (layer0_outputs(2285)));
    outputs(3470) <= layer0_outputs(3965);
    outputs(3471) <= (layer0_outputs(5023)) xor (layer0_outputs(133));
    outputs(3472) <= (layer0_outputs(4471)) and not (layer0_outputs(4182));
    outputs(3473) <= not((layer0_outputs(4690)) or (layer0_outputs(4606)));
    outputs(3474) <= not((layer0_outputs(1097)) xor (layer0_outputs(4832)));
    outputs(3475) <= (layer0_outputs(617)) and not (layer0_outputs(2443));
    outputs(3476) <= (layer0_outputs(1658)) and (layer0_outputs(2581));
    outputs(3477) <= not(layer0_outputs(1901));
    outputs(3478) <= (layer0_outputs(1194)) and not (layer0_outputs(4472));
    outputs(3479) <= not(layer0_outputs(3982));
    outputs(3480) <= not((layer0_outputs(1196)) xor (layer0_outputs(1799)));
    outputs(3481) <= not((layer0_outputs(4020)) xor (layer0_outputs(2715)));
    outputs(3482) <= layer0_outputs(657);
    outputs(3483) <= not(layer0_outputs(3251));
    outputs(3484) <= not(layer0_outputs(3392));
    outputs(3485) <= layer0_outputs(1846);
    outputs(3486) <= not((layer0_outputs(672)) and (layer0_outputs(1782)));
    outputs(3487) <= not(layer0_outputs(2653));
    outputs(3488) <= (layer0_outputs(1894)) and (layer0_outputs(1958));
    outputs(3489) <= not(layer0_outputs(3823));
    outputs(3490) <= not((layer0_outputs(3206)) or (layer0_outputs(3181)));
    outputs(3491) <= (layer0_outputs(357)) xor (layer0_outputs(4097));
    outputs(3492) <= not((layer0_outputs(2590)) or (layer0_outputs(1691)));
    outputs(3493) <= layer0_outputs(5081);
    outputs(3494) <= layer0_outputs(4065);
    outputs(3495) <= layer0_outputs(3978);
    outputs(3496) <= not(layer0_outputs(4313));
    outputs(3497) <= layer0_outputs(1295);
    outputs(3498) <= not(layer0_outputs(1234));
    outputs(3499) <= not(layer0_outputs(2305));
    outputs(3500) <= layer0_outputs(1514);
    outputs(3501) <= not(layer0_outputs(318));
    outputs(3502) <= layer0_outputs(900);
    outputs(3503) <= layer0_outputs(1751);
    outputs(3504) <= not(layer0_outputs(4076));
    outputs(3505) <= not(layer0_outputs(1266));
    outputs(3506) <= (layer0_outputs(1728)) xor (layer0_outputs(4253));
    outputs(3507) <= layer0_outputs(948);
    outputs(3508) <= layer0_outputs(211);
    outputs(3509) <= not(layer0_outputs(2584));
    outputs(3510) <= (layer0_outputs(461)) and not (layer0_outputs(1409));
    outputs(3511) <= layer0_outputs(1262);
    outputs(3512) <= (layer0_outputs(1874)) and not (layer0_outputs(3550));
    outputs(3513) <= (layer0_outputs(4283)) and not (layer0_outputs(2973));
    outputs(3514) <= (layer0_outputs(2104)) and not (layer0_outputs(3657));
    outputs(3515) <= (layer0_outputs(1681)) and not (layer0_outputs(2647));
    outputs(3516) <= (layer0_outputs(2222)) or (layer0_outputs(4263));
    outputs(3517) <= (layer0_outputs(915)) or (layer0_outputs(1057));
    outputs(3518) <= layer0_outputs(3622);
    outputs(3519) <= layer0_outputs(3545);
    outputs(3520) <= (layer0_outputs(2456)) and not (layer0_outputs(4664));
    outputs(3521) <= layer0_outputs(3279);
    outputs(3522) <= layer0_outputs(1861);
    outputs(3523) <= layer0_outputs(3123);
    outputs(3524) <= (layer0_outputs(4397)) xor (layer0_outputs(3891));
    outputs(3525) <= layer0_outputs(3040);
    outputs(3526) <= (layer0_outputs(2336)) or (layer0_outputs(3711));
    outputs(3527) <= layer0_outputs(4094);
    outputs(3528) <= layer0_outputs(3236);
    outputs(3529) <= not(layer0_outputs(4103)) or (layer0_outputs(3789));
    outputs(3530) <= layer0_outputs(2859);
    outputs(3531) <= (layer0_outputs(195)) xor (layer0_outputs(1990));
    outputs(3532) <= not((layer0_outputs(4867)) or (layer0_outputs(4464)));
    outputs(3533) <= layer0_outputs(3763);
    outputs(3534) <= (layer0_outputs(4850)) xor (layer0_outputs(1153));
    outputs(3535) <= (layer0_outputs(4282)) and (layer0_outputs(45));
    outputs(3536) <= layer0_outputs(4840);
    outputs(3537) <= not((layer0_outputs(4403)) xor (layer0_outputs(4829)));
    outputs(3538) <= (layer0_outputs(3074)) and (layer0_outputs(2110));
    outputs(3539) <= not(layer0_outputs(3113));
    outputs(3540) <= not(layer0_outputs(4097));
    outputs(3541) <= not(layer0_outputs(4260));
    outputs(3542) <= (layer0_outputs(111)) xor (layer0_outputs(2013));
    outputs(3543) <= not((layer0_outputs(947)) xor (layer0_outputs(2719)));
    outputs(3544) <= (layer0_outputs(1666)) or (layer0_outputs(3279));
    outputs(3545) <= not((layer0_outputs(3001)) and (layer0_outputs(4265)));
    outputs(3546) <= not(layer0_outputs(1913));
    outputs(3547) <= layer0_outputs(4830);
    outputs(3548) <= not(layer0_outputs(519));
    outputs(3549) <= not(layer0_outputs(894));
    outputs(3550) <= layer0_outputs(3267);
    outputs(3551) <= not(layer0_outputs(1128));
    outputs(3552) <= not((layer0_outputs(1988)) xor (layer0_outputs(1391)));
    outputs(3553) <= not(layer0_outputs(1440));
    outputs(3554) <= layer0_outputs(1806);
    outputs(3555) <= not(layer0_outputs(4963)) or (layer0_outputs(1227));
    outputs(3556) <= layer0_outputs(2924);
    outputs(3557) <= (layer0_outputs(4687)) and not (layer0_outputs(1998));
    outputs(3558) <= (layer0_outputs(4386)) xor (layer0_outputs(1043));
    outputs(3559) <= not((layer0_outputs(2656)) or (layer0_outputs(4014)));
    outputs(3560) <= not((layer0_outputs(2172)) xor (layer0_outputs(3444)));
    outputs(3561) <= layer0_outputs(428);
    outputs(3562) <= not(layer0_outputs(3523)) or (layer0_outputs(3849));
    outputs(3563) <= not(layer0_outputs(4546));
    outputs(3564) <= not(layer0_outputs(3));
    outputs(3565) <= (layer0_outputs(4309)) and (layer0_outputs(1974));
    outputs(3566) <= not(layer0_outputs(1037));
    outputs(3567) <= (layer0_outputs(4018)) and not (layer0_outputs(2776));
    outputs(3568) <= (layer0_outputs(1209)) and (layer0_outputs(2402));
    outputs(3569) <= (layer0_outputs(3461)) and not (layer0_outputs(2933));
    outputs(3570) <= not(layer0_outputs(3208));
    outputs(3571) <= not(layer0_outputs(2221));
    outputs(3572) <= not(layer0_outputs(3602));
    outputs(3573) <= not(layer0_outputs(2486)) or (layer0_outputs(3831));
    outputs(3574) <= not(layer0_outputs(480)) or (layer0_outputs(1450));
    outputs(3575) <= '0';
    outputs(3576) <= (layer0_outputs(4708)) xor (layer0_outputs(3693));
    outputs(3577) <= not(layer0_outputs(30));
    outputs(3578) <= not((layer0_outputs(4617)) xor (layer0_outputs(4)));
    outputs(3579) <= (layer0_outputs(2230)) or (layer0_outputs(1779));
    outputs(3580) <= layer0_outputs(273);
    outputs(3581) <= not(layer0_outputs(2554));
    outputs(3582) <= not((layer0_outputs(1189)) or (layer0_outputs(4028)));
    outputs(3583) <= not((layer0_outputs(217)) xor (layer0_outputs(1852)));
    outputs(3584) <= (layer0_outputs(1407)) or (layer0_outputs(3953));
    outputs(3585) <= not((layer0_outputs(4361)) and (layer0_outputs(4402)));
    outputs(3586) <= not(layer0_outputs(3534));
    outputs(3587) <= not(layer0_outputs(3506)) or (layer0_outputs(4799));
    outputs(3588) <= not((layer0_outputs(3782)) xor (layer0_outputs(4384)));
    outputs(3589) <= (layer0_outputs(512)) and not (layer0_outputs(1115));
    outputs(3590) <= not(layer0_outputs(2822)) or (layer0_outputs(2897));
    outputs(3591) <= not(layer0_outputs(4644));
    outputs(3592) <= not(layer0_outputs(2128));
    outputs(3593) <= not((layer0_outputs(4644)) or (layer0_outputs(915)));
    outputs(3594) <= not(layer0_outputs(4739));
    outputs(3595) <= not((layer0_outputs(4436)) xor (layer0_outputs(4160)));
    outputs(3596) <= not((layer0_outputs(762)) xor (layer0_outputs(4063)));
    outputs(3597) <= (layer0_outputs(4074)) and not (layer0_outputs(1831));
    outputs(3598) <= not((layer0_outputs(4841)) xor (layer0_outputs(1993)));
    outputs(3599) <= not((layer0_outputs(2978)) xor (layer0_outputs(2269)));
    outputs(3600) <= layer0_outputs(2673);
    outputs(3601) <= not((layer0_outputs(4493)) or (layer0_outputs(494)));
    outputs(3602) <= layer0_outputs(3868);
    outputs(3603) <= layer0_outputs(3133);
    outputs(3604) <= not(layer0_outputs(1044));
    outputs(3605) <= (layer0_outputs(1250)) xor (layer0_outputs(861));
    outputs(3606) <= not((layer0_outputs(4029)) and (layer0_outputs(4265)));
    outputs(3607) <= not((layer0_outputs(200)) xor (layer0_outputs(2605)));
    outputs(3608) <= (layer0_outputs(2058)) and not (layer0_outputs(1544));
    outputs(3609) <= (layer0_outputs(3762)) xor (layer0_outputs(4867));
    outputs(3610) <= (layer0_outputs(1178)) and not (layer0_outputs(2538));
    outputs(3611) <= (layer0_outputs(4802)) and not (layer0_outputs(1415));
    outputs(3612) <= layer0_outputs(1662);
    outputs(3613) <= (layer0_outputs(3612)) and not (layer0_outputs(3578));
    outputs(3614) <= not(layer0_outputs(1709));
    outputs(3615) <= layer0_outputs(905);
    outputs(3616) <= not(layer0_outputs(2608));
    outputs(3617) <= not(layer0_outputs(1349));
    outputs(3618) <= (layer0_outputs(361)) xor (layer0_outputs(2018));
    outputs(3619) <= not((layer0_outputs(1876)) xor (layer0_outputs(1388)));
    outputs(3620) <= (layer0_outputs(2133)) and not (layer0_outputs(3547));
    outputs(3621) <= (layer0_outputs(58)) xor (layer0_outputs(4463));
    outputs(3622) <= (layer0_outputs(85)) and (layer0_outputs(3723));
    outputs(3623) <= (layer0_outputs(4260)) and not (layer0_outputs(2071));
    outputs(3624) <= not(layer0_outputs(2380)) or (layer0_outputs(3465));
    outputs(3625) <= layer0_outputs(4490);
    outputs(3626) <= (layer0_outputs(1279)) and not (layer0_outputs(699));
    outputs(3627) <= layer0_outputs(993);
    outputs(3628) <= (layer0_outputs(3686)) and not (layer0_outputs(4021));
    outputs(3629) <= layer0_outputs(4379);
    outputs(3630) <= not(layer0_outputs(2431)) or (layer0_outputs(3058));
    outputs(3631) <= (layer0_outputs(3235)) and (layer0_outputs(4339));
    outputs(3632) <= (layer0_outputs(53)) and not (layer0_outputs(3100));
    outputs(3633) <= (layer0_outputs(429)) and not (layer0_outputs(912));
    outputs(3634) <= (layer0_outputs(4819)) xor (layer0_outputs(2392));
    outputs(3635) <= layer0_outputs(987);
    outputs(3636) <= not((layer0_outputs(4310)) xor (layer0_outputs(2502)));
    outputs(3637) <= layer0_outputs(4345);
    outputs(3638) <= (layer0_outputs(787)) and (layer0_outputs(5110));
    outputs(3639) <= layer0_outputs(3041);
    outputs(3640) <= (layer0_outputs(486)) xor (layer0_outputs(3356));
    outputs(3641) <= (layer0_outputs(4082)) and not (layer0_outputs(2041));
    outputs(3642) <= (layer0_outputs(1792)) and (layer0_outputs(4842));
    outputs(3643) <= (layer0_outputs(2316)) xor (layer0_outputs(45));
    outputs(3644) <= not((layer0_outputs(2484)) xor (layer0_outputs(3785)));
    outputs(3645) <= layer0_outputs(1873);
    outputs(3646) <= not(layer0_outputs(3852));
    outputs(3647) <= (layer0_outputs(2779)) and (layer0_outputs(1101));
    outputs(3648) <= layer0_outputs(4327);
    outputs(3649) <= (layer0_outputs(2365)) and not (layer0_outputs(4267));
    outputs(3650) <= layer0_outputs(4700);
    outputs(3651) <= layer0_outputs(4967);
    outputs(3652) <= not(layer0_outputs(2236));
    outputs(3653) <= layer0_outputs(2589);
    outputs(3654) <= not((layer0_outputs(3488)) or (layer0_outputs(4390)));
    outputs(3655) <= layer0_outputs(3434);
    outputs(3656) <= not(layer0_outputs(4835));
    outputs(3657) <= not((layer0_outputs(3022)) xor (layer0_outputs(4985)));
    outputs(3658) <= (layer0_outputs(3019)) and not (layer0_outputs(248));
    outputs(3659) <= not((layer0_outputs(5043)) xor (layer0_outputs(134)));
    outputs(3660) <= not(layer0_outputs(1124));
    outputs(3661) <= not(layer0_outputs(2687));
    outputs(3662) <= (layer0_outputs(3643)) and (layer0_outputs(4326));
    outputs(3663) <= not(layer0_outputs(4364));
    outputs(3664) <= not((layer0_outputs(664)) or (layer0_outputs(3409)));
    outputs(3665) <= not((layer0_outputs(1358)) or (layer0_outputs(4434)));
    outputs(3666) <= not(layer0_outputs(1483));
    outputs(3667) <= (layer0_outputs(863)) xor (layer0_outputs(2311));
    outputs(3668) <= not((layer0_outputs(1052)) and (layer0_outputs(2057)));
    outputs(3669) <= layer0_outputs(2289);
    outputs(3670) <= (layer0_outputs(4377)) and not (layer0_outputs(398));
    outputs(3671) <= not(layer0_outputs(1824));
    outputs(3672) <= not(layer0_outputs(942));
    outputs(3673) <= not(layer0_outputs(219));
    outputs(3674) <= (layer0_outputs(4025)) and not (layer0_outputs(4898));
    outputs(3675) <= (layer0_outputs(1060)) and not (layer0_outputs(717));
    outputs(3676) <= not(layer0_outputs(2956));
    outputs(3677) <= (layer0_outputs(3634)) and not (layer0_outputs(1929));
    outputs(3678) <= not((layer0_outputs(2003)) xor (layer0_outputs(1343)));
    outputs(3679) <= (layer0_outputs(966)) and not (layer0_outputs(4361));
    outputs(3680) <= (layer0_outputs(1935)) and not (layer0_outputs(3009));
    outputs(3681) <= not((layer0_outputs(1242)) xor (layer0_outputs(954)));
    outputs(3682) <= not(layer0_outputs(331));
    outputs(3683) <= layer0_outputs(4570);
    outputs(3684) <= not(layer0_outputs(2000));
    outputs(3685) <= layer0_outputs(450);
    outputs(3686) <= (layer0_outputs(2093)) and not (layer0_outputs(2986));
    outputs(3687) <= not((layer0_outputs(3063)) xor (layer0_outputs(1599)));
    outputs(3688) <= (layer0_outputs(1247)) xor (layer0_outputs(2358));
    outputs(3689) <= (layer0_outputs(9)) xor (layer0_outputs(1289));
    outputs(3690) <= not((layer0_outputs(1981)) xor (layer0_outputs(551)));
    outputs(3691) <= (layer0_outputs(4559)) xor (layer0_outputs(500));
    outputs(3692) <= (layer0_outputs(1627)) xor (layer0_outputs(3240));
    outputs(3693) <= (layer0_outputs(614)) and (layer0_outputs(1344));
    outputs(3694) <= not((layer0_outputs(3165)) or (layer0_outputs(3888)));
    outputs(3695) <= layer0_outputs(2722);
    outputs(3696) <= layer0_outputs(2246);
    outputs(3697) <= not(layer0_outputs(3471));
    outputs(3698) <= (layer0_outputs(2809)) and not (layer0_outputs(2566));
    outputs(3699) <= layer0_outputs(1368);
    outputs(3700) <= (layer0_outputs(3511)) and (layer0_outputs(90));
    outputs(3701) <= (layer0_outputs(2815)) and not (layer0_outputs(1624));
    outputs(3702) <= layer0_outputs(2723);
    outputs(3703) <= (layer0_outputs(4509)) and not (layer0_outputs(126));
    outputs(3704) <= not(layer0_outputs(98));
    outputs(3705) <= (layer0_outputs(3096)) and (layer0_outputs(656));
    outputs(3706) <= not((layer0_outputs(3742)) or (layer0_outputs(1148)));
    outputs(3707) <= not((layer0_outputs(674)) xor (layer0_outputs(4485)));
    outputs(3708) <= (layer0_outputs(4896)) and not (layer0_outputs(2354));
    outputs(3709) <= layer0_outputs(665);
    outputs(3710) <= (layer0_outputs(4576)) and (layer0_outputs(270));
    outputs(3711) <= (layer0_outputs(4686)) or (layer0_outputs(3838));
    outputs(3712) <= layer0_outputs(1608);
    outputs(3713) <= (layer0_outputs(4376)) and not (layer0_outputs(2816));
    outputs(3714) <= '0';
    outputs(3715) <= layer0_outputs(3979);
    outputs(3716) <= not((layer0_outputs(2408)) or (layer0_outputs(5060)));
    outputs(3717) <= (layer0_outputs(2387)) and not (layer0_outputs(3323));
    outputs(3718) <= (layer0_outputs(3684)) and not (layer0_outputs(4124));
    outputs(3719) <= layer0_outputs(2343);
    outputs(3720) <= not(layer0_outputs(4199));
    outputs(3721) <= not(layer0_outputs(1433));
    outputs(3722) <= layer0_outputs(3857);
    outputs(3723) <= not(layer0_outputs(3044));
    outputs(3724) <= (layer0_outputs(3379)) and (layer0_outputs(294));
    outputs(3725) <= (layer0_outputs(1371)) and not (layer0_outputs(1705));
    outputs(3726) <= not(layer0_outputs(3397)) or (layer0_outputs(420));
    outputs(3727) <= layer0_outputs(2156);
    outputs(3728) <= layer0_outputs(1006);
    outputs(3729) <= not(layer0_outputs(3557));
    outputs(3730) <= (layer0_outputs(884)) and not (layer0_outputs(4633));
    outputs(3731) <= layer0_outputs(637);
    outputs(3732) <= not((layer0_outputs(4916)) or (layer0_outputs(1221)));
    outputs(3733) <= not(layer0_outputs(180)) or (layer0_outputs(58));
    outputs(3734) <= layer0_outputs(4621);
    outputs(3735) <= not(layer0_outputs(2295));
    outputs(3736) <= (layer0_outputs(1519)) xor (layer0_outputs(4453));
    outputs(3737) <= not(layer0_outputs(4812));
    outputs(3738) <= (layer0_outputs(4315)) and not (layer0_outputs(4668));
    outputs(3739) <= not(layer0_outputs(7));
    outputs(3740) <= not((layer0_outputs(4332)) xor (layer0_outputs(4821)));
    outputs(3741) <= layer0_outputs(2998);
    outputs(3742) <= layer0_outputs(2696);
    outputs(3743) <= not(layer0_outputs(4614));
    outputs(3744) <= not(layer0_outputs(875));
    outputs(3745) <= layer0_outputs(344);
    outputs(3746) <= not((layer0_outputs(3645)) xor (layer0_outputs(4400)));
    outputs(3747) <= not(layer0_outputs(375)) or (layer0_outputs(2138));
    outputs(3748) <= (layer0_outputs(559)) and not (layer0_outputs(856));
    outputs(3749) <= (layer0_outputs(3996)) xor (layer0_outputs(2540));
    outputs(3750) <= (layer0_outputs(3323)) xor (layer0_outputs(1533));
    outputs(3751) <= not((layer0_outputs(4217)) xor (layer0_outputs(1477)));
    outputs(3752) <= (layer0_outputs(4181)) xor (layer0_outputs(1007));
    outputs(3753) <= (layer0_outputs(4544)) or (layer0_outputs(346));
    outputs(3754) <= (layer0_outputs(1992)) and not (layer0_outputs(2333));
    outputs(3755) <= (layer0_outputs(4531)) and (layer0_outputs(3412));
    outputs(3756) <= layer0_outputs(4389);
    outputs(3757) <= not((layer0_outputs(1289)) and (layer0_outputs(1394)));
    outputs(3758) <= '0';
    outputs(3759) <= layer0_outputs(4565);
    outputs(3760) <= not(layer0_outputs(4385));
    outputs(3761) <= (layer0_outputs(1580)) and (layer0_outputs(5069));
    outputs(3762) <= not((layer0_outputs(618)) xor (layer0_outputs(3941)));
    outputs(3763) <= (layer0_outputs(247)) and not (layer0_outputs(1267));
    outputs(3764) <= (layer0_outputs(2754)) xor (layer0_outputs(3524));
    outputs(3765) <= layer0_outputs(4132);
    outputs(3766) <= (layer0_outputs(4251)) and (layer0_outputs(575));
    outputs(3767) <= (layer0_outputs(1150)) and not (layer0_outputs(498));
    outputs(3768) <= not(layer0_outputs(2459));
    outputs(3769) <= layer0_outputs(788);
    outputs(3770) <= layer0_outputs(973);
    outputs(3771) <= not((layer0_outputs(2670)) xor (layer0_outputs(4345)));
    outputs(3772) <= (layer0_outputs(4588)) or (layer0_outputs(2331));
    outputs(3773) <= not((layer0_outputs(4608)) or (layer0_outputs(2841)));
    outputs(3774) <= not((layer0_outputs(1613)) or (layer0_outputs(100)));
    outputs(3775) <= not(layer0_outputs(2369));
    outputs(3776) <= layer0_outputs(451);
    outputs(3777) <= not((layer0_outputs(2433)) or (layer0_outputs(2794)));
    outputs(3778) <= not(layer0_outputs(3039));
    outputs(3779) <= not((layer0_outputs(3385)) or (layer0_outputs(4613)));
    outputs(3780) <= layer0_outputs(4184);
    outputs(3781) <= (layer0_outputs(4340)) and (layer0_outputs(2952));
    outputs(3782) <= (layer0_outputs(2425)) and (layer0_outputs(3840));
    outputs(3783) <= not(layer0_outputs(4474)) or (layer0_outputs(2334));
    outputs(3784) <= not(layer0_outputs(2888));
    outputs(3785) <= not(layer0_outputs(4253));
    outputs(3786) <= (layer0_outputs(1600)) and not (layer0_outputs(1326));
    outputs(3787) <= (layer0_outputs(4598)) xor (layer0_outputs(2969));
    outputs(3788) <= layer0_outputs(4735);
    outputs(3789) <= (layer0_outputs(138)) xor (layer0_outputs(2946));
    outputs(3790) <= (layer0_outputs(1083)) and (layer0_outputs(2021));
    outputs(3791) <= (layer0_outputs(256)) and not (layer0_outputs(2275));
    outputs(3792) <= (layer0_outputs(2578)) xor (layer0_outputs(4688));
    outputs(3793) <= not((layer0_outputs(376)) or (layer0_outputs(2411)));
    outputs(3794) <= layer0_outputs(685);
    outputs(3795) <= not(layer0_outputs(3145));
    outputs(3796) <= not(layer0_outputs(1996)) or (layer0_outputs(407));
    outputs(3797) <= (layer0_outputs(264)) and not (layer0_outputs(4167));
    outputs(3798) <= (layer0_outputs(510)) and not (layer0_outputs(2695));
    outputs(3799) <= not(layer0_outputs(147));
    outputs(3800) <= not((layer0_outputs(1708)) xor (layer0_outputs(4738)));
    outputs(3801) <= not(layer0_outputs(3160));
    outputs(3802) <= not((layer0_outputs(2597)) or (layer0_outputs(4835)));
    outputs(3803) <= layer0_outputs(4792);
    outputs(3804) <= not(layer0_outputs(2350));
    outputs(3805) <= not(layer0_outputs(4388));
    outputs(3806) <= not(layer0_outputs(640)) or (layer0_outputs(114));
    outputs(3807) <= (layer0_outputs(251)) and not (layer0_outputs(1704));
    outputs(3808) <= not(layer0_outputs(4561));
    outputs(3809) <= (layer0_outputs(964)) and (layer0_outputs(934));
    outputs(3810) <= layer0_outputs(1258);
    outputs(3811) <= not((layer0_outputs(1923)) xor (layer0_outputs(3619)));
    outputs(3812) <= (layer0_outputs(2421)) and not (layer0_outputs(5076));
    outputs(3813) <= (layer0_outputs(3271)) and (layer0_outputs(892));
    outputs(3814) <= not((layer0_outputs(2123)) xor (layer0_outputs(832)));
    outputs(3815) <= not((layer0_outputs(3797)) xor (layer0_outputs(1763)));
    outputs(3816) <= not((layer0_outputs(2376)) xor (layer0_outputs(2426)));
    outputs(3817) <= not((layer0_outputs(4189)) xor (layer0_outputs(3981)));
    outputs(3818) <= (layer0_outputs(4064)) xor (layer0_outputs(4298));
    outputs(3819) <= not(layer0_outputs(1056));
    outputs(3820) <= layer0_outputs(3584);
    outputs(3821) <= (layer0_outputs(1064)) and (layer0_outputs(4421));
    outputs(3822) <= not((layer0_outputs(2680)) xor (layer0_outputs(474)));
    outputs(3823) <= not(layer0_outputs(3357));
    outputs(3824) <= (layer0_outputs(3673)) and (layer0_outputs(4357));
    outputs(3825) <= not((layer0_outputs(3965)) or (layer0_outputs(3556)));
    outputs(3826) <= (layer0_outputs(1713)) xor (layer0_outputs(4643));
    outputs(3827) <= (layer0_outputs(3755)) xor (layer0_outputs(3413));
    outputs(3828) <= (layer0_outputs(2774)) and not (layer0_outputs(3664));
    outputs(3829) <= (layer0_outputs(2606)) and not (layer0_outputs(3321));
    outputs(3830) <= (layer0_outputs(4085)) xor (layer0_outputs(3443));
    outputs(3831) <= not((layer0_outputs(4445)) or (layer0_outputs(3722)));
    outputs(3832) <= not(layer0_outputs(4931));
    outputs(3833) <= (layer0_outputs(2410)) xor (layer0_outputs(3378));
    outputs(3834) <= layer0_outputs(451);
    outputs(3835) <= layer0_outputs(420);
    outputs(3836) <= not(layer0_outputs(1764));
    outputs(3837) <= (layer0_outputs(4626)) xor (layer0_outputs(3823));
    outputs(3838) <= (layer0_outputs(527)) xor (layer0_outputs(2184));
    outputs(3839) <= not(layer0_outputs(1899)) or (layer0_outputs(3378));
    outputs(3840) <= (layer0_outputs(561)) or (layer0_outputs(3692));
    outputs(3841) <= layer0_outputs(3498);
    outputs(3842) <= layer0_outputs(2359);
    outputs(3843) <= not((layer0_outputs(1966)) xor (layer0_outputs(1094)));
    outputs(3844) <= not(layer0_outputs(749));
    outputs(3845) <= (layer0_outputs(2007)) xor (layer0_outputs(4181));
    outputs(3846) <= layer0_outputs(1126);
    outputs(3847) <= layer0_outputs(800);
    outputs(3848) <= not((layer0_outputs(495)) and (layer0_outputs(4325)));
    outputs(3849) <= (layer0_outputs(365)) and (layer0_outputs(1114));
    outputs(3850) <= (layer0_outputs(4823)) xor (layer0_outputs(4993));
    outputs(3851) <= (layer0_outputs(4362)) and not (layer0_outputs(3853));
    outputs(3852) <= not(layer0_outputs(3036));
    outputs(3853) <= not(layer0_outputs(701));
    outputs(3854) <= (layer0_outputs(3766)) and not (layer0_outputs(244));
    outputs(3855) <= not((layer0_outputs(4566)) or (layer0_outputs(2293)));
    outputs(3856) <= (layer0_outputs(66)) or (layer0_outputs(4951));
    outputs(3857) <= (layer0_outputs(3197)) and not (layer0_outputs(574));
    outputs(3858) <= layer0_outputs(218);
    outputs(3859) <= layer0_outputs(933);
    outputs(3860) <= not((layer0_outputs(3496)) xor (layer0_outputs(74)));
    outputs(3861) <= not((layer0_outputs(4252)) xor (layer0_outputs(4975)));
    outputs(3862) <= (layer0_outputs(3127)) or (layer0_outputs(2196));
    outputs(3863) <= (layer0_outputs(1040)) xor (layer0_outputs(2850));
    outputs(3864) <= not((layer0_outputs(3707)) or (layer0_outputs(870)));
    outputs(3865) <= (layer0_outputs(692)) and not (layer0_outputs(4921));
    outputs(3866) <= layer0_outputs(3071);
    outputs(3867) <= not(layer0_outputs(2716));
    outputs(3868) <= (layer0_outputs(4697)) and (layer0_outputs(4251));
    outputs(3869) <= not(layer0_outputs(2549));
    outputs(3870) <= layer0_outputs(1808);
    outputs(3871) <= layer0_outputs(3779);
    outputs(3872) <= (layer0_outputs(265)) and not (layer0_outputs(412));
    outputs(3873) <= not(layer0_outputs(3726));
    outputs(3874) <= (layer0_outputs(4117)) and not (layer0_outputs(2485));
    outputs(3875) <= not(layer0_outputs(1184)) or (layer0_outputs(502));
    outputs(3876) <= (layer0_outputs(4279)) and not (layer0_outputs(1648));
    outputs(3877) <= not((layer0_outputs(4393)) or (layer0_outputs(27)));
    outputs(3878) <= not(layer0_outputs(3456)) or (layer0_outputs(2089));
    outputs(3879) <= (layer0_outputs(1298)) xor (layer0_outputs(2462));
    outputs(3880) <= not((layer0_outputs(4987)) xor (layer0_outputs(1414)));
    outputs(3881) <= not(layer0_outputs(3256));
    outputs(3882) <= not((layer0_outputs(1741)) xor (layer0_outputs(71)));
    outputs(3883) <= not(layer0_outputs(4174));
    outputs(3884) <= layer0_outputs(2629);
    outputs(3885) <= (layer0_outputs(5058)) xor (layer0_outputs(4031));
    outputs(3886) <= not((layer0_outputs(1782)) xor (layer0_outputs(1523)));
    outputs(3887) <= layer0_outputs(409);
    outputs(3888) <= (layer0_outputs(2627)) and not (layer0_outputs(2718));
    outputs(3889) <= (layer0_outputs(123)) xor (layer0_outputs(2594));
    outputs(3890) <= layer0_outputs(1355);
    outputs(3891) <= not(layer0_outputs(1597));
    outputs(3892) <= (layer0_outputs(382)) and (layer0_outputs(2811));
    outputs(3893) <= layer0_outputs(1997);
    outputs(3894) <= not((layer0_outputs(904)) or (layer0_outputs(1192)));
    outputs(3895) <= layer0_outputs(4511);
    outputs(3896) <= not((layer0_outputs(2413)) or (layer0_outputs(3529)));
    outputs(3897) <= (layer0_outputs(4869)) and (layer0_outputs(265));
    outputs(3898) <= (layer0_outputs(5028)) xor (layer0_outputs(3447));
    outputs(3899) <= not(layer0_outputs(155));
    outputs(3900) <= not(layer0_outputs(1334));
    outputs(3901) <= (layer0_outputs(1993)) xor (layer0_outputs(2060));
    outputs(3902) <= layer0_outputs(261);
    outputs(3903) <= layer0_outputs(2266);
    outputs(3904) <= not((layer0_outputs(4236)) or (layer0_outputs(4102)));
    outputs(3905) <= not(layer0_outputs(1985)) or (layer0_outputs(3873));
    outputs(3906) <= not(layer0_outputs(4890));
    outputs(3907) <= layer0_outputs(3304);
    outputs(3908) <= (layer0_outputs(1890)) xor (layer0_outputs(4187));
    outputs(3909) <= layer0_outputs(40);
    outputs(3910) <= layer0_outputs(3449);
    outputs(3911) <= layer0_outputs(4333);
    outputs(3912) <= (layer0_outputs(3218)) and not (layer0_outputs(3885));
    outputs(3913) <= layer0_outputs(2101);
    outputs(3914) <= (layer0_outputs(5015)) and not (layer0_outputs(2676));
    outputs(3915) <= (layer0_outputs(755)) and not (layer0_outputs(4845));
    outputs(3916) <= not(layer0_outputs(1717));
    outputs(3917) <= layer0_outputs(2647);
    outputs(3918) <= (layer0_outputs(4926)) and (layer0_outputs(413));
    outputs(3919) <= layer0_outputs(2396);
    outputs(3920) <= layer0_outputs(1934);
    outputs(3921) <= not(layer0_outputs(2215));
    outputs(3922) <= (layer0_outputs(1863)) xor (layer0_outputs(1008));
    outputs(3923) <= not(layer0_outputs(3783));
    outputs(3924) <= (layer0_outputs(1560)) and not (layer0_outputs(2587));
    outputs(3925) <= not(layer0_outputs(2172)) or (layer0_outputs(4070));
    outputs(3926) <= (layer0_outputs(4752)) and not (layer0_outputs(389));
    outputs(3927) <= (layer0_outputs(4320)) and not (layer0_outputs(2503));
    outputs(3928) <= not(layer0_outputs(4408));
    outputs(3929) <= not(layer0_outputs(215));
    outputs(3930) <= (layer0_outputs(2196)) or (layer0_outputs(4810));
    outputs(3931) <= (layer0_outputs(2518)) and (layer0_outputs(3975));
    outputs(3932) <= (layer0_outputs(3630)) and not (layer0_outputs(3038));
    outputs(3933) <= not(layer0_outputs(4081)) or (layer0_outputs(2010));
    outputs(3934) <= (layer0_outputs(3689)) xor (layer0_outputs(4575));
    outputs(3935) <= layer0_outputs(4195);
    outputs(3936) <= not((layer0_outputs(535)) xor (layer0_outputs(959)));
    outputs(3937) <= not(layer0_outputs(781));
    outputs(3938) <= not((layer0_outputs(3015)) or (layer0_outputs(2469)));
    outputs(3939) <= (layer0_outputs(1555)) xor (layer0_outputs(3309));
    outputs(3940) <= not((layer0_outputs(2524)) or (layer0_outputs(76)));
    outputs(3941) <= (layer0_outputs(1207)) and not (layer0_outputs(3207));
    outputs(3942) <= not((layer0_outputs(2179)) or (layer0_outputs(780)));
    outputs(3943) <= not((layer0_outputs(3168)) xor (layer0_outputs(1026)));
    outputs(3944) <= (layer0_outputs(1629)) xor (layer0_outputs(2085));
    outputs(3945) <= layer0_outputs(4242);
    outputs(3946) <= (layer0_outputs(3495)) and not (layer0_outputs(4194));
    outputs(3947) <= (layer0_outputs(1257)) xor (layer0_outputs(1196));
    outputs(3948) <= (layer0_outputs(2533)) and (layer0_outputs(2926));
    outputs(3949) <= layer0_outputs(4947);
    outputs(3950) <= (layer0_outputs(3603)) and not (layer0_outputs(4174));
    outputs(3951) <= (layer0_outputs(395)) and (layer0_outputs(4522));
    outputs(3952) <= not((layer0_outputs(3459)) xor (layer0_outputs(3255)));
    outputs(3953) <= (layer0_outputs(3630)) xor (layer0_outputs(2137));
    outputs(3954) <= (layer0_outputs(3458)) and not (layer0_outputs(415));
    outputs(3955) <= (layer0_outputs(4216)) and not (layer0_outputs(5114));
    outputs(3956) <= not(layer0_outputs(913));
    outputs(3957) <= '0';
    outputs(3958) <= not(layer0_outputs(3688));
    outputs(3959) <= layer0_outputs(1861);
    outputs(3960) <= (layer0_outputs(3835)) and (layer0_outputs(4235));
    outputs(3961) <= not((layer0_outputs(3242)) xor (layer0_outputs(2821)));
    outputs(3962) <= not((layer0_outputs(3048)) xor (layer0_outputs(2470)));
    outputs(3963) <= not(layer0_outputs(2634));
    outputs(3964) <= not((layer0_outputs(2248)) xor (layer0_outputs(4564)));
    outputs(3965) <= (layer0_outputs(4192)) xor (layer0_outputs(2443));
    outputs(3966) <= layer0_outputs(3618);
    outputs(3967) <= layer0_outputs(2975);
    outputs(3968) <= not((layer0_outputs(2032)) xor (layer0_outputs(3739)));
    outputs(3969) <= not(layer0_outputs(2292));
    outputs(3970) <= layer0_outputs(93);
    outputs(3971) <= not((layer0_outputs(625)) xor (layer0_outputs(1205)));
    outputs(3972) <= (layer0_outputs(4777)) and (layer0_outputs(1303));
    outputs(3973) <= not((layer0_outputs(3162)) xor (layer0_outputs(4026)));
    outputs(3974) <= not(layer0_outputs(1912));
    outputs(3975) <= layer0_outputs(744);
    outputs(3976) <= not(layer0_outputs(4058));
    outputs(3977) <= (layer0_outputs(1222)) and not (layer0_outputs(5071));
    outputs(3978) <= not(layer0_outputs(3578)) or (layer0_outputs(2590));
    outputs(3979) <= not(layer0_outputs(4942));
    outputs(3980) <= not(layer0_outputs(540));
    outputs(3981) <= layer0_outputs(1758);
    outputs(3982) <= not((layer0_outputs(1652)) and (layer0_outputs(1193)));
    outputs(3983) <= not(layer0_outputs(5033));
    outputs(3984) <= not((layer0_outputs(2287)) xor (layer0_outputs(3159)));
    outputs(3985) <= not(layer0_outputs(1268)) or (layer0_outputs(70));
    outputs(3986) <= (layer0_outputs(1682)) xor (layer0_outputs(320));
    outputs(3987) <= layer0_outputs(3796);
    outputs(3988) <= not(layer0_outputs(1565));
    outputs(3989) <= not(layer0_outputs(4434));
    outputs(3990) <= layer0_outputs(3079);
    outputs(3991) <= (layer0_outputs(3943)) and not (layer0_outputs(5032));
    outputs(3992) <= not(layer0_outputs(4168));
    outputs(3993) <= (layer0_outputs(5009)) and (layer0_outputs(232));
    outputs(3994) <= layer0_outputs(2675);
    outputs(3995) <= (layer0_outputs(4446)) and not (layer0_outputs(2335));
    outputs(3996) <= not((layer0_outputs(543)) xor (layer0_outputs(5028)));
    outputs(3997) <= not(layer0_outputs(3268));
    outputs(3998) <= layer0_outputs(1698);
    outputs(3999) <= (layer0_outputs(2496)) xor (layer0_outputs(3738));
    outputs(4000) <= layer0_outputs(1282);
    outputs(4001) <= not((layer0_outputs(4377)) xor (layer0_outputs(3438)));
    outputs(4002) <= (layer0_outputs(2808)) and (layer0_outputs(4373));
    outputs(4003) <= (layer0_outputs(2255)) and not (layer0_outputs(4966));
    outputs(4004) <= layer0_outputs(299);
    outputs(4005) <= not(layer0_outputs(901));
    outputs(4006) <= not(layer0_outputs(2105));
    outputs(4007) <= (layer0_outputs(3839)) xor (layer0_outputs(2384));
    outputs(4008) <= (layer0_outputs(3804)) xor (layer0_outputs(1291));
    outputs(4009) <= (layer0_outputs(3356)) xor (layer0_outputs(3833));
    outputs(4010) <= not((layer0_outputs(1304)) or (layer0_outputs(4155)));
    outputs(4011) <= not((layer0_outputs(2092)) or (layer0_outputs(1359)));
    outputs(4012) <= (layer0_outputs(4442)) and not (layer0_outputs(2039));
    outputs(4013) <= not(layer0_outputs(458));
    outputs(4014) <= not((layer0_outputs(4709)) xor (layer0_outputs(1412)));
    outputs(4015) <= (layer0_outputs(3274)) and not (layer0_outputs(1702));
    outputs(4016) <= not(layer0_outputs(1022));
    outputs(4017) <= (layer0_outputs(4281)) and not (layer0_outputs(955));
    outputs(4018) <= layer0_outputs(4379);
    outputs(4019) <= (layer0_outputs(2243)) xor (layer0_outputs(2065));
    outputs(4020) <= not(layer0_outputs(4594));
    outputs(4021) <= not(layer0_outputs(2612));
    outputs(4022) <= not(layer0_outputs(862));
    outputs(4023) <= (layer0_outputs(4960)) and not (layer0_outputs(5098));
    outputs(4024) <= not((layer0_outputs(513)) and (layer0_outputs(5073)));
    outputs(4025) <= layer0_outputs(3656);
    outputs(4026) <= (layer0_outputs(4221)) xor (layer0_outputs(1593));
    outputs(4027) <= (layer0_outputs(923)) and (layer0_outputs(2119));
    outputs(4028) <= (layer0_outputs(2217)) and (layer0_outputs(4222));
    outputs(4029) <= not(layer0_outputs(4461));
    outputs(4030) <= not((layer0_outputs(1670)) or (layer0_outputs(3516)));
    outputs(4031) <= not(layer0_outputs(2515)) or (layer0_outputs(2904));
    outputs(4032) <= layer0_outputs(2210);
    outputs(4033) <= layer0_outputs(1424);
    outputs(4034) <= not((layer0_outputs(4688)) xor (layer0_outputs(4674)));
    outputs(4035) <= layer0_outputs(1361);
    outputs(4036) <= layer0_outputs(80);
    outputs(4037) <= (layer0_outputs(1692)) and not (layer0_outputs(3208));
    outputs(4038) <= not(layer0_outputs(5099));
    outputs(4039) <= (layer0_outputs(1010)) and not (layer0_outputs(1750));
    outputs(4040) <= '0';
    outputs(4041) <= not(layer0_outputs(1511));
    outputs(4042) <= layer0_outputs(5103);
    outputs(4043) <= not((layer0_outputs(4770)) or (layer0_outputs(2799)));
    outputs(4044) <= not((layer0_outputs(2967)) xor (layer0_outputs(1192)));
    outputs(4045) <= (layer0_outputs(1658)) and not (layer0_outputs(4633));
    outputs(4046) <= layer0_outputs(3386);
    outputs(4047) <= not(layer0_outputs(1855));
    outputs(4048) <= not(layer0_outputs(4190));
    outputs(4049) <= not(layer0_outputs(2710)) or (layer0_outputs(653));
    outputs(4050) <= (layer0_outputs(744)) and (layer0_outputs(3972));
    outputs(4051) <= (layer0_outputs(4619)) and (layer0_outputs(4593));
    outputs(4052) <= layer0_outputs(4467);
    outputs(4053) <= not(layer0_outputs(1541));
    outputs(4054) <= not(layer0_outputs(3328));
    outputs(4055) <= not((layer0_outputs(797)) xor (layer0_outputs(2933)));
    outputs(4056) <= '0';
    outputs(4057) <= layer0_outputs(1510);
    outputs(4058) <= (layer0_outputs(1759)) or (layer0_outputs(1632));
    outputs(4059) <= layer0_outputs(3807);
    outputs(4060) <= (layer0_outputs(1601)) and not (layer0_outputs(1322));
    outputs(4061) <= not(layer0_outputs(778));
    outputs(4062) <= (layer0_outputs(3013)) and not (layer0_outputs(3107));
    outputs(4063) <= not(layer0_outputs(3817));
    outputs(4064) <= layer0_outputs(2887);
    outputs(4065) <= (layer0_outputs(731)) xor (layer0_outputs(1778));
    outputs(4066) <= not(layer0_outputs(2599));
    outputs(4067) <= not((layer0_outputs(4973)) and (layer0_outputs(5000)));
    outputs(4068) <= (layer0_outputs(1547)) xor (layer0_outputs(4995));
    outputs(4069) <= (layer0_outputs(2158)) and not (layer0_outputs(250));
    outputs(4070) <= not((layer0_outputs(280)) xor (layer0_outputs(2940)));
    outputs(4071) <= layer0_outputs(1570);
    outputs(4072) <= layer0_outputs(1145);
    outputs(4073) <= (layer0_outputs(4950)) and (layer0_outputs(2142));
    outputs(4074) <= not(layer0_outputs(521));
    outputs(4075) <= not(layer0_outputs(3368));
    outputs(4076) <= not(layer0_outputs(1069));
    outputs(4077) <= not((layer0_outputs(4542)) or (layer0_outputs(3785)));
    outputs(4078) <= not((layer0_outputs(2786)) or (layer0_outputs(4270)));
    outputs(4079) <= layer0_outputs(2396);
    outputs(4080) <= (layer0_outputs(3059)) and not (layer0_outputs(2660));
    outputs(4081) <= not(layer0_outputs(252));
    outputs(4082) <= not((layer0_outputs(1434)) or (layer0_outputs(1013)));
    outputs(4083) <= not(layer0_outputs(3896)) or (layer0_outputs(4999));
    outputs(4084) <= not(layer0_outputs(329));
    outputs(4085) <= layer0_outputs(3906);
    outputs(4086) <= (layer0_outputs(13)) xor (layer0_outputs(2285));
    outputs(4087) <= not((layer0_outputs(4540)) xor (layer0_outputs(116)));
    outputs(4088) <= layer0_outputs(163);
    outputs(4089) <= (layer0_outputs(3580)) and not (layer0_outputs(147));
    outputs(4090) <= (layer0_outputs(506)) or (layer0_outputs(1545));
    outputs(4091) <= not((layer0_outputs(411)) or (layer0_outputs(3519)));
    outputs(4092) <= (layer0_outputs(2244)) and (layer0_outputs(3956));
    outputs(4093) <= layer0_outputs(1630);
    outputs(4094) <= not((layer0_outputs(4010)) or (layer0_outputs(4023)));
    outputs(4095) <= (layer0_outputs(4963)) and (layer0_outputs(1585));
    outputs(4096) <= not((layer0_outputs(5067)) or (layer0_outputs(3829)));
    outputs(4097) <= not(layer0_outputs(1134));
    outputs(4098) <= (layer0_outputs(5)) and not (layer0_outputs(481));
    outputs(4099) <= not(layer0_outputs(954));
    outputs(4100) <= layer0_outputs(351);
    outputs(4101) <= not(layer0_outputs(4825));
    outputs(4102) <= layer0_outputs(2488);
    outputs(4103) <= (layer0_outputs(4905)) xor (layer0_outputs(1889));
    outputs(4104) <= not(layer0_outputs(3950));
    outputs(4105) <= not((layer0_outputs(4294)) xor (layer0_outputs(1309)));
    outputs(4106) <= layer0_outputs(2073);
    outputs(4107) <= (layer0_outputs(2979)) and not (layer0_outputs(752));
    outputs(4108) <= not((layer0_outputs(1914)) xor (layer0_outputs(4533)));
    outputs(4109) <= (layer0_outputs(3654)) or (layer0_outputs(1680));
    outputs(4110) <= (layer0_outputs(229)) and not (layer0_outputs(2386));
    outputs(4111) <= not(layer0_outputs(4543)) or (layer0_outputs(3789));
    outputs(4112) <= not(layer0_outputs(4438)) or (layer0_outputs(3319));
    outputs(4113) <= (layer0_outputs(2085)) and not (layer0_outputs(4405));
    outputs(4114) <= not(layer0_outputs(4933)) or (layer0_outputs(3078));
    outputs(4115) <= not(layer0_outputs(4247));
    outputs(4116) <= (layer0_outputs(1346)) or (layer0_outputs(3635));
    outputs(4117) <= not(layer0_outputs(3983));
    outputs(4118) <= (layer0_outputs(3874)) and not (layer0_outputs(870));
    outputs(4119) <= (layer0_outputs(4338)) and (layer0_outputs(3340));
    outputs(4120) <= layer0_outputs(2006);
    outputs(4121) <= not(layer0_outputs(4534));
    outputs(4122) <= not(layer0_outputs(707));
    outputs(4123) <= (layer0_outputs(4694)) xor (layer0_outputs(4463));
    outputs(4124) <= (layer0_outputs(3452)) or (layer0_outputs(3143));
    outputs(4125) <= (layer0_outputs(1765)) and (layer0_outputs(2507));
    outputs(4126) <= not((layer0_outputs(3120)) xor (layer0_outputs(1435)));
    outputs(4127) <= not(layer0_outputs(4712));
    outputs(4128) <= (layer0_outputs(2784)) and (layer0_outputs(1012));
    outputs(4129) <= not(layer0_outputs(646));
    outputs(4130) <= layer0_outputs(421);
    outputs(4131) <= not(layer0_outputs(2668));
    outputs(4132) <= (layer0_outputs(1804)) xor (layer0_outputs(1677));
    outputs(4133) <= not(layer0_outputs(981)) or (layer0_outputs(1986));
    outputs(4134) <= (layer0_outputs(71)) or (layer0_outputs(2875));
    outputs(4135) <= '1';
    outputs(4136) <= layer0_outputs(3469);
    outputs(4137) <= not(layer0_outputs(1352));
    outputs(4138) <= not(layer0_outputs(881)) or (layer0_outputs(2970));
    outputs(4139) <= not((layer0_outputs(396)) and (layer0_outputs(1677)));
    outputs(4140) <= (layer0_outputs(644)) or (layer0_outputs(3911));
    outputs(4141) <= not(layer0_outputs(815));
    outputs(4142) <= (layer0_outputs(1204)) and not (layer0_outputs(4323));
    outputs(4143) <= layer0_outputs(4607);
    outputs(4144) <= not(layer0_outputs(4853)) or (layer0_outputs(3651));
    outputs(4145) <= not(layer0_outputs(638));
    outputs(4146) <= layer0_outputs(1266);
    outputs(4147) <= not((layer0_outputs(1916)) xor (layer0_outputs(3959)));
    outputs(4148) <= not(layer0_outputs(4961));
    outputs(4149) <= layer0_outputs(4331);
    outputs(4150) <= layer0_outputs(443);
    outputs(4151) <= '1';
    outputs(4152) <= layer0_outputs(2909);
    outputs(4153) <= (layer0_outputs(33)) and (layer0_outputs(1091));
    outputs(4154) <= not(layer0_outputs(1840)) or (layer0_outputs(3275));
    outputs(4155) <= not(layer0_outputs(2951)) or (layer0_outputs(2000));
    outputs(4156) <= not(layer0_outputs(5088)) or (layer0_outputs(680));
    outputs(4157) <= not((layer0_outputs(634)) or (layer0_outputs(1830)));
    outputs(4158) <= not((layer0_outputs(4606)) xor (layer0_outputs(4997)));
    outputs(4159) <= not(layer0_outputs(3374)) or (layer0_outputs(2475));
    outputs(4160) <= layer0_outputs(2415);
    outputs(4161) <= not(layer0_outputs(2287));
    outputs(4162) <= not(layer0_outputs(2629));
    outputs(4163) <= (layer0_outputs(4156)) and not (layer0_outputs(202));
    outputs(4164) <= not((layer0_outputs(3047)) or (layer0_outputs(391)));
    outputs(4165) <= not(layer0_outputs(1501)) or (layer0_outputs(2733));
    outputs(4166) <= (layer0_outputs(695)) xor (layer0_outputs(5098));
    outputs(4167) <= not((layer0_outputs(3228)) or (layer0_outputs(2290)));
    outputs(4168) <= (layer0_outputs(924)) or (layer0_outputs(2768));
    outputs(4169) <= not(layer0_outputs(305));
    outputs(4170) <= (layer0_outputs(2432)) and not (layer0_outputs(1434));
    outputs(4171) <= layer0_outputs(2749);
    outputs(4172) <= (layer0_outputs(1564)) and (layer0_outputs(1542));
    outputs(4173) <= layer0_outputs(1116);
    outputs(4174) <= (layer0_outputs(4741)) xor (layer0_outputs(3364));
    outputs(4175) <= (layer0_outputs(1866)) and (layer0_outputs(1395));
    outputs(4176) <= not((layer0_outputs(3217)) xor (layer0_outputs(3399)));
    outputs(4177) <= layer0_outputs(4766);
    outputs(4178) <= not((layer0_outputs(891)) xor (layer0_outputs(4791)));
    outputs(4179) <= not(layer0_outputs(3004));
    outputs(4180) <= not((layer0_outputs(735)) xor (layer0_outputs(1977)));
    outputs(4181) <= (layer0_outputs(2573)) and not (layer0_outputs(4062));
    outputs(4182) <= not((layer0_outputs(4715)) or (layer0_outputs(419)));
    outputs(4183) <= (layer0_outputs(1868)) xor (layer0_outputs(4534));
    outputs(4184) <= layer0_outputs(1714);
    outputs(4185) <= layer0_outputs(4353);
    outputs(4186) <= not((layer0_outputs(4149)) or (layer0_outputs(4203)));
    outputs(4187) <= (layer0_outputs(2964)) or (layer0_outputs(276));
    outputs(4188) <= layer0_outputs(289);
    outputs(4189) <= layer0_outputs(3055);
    outputs(4190) <= (layer0_outputs(768)) and not (layer0_outputs(4275));
    outputs(4191) <= (layer0_outputs(2100)) xor (layer0_outputs(16));
    outputs(4192) <= not((layer0_outputs(1767)) xor (layer0_outputs(2604)));
    outputs(4193) <= layer0_outputs(1432);
    outputs(4194) <= layer0_outputs(142);
    outputs(4195) <= not(layer0_outputs(2792));
    outputs(4196) <= layer0_outputs(4336);
    outputs(4197) <= layer0_outputs(378);
    outputs(4198) <= not(layer0_outputs(2871));
    outputs(4199) <= not(layer0_outputs(3051)) or (layer0_outputs(194));
    outputs(4200) <= not((layer0_outputs(911)) and (layer0_outputs(5074)));
    outputs(4201) <= (layer0_outputs(2807)) and not (layer0_outputs(3361));
    outputs(4202) <= layer0_outputs(10);
    outputs(4203) <= not(layer0_outputs(647));
    outputs(4204) <= not(layer0_outputs(2504)) or (layer0_outputs(3441));
    outputs(4205) <= not(layer0_outputs(4140)) or (layer0_outputs(2702));
    outputs(4206) <= layer0_outputs(3855);
    outputs(4207) <= not(layer0_outputs(5113));
    outputs(4208) <= layer0_outputs(2075);
    outputs(4209) <= (layer0_outputs(1964)) and (layer0_outputs(150));
    outputs(4210) <= (layer0_outputs(1296)) xor (layer0_outputs(2292));
    outputs(4211) <= (layer0_outputs(1620)) and not (layer0_outputs(4601));
    outputs(4212) <= (layer0_outputs(2936)) xor (layer0_outputs(4371));
    outputs(4213) <= layer0_outputs(115);
    outputs(4214) <= not((layer0_outputs(1265)) and (layer0_outputs(3513)));
    outputs(4215) <= layer0_outputs(3795);
    outputs(4216) <= not(layer0_outputs(2789));
    outputs(4217) <= (layer0_outputs(5094)) xor (layer0_outputs(3454));
    outputs(4218) <= not((layer0_outputs(4019)) and (layer0_outputs(442)));
    outputs(4219) <= not(layer0_outputs(865));
    outputs(4220) <= (layer0_outputs(2593)) or (layer0_outputs(3624));
    outputs(4221) <= layer0_outputs(1155);
    outputs(4222) <= not((layer0_outputs(2450)) and (layer0_outputs(991)));
    outputs(4223) <= not((layer0_outputs(2229)) xor (layer0_outputs(2339)));
    outputs(4224) <= not(layer0_outputs(2492)) or (layer0_outputs(4737));
    outputs(4225) <= not(layer0_outputs(2505));
    outputs(4226) <= layer0_outputs(2596);
    outputs(4227) <= not(layer0_outputs(4575));
    outputs(4228) <= not(layer0_outputs(112)) or (layer0_outputs(1922));
    outputs(4229) <= (layer0_outputs(1863)) or (layer0_outputs(4415));
    outputs(4230) <= not(layer0_outputs(2107));
    outputs(4231) <= layer0_outputs(55);
    outputs(4232) <= layer0_outputs(1097);
    outputs(4233) <= layer0_outputs(198);
    outputs(4234) <= not(layer0_outputs(4152));
    outputs(4235) <= layer0_outputs(3732);
    outputs(4236) <= layer0_outputs(4984);
    outputs(4237) <= not(layer0_outputs(2606));
    outputs(4238) <= layer0_outputs(273);
    outputs(4239) <= layer0_outputs(4477);
    outputs(4240) <= layer0_outputs(789);
    outputs(4241) <= not((layer0_outputs(4004)) and (layer0_outputs(1942)));
    outputs(4242) <= not(layer0_outputs(166));
    outputs(4243) <= not(layer0_outputs(3264));
    outputs(4244) <= not((layer0_outputs(2603)) and (layer0_outputs(3558)));
    outputs(4245) <= not(layer0_outputs(783));
    outputs(4246) <= not(layer0_outputs(1873));
    outputs(4247) <= not(layer0_outputs(3248));
    outputs(4248) <= (layer0_outputs(3053)) xor (layer0_outputs(1609));
    outputs(4249) <= not((layer0_outputs(4634)) or (layer0_outputs(3501)));
    outputs(4250) <= (layer0_outputs(2667)) xor (layer0_outputs(33));
    outputs(4251) <= not(layer0_outputs(1027));
    outputs(4252) <= not(layer0_outputs(889)) or (layer0_outputs(3414));
    outputs(4253) <= (layer0_outputs(2851)) or (layer0_outputs(1579));
    outputs(4254) <= not((layer0_outputs(594)) or (layer0_outputs(458)));
    outputs(4255) <= not((layer0_outputs(2136)) and (layer0_outputs(932)));
    outputs(4256) <= layer0_outputs(1122);
    outputs(4257) <= layer0_outputs(1940);
    outputs(4258) <= not((layer0_outputs(3314)) xor (layer0_outputs(4700)));
    outputs(4259) <= layer0_outputs(5093);
    outputs(4260) <= layer0_outputs(3272);
    outputs(4261) <= layer0_outputs(4084);
    outputs(4262) <= (layer0_outputs(1504)) and not (layer0_outputs(4957));
    outputs(4263) <= layer0_outputs(183);
    outputs(4264) <= (layer0_outputs(3909)) xor (layer0_outputs(389));
    outputs(4265) <= not((layer0_outputs(122)) xor (layer0_outputs(2848)));
    outputs(4266) <= layer0_outputs(4934);
    outputs(4267) <= not(layer0_outputs(245)) or (layer0_outputs(5096));
    outputs(4268) <= not(layer0_outputs(2294));
    outputs(4269) <= layer0_outputs(3172);
    outputs(4270) <= (layer0_outputs(3278)) xor (layer0_outputs(4480));
    outputs(4271) <= not(layer0_outputs(577));
    outputs(4272) <= (layer0_outputs(345)) xor (layer0_outputs(3689));
    outputs(4273) <= not(layer0_outputs(3622)) or (layer0_outputs(1370));
    outputs(4274) <= (layer0_outputs(3966)) and not (layer0_outputs(4086));
    outputs(4275) <= layer0_outputs(4215);
    outputs(4276) <= (layer0_outputs(4067)) xor (layer0_outputs(3146));
    outputs(4277) <= (layer0_outputs(331)) and (layer0_outputs(1972));
    outputs(4278) <= not(layer0_outputs(640));
    outputs(4279) <= layer0_outputs(828);
    outputs(4280) <= (layer0_outputs(34)) xor (layer0_outputs(1038));
    outputs(4281) <= not((layer0_outputs(3405)) and (layer0_outputs(2966)));
    outputs(4282) <= not(layer0_outputs(2870));
    outputs(4283) <= not(layer0_outputs(3347));
    outputs(4284) <= layer0_outputs(3646);
    outputs(4285) <= (layer0_outputs(4095)) xor (layer0_outputs(2244));
    outputs(4286) <= (layer0_outputs(4629)) or (layer0_outputs(4272));
    outputs(4287) <= layer0_outputs(59);
    outputs(4288) <= not(layer0_outputs(262)) or (layer0_outputs(3233));
    outputs(4289) <= not(layer0_outputs(3639));
    outputs(4290) <= not(layer0_outputs(4444));
    outputs(4291) <= not((layer0_outputs(1377)) xor (layer0_outputs(1747)));
    outputs(4292) <= layer0_outputs(789);
    outputs(4293) <= layer0_outputs(1433);
    outputs(4294) <= (layer0_outputs(953)) or (layer0_outputs(3187));
    outputs(4295) <= (layer0_outputs(4309)) xor (layer0_outputs(4316));
    outputs(4296) <= (layer0_outputs(2126)) xor (layer0_outputs(2016));
    outputs(4297) <= layer0_outputs(1284);
    outputs(4298) <= not(layer0_outputs(4717));
    outputs(4299) <= layer0_outputs(5083);
    outputs(4300) <= not(layer0_outputs(4486));
    outputs(4301) <= not((layer0_outputs(903)) xor (layer0_outputs(1727)));
    outputs(4302) <= (layer0_outputs(3508)) and not (layer0_outputs(3032));
    outputs(4303) <= (layer0_outputs(3872)) or (layer0_outputs(2194));
    outputs(4304) <= not((layer0_outputs(1269)) xor (layer0_outputs(622)));
    outputs(4305) <= not(layer0_outputs(22));
    outputs(4306) <= (layer0_outputs(1226)) xor (layer0_outputs(2034));
    outputs(4307) <= not(layer0_outputs(846));
    outputs(4308) <= (layer0_outputs(3909)) and not (layer0_outputs(2133));
    outputs(4309) <= (layer0_outputs(2274)) or (layer0_outputs(4866));
    outputs(4310) <= layer0_outputs(3411);
    outputs(4311) <= not((layer0_outputs(4875)) and (layer0_outputs(439)));
    outputs(4312) <= layer0_outputs(3802);
    outputs(4313) <= not(layer0_outputs(2821)) or (layer0_outputs(1556));
    outputs(4314) <= (layer0_outputs(4094)) and not (layer0_outputs(1785));
    outputs(4315) <= (layer0_outputs(4788)) and not (layer0_outputs(4716));
    outputs(4316) <= (layer0_outputs(967)) and not (layer0_outputs(423));
    outputs(4317) <= not(layer0_outputs(4677));
    outputs(4318) <= not((layer0_outputs(3918)) xor (layer0_outputs(4041)));
    outputs(4319) <= layer0_outputs(4107);
    outputs(4320) <= not((layer0_outputs(1563)) or (layer0_outputs(2544)));
    outputs(4321) <= not((layer0_outputs(1839)) xor (layer0_outputs(3786)));
    outputs(4322) <= layer0_outputs(1179);
    outputs(4323) <= (layer0_outputs(362)) and not (layer0_outputs(4360));
    outputs(4324) <= not((layer0_outputs(2068)) and (layer0_outputs(3838)));
    outputs(4325) <= not(layer0_outputs(3462)) or (layer0_outputs(1340));
    outputs(4326) <= layer0_outputs(2814);
    outputs(4327) <= (layer0_outputs(3775)) and (layer0_outputs(2291));
    outputs(4328) <= not(layer0_outputs(1498));
    outputs(4329) <= not(layer0_outputs(4489));
    outputs(4330) <= layer0_outputs(4465);
    outputs(4331) <= layer0_outputs(3567);
    outputs(4332) <= not(layer0_outputs(4504)) or (layer0_outputs(890));
    outputs(4333) <= '1';
    outputs(4334) <= not(layer0_outputs(303));
    outputs(4335) <= (layer0_outputs(2029)) xor (layer0_outputs(929));
    outputs(4336) <= not(layer0_outputs(1347));
    outputs(4337) <= (layer0_outputs(4924)) or (layer0_outputs(4128));
    outputs(4338) <= not(layer0_outputs(4888));
    outputs(4339) <= (layer0_outputs(3393)) or (layer0_outputs(4877));
    outputs(4340) <= layer0_outputs(131);
    outputs(4341) <= layer0_outputs(755);
    outputs(4342) <= not((layer0_outputs(4068)) xor (layer0_outputs(2690)));
    outputs(4343) <= not(layer0_outputs(4271));
    outputs(4344) <= (layer0_outputs(1644)) and not (layer0_outputs(3353));
    outputs(4345) <= not((layer0_outputs(2466)) xor (layer0_outputs(2805)));
    outputs(4346) <= not(layer0_outputs(2571));
    outputs(4347) <= (layer0_outputs(2848)) xor (layer0_outputs(1096));
    outputs(4348) <= not(layer0_outputs(4032)) or (layer0_outputs(2127));
    outputs(4349) <= layer0_outputs(1473);
    outputs(4350) <= not(layer0_outputs(2697)) or (layer0_outputs(2417));
    outputs(4351) <= not(layer0_outputs(1756)) or (layer0_outputs(2651));
    outputs(4352) <= (layer0_outputs(2499)) and not (layer0_outputs(726));
    outputs(4353) <= not(layer0_outputs(2729));
    outputs(4354) <= layer0_outputs(1095);
    outputs(4355) <= not((layer0_outputs(4053)) or (layer0_outputs(864)));
    outputs(4356) <= (layer0_outputs(1865)) xor (layer0_outputs(4311));
    outputs(4357) <= not(layer0_outputs(3758));
    outputs(4358) <= layer0_outputs(4484);
    outputs(4359) <= (layer0_outputs(4755)) xor (layer0_outputs(2637));
    outputs(4360) <= not((layer0_outputs(797)) and (layer0_outputs(1643)));
    outputs(4361) <= (layer0_outputs(5013)) xor (layer0_outputs(4270));
    outputs(4362) <= not(layer0_outputs(2208));
    outputs(4363) <= (layer0_outputs(3803)) and not (layer0_outputs(191));
    outputs(4364) <= layer0_outputs(1095);
    outputs(4365) <= not(layer0_outputs(4073));
    outputs(4366) <= layer0_outputs(1969);
    outputs(4367) <= (layer0_outputs(1984)) and (layer0_outputs(1868));
    outputs(4368) <= not(layer0_outputs(3132)) or (layer0_outputs(3318));
    outputs(4369) <= not((layer0_outputs(2921)) or (layer0_outputs(4728)));
    outputs(4370) <= (layer0_outputs(3930)) or (layer0_outputs(4430));
    outputs(4371) <= not(layer0_outputs(2845));
    outputs(4372) <= not(layer0_outputs(4970)) or (layer0_outputs(3016));
    outputs(4373) <= not((layer0_outputs(4623)) xor (layer0_outputs(3330)));
    outputs(4374) <= (layer0_outputs(3254)) or (layer0_outputs(1738));
    outputs(4375) <= layer0_outputs(1641);
    outputs(4376) <= layer0_outputs(54);
    outputs(4377) <= not((layer0_outputs(497)) or (layer0_outputs(996)));
    outputs(4378) <= (layer0_outputs(192)) and (layer0_outputs(4909));
    outputs(4379) <= not((layer0_outputs(4708)) and (layer0_outputs(3536)));
    outputs(4380) <= not((layer0_outputs(2871)) xor (layer0_outputs(3325)));
    outputs(4381) <= not((layer0_outputs(3922)) xor (layer0_outputs(1300)));
    outputs(4382) <= layer0_outputs(1044);
    outputs(4383) <= layer0_outputs(785);
    outputs(4384) <= not(layer0_outputs(1973));
    outputs(4385) <= layer0_outputs(4886);
    outputs(4386) <= not(layer0_outputs(2390));
    outputs(4387) <= layer0_outputs(3648);
    outputs(4388) <= not(layer0_outputs(2111)) or (layer0_outputs(3895));
    outputs(4389) <= not(layer0_outputs(384)) or (layer0_outputs(2823));
    outputs(4390) <= not(layer0_outputs(2357)) or (layer0_outputs(1506));
    outputs(4391) <= (layer0_outputs(1015)) and not (layer0_outputs(558));
    outputs(4392) <= not(layer0_outputs(3097));
    outputs(4393) <= (layer0_outputs(4501)) or (layer0_outputs(4653));
    outputs(4394) <= '1';
    outputs(4395) <= (layer0_outputs(2532)) and (layer0_outputs(3713));
    outputs(4396) <= layer0_outputs(2879);
    outputs(4397) <= not((layer0_outputs(946)) xor (layer0_outputs(854)));
    outputs(4398) <= not(layer0_outputs(172));
    outputs(4399) <= layer0_outputs(235);
    outputs(4400) <= not(layer0_outputs(2304));
    outputs(4401) <= layer0_outputs(1881);
    outputs(4402) <= (layer0_outputs(5086)) and (layer0_outputs(3730));
    outputs(4403) <= layer0_outputs(729);
    outputs(4404) <= (layer0_outputs(3787)) xor (layer0_outputs(326));
    outputs(4405) <= not(layer0_outputs(4320)) or (layer0_outputs(3306));
    outputs(4406) <= layer0_outputs(4335);
    outputs(4407) <= not(layer0_outputs(4053));
    outputs(4408) <= layer0_outputs(2793);
    outputs(4409) <= (layer0_outputs(2432)) and (layer0_outputs(3546));
    outputs(4410) <= not(layer0_outputs(1034));
    outputs(4411) <= (layer0_outputs(472)) and not (layer0_outputs(2461));
    outputs(4412) <= not((layer0_outputs(1686)) and (layer0_outputs(688)));
    outputs(4413) <= layer0_outputs(2424);
    outputs(4414) <= layer0_outputs(86);
    outputs(4415) <= (layer0_outputs(3331)) and not (layer0_outputs(4191));
    outputs(4416) <= not(layer0_outputs(2379)) or (layer0_outputs(1142));
    outputs(4417) <= (layer0_outputs(2623)) or (layer0_outputs(1952));
    outputs(4418) <= layer0_outputs(4187);
    outputs(4419) <= (layer0_outputs(3044)) xor (layer0_outputs(580));
    outputs(4420) <= not(layer0_outputs(3282)) or (layer0_outputs(1975));
    outputs(4421) <= (layer0_outputs(4189)) and not (layer0_outputs(3475));
    outputs(4422) <= layer0_outputs(105);
    outputs(4423) <= layer0_outputs(3117);
    outputs(4424) <= not(layer0_outputs(1302));
    outputs(4425) <= not((layer0_outputs(975)) xor (layer0_outputs(1943)));
    outputs(4426) <= layer0_outputs(1443);
    outputs(4427) <= (layer0_outputs(1601)) xor (layer0_outputs(3290));
    outputs(4428) <= not((layer0_outputs(3919)) xor (layer0_outputs(1475)));
    outputs(4429) <= not(layer0_outputs(2445));
    outputs(4430) <= (layer0_outputs(2236)) xor (layer0_outputs(929));
    outputs(4431) <= (layer0_outputs(4863)) or (layer0_outputs(4668));
    outputs(4432) <= (layer0_outputs(4976)) and (layer0_outputs(2170));
    outputs(4433) <= not(layer0_outputs(2930));
    outputs(4434) <= not((layer0_outputs(2240)) and (layer0_outputs(935)));
    outputs(4435) <= layer0_outputs(712);
    outputs(4436) <= not(layer0_outputs(3425));
    outputs(4437) <= (layer0_outputs(3346)) xor (layer0_outputs(1243));
    outputs(4438) <= not((layer0_outputs(2367)) xor (layer0_outputs(448)));
    outputs(4439) <= (layer0_outputs(490)) xor (layer0_outputs(4363));
    outputs(4440) <= layer0_outputs(4353);
    outputs(4441) <= not(layer0_outputs(4035));
    outputs(4442) <= not((layer0_outputs(3389)) and (layer0_outputs(1114)));
    outputs(4443) <= (layer0_outputs(4376)) and not (layer0_outputs(722));
    outputs(4444) <= not(layer0_outputs(4940));
    outputs(4445) <= layer0_outputs(4113);
    outputs(4446) <= not(layer0_outputs(396));
    outputs(4447) <= not(layer0_outputs(2319));
    outputs(4448) <= layer0_outputs(2992);
    outputs(4449) <= not(layer0_outputs(2565)) or (layer0_outputs(547));
    outputs(4450) <= not((layer0_outputs(2037)) xor (layer0_outputs(2490)));
    outputs(4451) <= (layer0_outputs(4285)) xor (layer0_outputs(3141));
    outputs(4452) <= (layer0_outputs(1612)) and not (layer0_outputs(1286));
    outputs(4453) <= not((layer0_outputs(1791)) xor (layer0_outputs(880)));
    outputs(4454) <= (layer0_outputs(1787)) and (layer0_outputs(3886));
    outputs(4455) <= not(layer0_outputs(2928));
    outputs(4456) <= not(layer0_outputs(3710));
    outputs(4457) <= (layer0_outputs(1825)) and not (layer0_outputs(4288));
    outputs(4458) <= layer0_outputs(4429);
    outputs(4459) <= layer0_outputs(3308);
    outputs(4460) <= (layer0_outputs(4824)) and (layer0_outputs(1787));
    outputs(4461) <= not(layer0_outputs(3472));
    outputs(4462) <= (layer0_outputs(1010)) and (layer0_outputs(1908));
    outputs(4463) <= layer0_outputs(3869);
    outputs(4464) <= layer0_outputs(2362);
    outputs(4465) <= layer0_outputs(828);
    outputs(4466) <= not(layer0_outputs(4996));
    outputs(4467) <= (layer0_outputs(1558)) xor (layer0_outputs(4657));
    outputs(4468) <= (layer0_outputs(1968)) and (layer0_outputs(1251));
    outputs(4469) <= layer0_outputs(587);
    outputs(4470) <= not(layer0_outputs(309)) or (layer0_outputs(3772));
    outputs(4471) <= not((layer0_outputs(3918)) xor (layer0_outputs(2082)));
    outputs(4472) <= not(layer0_outputs(1687)) or (layer0_outputs(3157));
    outputs(4473) <= not(layer0_outputs(1176));
    outputs(4474) <= (layer0_outputs(535)) xor (layer0_outputs(2517));
    outputs(4475) <= not((layer0_outputs(3683)) or (layer0_outputs(3257)));
    outputs(4476) <= not(layer0_outputs(3695));
    outputs(4477) <= layer0_outputs(609);
    outputs(4478) <= not(layer0_outputs(139));
    outputs(4479) <= layer0_outputs(3764);
    outputs(4480) <= layer0_outputs(4805);
    outputs(4481) <= not((layer0_outputs(202)) or (layer0_outputs(1276)));
    outputs(4482) <= layer0_outputs(578);
    outputs(4483) <= not(layer0_outputs(5044)) or (layer0_outputs(3478));
    outputs(4484) <= not(layer0_outputs(5008));
    outputs(4485) <= not(layer0_outputs(4213));
    outputs(4486) <= (layer0_outputs(4683)) and not (layer0_outputs(3006));
    outputs(4487) <= (layer0_outputs(2006)) or (layer0_outputs(3115));
    outputs(4488) <= not((layer0_outputs(1571)) xor (layer0_outputs(1387)));
    outputs(4489) <= layer0_outputs(3803);
    outputs(4490) <= (layer0_outputs(985)) xor (layer0_outputs(1721));
    outputs(4491) <= (layer0_outputs(2847)) and (layer0_outputs(601));
    outputs(4492) <= layer0_outputs(1970);
    outputs(4493) <= (layer0_outputs(1205)) xor (layer0_outputs(856));
    outputs(4494) <= not(layer0_outputs(2158));
    outputs(4495) <= (layer0_outputs(4011)) xor (layer0_outputs(1318));
    outputs(4496) <= not(layer0_outputs(3763)) or (layer0_outputs(408));
    outputs(4497) <= layer0_outputs(1392);
    outputs(4498) <= not((layer0_outputs(850)) xor (layer0_outputs(1976)));
    outputs(4499) <= not(layer0_outputs(2873));
    outputs(4500) <= not(layer0_outputs(2192)) or (layer0_outputs(99));
    outputs(4501) <= not(layer0_outputs(3370));
    outputs(4502) <= (layer0_outputs(1297)) and not (layer0_outputs(4656));
    outputs(4503) <= (layer0_outputs(4545)) or (layer0_outputs(2493));
    outputs(4504) <= (layer0_outputs(4705)) or (layer0_outputs(1834));
    outputs(4505) <= (layer0_outputs(4732)) xor (layer0_outputs(2280));
    outputs(4506) <= (layer0_outputs(2756)) or (layer0_outputs(3320));
    outputs(4507) <= (layer0_outputs(1746)) and (layer0_outputs(3380));
    outputs(4508) <= layer0_outputs(1639);
    outputs(4509) <= (layer0_outputs(3308)) and not (layer0_outputs(2902));
    outputs(4510) <= (layer0_outputs(4095)) or (layer0_outputs(1489));
    outputs(4511) <= not(layer0_outputs(2164));
    outputs(4512) <= not(layer0_outputs(1190));
    outputs(4513) <= (layer0_outputs(1681)) and (layer0_outputs(1431));
    outputs(4514) <= (layer0_outputs(5083)) and not (layer0_outputs(3349));
    outputs(4515) <= not(layer0_outputs(3376));
    outputs(4516) <= '1';
    outputs(4517) <= layer0_outputs(370);
    outputs(4518) <= not((layer0_outputs(4437)) xor (layer0_outputs(4744)));
    outputs(4519) <= layer0_outputs(3260);
    outputs(4520) <= not((layer0_outputs(4904)) xor (layer0_outputs(484)));
    outputs(4521) <= not(layer0_outputs(1903));
    outputs(4522) <= not(layer0_outputs(4136));
    outputs(4523) <= (layer0_outputs(2182)) or (layer0_outputs(3486));
    outputs(4524) <= not((layer0_outputs(4596)) or (layer0_outputs(1446)));
    outputs(4525) <= not(layer0_outputs(470));
    outputs(4526) <= not(layer0_outputs(2643));
    outputs(4527) <= not((layer0_outputs(2467)) and (layer0_outputs(555)));
    outputs(4528) <= (layer0_outputs(3509)) xor (layer0_outputs(3913));
    outputs(4529) <= layer0_outputs(2353);
    outputs(4530) <= not(layer0_outputs(2643));
    outputs(4531) <= layer0_outputs(3144);
    outputs(4532) <= (layer0_outputs(2195)) and (layer0_outputs(1239));
    outputs(4533) <= layer0_outputs(3737);
    outputs(4534) <= not((layer0_outputs(718)) xor (layer0_outputs(816)));
    outputs(4535) <= not(layer0_outputs(4573));
    outputs(4536) <= not((layer0_outputs(3546)) xor (layer0_outputs(3933)));
    outputs(4537) <= (layer0_outputs(4669)) xor (layer0_outputs(1656));
    outputs(4538) <= layer0_outputs(3391);
    outputs(4539) <= not(layer0_outputs(2563));
    outputs(4540) <= (layer0_outputs(3252)) and (layer0_outputs(4554));
    outputs(4541) <= not((layer0_outputs(1492)) xor (layer0_outputs(697)));
    outputs(4542) <= not((layer0_outputs(1669)) xor (layer0_outputs(4545)));
    outputs(4543) <= not(layer0_outputs(559));
    outputs(4544) <= not(layer0_outputs(4945)) or (layer0_outputs(4808));
    outputs(4545) <= not(layer0_outputs(1757));
    outputs(4546) <= (layer0_outputs(2736)) and not (layer0_outputs(4597));
    outputs(4547) <= not((layer0_outputs(1562)) or (layer0_outputs(722)));
    outputs(4548) <= layer0_outputs(3605);
    outputs(4549) <= (layer0_outputs(971)) and not (layer0_outputs(3862));
    outputs(4550) <= not((layer0_outputs(1080)) xor (layer0_outputs(1045)));
    outputs(4551) <= not((layer0_outputs(2914)) xor (layer0_outputs(2949)));
    outputs(4552) <= not((layer0_outputs(3520)) xor (layer0_outputs(643)));
    outputs(4553) <= layer0_outputs(2317);
    outputs(4554) <= (layer0_outputs(4085)) and (layer0_outputs(2394));
    outputs(4555) <= layer0_outputs(1077);
    outputs(4556) <= not((layer0_outputs(4504)) and (layer0_outputs(2337)));
    outputs(4557) <= not((layer0_outputs(2042)) xor (layer0_outputs(2803)));
    outputs(4558) <= not((layer0_outputs(3474)) xor (layer0_outputs(4093)));
    outputs(4559) <= layer0_outputs(1212);
    outputs(4560) <= not(layer0_outputs(4892)) or (layer0_outputs(4948));
    outputs(4561) <= not(layer0_outputs(193));
    outputs(4562) <= not(layer0_outputs(2564));
    outputs(4563) <= (layer0_outputs(1456)) xor (layer0_outputs(1317));
    outputs(4564) <= (layer0_outputs(517)) xor (layer0_outputs(3525));
    outputs(4565) <= layer0_outputs(5034);
    outputs(4566) <= layer0_outputs(2597);
    outputs(4567) <= (layer0_outputs(525)) and not (layer0_outputs(5021));
    outputs(4568) <= not(layer0_outputs(1487)) or (layer0_outputs(739));
    outputs(4569) <= not(layer0_outputs(3212));
    outputs(4570) <= not(layer0_outputs(3584));
    outputs(4571) <= (layer0_outputs(2033)) and not (layer0_outputs(320));
    outputs(4572) <= layer0_outputs(2974);
    outputs(4573) <= not(layer0_outputs(4435));
    outputs(4574) <= not(layer0_outputs(104)) or (layer0_outputs(2545));
    outputs(4575) <= not((layer0_outputs(2705)) xor (layer0_outputs(5102)));
    outputs(4576) <= not((layer0_outputs(272)) xor (layer0_outputs(2859)));
    outputs(4577) <= (layer0_outputs(211)) xor (layer0_outputs(1415));
    outputs(4578) <= layer0_outputs(1694);
    outputs(4579) <= (layer0_outputs(4843)) and not (layer0_outputs(4087));
    outputs(4580) <= (layer0_outputs(1383)) or (layer0_outputs(321));
    outputs(4581) <= not((layer0_outputs(3318)) and (layer0_outputs(118)));
    outputs(4582) <= layer0_outputs(3942);
    outputs(4583) <= not(layer0_outputs(1830));
    outputs(4584) <= (layer0_outputs(2416)) or (layer0_outputs(3881));
    outputs(4585) <= (layer0_outputs(4009)) xor (layer0_outputs(792));
    outputs(4586) <= not(layer0_outputs(314));
    outputs(4587) <= layer0_outputs(4319);
    outputs(4588) <= not(layer0_outputs(3615));
    outputs(4589) <= (layer0_outputs(2252)) xor (layer0_outputs(3522));
    outputs(4590) <= layer0_outputs(3708);
    outputs(4591) <= layer0_outputs(1223);
    outputs(4592) <= layer0_outputs(2502);
    outputs(4593) <= not(layer0_outputs(4765));
    outputs(4594) <= not(layer0_outputs(1072));
    outputs(4595) <= not(layer0_outputs(606));
    outputs(4596) <= not(layer0_outputs(373));
    outputs(4597) <= not(layer0_outputs(4367));
    outputs(4598) <= not(layer0_outputs(3397)) or (layer0_outputs(2375));
    outputs(4599) <= not(layer0_outputs(2971));
    outputs(4600) <= (layer0_outputs(5077)) or (layer0_outputs(3302));
    outputs(4601) <= (layer0_outputs(1163)) and (layer0_outputs(2809));
    outputs(4602) <= not(layer0_outputs(433));
    outputs(4603) <= not(layer0_outputs(4047));
    outputs(4604) <= not(layer0_outputs(4183));
    outputs(4605) <= not((layer0_outputs(1057)) and (layer0_outputs(3025)));
    outputs(4606) <= not(layer0_outputs(647));
    outputs(4607) <= layer0_outputs(2612);
    outputs(4608) <= not((layer0_outputs(4143)) xor (layer0_outputs(969)));
    outputs(4609) <= (layer0_outputs(3524)) xor (layer0_outputs(1906));
    outputs(4610) <= (layer0_outputs(1506)) xor (layer0_outputs(2062));
    outputs(4611) <= (layer0_outputs(3975)) and (layer0_outputs(4516));
    outputs(4612) <= not(layer0_outputs(1675)) or (layer0_outputs(1944));
    outputs(4613) <= (layer0_outputs(3001)) and (layer0_outputs(1325));
    outputs(4614) <= (layer0_outputs(4417)) xor (layer0_outputs(4859));
    outputs(4615) <= not((layer0_outputs(446)) xor (layer0_outputs(3543)));
    outputs(4616) <= not(layer0_outputs(2615));
    outputs(4617) <= layer0_outputs(4195);
    outputs(4618) <= not((layer0_outputs(1616)) xor (layer0_outputs(4439)));
    outputs(4619) <= (layer0_outputs(288)) and not (layer0_outputs(3447));
    outputs(4620) <= not((layer0_outputs(5056)) xor (layer0_outputs(4562)));
    outputs(4621) <= not((layer0_outputs(749)) and (layer0_outputs(4340)));
    outputs(4622) <= (layer0_outputs(539)) and not (layer0_outputs(871));
    outputs(4623) <= (layer0_outputs(3582)) xor (layer0_outputs(2837));
    outputs(4624) <= (layer0_outputs(922)) and not (layer0_outputs(1292));
    outputs(4625) <= not(layer0_outputs(257)) or (layer0_outputs(2301));
    outputs(4626) <= layer0_outputs(1849);
    outputs(4627) <= not(layer0_outputs(3479));
    outputs(4628) <= (layer0_outputs(3092)) and not (layer0_outputs(1043));
    outputs(4629) <= '0';
    outputs(4630) <= not((layer0_outputs(1835)) xor (layer0_outputs(339)));
    outputs(4631) <= layer0_outputs(2117);
    outputs(4632) <= not((layer0_outputs(308)) or (layer0_outputs(334)));
    outputs(4633) <= not((layer0_outputs(2449)) xor (layer0_outputs(605)));
    outputs(4634) <= (layer0_outputs(1878)) and not (layer0_outputs(1036));
    outputs(4635) <= (layer0_outputs(4411)) and not (layer0_outputs(343));
    outputs(4636) <= (layer0_outputs(5047)) xor (layer0_outputs(222));
    outputs(4637) <= not(layer0_outputs(2465));
    outputs(4638) <= (layer0_outputs(4160)) and not (layer0_outputs(2350));
    outputs(4639) <= layer0_outputs(2501);
    outputs(4640) <= not((layer0_outputs(3374)) xor (layer0_outputs(1220)));
    outputs(4641) <= not(layer0_outputs(765));
    outputs(4642) <= (layer0_outputs(4016)) and not (layer0_outputs(1487));
    outputs(4643) <= not(layer0_outputs(4975));
    outputs(4644) <= layer0_outputs(413);
    outputs(4645) <= layer0_outputs(1722);
    outputs(4646) <= layer0_outputs(4079);
    outputs(4647) <= not((layer0_outputs(1280)) or (layer0_outputs(4144)));
    outputs(4648) <= not(layer0_outputs(848));
    outputs(4649) <= (layer0_outputs(2954)) and not (layer0_outputs(2002));
    outputs(4650) <= not(layer0_outputs(78));
    outputs(4651) <= not(layer0_outputs(604));
    outputs(4652) <= not((layer0_outputs(1046)) or (layer0_outputs(426)));
    outputs(4653) <= (layer0_outputs(740)) or (layer0_outputs(1299));
    outputs(4654) <= (layer0_outputs(2177)) xor (layer0_outputs(110));
    outputs(4655) <= (layer0_outputs(1559)) and not (layer0_outputs(4992));
    outputs(4656) <= layer0_outputs(3193);
    outputs(4657) <= (layer0_outputs(4495)) and (layer0_outputs(3768));
    outputs(4658) <= not((layer0_outputs(197)) or (layer0_outputs(910)));
    outputs(4659) <= layer0_outputs(4837);
    outputs(4660) <= not(layer0_outputs(2868));
    outputs(4661) <= (layer0_outputs(231)) and not (layer0_outputs(2645));
    outputs(4662) <= (layer0_outputs(192)) xor (layer0_outputs(2791));
    outputs(4663) <= (layer0_outputs(3963)) and not (layer0_outputs(3944));
    outputs(4664) <= not((layer0_outputs(2383)) xor (layer0_outputs(3422)));
    outputs(4665) <= (layer0_outputs(3646)) and (layer0_outputs(4620));
    outputs(4666) <= (layer0_outputs(3241)) xor (layer0_outputs(3421));
    outputs(4667) <= (layer0_outputs(641)) or (layer0_outputs(2965));
    outputs(4668) <= (layer0_outputs(1374)) and not (layer0_outputs(595));
    outputs(4669) <= layer0_outputs(581);
    outputs(4670) <= not((layer0_outputs(124)) or (layer0_outputs(3426)));
    outputs(4671) <= not(layer0_outputs(3463)) or (layer0_outputs(803));
    outputs(4672) <= not(layer0_outputs(4058));
    outputs(4673) <= not(layer0_outputs(2125));
    outputs(4674) <= not(layer0_outputs(1495)) or (layer0_outputs(2262));
    outputs(4675) <= (layer0_outputs(4712)) or (layer0_outputs(4704));
    outputs(4676) <= (layer0_outputs(4401)) and not (layer0_outputs(4011));
    outputs(4677) <= (layer0_outputs(5078)) xor (layer0_outputs(4938));
    outputs(4678) <= layer0_outputs(352);
    outputs(4679) <= not(layer0_outputs(4013));
    outputs(4680) <= (layer0_outputs(2989)) and not (layer0_outputs(3565));
    outputs(4681) <= not((layer0_outputs(3018)) xor (layer0_outputs(1130)));
    outputs(4682) <= (layer0_outputs(379)) and not (layer0_outputs(3865));
    outputs(4683) <= not(layer0_outputs(1281));
    outputs(4684) <= not(layer0_outputs(2850)) or (layer0_outputs(2642));
    outputs(4685) <= (layer0_outputs(342)) xor (layer0_outputs(143));
    outputs(4686) <= (layer0_outputs(330)) and not (layer0_outputs(3227));
    outputs(4687) <= layer0_outputs(3683);
    outputs(4688) <= '1';
    outputs(4689) <= (layer0_outputs(2393)) and (layer0_outputs(4164));
    outputs(4690) <= not(layer0_outputs(2082));
    outputs(4691) <= (layer0_outputs(3362)) xor (layer0_outputs(3099));
    outputs(4692) <= (layer0_outputs(3657)) xor (layer0_outputs(2387));
    outputs(4693) <= (layer0_outputs(4171)) and (layer0_outputs(3714));
    outputs(4694) <= not(layer0_outputs(3954));
    outputs(4695) <= (layer0_outputs(2241)) and not (layer0_outputs(3142));
    outputs(4696) <= not((layer0_outputs(1493)) or (layer0_outputs(1820)));
    outputs(4697) <= (layer0_outputs(2724)) and not (layer0_outputs(1252));
    outputs(4698) <= not(layer0_outputs(3677));
    outputs(4699) <= not(layer0_outputs(4369));
    outputs(4700) <= (layer0_outputs(1754)) xor (layer0_outputs(1568));
    outputs(4701) <= layer0_outputs(3396);
    outputs(4702) <= not(layer0_outputs(4530));
    outputs(4703) <= not(layer0_outputs(4078));
    outputs(4704) <= layer0_outputs(1867);
    outputs(4705) <= (layer0_outputs(623)) xor (layer0_outputs(3710));
    outputs(4706) <= (layer0_outputs(845)) and not (layer0_outputs(5111));
    outputs(4707) <= not((layer0_outputs(1084)) or (layer0_outputs(4706)));
    outputs(4708) <= not((layer0_outputs(1503)) or (layer0_outputs(1080)));
    outputs(4709) <= not(layer0_outputs(1042));
    outputs(4710) <= layer0_outputs(1363);
    outputs(4711) <= (layer0_outputs(2774)) and not (layer0_outputs(1140));
    outputs(4712) <= (layer0_outputs(4689)) and not (layer0_outputs(3589));
    outputs(4713) <= layer0_outputs(3433);
    outputs(4714) <= layer0_outputs(2052);
    outputs(4715) <= not(layer0_outputs(371));
    outputs(4716) <= layer0_outputs(169);
    outputs(4717) <= layer0_outputs(3593);
    outputs(4718) <= (layer0_outputs(928)) and (layer0_outputs(3694));
    outputs(4719) <= layer0_outputs(4413);
    outputs(4720) <= layer0_outputs(2012);
    outputs(4721) <= layer0_outputs(121);
    outputs(4722) <= (layer0_outputs(1739)) and not (layer0_outputs(2692));
    outputs(4723) <= not((layer0_outputs(2481)) xor (layer0_outputs(3223)));
    outputs(4724) <= (layer0_outputs(5106)) and (layer0_outputs(5043));
    outputs(4725) <= layer0_outputs(2907);
    outputs(4726) <= (layer0_outputs(3870)) and not (layer0_outputs(2500));
    outputs(4727) <= (layer0_outputs(3570)) and not (layer0_outputs(4502));
    outputs(4728) <= (layer0_outputs(1045)) xor (layer0_outputs(2759));
    outputs(4729) <= layer0_outputs(468);
    outputs(4730) <= not(layer0_outputs(998));
    outputs(4731) <= (layer0_outputs(82)) and not (layer0_outputs(4663));
    outputs(4732) <= (layer0_outputs(3735)) xor (layer0_outputs(3230));
    outputs(4733) <= (layer0_outputs(4819)) xor (layer0_outputs(4114));
    outputs(4734) <= (layer0_outputs(3827)) xor (layer0_outputs(4910));
    outputs(4735) <= (layer0_outputs(1382)) and not (layer0_outputs(3717));
    outputs(4736) <= layer0_outputs(4247);
    outputs(4737) <= not(layer0_outputs(2078));
    outputs(4738) <= (layer0_outputs(4979)) and not (layer0_outputs(4833));
    outputs(4739) <= (layer0_outputs(916)) and not (layer0_outputs(1576));
    outputs(4740) <= not((layer0_outputs(2410)) or (layer0_outputs(1050)));
    outputs(4741) <= not(layer0_outputs(3937)) or (layer0_outputs(2961));
    outputs(4742) <= (layer0_outputs(1918)) and not (layer0_outputs(3210));
    outputs(4743) <= layer0_outputs(3028);
    outputs(4744) <= layer0_outputs(52);
    outputs(4745) <= not(layer0_outputs(4008));
    outputs(4746) <= (layer0_outputs(1989)) xor (layer0_outputs(260));
    outputs(4747) <= layer0_outputs(1152);
    outputs(4748) <= (layer0_outputs(5101)) and not (layer0_outputs(1223));
    outputs(4749) <= not(layer0_outputs(4059));
    outputs(4750) <= not((layer0_outputs(1087)) or (layer0_outputs(4348)));
    outputs(4751) <= (layer0_outputs(3650)) xor (layer0_outputs(3338));
    outputs(4752) <= (layer0_outputs(1827)) xor (layer0_outputs(4046));
    outputs(4753) <= (layer0_outputs(536)) and (layer0_outputs(223));
    outputs(4754) <= (layer0_outputs(4172)) and not (layer0_outputs(3903));
    outputs(4755) <= (layer0_outputs(4812)) xor (layer0_outputs(633));
    outputs(4756) <= not((layer0_outputs(4510)) or (layer0_outputs(3326)));
    outputs(4757) <= not(layer0_outputs(4786));
    outputs(4758) <= not(layer0_outputs(1850));
    outputs(4759) <= layer0_outputs(1234);
    outputs(4760) <= not((layer0_outputs(1383)) xor (layer0_outputs(1238)));
    outputs(4761) <= not((layer0_outputs(1954)) and (layer0_outputs(4163)));
    outputs(4762) <= (layer0_outputs(2570)) xor (layer0_outputs(3814));
    outputs(4763) <= layer0_outputs(3037);
    outputs(4764) <= layer0_outputs(2016);
    outputs(4765) <= not((layer0_outputs(3833)) xor (layer0_outputs(3675)));
    outputs(4766) <= layer0_outputs(314);
    outputs(4767) <= (layer0_outputs(3244)) xor (layer0_outputs(1877));
    outputs(4768) <= not((layer0_outputs(2962)) xor (layer0_outputs(1773)));
    outputs(4769) <= (layer0_outputs(1862)) or (layer0_outputs(1848));
    outputs(4770) <= not((layer0_outputs(2160)) or (layer0_outputs(199)));
    outputs(4771) <= not(layer0_outputs(2066));
    outputs(4772) <= (layer0_outputs(1117)) and not (layer0_outputs(1466));
    outputs(4773) <= (layer0_outputs(1853)) xor (layer0_outputs(1074));
    outputs(4774) <= layer0_outputs(4002);
    outputs(4775) <= not((layer0_outputs(4711)) xor (layer0_outputs(3759)));
    outputs(4776) <= layer0_outputs(5045);
    outputs(4777) <= (layer0_outputs(1722)) and not (layer0_outputs(4486));
    outputs(4778) <= layer0_outputs(1563);
    outputs(4779) <= (layer0_outputs(1187)) and not (layer0_outputs(170));
    outputs(4780) <= not(layer0_outputs(4916));
    outputs(4781) <= not((layer0_outputs(4175)) or (layer0_outputs(2064)));
    outputs(4782) <= layer0_outputs(851);
    outputs(4783) <= layer0_outputs(3274);
    outputs(4784) <= not((layer0_outputs(1949)) xor (layer0_outputs(1137)));
    outputs(4785) <= layer0_outputs(3105);
    outputs(4786) <= not(layer0_outputs(921)) or (layer0_outputs(1635));
    outputs(4787) <= layer0_outputs(962);
    outputs(4788) <= layer0_outputs(3777);
    outputs(4789) <= not(layer0_outputs(2348));
    outputs(4790) <= not(layer0_outputs(1952));
    outputs(4791) <= not((layer0_outputs(3229)) xor (layer0_outputs(3367)));
    outputs(4792) <= not(layer0_outputs(3163));
    outputs(4793) <= not(layer0_outputs(3516));
    outputs(4794) <= not(layer0_outputs(2099)) or (layer0_outputs(237));
    outputs(4795) <= not(layer0_outputs(1046));
    outputs(4796) <= not(layer0_outputs(246));
    outputs(4797) <= layer0_outputs(1946);
    outputs(4798) <= layer0_outputs(1368);
    outputs(4799) <= not(layer0_outputs(4328));
    outputs(4800) <= not(layer0_outputs(3902));
    outputs(4801) <= (layer0_outputs(1739)) and not (layer0_outputs(6));
    outputs(4802) <= layer0_outputs(3950);
    outputs(4803) <= not((layer0_outputs(3712)) and (layer0_outputs(3551)));
    outputs(4804) <= not((layer0_outputs(4399)) xor (layer0_outputs(4711)));
    outputs(4805) <= (layer0_outputs(731)) or (layer0_outputs(3015));
    outputs(4806) <= layer0_outputs(4307);
    outputs(4807) <= (layer0_outputs(1371)) and (layer0_outputs(2135));
    outputs(4808) <= layer0_outputs(4298);
    outputs(4809) <= (layer0_outputs(2829)) and (layer0_outputs(1717));
    outputs(4810) <= layer0_outputs(4913);
    outputs(4811) <= (layer0_outputs(4356)) and not (layer0_outputs(822));
    outputs(4812) <= not((layer0_outputs(2555)) or (layer0_outputs(1147)));
    outputs(4813) <= (layer0_outputs(2010)) or (layer0_outputs(3004));
    outputs(4814) <= not((layer0_outputs(527)) or (layer0_outputs(2833)));
    outputs(4815) <= (layer0_outputs(4727)) and not (layer0_outputs(770));
    outputs(4816) <= layer0_outputs(1548);
    outputs(4817) <= not(layer0_outputs(3375)) or (layer0_outputs(2858));
    outputs(4818) <= not((layer0_outputs(1444)) or (layer0_outputs(2795)));
    outputs(4819) <= layer0_outputs(115);
    outputs(4820) <= layer0_outputs(2665);
    outputs(4821) <= not(layer0_outputs(3774));
    outputs(4822) <= layer0_outputs(1358);
    outputs(4823) <= (layer0_outputs(3678)) xor (layer0_outputs(3821));
    outputs(4824) <= (layer0_outputs(2787)) and (layer0_outputs(2589));
    outputs(4825) <= not(layer0_outputs(3548));
    outputs(4826) <= layer0_outputs(2205);
    outputs(4827) <= (layer0_outputs(721)) and (layer0_outputs(1980));
    outputs(4828) <= layer0_outputs(4367);
    outputs(4829) <= (layer0_outputs(2701)) and (layer0_outputs(684));
    outputs(4830) <= layer0_outputs(3124);
    outputs(4831) <= (layer0_outputs(768)) and not (layer0_outputs(978));
    outputs(4832) <= layer0_outputs(3255);
    outputs(4833) <= layer0_outputs(154);
    outputs(4834) <= not(layer0_outputs(3614));
    outputs(4835) <= (layer0_outputs(1149)) xor (layer0_outputs(2876));
    outputs(4836) <= (layer0_outputs(1882)) and not (layer0_outputs(799));
    outputs(4837) <= (layer0_outputs(3024)) and not (layer0_outputs(4419));
    outputs(4838) <= layer0_outputs(4607);
    outputs(4839) <= (layer0_outputs(1225)) and (layer0_outputs(166));
    outputs(4840) <= layer0_outputs(695);
    outputs(4841) <= (layer0_outputs(1991)) and not (layer0_outputs(3479));
    outputs(4842) <= not(layer0_outputs(2849));
    outputs(4843) <= not((layer0_outputs(2965)) or (layer0_outputs(2843)));
    outputs(4844) <= not((layer0_outputs(568)) or (layer0_outputs(562)));
    outputs(4845) <= not(layer0_outputs(4922));
    outputs(4846) <= (layer0_outputs(5019)) xor (layer0_outputs(1763));
    outputs(4847) <= layer0_outputs(3582);
    outputs(4848) <= (layer0_outputs(1943)) and not (layer0_outputs(996));
    outputs(4849) <= (layer0_outputs(1556)) xor (layer0_outputs(3586));
    outputs(4850) <= layer0_outputs(2653);
    outputs(4851) <= not(layer0_outputs(4572));
    outputs(4852) <= (layer0_outputs(3453)) and not (layer0_outputs(538));
    outputs(4853) <= not((layer0_outputs(426)) xor (layer0_outputs(2947)));
    outputs(4854) <= (layer0_outputs(57)) xor (layer0_outputs(2103));
    outputs(4855) <= not(layer0_outputs(8));
    outputs(4856) <= (layer0_outputs(4045)) and not (layer0_outputs(1592));
    outputs(4857) <= (layer0_outputs(4852)) and (layer0_outputs(5075));
    outputs(4858) <= not(layer0_outputs(146));
    outputs(4859) <= not(layer0_outputs(3497));
    outputs(4860) <= (layer0_outputs(909)) and (layer0_outputs(1913));
    outputs(4861) <= not(layer0_outputs(813));
    outputs(4862) <= (layer0_outputs(2454)) and (layer0_outputs(2852));
    outputs(4863) <= (layer0_outputs(1083)) and not (layer0_outputs(2422));
    outputs(4864) <= (layer0_outputs(4074)) and (layer0_outputs(3470));
    outputs(4865) <= not(layer0_outputs(4551));
    outputs(4866) <= not((layer0_outputs(4973)) xor (layer0_outputs(1540)));
    outputs(4867) <= layer0_outputs(3751);
    outputs(4868) <= layer0_outputs(4409);
    outputs(4869) <= not((layer0_outputs(1618)) or (layer0_outputs(3747)));
    outputs(4870) <= not((layer0_outputs(4691)) xor (layer0_outputs(3542)));
    outputs(4871) <= (layer0_outputs(2253)) and not (layer0_outputs(3556));
    outputs(4872) <= (layer0_outputs(1553)) and not (layer0_outputs(408));
    outputs(4873) <= (layer0_outputs(2631)) and (layer0_outputs(2746));
    outputs(4874) <= (layer0_outputs(1723)) xor (layer0_outputs(1270));
    outputs(4875) <= not((layer0_outputs(952)) or (layer0_outputs(1874)));
    outputs(4876) <= (layer0_outputs(771)) and not (layer0_outputs(1200));
    outputs(4877) <= (layer0_outputs(2704)) xor (layer0_outputs(3151));
    outputs(4878) <= not((layer0_outputs(3996)) or (layer0_outputs(490)));
    outputs(4879) <= (layer0_outputs(1620)) xor (layer0_outputs(4664));
    outputs(4880) <= not(layer0_outputs(657));
    outputs(4881) <= (layer0_outputs(318)) and not (layer0_outputs(1194));
    outputs(4882) <= layer0_outputs(2251);
    outputs(4883) <= (layer0_outputs(620)) xor (layer0_outputs(1250));
    outputs(4884) <= layer0_outputs(1656);
    outputs(4885) <= (layer0_outputs(3204)) or (layer0_outputs(5080));
    outputs(4886) <= (layer0_outputs(1543)) and (layer0_outputs(2159));
    outputs(4887) <= (layer0_outputs(2511)) and (layer0_outputs(845));
    outputs(4888) <= (layer0_outputs(5013)) or (layer0_outputs(3836));
    outputs(4889) <= not((layer0_outputs(1112)) or (layer0_outputs(28)));
    outputs(4890) <= not(layer0_outputs(1699));
    outputs(4891) <= layer0_outputs(3033);
    outputs(4892) <= layer0_outputs(4943);
    outputs(4893) <= not((layer0_outputs(3991)) or (layer0_outputs(571)));
    outputs(4894) <= layer0_outputs(3037);
    outputs(4895) <= not((layer0_outputs(145)) xor (layer0_outputs(1312)));
    outputs(4896) <= not(layer0_outputs(1356)) or (layer0_outputs(3664));
    outputs(4897) <= (layer0_outputs(4273)) and not (layer0_outputs(2760));
    outputs(4898) <= (layer0_outputs(1278)) xor (layer0_outputs(2981));
    outputs(4899) <= not(layer0_outputs(1307)) or (layer0_outputs(4881));
    outputs(4900) <= (layer0_outputs(1570)) and (layer0_outputs(1871));
    outputs(4901) <= (layer0_outputs(1088)) and (layer0_outputs(1306));
    outputs(4902) <= not(layer0_outputs(4929));
    outputs(4903) <= (layer0_outputs(3743)) xor (layer0_outputs(1856));
    outputs(4904) <= layer0_outputs(1884);
    outputs(4905) <= (layer0_outputs(4658)) and (layer0_outputs(3865));
    outputs(4906) <= layer0_outputs(1865);
    outputs(4907) <= (layer0_outputs(3416)) and not (layer0_outputs(927));
    outputs(4908) <= not(layer0_outputs(806));
    outputs(4909) <= not(layer0_outputs(269));
    outputs(4910) <= (layer0_outputs(1256)) xor (layer0_outputs(4920));
    outputs(4911) <= layer0_outputs(930);
    outputs(4912) <= layer0_outputs(1230);
    outputs(4913) <= not((layer0_outputs(4065)) or (layer0_outputs(1537)));
    outputs(4914) <= (layer0_outputs(2935)) xor (layer0_outputs(3736));
    outputs(4915) <= not(layer0_outputs(4856)) or (layer0_outputs(2583));
    outputs(4916) <= not(layer0_outputs(2300));
    outputs(4917) <= not(layer0_outputs(3987));
    outputs(4918) <= (layer0_outputs(2872)) and not (layer0_outputs(4538));
    outputs(4919) <= layer0_outputs(189);
    outputs(4920) <= (layer0_outputs(4162)) xor (layer0_outputs(4661));
    outputs(4921) <= not(layer0_outputs(3406));
    outputs(4922) <= not(layer0_outputs(2050));
    outputs(4923) <= layer0_outputs(2420);
    outputs(4924) <= layer0_outputs(4803);
    outputs(4925) <= not(layer0_outputs(719)) or (layer0_outputs(4690));
    outputs(4926) <= not(layer0_outputs(3567));
    outputs(4927) <= (layer0_outputs(1393)) and (layer0_outputs(23));
    outputs(4928) <= (layer0_outputs(916)) and (layer0_outputs(5062));
    outputs(4929) <= layer0_outputs(3050);
    outputs(4930) <= not((layer0_outputs(2942)) or (layer0_outputs(1039)));
    outputs(4931) <= not((layer0_outputs(3243)) and (layer0_outputs(1350)));
    outputs(4932) <= not(layer0_outputs(4517));
    outputs(4933) <= not((layer0_outputs(2990)) and (layer0_outputs(4974)));
    outputs(4934) <= not((layer0_outputs(2888)) or (layer0_outputs(3911)));
    outputs(4935) <= not((layer0_outputs(4389)) xor (layer0_outputs(2611)));
    outputs(4936) <= not(layer0_outputs(1158));
    outputs(4937) <= not(layer0_outputs(919));
    outputs(4938) <= (layer0_outputs(1732)) xor (layer0_outputs(190));
    outputs(4939) <= layer0_outputs(4560);
    outputs(4940) <= not((layer0_outputs(2250)) or (layer0_outputs(972)));
    outputs(4941) <= not(layer0_outputs(3328));
    outputs(4942) <= (layer0_outputs(5016)) and (layer0_outputs(2351));
    outputs(4943) <= (layer0_outputs(1950)) and not (layer0_outputs(3347));
    outputs(4944) <= not((layer0_outputs(1486)) or (layer0_outputs(3531)));
    outputs(4945) <= layer0_outputs(1883);
    outputs(4946) <= not((layer0_outputs(3900)) and (layer0_outputs(2278)));
    outputs(4947) <= not((layer0_outputs(4088)) and (layer0_outputs(2953)));
    outputs(4948) <= layer0_outputs(1987);
    outputs(4949) <= layer0_outputs(31);
    outputs(4950) <= (layer0_outputs(5082)) and (layer0_outputs(1673));
    outputs(4951) <= layer0_outputs(51);
    outputs(4952) <= not(layer0_outputs(4365));
    outputs(4953) <= (layer0_outputs(2811)) and not (layer0_outputs(3885));
    outputs(4954) <= not(layer0_outputs(819));
    outputs(4955) <= (layer0_outputs(1674)) xor (layer0_outputs(682));
    outputs(4956) <= not((layer0_outputs(3954)) or (layer0_outputs(1807)));
    outputs(4957) <= (layer0_outputs(3853)) xor (layer0_outputs(3986));
    outputs(4958) <= not(layer0_outputs(2310));
    outputs(4959) <= not(layer0_outputs(3062));
    outputs(4960) <= (layer0_outputs(847)) xor (layer0_outputs(132));
    outputs(4961) <= not((layer0_outputs(3969)) xor (layer0_outputs(740)));
    outputs(4962) <= layer0_outputs(4355);
    outputs(4963) <= layer0_outputs(1674);
    outputs(4964) <= not(layer0_outputs(2801));
    outputs(4965) <= layer0_outputs(3050);
    outputs(4966) <= (layer0_outputs(234)) and not (layer0_outputs(1734));
    outputs(4967) <= not((layer0_outputs(1696)) or (layer0_outputs(547)));
    outputs(4968) <= layer0_outputs(4722);
    outputs(4969) <= layer0_outputs(877);
    outputs(4970) <= (layer0_outputs(1263)) and not (layer0_outputs(2476));
    outputs(4971) <= (layer0_outputs(2077)) xor (layer0_outputs(4070));
    outputs(4972) <= layer0_outputs(4505);
    outputs(4973) <= layer0_outputs(4387);
    outputs(4974) <= not((layer0_outputs(3970)) xor (layer0_outputs(4008)));
    outputs(4975) <= layer0_outputs(1033);
    outputs(4976) <= not(layer0_outputs(3743));
    outputs(4977) <= (layer0_outputs(1887)) and not (layer0_outputs(4033));
    outputs(4978) <= (layer0_outputs(1699)) xor (layer0_outputs(2213));
    outputs(4979) <= not((layer0_outputs(2381)) and (layer0_outputs(3830)));
    outputs(4980) <= (layer0_outputs(2376)) and not (layer0_outputs(149));
    outputs(4981) <= (layer0_outputs(821)) and not (layer0_outputs(4153));
    outputs(4982) <= (layer0_outputs(4869)) and not (layer0_outputs(1446));
    outputs(4983) <= not(layer0_outputs(2329));
    outputs(4984) <= not((layer0_outputs(1104)) or (layer0_outputs(369)));
    outputs(4985) <= (layer0_outputs(210)) xor (layer0_outputs(4204));
    outputs(4986) <= (layer0_outputs(3873)) and not (layer0_outputs(2256));
    outputs(4987) <= not(layer0_outputs(124));
    outputs(4988) <= not(layer0_outputs(4304));
    outputs(4989) <= (layer0_outputs(1072)) xor (layer0_outputs(142));
    outputs(4990) <= not((layer0_outputs(2883)) xor (layer0_outputs(2980)));
    outputs(4991) <= (layer0_outputs(2)) and (layer0_outputs(4448));
    outputs(4992) <= not(layer0_outputs(2687));
    outputs(4993) <= not((layer0_outputs(681)) xor (layer0_outputs(1645)));
    outputs(4994) <= (layer0_outputs(302)) and not (layer0_outputs(3769));
    outputs(4995) <= (layer0_outputs(732)) and not (layer0_outputs(3907));
    outputs(4996) <= layer0_outputs(1686);
    outputs(4997) <= layer0_outputs(1463);
    outputs(4998) <= (layer0_outputs(4747)) and (layer0_outputs(1857));
    outputs(4999) <= not(layer0_outputs(96)) or (layer0_outputs(3386));
    outputs(5000) <= not(layer0_outputs(333));
    outputs(5001) <= (layer0_outputs(2671)) and (layer0_outputs(4546));
    outputs(5002) <= not((layer0_outputs(713)) xor (layer0_outputs(3928)));
    outputs(5003) <= not(layer0_outputs(1649));
    outputs(5004) <= (layer0_outputs(2582)) and not (layer0_outputs(2951));
    outputs(5005) <= (layer0_outputs(592)) and not (layer0_outputs(5027));
    outputs(5006) <= not(layer0_outputs(4352));
    outputs(5007) <= (layer0_outputs(425)) xor (layer0_outputs(936));
    outputs(5008) <= not(layer0_outputs(4365));
    outputs(5009) <= (layer0_outputs(1956)) and (layer0_outputs(2407));
    outputs(5010) <= (layer0_outputs(1213)) xor (layer0_outputs(4096));
    outputs(5011) <= layer0_outputs(3105);
    outputs(5012) <= not(layer0_outputs(2814));
    outputs(5013) <= (layer0_outputs(3771)) and not (layer0_outputs(2492));
    outputs(5014) <= (layer0_outputs(1626)) and not (layer0_outputs(564));
    outputs(5015) <= (layer0_outputs(1762)) xor (layer0_outputs(4863));
    outputs(5016) <= not(layer0_outputs(4900));
    outputs(5017) <= not(layer0_outputs(1917)) or (layer0_outputs(4245));
    outputs(5018) <= not(layer0_outputs(3210));
    outputs(5019) <= not((layer0_outputs(4112)) or (layer0_outputs(3856)));
    outputs(5020) <= not(layer0_outputs(1793)) or (layer0_outputs(2224));
    outputs(5021) <= (layer0_outputs(4431)) and not (layer0_outputs(3177));
    outputs(5022) <= (layer0_outputs(1019)) and not (layer0_outputs(2500));
    outputs(5023) <= not((layer0_outputs(949)) and (layer0_outputs(2422)));
    outputs(5024) <= not(layer0_outputs(2459));
    outputs(5025) <= (layer0_outputs(824)) xor (layer0_outputs(2235));
    outputs(5026) <= not((layer0_outputs(941)) and (layer0_outputs(4972)));
    outputs(5027) <= (layer0_outputs(2197)) and (layer0_outputs(3780));
    outputs(5028) <= (layer0_outputs(667)) or (layer0_outputs(4764));
    outputs(5029) <= layer0_outputs(4638);
    outputs(5030) <= (layer0_outputs(1798)) and not (layer0_outputs(899));
    outputs(5031) <= (layer0_outputs(672)) and not (layer0_outputs(629));
    outputs(5032) <= not((layer0_outputs(5096)) or (layer0_outputs(1249)));
    outputs(5033) <= not(layer0_outputs(2775));
    outputs(5034) <= (layer0_outputs(1669)) and (layer0_outputs(4051));
    outputs(5035) <= (layer0_outputs(2037)) xor (layer0_outputs(767));
    outputs(5036) <= not(layer0_outputs(557));
    outputs(5037) <= not((layer0_outputs(2303)) xor (layer0_outputs(885)));
    outputs(5038) <= layer0_outputs(2907);
    outputs(5039) <= (layer0_outputs(4878)) or (layer0_outputs(2294));
    outputs(5040) <= layer0_outputs(2533);
    outputs(5041) <= (layer0_outputs(4208)) and not (layer0_outputs(1419));
    outputs(5042) <= not((layer0_outputs(4781)) xor (layer0_outputs(994)));
    outputs(5043) <= (layer0_outputs(2048)) and (layer0_outputs(1090));
    outputs(5044) <= not((layer0_outputs(422)) or (layer0_outputs(1116)));
    outputs(5045) <= (layer0_outputs(4625)) and not (layer0_outputs(136));
    outputs(5046) <= (layer0_outputs(1255)) or (layer0_outputs(1737));
    outputs(5047) <= not((layer0_outputs(1578)) or (layer0_outputs(1068)));
    outputs(5048) <= not(layer0_outputs(2620));
    outputs(5049) <= (layer0_outputs(3305)) and (layer0_outputs(3064));
    outputs(5050) <= (layer0_outputs(2941)) and not (layer0_outputs(1359));
    outputs(5051) <= layer0_outputs(460);
    outputs(5052) <= (layer0_outputs(4897)) and (layer0_outputs(2777));
    outputs(5053) <= layer0_outputs(4721);
    outputs(5054) <= (layer0_outputs(3364)) and not (layer0_outputs(75));
    outputs(5055) <= layer0_outputs(4557);
    outputs(5056) <= not((layer0_outputs(2345)) xor (layer0_outputs(3880)));
    outputs(5057) <= not((layer0_outputs(5049)) or (layer0_outputs(2174)));
    outputs(5058) <= not((layer0_outputs(597)) xor (layer0_outputs(4897)));
    outputs(5059) <= not(layer0_outputs(1353));
    outputs(5060) <= not((layer0_outputs(4311)) or (layer0_outputs(861)));
    outputs(5061) <= (layer0_outputs(646)) and not (layer0_outputs(1274));
    outputs(5062) <= (layer0_outputs(831)) and not (layer0_outputs(3902));
    outputs(5063) <= not(layer0_outputs(4581)) or (layer0_outputs(1183));
    outputs(5064) <= (layer0_outputs(2945)) and not (layer0_outputs(3462));
    outputs(5065) <= layer0_outputs(2412);
    outputs(5066) <= (layer0_outputs(917)) and not (layer0_outputs(1859));
    outputs(5067) <= not((layer0_outputs(1796)) or (layer0_outputs(482)));
    outputs(5068) <= not((layer0_outputs(2165)) and (layer0_outputs(3070)));
    outputs(5069) <= not(layer0_outputs(4077)) or (layer0_outputs(3269));
    outputs(5070) <= (layer0_outputs(2864)) and (layer0_outputs(3023));
    outputs(5071) <= (layer0_outputs(1911)) and not (layer0_outputs(1376));
    outputs(5072) <= (layer0_outputs(1155)) and (layer0_outputs(4330));
    outputs(5073) <= (layer0_outputs(3751)) and (layer0_outputs(4978));
    outputs(5074) <= (layer0_outputs(2609)) xor (layer0_outputs(1485));
    outputs(5075) <= layer0_outputs(2970);
    outputs(5076) <= not((layer0_outputs(2833)) or (layer0_outputs(4473)));
    outputs(5077) <= layer0_outputs(4438);
    outputs(5078) <= layer0_outputs(4986);
    outputs(5079) <= not((layer0_outputs(4861)) and (layer0_outputs(3121)));
    outputs(5080) <= not((layer0_outputs(4675)) xor (layer0_outputs(2181)));
    outputs(5081) <= layer0_outputs(2164);
    outputs(5082) <= layer0_outputs(3183);
    outputs(5083) <= not(layer0_outputs(605));
    outputs(5084) <= (layer0_outputs(2255)) and not (layer0_outputs(4616));
    outputs(5085) <= layer0_outputs(874);
    outputs(5086) <= (layer0_outputs(809)) xor (layer0_outputs(2626));
    outputs(5087) <= (layer0_outputs(3066)) xor (layer0_outputs(3166));
    outputs(5088) <= not((layer0_outputs(3616)) or (layer0_outputs(334)));
    outputs(5089) <= layer0_outputs(530);
    outputs(5090) <= layer0_outputs(84);
    outputs(5091) <= not((layer0_outputs(1539)) and (layer0_outputs(3070)));
    outputs(5092) <= not((layer0_outputs(5046)) xor (layer0_outputs(372)));
    outputs(5093) <= (layer0_outputs(4269)) and not (layer0_outputs(4469));
    outputs(5094) <= not((layer0_outputs(3191)) xor (layer0_outputs(681)));
    outputs(5095) <= layer0_outputs(2288);
    outputs(5096) <= (layer0_outputs(4220)) and not (layer0_outputs(3768));
    outputs(5097) <= (layer0_outputs(1181)) and not (layer0_outputs(4603));
    outputs(5098) <= (layer0_outputs(2553)) and not (layer0_outputs(1310));
    outputs(5099) <= layer0_outputs(802);
    outputs(5100) <= not(layer0_outputs(3036));
    outputs(5101) <= layer0_outputs(2572);
    outputs(5102) <= not((layer0_outputs(2474)) xor (layer0_outputs(1278)));
    outputs(5103) <= (layer0_outputs(1315)) and (layer0_outputs(4296));
    outputs(5104) <= not((layer0_outputs(908)) or (layer0_outputs(2832)));
    outputs(5105) <= layer0_outputs(1653);
    outputs(5106) <= layer0_outputs(2438);
    outputs(5107) <= (layer0_outputs(3777)) xor (layer0_outputs(581));
    outputs(5108) <= not((layer0_outputs(3828)) xor (layer0_outputs(4417)));
    outputs(5109) <= not((layer0_outputs(565)) or (layer0_outputs(1704)));
    outputs(5110) <= (layer0_outputs(2755)) xor (layer0_outputs(2118));
    outputs(5111) <= not((layer0_outputs(2115)) and (layer0_outputs(4790)));
    outputs(5112) <= (layer0_outputs(645)) xor (layer0_outputs(4062));
    outputs(5113) <= '0';
    outputs(5114) <= not((layer0_outputs(2537)) or (layer0_outputs(359)));
    outputs(5115) <= layer0_outputs(2402);
    outputs(5116) <= (layer0_outputs(4088)) and not (layer0_outputs(3512));
    outputs(5117) <= (layer0_outputs(2497)) and not (layer0_outputs(4928));
    outputs(5118) <= (layer0_outputs(1517)) and not (layer0_outputs(4663));
    outputs(5119) <= (layer0_outputs(3017)) and not (layer0_outputs(3599));

end Behavioral;
