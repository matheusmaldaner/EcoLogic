library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(2559 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(2559 downto 0);

begin

    layer0_outputs(0) <= not(inputs(13));
    layer0_outputs(1) <= (inputs(215)) and not (inputs(225));
    layer0_outputs(2) <= not((inputs(248)) or (inputs(239)));
    layer0_outputs(3) <= not((inputs(180)) xor (inputs(193)));
    layer0_outputs(4) <= not(inputs(24)) or (inputs(254));
    layer0_outputs(5) <= not((inputs(204)) or (inputs(61)));
    layer0_outputs(6) <= (inputs(41)) or (inputs(96));
    layer0_outputs(7) <= (inputs(120)) and not (inputs(178));
    layer0_outputs(8) <= '1';
    layer0_outputs(9) <= not((inputs(142)) or (inputs(55)));
    layer0_outputs(10) <= (inputs(222)) or (inputs(117));
    layer0_outputs(11) <= (inputs(136)) or (inputs(254));
    layer0_outputs(12) <= not((inputs(45)) or (inputs(176)));
    layer0_outputs(13) <= '1';
    layer0_outputs(14) <= inputs(239);
    layer0_outputs(15) <= '0';
    layer0_outputs(16) <= inputs(18);
    layer0_outputs(17) <= (inputs(186)) and not (inputs(71));
    layer0_outputs(18) <= not((inputs(246)) and (inputs(111)));
    layer0_outputs(19) <= not(inputs(136));
    layer0_outputs(20) <= (inputs(47)) or (inputs(24));
    layer0_outputs(21) <= not(inputs(41)) or (inputs(149));
    layer0_outputs(22) <= inputs(47);
    layer0_outputs(23) <= (inputs(149)) and not (inputs(15));
    layer0_outputs(24) <= inputs(57);
    layer0_outputs(25) <= not(inputs(24)) or (inputs(239));
    layer0_outputs(26) <= not(inputs(60)) or (inputs(32));
    layer0_outputs(27) <= not(inputs(211));
    layer0_outputs(28) <= not(inputs(253));
    layer0_outputs(29) <= not(inputs(29)) or (inputs(179));
    layer0_outputs(30) <= (inputs(210)) and not (inputs(2));
    layer0_outputs(31) <= inputs(100);
    layer0_outputs(32) <= (inputs(21)) or (inputs(5));
    layer0_outputs(33) <= not(inputs(246));
    layer0_outputs(34) <= not((inputs(111)) and (inputs(17)));
    layer0_outputs(35) <= not(inputs(85));
    layer0_outputs(36) <= inputs(100);
    layer0_outputs(37) <= inputs(179);
    layer0_outputs(38) <= (inputs(140)) or (inputs(2));
    layer0_outputs(39) <= inputs(178);
    layer0_outputs(40) <= not(inputs(196)) or (inputs(101));
    layer0_outputs(41) <= not(inputs(29));
    layer0_outputs(42) <= not(inputs(196));
    layer0_outputs(43) <= (inputs(49)) xor (inputs(47));
    layer0_outputs(44) <= not((inputs(99)) or (inputs(97)));
    layer0_outputs(45) <= inputs(111);
    layer0_outputs(46) <= not(inputs(105));
    layer0_outputs(47) <= inputs(127);
    layer0_outputs(48) <= inputs(92);
    layer0_outputs(49) <= inputs(105);
    layer0_outputs(50) <= not(inputs(42));
    layer0_outputs(51) <= not(inputs(169)) or (inputs(31));
    layer0_outputs(52) <= not(inputs(136)) or (inputs(180));
    layer0_outputs(53) <= not(inputs(62));
    layer0_outputs(54) <= not(inputs(67));
    layer0_outputs(55) <= '0';
    layer0_outputs(56) <= not(inputs(117));
    layer0_outputs(57) <= not(inputs(10)) or (inputs(227));
    layer0_outputs(58) <= (inputs(123)) and not (inputs(94));
    layer0_outputs(59) <= not(inputs(59));
    layer0_outputs(60) <= (inputs(212)) or (inputs(86));
    layer0_outputs(61) <= not(inputs(191)) or (inputs(156));
    layer0_outputs(62) <= not(inputs(228));
    layer0_outputs(63) <= inputs(109);
    layer0_outputs(64) <= (inputs(55)) and not (inputs(75));
    layer0_outputs(65) <= not(inputs(114));
    layer0_outputs(66) <= inputs(175);
    layer0_outputs(67) <= not((inputs(0)) or (inputs(63)));
    layer0_outputs(68) <= inputs(146);
    layer0_outputs(69) <= not((inputs(21)) or (inputs(234)));
    layer0_outputs(70) <= not(inputs(55));
    layer0_outputs(71) <= not(inputs(241)) or (inputs(199));
    layer0_outputs(72) <= not(inputs(107));
    layer0_outputs(73) <= not((inputs(184)) or (inputs(237)));
    layer0_outputs(74) <= not((inputs(72)) or (inputs(84)));
    layer0_outputs(75) <= not((inputs(180)) or (inputs(59)));
    layer0_outputs(76) <= (inputs(160)) or (inputs(94));
    layer0_outputs(77) <= '1';
    layer0_outputs(78) <= not(inputs(66));
    layer0_outputs(79) <= not(inputs(145)) or (inputs(112));
    layer0_outputs(80) <= inputs(226);
    layer0_outputs(81) <= not(inputs(110));
    layer0_outputs(82) <= (inputs(14)) or (inputs(136));
    layer0_outputs(83) <= not(inputs(189)) or (inputs(129));
    layer0_outputs(84) <= (inputs(71)) and not (inputs(91));
    layer0_outputs(85) <= not(inputs(27)) or (inputs(170));
    layer0_outputs(86) <= not(inputs(234));
    layer0_outputs(87) <= (inputs(193)) or (inputs(213));
    layer0_outputs(88) <= (inputs(173)) and not (inputs(152));
    layer0_outputs(89) <= not((inputs(240)) or (inputs(224)));
    layer0_outputs(90) <= (inputs(64)) or (inputs(177));
    layer0_outputs(91) <= not(inputs(237));
    layer0_outputs(92) <= (inputs(48)) and not (inputs(12));
    layer0_outputs(93) <= not((inputs(236)) or (inputs(174)));
    layer0_outputs(94) <= '1';
    layer0_outputs(95) <= inputs(196);
    layer0_outputs(96) <= not(inputs(186)) or (inputs(13));
    layer0_outputs(97) <= (inputs(51)) or (inputs(13));
    layer0_outputs(98) <= (inputs(117)) or (inputs(149));
    layer0_outputs(99) <= inputs(175);
    layer0_outputs(100) <= inputs(5);
    layer0_outputs(101) <= not(inputs(195)) or (inputs(28));
    layer0_outputs(102) <= '0';
    layer0_outputs(103) <= not(inputs(237));
    layer0_outputs(104) <= (inputs(60)) and not (inputs(160));
    layer0_outputs(105) <= (inputs(204)) and not (inputs(1));
    layer0_outputs(106) <= '1';
    layer0_outputs(107) <= (inputs(153)) or (inputs(200));
    layer0_outputs(108) <= not(inputs(135));
    layer0_outputs(109) <= inputs(164);
    layer0_outputs(110) <= not((inputs(113)) xor (inputs(147)));
    layer0_outputs(111) <= inputs(43);
    layer0_outputs(112) <= not(inputs(189)) or (inputs(253));
    layer0_outputs(113) <= not((inputs(1)) or (inputs(205)));
    layer0_outputs(114) <= inputs(131);
    layer0_outputs(115) <= not(inputs(146));
    layer0_outputs(116) <= not((inputs(110)) or (inputs(116)));
    layer0_outputs(117) <= (inputs(118)) or (inputs(0));
    layer0_outputs(118) <= inputs(126);
    layer0_outputs(119) <= (inputs(25)) and not (inputs(159));
    layer0_outputs(120) <= inputs(36);
    layer0_outputs(121) <= (inputs(31)) or (inputs(246));
    layer0_outputs(122) <= (inputs(254)) or (inputs(121));
    layer0_outputs(123) <= not((inputs(191)) or (inputs(215)));
    layer0_outputs(124) <= (inputs(151)) and not (inputs(126));
    layer0_outputs(125) <= not((inputs(53)) and (inputs(49)));
    layer0_outputs(126) <= not(inputs(166));
    layer0_outputs(127) <= inputs(111);
    layer0_outputs(128) <= inputs(182);
    layer0_outputs(129) <= (inputs(186)) and not (inputs(208));
    layer0_outputs(130) <= not(inputs(178));
    layer0_outputs(131) <= not((inputs(88)) or (inputs(173)));
    layer0_outputs(132) <= not(inputs(100));
    layer0_outputs(133) <= (inputs(152)) and not (inputs(189));
    layer0_outputs(134) <= (inputs(209)) or (inputs(220));
    layer0_outputs(135) <= inputs(124);
    layer0_outputs(136) <= inputs(14);
    layer0_outputs(137) <= not((inputs(121)) or (inputs(33)));
    layer0_outputs(138) <= not((inputs(233)) and (inputs(197)));
    layer0_outputs(139) <= inputs(120);
    layer0_outputs(140) <= not(inputs(6));
    layer0_outputs(141) <= inputs(157);
    layer0_outputs(142) <= not((inputs(183)) and (inputs(189)));
    layer0_outputs(143) <= inputs(176);
    layer0_outputs(144) <= not((inputs(109)) or (inputs(254)));
    layer0_outputs(145) <= not((inputs(98)) or (inputs(14)));
    layer0_outputs(146) <= not(inputs(137)) or (inputs(4));
    layer0_outputs(147) <= not((inputs(6)) or (inputs(32)));
    layer0_outputs(148) <= (inputs(160)) and not (inputs(241));
    layer0_outputs(149) <= (inputs(156)) or (inputs(125));
    layer0_outputs(150) <= inputs(146);
    layer0_outputs(151) <= inputs(133);
    layer0_outputs(152) <= (inputs(76)) or (inputs(193));
    layer0_outputs(153) <= (inputs(40)) and not (inputs(40));
    layer0_outputs(154) <= not(inputs(26)) or (inputs(64));
    layer0_outputs(155) <= (inputs(94)) or (inputs(238));
    layer0_outputs(156) <= (inputs(23)) and not (inputs(184));
    layer0_outputs(157) <= not((inputs(131)) or (inputs(142)));
    layer0_outputs(158) <= not(inputs(99));
    layer0_outputs(159) <= inputs(103);
    layer0_outputs(160) <= (inputs(125)) xor (inputs(61));
    layer0_outputs(161) <= inputs(247);
    layer0_outputs(162) <= (inputs(2)) or (inputs(136));
    layer0_outputs(163) <= not(inputs(53));
    layer0_outputs(164) <= not((inputs(25)) or (inputs(192)));
    layer0_outputs(165) <= (inputs(151)) and not (inputs(78));
    layer0_outputs(166) <= not(inputs(145));
    layer0_outputs(167) <= (inputs(68)) and not (inputs(95));
    layer0_outputs(168) <= (inputs(44)) and not (inputs(158));
    layer0_outputs(169) <= '1';
    layer0_outputs(170) <= not(inputs(90));
    layer0_outputs(171) <= '0';
    layer0_outputs(172) <= not((inputs(9)) or (inputs(26)));
    layer0_outputs(173) <= inputs(106);
    layer0_outputs(174) <= inputs(103);
    layer0_outputs(175) <= (inputs(163)) or (inputs(99));
    layer0_outputs(176) <= (inputs(205)) and (inputs(200));
    layer0_outputs(177) <= (inputs(228)) or (inputs(208));
    layer0_outputs(178) <= not(inputs(121));
    layer0_outputs(179) <= inputs(59);
    layer0_outputs(180) <= '1';
    layer0_outputs(181) <= '1';
    layer0_outputs(182) <= inputs(118);
    layer0_outputs(183) <= not(inputs(104));
    layer0_outputs(184) <= not((inputs(31)) or (inputs(30)));
    layer0_outputs(185) <= not(inputs(71)) or (inputs(142));
    layer0_outputs(186) <= (inputs(181)) or (inputs(225));
    layer0_outputs(187) <= (inputs(27)) or (inputs(94));
    layer0_outputs(188) <= not(inputs(197)) or (inputs(45));
    layer0_outputs(189) <= (inputs(5)) and not (inputs(133));
    layer0_outputs(190) <= inputs(247);
    layer0_outputs(191) <= inputs(164);
    layer0_outputs(192) <= not((inputs(143)) or (inputs(166)));
    layer0_outputs(193) <= not((inputs(168)) and (inputs(5)));
    layer0_outputs(194) <= (inputs(59)) xor (inputs(22));
    layer0_outputs(195) <= not((inputs(15)) or (inputs(225)));
    layer0_outputs(196) <= (inputs(172)) xor (inputs(76));
    layer0_outputs(197) <= not(inputs(216)) or (inputs(61));
    layer0_outputs(198) <= (inputs(38)) and not (inputs(234));
    layer0_outputs(199) <= not(inputs(51)) or (inputs(157));
    layer0_outputs(200) <= (inputs(34)) or (inputs(46));
    layer0_outputs(201) <= inputs(85);
    layer0_outputs(202) <= not((inputs(9)) and (inputs(89)));
    layer0_outputs(203) <= not((inputs(187)) or (inputs(253)));
    layer0_outputs(204) <= not(inputs(98));
    layer0_outputs(205) <= not(inputs(76));
    layer0_outputs(206) <= not(inputs(142)) or (inputs(0));
    layer0_outputs(207) <= not(inputs(130));
    layer0_outputs(208) <= (inputs(221)) and (inputs(238));
    layer0_outputs(209) <= not(inputs(243));
    layer0_outputs(210) <= (inputs(174)) and not (inputs(115));
    layer0_outputs(211) <= (inputs(106)) or (inputs(93));
    layer0_outputs(212) <= not(inputs(152)) or (inputs(66));
    layer0_outputs(213) <= (inputs(191)) and not (inputs(95));
    layer0_outputs(214) <= not((inputs(171)) xor (inputs(120)));
    layer0_outputs(215) <= not(inputs(41)) or (inputs(165));
    layer0_outputs(216) <= (inputs(232)) and not (inputs(13));
    layer0_outputs(217) <= not(inputs(217)) or (inputs(45));
    layer0_outputs(218) <= (inputs(104)) and not (inputs(48));
    layer0_outputs(219) <= (inputs(84)) and not (inputs(48));
    layer0_outputs(220) <= not(inputs(38)) or (inputs(139));
    layer0_outputs(221) <= not((inputs(230)) xor (inputs(38)));
    layer0_outputs(222) <= not((inputs(205)) or (inputs(18)));
    layer0_outputs(223) <= (inputs(32)) or (inputs(30));
    layer0_outputs(224) <= inputs(124);
    layer0_outputs(225) <= inputs(66);
    layer0_outputs(226) <= inputs(74);
    layer0_outputs(227) <= not(inputs(195));
    layer0_outputs(228) <= not(inputs(155));
    layer0_outputs(229) <= not(inputs(245));
    layer0_outputs(230) <= inputs(121);
    layer0_outputs(231) <= not((inputs(170)) or (inputs(4)));
    layer0_outputs(232) <= not((inputs(112)) or (inputs(123)));
    layer0_outputs(233) <= not(inputs(116)) or (inputs(14));
    layer0_outputs(234) <= not(inputs(154)) or (inputs(26));
    layer0_outputs(235) <= inputs(196);
    layer0_outputs(236) <= not(inputs(158)) or (inputs(238));
    layer0_outputs(237) <= '1';
    layer0_outputs(238) <= (inputs(216)) and not (inputs(145));
    layer0_outputs(239) <= not(inputs(199));
    layer0_outputs(240) <= (inputs(173)) or (inputs(180));
    layer0_outputs(241) <= inputs(120);
    layer0_outputs(242) <= not(inputs(141));
    layer0_outputs(243) <= not((inputs(206)) and (inputs(206)));
    layer0_outputs(244) <= inputs(119);
    layer0_outputs(245) <= not(inputs(53)) or (inputs(42));
    layer0_outputs(246) <= not(inputs(39));
    layer0_outputs(247) <= (inputs(113)) xor (inputs(55));
    layer0_outputs(248) <= not(inputs(42));
    layer0_outputs(249) <= inputs(183);
    layer0_outputs(250) <= inputs(132);
    layer0_outputs(251) <= inputs(121);
    layer0_outputs(252) <= not(inputs(36));
    layer0_outputs(253) <= not(inputs(152));
    layer0_outputs(254) <= '1';
    layer0_outputs(255) <= (inputs(211)) and not (inputs(81));
    layer0_outputs(256) <= '1';
    layer0_outputs(257) <= not(inputs(232));
    layer0_outputs(258) <= inputs(115);
    layer0_outputs(259) <= (inputs(54)) and not (inputs(47));
    layer0_outputs(260) <= (inputs(222)) or (inputs(174));
    layer0_outputs(261) <= not((inputs(189)) or (inputs(54)));
    layer0_outputs(262) <= not(inputs(106)) or (inputs(17));
    layer0_outputs(263) <= inputs(121);
    layer0_outputs(264) <= not(inputs(123));
    layer0_outputs(265) <= (inputs(204)) and not (inputs(15));
    layer0_outputs(266) <= inputs(47);
    layer0_outputs(267) <= not(inputs(130));
    layer0_outputs(268) <= not(inputs(152));
    layer0_outputs(269) <= not((inputs(189)) or (inputs(125)));
    layer0_outputs(270) <= inputs(223);
    layer0_outputs(271) <= not((inputs(4)) xor (inputs(160)));
    layer0_outputs(272) <= not((inputs(152)) or (inputs(236)));
    layer0_outputs(273) <= not(inputs(188)) or (inputs(240));
    layer0_outputs(274) <= not((inputs(131)) or (inputs(124)));
    layer0_outputs(275) <= not(inputs(138));
    layer0_outputs(276) <= inputs(124);
    layer0_outputs(277) <= (inputs(19)) or (inputs(158));
    layer0_outputs(278) <= not(inputs(164));
    layer0_outputs(279) <= (inputs(173)) or (inputs(158));
    layer0_outputs(280) <= not((inputs(2)) or (inputs(177)));
    layer0_outputs(281) <= (inputs(174)) and not (inputs(251));
    layer0_outputs(282) <= not(inputs(121));
    layer0_outputs(283) <= (inputs(202)) or (inputs(136));
    layer0_outputs(284) <= inputs(216);
    layer0_outputs(285) <= (inputs(138)) or (inputs(198));
    layer0_outputs(286) <= not((inputs(85)) or (inputs(143)));
    layer0_outputs(287) <= (inputs(255)) or (inputs(83));
    layer0_outputs(288) <= (inputs(83)) or (inputs(158));
    layer0_outputs(289) <= inputs(206);
    layer0_outputs(290) <= not(inputs(85));
    layer0_outputs(291) <= not(inputs(230)) or (inputs(29));
    layer0_outputs(292) <= not(inputs(27));
    layer0_outputs(293) <= (inputs(77)) or (inputs(143));
    layer0_outputs(294) <= not((inputs(176)) or (inputs(177)));
    layer0_outputs(295) <= not(inputs(119)) or (inputs(207));
    layer0_outputs(296) <= (inputs(177)) or (inputs(89));
    layer0_outputs(297) <= not(inputs(44));
    layer0_outputs(298) <= (inputs(216)) and (inputs(240));
    layer0_outputs(299) <= not((inputs(150)) or (inputs(13)));
    layer0_outputs(300) <= inputs(167);
    layer0_outputs(301) <= inputs(149);
    layer0_outputs(302) <= (inputs(255)) xor (inputs(44));
    layer0_outputs(303) <= inputs(115);
    layer0_outputs(304) <= not(inputs(26)) or (inputs(190));
    layer0_outputs(305) <= not(inputs(185)) or (inputs(81));
    layer0_outputs(306) <= not(inputs(84));
    layer0_outputs(307) <= (inputs(103)) or (inputs(117));
    layer0_outputs(308) <= (inputs(114)) or (inputs(135));
    layer0_outputs(309) <= (inputs(199)) and not (inputs(207));
    layer0_outputs(310) <= inputs(103);
    layer0_outputs(311) <= (inputs(236)) or (inputs(215));
    layer0_outputs(312) <= inputs(9);
    layer0_outputs(313) <= (inputs(249)) or (inputs(76));
    layer0_outputs(314) <= (inputs(242)) xor (inputs(235));
    layer0_outputs(315) <= not(inputs(172));
    layer0_outputs(316) <= inputs(75);
    layer0_outputs(317) <= (inputs(108)) or (inputs(52));
    layer0_outputs(318) <= not(inputs(88));
    layer0_outputs(319) <= not(inputs(235));
    layer0_outputs(320) <= not((inputs(141)) xor (inputs(121)));
    layer0_outputs(321) <= inputs(152);
    layer0_outputs(322) <= (inputs(182)) xor (inputs(77));
    layer0_outputs(323) <= (inputs(91)) or (inputs(60));
    layer0_outputs(324) <= not(inputs(182));
    layer0_outputs(325) <= (inputs(122)) and not (inputs(12));
    layer0_outputs(326) <= not(inputs(180));
    layer0_outputs(327) <= inputs(183);
    layer0_outputs(328) <= not(inputs(91));
    layer0_outputs(329) <= (inputs(26)) and not (inputs(222));
    layer0_outputs(330) <= (inputs(51)) or (inputs(42));
    layer0_outputs(331) <= (inputs(251)) or (inputs(254));
    layer0_outputs(332) <= (inputs(122)) and not (inputs(10));
    layer0_outputs(333) <= not((inputs(49)) xor (inputs(110)));
    layer0_outputs(334) <= not(inputs(50)) or (inputs(173));
    layer0_outputs(335) <= (inputs(192)) and not (inputs(158));
    layer0_outputs(336) <= not(inputs(115));
    layer0_outputs(337) <= not((inputs(203)) or (inputs(193)));
    layer0_outputs(338) <= not(inputs(102));
    layer0_outputs(339) <= not(inputs(88));
    layer0_outputs(340) <= (inputs(102)) or (inputs(130));
    layer0_outputs(341) <= not(inputs(151));
    layer0_outputs(342) <= not((inputs(126)) xor (inputs(180)));
    layer0_outputs(343) <= (inputs(94)) xor (inputs(63));
    layer0_outputs(344) <= not((inputs(146)) or (inputs(169)));
    layer0_outputs(345) <= (inputs(196)) and not (inputs(107));
    layer0_outputs(346) <= not(inputs(195)) or (inputs(121));
    layer0_outputs(347) <= not(inputs(133)) or (inputs(63));
    layer0_outputs(348) <= not(inputs(67)) or (inputs(211));
    layer0_outputs(349) <= '0';
    layer0_outputs(350) <= not(inputs(35));
    layer0_outputs(351) <= (inputs(43)) and not (inputs(72));
    layer0_outputs(352) <= (inputs(143)) or (inputs(133));
    layer0_outputs(353) <= not(inputs(205));
    layer0_outputs(354) <= (inputs(223)) xor (inputs(180));
    layer0_outputs(355) <= inputs(120);
    layer0_outputs(356) <= (inputs(237)) and not (inputs(80));
    layer0_outputs(357) <= inputs(97);
    layer0_outputs(358) <= not(inputs(126));
    layer0_outputs(359) <= (inputs(79)) or (inputs(58));
    layer0_outputs(360) <= (inputs(105)) and not (inputs(172));
    layer0_outputs(361) <= not((inputs(162)) or (inputs(122)));
    layer0_outputs(362) <= (inputs(86)) or (inputs(190));
    layer0_outputs(363) <= not(inputs(72));
    layer0_outputs(364) <= not(inputs(56));
    layer0_outputs(365) <= '0';
    layer0_outputs(366) <= (inputs(187)) and not (inputs(97));
    layer0_outputs(367) <= not(inputs(57));
    layer0_outputs(368) <= not((inputs(118)) or (inputs(85)));
    layer0_outputs(369) <= not(inputs(211)) or (inputs(95));
    layer0_outputs(370) <= not(inputs(235));
    layer0_outputs(371) <= (inputs(17)) and not (inputs(189));
    layer0_outputs(372) <= inputs(161);
    layer0_outputs(373) <= (inputs(229)) and not (inputs(88));
    layer0_outputs(374) <= not(inputs(165));
    layer0_outputs(375) <= not((inputs(4)) or (inputs(52)));
    layer0_outputs(376) <= not((inputs(163)) or (inputs(111)));
    layer0_outputs(377) <= not((inputs(118)) or (inputs(31)));
    layer0_outputs(378) <= (inputs(200)) or (inputs(238));
    layer0_outputs(379) <= inputs(63);
    layer0_outputs(380) <= not(inputs(203)) or (inputs(225));
    layer0_outputs(381) <= not(inputs(25)) or (inputs(134));
    layer0_outputs(382) <= not(inputs(132));
    layer0_outputs(383) <= not((inputs(175)) or (inputs(68)));
    layer0_outputs(384) <= not(inputs(28)) or (inputs(16));
    layer0_outputs(385) <= not((inputs(139)) and (inputs(109)));
    layer0_outputs(386) <= not((inputs(147)) xor (inputs(100)));
    layer0_outputs(387) <= not(inputs(234)) or (inputs(127));
    layer0_outputs(388) <= not((inputs(178)) or (inputs(195)));
    layer0_outputs(389) <= not(inputs(102)) or (inputs(33));
    layer0_outputs(390) <= (inputs(121)) and not (inputs(251));
    layer0_outputs(391) <= (inputs(162)) or (inputs(58));
    layer0_outputs(392) <= inputs(227);
    layer0_outputs(393) <= (inputs(182)) or (inputs(98));
    layer0_outputs(394) <= '0';
    layer0_outputs(395) <= not(inputs(87));
    layer0_outputs(396) <= inputs(103);
    layer0_outputs(397) <= not(inputs(191)) or (inputs(44));
    layer0_outputs(398) <= not(inputs(63));
    layer0_outputs(399) <= not(inputs(21));
    layer0_outputs(400) <= not(inputs(91));
    layer0_outputs(401) <= not(inputs(20));
    layer0_outputs(402) <= not(inputs(135));
    layer0_outputs(403) <= not(inputs(153));
    layer0_outputs(404) <= not(inputs(73)) or (inputs(225));
    layer0_outputs(405) <= (inputs(188)) and not (inputs(109));
    layer0_outputs(406) <= not(inputs(135));
    layer0_outputs(407) <= not((inputs(24)) and (inputs(243)));
    layer0_outputs(408) <= not(inputs(89));
    layer0_outputs(409) <= inputs(67);
    layer0_outputs(410) <= (inputs(22)) and (inputs(232));
    layer0_outputs(411) <= (inputs(151)) and not (inputs(221));
    layer0_outputs(412) <= inputs(144);
    layer0_outputs(413) <= inputs(202);
    layer0_outputs(414) <= inputs(85);
    layer0_outputs(415) <= (inputs(126)) or (inputs(137));
    layer0_outputs(416) <= inputs(171);
    layer0_outputs(417) <= inputs(137);
    layer0_outputs(418) <= inputs(196);
    layer0_outputs(419) <= inputs(213);
    layer0_outputs(420) <= not(inputs(1));
    layer0_outputs(421) <= not((inputs(220)) or (inputs(190)));
    layer0_outputs(422) <= inputs(15);
    layer0_outputs(423) <= (inputs(214)) or (inputs(207));
    layer0_outputs(424) <= not((inputs(41)) and (inputs(42)));
    layer0_outputs(425) <= (inputs(65)) and not (inputs(158));
    layer0_outputs(426) <= (inputs(85)) and not (inputs(223));
    layer0_outputs(427) <= '0';
    layer0_outputs(428) <= not(inputs(35));
    layer0_outputs(429) <= inputs(117);
    layer0_outputs(430) <= (inputs(226)) and not (inputs(129));
    layer0_outputs(431) <= inputs(96);
    layer0_outputs(432) <= inputs(247);
    layer0_outputs(433) <= (inputs(190)) or (inputs(194));
    layer0_outputs(434) <= (inputs(131)) xor (inputs(159));
    layer0_outputs(435) <= not((inputs(27)) or (inputs(33)));
    layer0_outputs(436) <= not(inputs(216));
    layer0_outputs(437) <= not((inputs(242)) and (inputs(27)));
    layer0_outputs(438) <= (inputs(195)) and not (inputs(113));
    layer0_outputs(439) <= not((inputs(84)) or (inputs(112)));
    layer0_outputs(440) <= not((inputs(177)) or (inputs(24)));
    layer0_outputs(441) <= inputs(248);
    layer0_outputs(442) <= not(inputs(128)) or (inputs(255));
    layer0_outputs(443) <= not((inputs(82)) or (inputs(64)));
    layer0_outputs(444) <= (inputs(209)) or (inputs(202));
    layer0_outputs(445) <= (inputs(31)) or (inputs(144));
    layer0_outputs(446) <= inputs(179);
    layer0_outputs(447) <= inputs(84);
    layer0_outputs(448) <= not(inputs(43)) or (inputs(241));
    layer0_outputs(449) <= inputs(37);
    layer0_outputs(450) <= inputs(120);
    layer0_outputs(451) <= inputs(179);
    layer0_outputs(452) <= inputs(230);
    layer0_outputs(453) <= (inputs(150)) and not (inputs(194));
    layer0_outputs(454) <= inputs(134);
    layer0_outputs(455) <= not(inputs(148)) or (inputs(187));
    layer0_outputs(456) <= not(inputs(24));
    layer0_outputs(457) <= (inputs(32)) or (inputs(168));
    layer0_outputs(458) <= not((inputs(229)) and (inputs(164)));
    layer0_outputs(459) <= not(inputs(87));
    layer0_outputs(460) <= inputs(118);
    layer0_outputs(461) <= not(inputs(219)) or (inputs(238));
    layer0_outputs(462) <= not(inputs(73));
    layer0_outputs(463) <= not(inputs(92)) or (inputs(143));
    layer0_outputs(464) <= (inputs(71)) and not (inputs(124));
    layer0_outputs(465) <= (inputs(59)) and not (inputs(87));
    layer0_outputs(466) <= inputs(83);
    layer0_outputs(467) <= not(inputs(174)) or (inputs(111));
    layer0_outputs(468) <= not((inputs(195)) or (inputs(213)));
    layer0_outputs(469) <= not((inputs(119)) and (inputs(94)));
    layer0_outputs(470) <= (inputs(128)) and (inputs(236));
    layer0_outputs(471) <= not(inputs(102));
    layer0_outputs(472) <= not(inputs(48)) or (inputs(160));
    layer0_outputs(473) <= (inputs(235)) xor (inputs(170));
    layer0_outputs(474) <= (inputs(87)) and not (inputs(64));
    layer0_outputs(475) <= (inputs(36)) and not (inputs(130));
    layer0_outputs(476) <= inputs(129);
    layer0_outputs(477) <= (inputs(2)) and not (inputs(129));
    layer0_outputs(478) <= not((inputs(246)) or (inputs(34)));
    layer0_outputs(479) <= inputs(170);
    layer0_outputs(480) <= (inputs(184)) and not (inputs(111));
    layer0_outputs(481) <= not((inputs(214)) or (inputs(191)));
    layer0_outputs(482) <= inputs(140);
    layer0_outputs(483) <= not((inputs(107)) xor (inputs(197)));
    layer0_outputs(484) <= not(inputs(166));
    layer0_outputs(485) <= inputs(78);
    layer0_outputs(486) <= inputs(84);
    layer0_outputs(487) <= not(inputs(232)) or (inputs(12));
    layer0_outputs(488) <= not(inputs(216));
    layer0_outputs(489) <= inputs(117);
    layer0_outputs(490) <= not((inputs(34)) or (inputs(241)));
    layer0_outputs(491) <= not(inputs(148)) or (inputs(92));
    layer0_outputs(492) <= (inputs(254)) or (inputs(163));
    layer0_outputs(493) <= not((inputs(60)) or (inputs(21)));
    layer0_outputs(494) <= not(inputs(187)) or (inputs(1));
    layer0_outputs(495) <= not((inputs(118)) xor (inputs(68)));
    layer0_outputs(496) <= not(inputs(148));
    layer0_outputs(497) <= inputs(153);
    layer0_outputs(498) <= not(inputs(63));
    layer0_outputs(499) <= inputs(5);
    layer0_outputs(500) <= (inputs(239)) or (inputs(126));
    layer0_outputs(501) <= (inputs(177)) xor (inputs(147));
    layer0_outputs(502) <= not((inputs(80)) or (inputs(147)));
    layer0_outputs(503) <= not((inputs(162)) or (inputs(216)));
    layer0_outputs(504) <= not(inputs(70)) or (inputs(121));
    layer0_outputs(505) <= inputs(67);
    layer0_outputs(506) <= (inputs(227)) and not (inputs(92));
    layer0_outputs(507) <= (inputs(250)) and (inputs(171));
    layer0_outputs(508) <= not(inputs(1));
    layer0_outputs(509) <= (inputs(199)) xor (inputs(225));
    layer0_outputs(510) <= not(inputs(162));
    layer0_outputs(511) <= not((inputs(214)) xor (inputs(111)));
    layer0_outputs(512) <= not((inputs(147)) or (inputs(132)));
    layer0_outputs(513) <= not(inputs(107));
    layer0_outputs(514) <= not(inputs(88));
    layer0_outputs(515) <= inputs(195);
    layer0_outputs(516) <= (inputs(47)) or (inputs(188));
    layer0_outputs(517) <= not((inputs(88)) or (inputs(218)));
    layer0_outputs(518) <= (inputs(98)) or (inputs(81));
    layer0_outputs(519) <= not(inputs(22));
    layer0_outputs(520) <= not((inputs(138)) or (inputs(235)));
    layer0_outputs(521) <= (inputs(60)) and (inputs(73));
    layer0_outputs(522) <= (inputs(245)) and not (inputs(153));
    layer0_outputs(523) <= not(inputs(185));
    layer0_outputs(524) <= not(inputs(52));
    layer0_outputs(525) <= inputs(54);
    layer0_outputs(526) <= inputs(192);
    layer0_outputs(527) <= not((inputs(226)) xor (inputs(62)));
    layer0_outputs(528) <= not(inputs(111));
    layer0_outputs(529) <= not(inputs(245));
    layer0_outputs(530) <= inputs(189);
    layer0_outputs(531) <= not(inputs(123));
    layer0_outputs(532) <= not(inputs(64)) or (inputs(96));
    layer0_outputs(533) <= not((inputs(227)) and (inputs(33)));
    layer0_outputs(534) <= not(inputs(93));
    layer0_outputs(535) <= inputs(100);
    layer0_outputs(536) <= (inputs(214)) and not (inputs(253));
    layer0_outputs(537) <= inputs(153);
    layer0_outputs(538) <= not(inputs(246));
    layer0_outputs(539) <= (inputs(63)) or (inputs(248));
    layer0_outputs(540) <= (inputs(216)) xor (inputs(249));
    layer0_outputs(541) <= (inputs(109)) or (inputs(18));
    layer0_outputs(542) <= (inputs(148)) and not (inputs(94));
    layer0_outputs(543) <= not(inputs(115));
    layer0_outputs(544) <= not(inputs(150));
    layer0_outputs(545) <= (inputs(30)) and (inputs(229));
    layer0_outputs(546) <= (inputs(19)) or (inputs(31));
    layer0_outputs(547) <= inputs(23);
    layer0_outputs(548) <= inputs(89);
    layer0_outputs(549) <= not(inputs(89));
    layer0_outputs(550) <= (inputs(169)) or (inputs(106));
    layer0_outputs(551) <= inputs(230);
    layer0_outputs(552) <= (inputs(223)) or (inputs(109));
    layer0_outputs(553) <= inputs(189);
    layer0_outputs(554) <= (inputs(9)) and not (inputs(113));
    layer0_outputs(555) <= not((inputs(6)) or (inputs(158)));
    layer0_outputs(556) <= (inputs(60)) and not (inputs(220));
    layer0_outputs(557) <= not(inputs(210));
    layer0_outputs(558) <= (inputs(62)) or (inputs(155));
    layer0_outputs(559) <= inputs(116);
    layer0_outputs(560) <= not(inputs(205));
    layer0_outputs(561) <= inputs(193);
    layer0_outputs(562) <= not((inputs(21)) and (inputs(29)));
    layer0_outputs(563) <= not((inputs(206)) or (inputs(213)));
    layer0_outputs(564) <= not(inputs(233));
    layer0_outputs(565) <= inputs(182);
    layer0_outputs(566) <= not(inputs(99));
    layer0_outputs(567) <= (inputs(83)) and not (inputs(54));
    layer0_outputs(568) <= (inputs(47)) or (inputs(23));
    layer0_outputs(569) <= not((inputs(191)) or (inputs(208)));
    layer0_outputs(570) <= (inputs(52)) and not (inputs(222));
    layer0_outputs(571) <= inputs(211);
    layer0_outputs(572) <= '1';
    layer0_outputs(573) <= not(inputs(75)) or (inputs(3));
    layer0_outputs(574) <= not(inputs(114));
    layer0_outputs(575) <= not((inputs(238)) or (inputs(16)));
    layer0_outputs(576) <= not(inputs(197));
    layer0_outputs(577) <= not((inputs(251)) xor (inputs(187)));
    layer0_outputs(578) <= inputs(174);
    layer0_outputs(579) <= not(inputs(83));
    layer0_outputs(580) <= not((inputs(193)) or (inputs(208)));
    layer0_outputs(581) <= not(inputs(133)) or (inputs(72));
    layer0_outputs(582) <= '1';
    layer0_outputs(583) <= (inputs(238)) or (inputs(245));
    layer0_outputs(584) <= not(inputs(174));
    layer0_outputs(585) <= (inputs(204)) and not (inputs(247));
    layer0_outputs(586) <= not((inputs(153)) or (inputs(220)));
    layer0_outputs(587) <= not((inputs(245)) and (inputs(227)));
    layer0_outputs(588) <= (inputs(78)) and not (inputs(15));
    layer0_outputs(589) <= (inputs(95)) and not (inputs(157));
    layer0_outputs(590) <= not(inputs(14));
    layer0_outputs(591) <= not(inputs(124)) or (inputs(129));
    layer0_outputs(592) <= not((inputs(83)) or (inputs(90)));
    layer0_outputs(593) <= not(inputs(230));
    layer0_outputs(594) <= not((inputs(197)) xor (inputs(65)));
    layer0_outputs(595) <= not(inputs(100));
    layer0_outputs(596) <= not((inputs(223)) xor (inputs(204)));
    layer0_outputs(597) <= (inputs(37)) and (inputs(12));
    layer0_outputs(598) <= inputs(228);
    layer0_outputs(599) <= not(inputs(39));
    layer0_outputs(600) <= (inputs(122)) and not (inputs(141));
    layer0_outputs(601) <= not(inputs(245));
    layer0_outputs(602) <= (inputs(33)) or (inputs(210));
    layer0_outputs(603) <= (inputs(173)) xor (inputs(204));
    layer0_outputs(604) <= (inputs(83)) or (inputs(151));
    layer0_outputs(605) <= inputs(157);
    layer0_outputs(606) <= not(inputs(244));
    layer0_outputs(607) <= '1';
    layer0_outputs(608) <= (inputs(90)) or (inputs(149));
    layer0_outputs(609) <= (inputs(138)) and not (inputs(179));
    layer0_outputs(610) <= not(inputs(251));
    layer0_outputs(611) <= not(inputs(162));
    layer0_outputs(612) <= not(inputs(209));
    layer0_outputs(613) <= not((inputs(177)) and (inputs(188)));
    layer0_outputs(614) <= not(inputs(1));
    layer0_outputs(615) <= inputs(84);
    layer0_outputs(616) <= not(inputs(75)) or (inputs(180));
    layer0_outputs(617) <= inputs(171);
    layer0_outputs(618) <= not((inputs(176)) or (inputs(202)));
    layer0_outputs(619) <= (inputs(248)) and not (inputs(76));
    layer0_outputs(620) <= not(inputs(68));
    layer0_outputs(621) <= inputs(91);
    layer0_outputs(622) <= not(inputs(180));
    layer0_outputs(623) <= not((inputs(154)) or (inputs(179)));
    layer0_outputs(624) <= not(inputs(157));
    layer0_outputs(625) <= inputs(114);
    layer0_outputs(626) <= (inputs(65)) xor (inputs(69));
    layer0_outputs(627) <= inputs(133);
    layer0_outputs(628) <= (inputs(227)) and not (inputs(125));
    layer0_outputs(629) <= '0';
    layer0_outputs(630) <= not((inputs(80)) or (inputs(178)));
    layer0_outputs(631) <= not((inputs(235)) or (inputs(141)));
    layer0_outputs(632) <= not(inputs(138)) or (inputs(196));
    layer0_outputs(633) <= (inputs(121)) and not (inputs(128));
    layer0_outputs(634) <= inputs(70);
    layer0_outputs(635) <= (inputs(130)) xor (inputs(113));
    layer0_outputs(636) <= inputs(217);
    layer0_outputs(637) <= inputs(101);
    layer0_outputs(638) <= not((inputs(193)) or (inputs(225)));
    layer0_outputs(639) <= inputs(253);
    layer0_outputs(640) <= inputs(101);
    layer0_outputs(641) <= not((inputs(224)) or (inputs(1)));
    layer0_outputs(642) <= (inputs(72)) and not (inputs(127));
    layer0_outputs(643) <= not(inputs(147));
    layer0_outputs(644) <= (inputs(123)) or (inputs(32));
    layer0_outputs(645) <= (inputs(16)) xor (inputs(44));
    layer0_outputs(646) <= not((inputs(60)) xor (inputs(71)));
    layer0_outputs(647) <= inputs(102);
    layer0_outputs(648) <= (inputs(204)) and not (inputs(238));
    layer0_outputs(649) <= not((inputs(123)) or (inputs(80)));
    layer0_outputs(650) <= inputs(82);
    layer0_outputs(651) <= (inputs(30)) or (inputs(59));
    layer0_outputs(652) <= not((inputs(203)) or (inputs(97)));
    layer0_outputs(653) <= inputs(98);
    layer0_outputs(654) <= not(inputs(97));
    layer0_outputs(655) <= not(inputs(39));
    layer0_outputs(656) <= (inputs(249)) or (inputs(244));
    layer0_outputs(657) <= not(inputs(13));
    layer0_outputs(658) <= not(inputs(231)) or (inputs(1));
    layer0_outputs(659) <= (inputs(13)) and not (inputs(76));
    layer0_outputs(660) <= (inputs(172)) and not (inputs(168));
    layer0_outputs(661) <= (inputs(215)) and not (inputs(252));
    layer0_outputs(662) <= (inputs(37)) or (inputs(95));
    layer0_outputs(663) <= not((inputs(141)) or (inputs(114)));
    layer0_outputs(664) <= inputs(98);
    layer0_outputs(665) <= (inputs(68)) xor (inputs(48));
    layer0_outputs(666) <= inputs(100);
    layer0_outputs(667) <= not(inputs(14));
    layer0_outputs(668) <= not((inputs(24)) xor (inputs(70)));
    layer0_outputs(669) <= (inputs(229)) and not (inputs(96));
    layer0_outputs(670) <= (inputs(219)) or (inputs(79));
    layer0_outputs(671) <= (inputs(182)) or (inputs(38));
    layer0_outputs(672) <= not(inputs(23)) or (inputs(77));
    layer0_outputs(673) <= not(inputs(103)) or (inputs(57));
    layer0_outputs(674) <= not((inputs(222)) or (inputs(254)));
    layer0_outputs(675) <= not(inputs(240));
    layer0_outputs(676) <= not(inputs(174));
    layer0_outputs(677) <= (inputs(63)) or (inputs(59));
    layer0_outputs(678) <= not((inputs(248)) and (inputs(28)));
    layer0_outputs(679) <= not(inputs(108));
    layer0_outputs(680) <= inputs(163);
    layer0_outputs(681) <= inputs(16);
    layer0_outputs(682) <= not(inputs(23)) or (inputs(212));
    layer0_outputs(683) <= inputs(68);
    layer0_outputs(684) <= not(inputs(21));
    layer0_outputs(685) <= inputs(209);
    layer0_outputs(686) <= (inputs(95)) and not (inputs(231));
    layer0_outputs(687) <= not((inputs(226)) or (inputs(163)));
    layer0_outputs(688) <= inputs(192);
    layer0_outputs(689) <= inputs(115);
    layer0_outputs(690) <= not((inputs(139)) or (inputs(222)));
    layer0_outputs(691) <= (inputs(240)) xor (inputs(74));
    layer0_outputs(692) <= inputs(94);
    layer0_outputs(693) <= inputs(219);
    layer0_outputs(694) <= not((inputs(107)) or (inputs(149)));
    layer0_outputs(695) <= not(inputs(172));
    layer0_outputs(696) <= (inputs(15)) or (inputs(201));
    layer0_outputs(697) <= not(inputs(169));
    layer0_outputs(698) <= not((inputs(194)) or (inputs(239)));
    layer0_outputs(699) <= not((inputs(96)) or (inputs(230)));
    layer0_outputs(700) <= (inputs(147)) xor (inputs(45));
    layer0_outputs(701) <= not(inputs(154));
    layer0_outputs(702) <= inputs(61);
    layer0_outputs(703) <= not((inputs(215)) and (inputs(70)));
    layer0_outputs(704) <= inputs(119);
    layer0_outputs(705) <= not(inputs(114));
    layer0_outputs(706) <= not((inputs(89)) or (inputs(48)));
    layer0_outputs(707) <= not(inputs(85));
    layer0_outputs(708) <= not(inputs(15));
    layer0_outputs(709) <= inputs(83);
    layer0_outputs(710) <= not((inputs(228)) or (inputs(33)));
    layer0_outputs(711) <= not((inputs(205)) or (inputs(202)));
    layer0_outputs(712) <= inputs(101);
    layer0_outputs(713) <= inputs(149);
    layer0_outputs(714) <= inputs(100);
    layer0_outputs(715) <= not((inputs(89)) and (inputs(57)));
    layer0_outputs(716) <= not(inputs(176));
    layer0_outputs(717) <= (inputs(131)) and not (inputs(207));
    layer0_outputs(718) <= inputs(136);
    layer0_outputs(719) <= (inputs(203)) and not (inputs(123));
    layer0_outputs(720) <= not(inputs(246));
    layer0_outputs(721) <= (inputs(186)) and (inputs(225));
    layer0_outputs(722) <= not((inputs(236)) or (inputs(221)));
    layer0_outputs(723) <= not(inputs(209)) or (inputs(33));
    layer0_outputs(724) <= not(inputs(11));
    layer0_outputs(725) <= not((inputs(234)) and (inputs(69)));
    layer0_outputs(726) <= not((inputs(127)) or (inputs(146)));
    layer0_outputs(727) <= not(inputs(179));
    layer0_outputs(728) <= inputs(226);
    layer0_outputs(729) <= not(inputs(49));
    layer0_outputs(730) <= inputs(233);
    layer0_outputs(731) <= not(inputs(203));
    layer0_outputs(732) <= (inputs(189)) and not (inputs(66));
    layer0_outputs(733) <= not(inputs(113));
    layer0_outputs(734) <= inputs(139);
    layer0_outputs(735) <= not((inputs(133)) or (inputs(140)));
    layer0_outputs(736) <= not((inputs(234)) or (inputs(36)));
    layer0_outputs(737) <= (inputs(138)) xor (inputs(58));
    layer0_outputs(738) <= not((inputs(57)) or (inputs(227)));
    layer0_outputs(739) <= inputs(181);
    layer0_outputs(740) <= (inputs(45)) or (inputs(17));
    layer0_outputs(741) <= inputs(204);
    layer0_outputs(742) <= inputs(168);
    layer0_outputs(743) <= inputs(35);
    layer0_outputs(744) <= (inputs(217)) or (inputs(158));
    layer0_outputs(745) <= (inputs(24)) and not (inputs(18));
    layer0_outputs(746) <= inputs(163);
    layer0_outputs(747) <= not(inputs(198)) or (inputs(239));
    layer0_outputs(748) <= (inputs(123)) and (inputs(67));
    layer0_outputs(749) <= not((inputs(137)) or (inputs(94)));
    layer0_outputs(750) <= inputs(104);
    layer0_outputs(751) <= not(inputs(141));
    layer0_outputs(752) <= '0';
    layer0_outputs(753) <= '0';
    layer0_outputs(754) <= (inputs(221)) or (inputs(219));
    layer0_outputs(755) <= (inputs(134)) and not (inputs(252));
    layer0_outputs(756) <= not((inputs(27)) and (inputs(100)));
    layer0_outputs(757) <= inputs(195);
    layer0_outputs(758) <= not((inputs(8)) or (inputs(208)));
    layer0_outputs(759) <= (inputs(106)) or (inputs(179));
    layer0_outputs(760) <= not(inputs(76));
    layer0_outputs(761) <= not(inputs(194));
    layer0_outputs(762) <= inputs(80);
    layer0_outputs(763) <= not((inputs(161)) or (inputs(142)));
    layer0_outputs(764) <= (inputs(131)) and not (inputs(237));
    layer0_outputs(765) <= not(inputs(197));
    layer0_outputs(766) <= not(inputs(123));
    layer0_outputs(767) <= not((inputs(176)) or (inputs(13)));
    layer0_outputs(768) <= not(inputs(230));
    layer0_outputs(769) <= inputs(206);
    layer0_outputs(770) <= not(inputs(39));
    layer0_outputs(771) <= not(inputs(34)) or (inputs(24));
    layer0_outputs(772) <= inputs(117);
    layer0_outputs(773) <= (inputs(102)) or (inputs(81));
    layer0_outputs(774) <= inputs(77);
    layer0_outputs(775) <= (inputs(91)) and not (inputs(2));
    layer0_outputs(776) <= not(inputs(116));
    layer0_outputs(777) <= inputs(218);
    layer0_outputs(778) <= not(inputs(13)) or (inputs(147));
    layer0_outputs(779) <= (inputs(142)) and not (inputs(9));
    layer0_outputs(780) <= (inputs(65)) or (inputs(26));
    layer0_outputs(781) <= not(inputs(232)) or (inputs(26));
    layer0_outputs(782) <= inputs(123);
    layer0_outputs(783) <= not(inputs(149)) or (inputs(241));
    layer0_outputs(784) <= not(inputs(21));
    layer0_outputs(785) <= not(inputs(129)) or (inputs(240));
    layer0_outputs(786) <= not(inputs(162)) or (inputs(170));
    layer0_outputs(787) <= not(inputs(153)) or (inputs(153));
    layer0_outputs(788) <= (inputs(231)) and not (inputs(150));
    layer0_outputs(789) <= inputs(162);
    layer0_outputs(790) <= not(inputs(21));
    layer0_outputs(791) <= not(inputs(218)) or (inputs(130));
    layer0_outputs(792) <= (inputs(138)) and not (inputs(165));
    layer0_outputs(793) <= not(inputs(118));
    layer0_outputs(794) <= not(inputs(97));
    layer0_outputs(795) <= not((inputs(198)) and (inputs(187)));
    layer0_outputs(796) <= not((inputs(81)) or (inputs(10)));
    layer0_outputs(797) <= not((inputs(243)) or (inputs(168)));
    layer0_outputs(798) <= (inputs(160)) and not (inputs(140));
    layer0_outputs(799) <= (inputs(242)) xor (inputs(76));
    layer0_outputs(800) <= (inputs(196)) or (inputs(223));
    layer0_outputs(801) <= not((inputs(69)) or (inputs(150)));
    layer0_outputs(802) <= (inputs(177)) or (inputs(7));
    layer0_outputs(803) <= not(inputs(40));
    layer0_outputs(804) <= inputs(247);
    layer0_outputs(805) <= (inputs(31)) or (inputs(65));
    layer0_outputs(806) <= inputs(218);
    layer0_outputs(807) <= inputs(11);
    layer0_outputs(808) <= not(inputs(203));
    layer0_outputs(809) <= (inputs(189)) and (inputs(141));
    layer0_outputs(810) <= (inputs(210)) or (inputs(246));
    layer0_outputs(811) <= (inputs(189)) and not (inputs(49));
    layer0_outputs(812) <= not(inputs(240)) or (inputs(148));
    layer0_outputs(813) <= not((inputs(165)) xor (inputs(145)));
    layer0_outputs(814) <= (inputs(72)) xor (inputs(96));
    layer0_outputs(815) <= not(inputs(75)) or (inputs(173));
    layer0_outputs(816) <= not((inputs(186)) or (inputs(204)));
    layer0_outputs(817) <= not(inputs(124)) or (inputs(163));
    layer0_outputs(818) <= (inputs(94)) or (inputs(197));
    layer0_outputs(819) <= not(inputs(73));
    layer0_outputs(820) <= not(inputs(135)) or (inputs(198));
    layer0_outputs(821) <= inputs(169);
    layer0_outputs(822) <= not((inputs(181)) or (inputs(195)));
    layer0_outputs(823) <= not((inputs(158)) or (inputs(141)));
    layer0_outputs(824) <= (inputs(160)) xor (inputs(95));
    layer0_outputs(825) <= not(inputs(105));
    layer0_outputs(826) <= not(inputs(115)) or (inputs(0));
    layer0_outputs(827) <= (inputs(41)) and not (inputs(129));
    layer0_outputs(828) <= inputs(157);
    layer0_outputs(829) <= (inputs(90)) or (inputs(77));
    layer0_outputs(830) <= not((inputs(127)) or (inputs(231)));
    layer0_outputs(831) <= (inputs(246)) or (inputs(255));
    layer0_outputs(832) <= not(inputs(173));
    layer0_outputs(833) <= (inputs(116)) or (inputs(220));
    layer0_outputs(834) <= not(inputs(137));
    layer0_outputs(835) <= not(inputs(227));
    layer0_outputs(836) <= (inputs(158)) or (inputs(172));
    layer0_outputs(837) <= '1';
    layer0_outputs(838) <= (inputs(69)) and not (inputs(175));
    layer0_outputs(839) <= (inputs(49)) or (inputs(22));
    layer0_outputs(840) <= not((inputs(22)) or (inputs(177)));
    layer0_outputs(841) <= (inputs(191)) or (inputs(95));
    layer0_outputs(842) <= inputs(198);
    layer0_outputs(843) <= not(inputs(42)) or (inputs(207));
    layer0_outputs(844) <= not((inputs(194)) or (inputs(30)));
    layer0_outputs(845) <= (inputs(187)) and not (inputs(226));
    layer0_outputs(846) <= not((inputs(141)) or (inputs(138)));
    layer0_outputs(847) <= inputs(122);
    layer0_outputs(848) <= not(inputs(24));
    layer0_outputs(849) <= not(inputs(78)) or (inputs(144));
    layer0_outputs(850) <= (inputs(66)) or (inputs(124));
    layer0_outputs(851) <= (inputs(91)) or (inputs(33));
    layer0_outputs(852) <= inputs(116);
    layer0_outputs(853) <= not((inputs(25)) and (inputs(168)));
    layer0_outputs(854) <= not(inputs(73));
    layer0_outputs(855) <= not(inputs(24)) or (inputs(167));
    layer0_outputs(856) <= (inputs(103)) or (inputs(147));
    layer0_outputs(857) <= (inputs(101)) xor (inputs(148));
    layer0_outputs(858) <= (inputs(161)) xor (inputs(60));
    layer0_outputs(859) <= not(inputs(13));
    layer0_outputs(860) <= inputs(166);
    layer0_outputs(861) <= not((inputs(159)) or (inputs(46)));
    layer0_outputs(862) <= not(inputs(75)) or (inputs(18));
    layer0_outputs(863) <= (inputs(2)) or (inputs(62));
    layer0_outputs(864) <= not(inputs(105)) or (inputs(157));
    layer0_outputs(865) <= (inputs(170)) or (inputs(147));
    layer0_outputs(866) <= not((inputs(135)) or (inputs(234)));
    layer0_outputs(867) <= (inputs(54)) or (inputs(206));
    layer0_outputs(868) <= not(inputs(149));
    layer0_outputs(869) <= not((inputs(86)) or (inputs(172)));
    layer0_outputs(870) <= not(inputs(64));
    layer0_outputs(871) <= (inputs(5)) and not (inputs(112));
    layer0_outputs(872) <= not(inputs(55));
    layer0_outputs(873) <= inputs(40);
    layer0_outputs(874) <= (inputs(197)) or (inputs(193));
    layer0_outputs(875) <= inputs(90);
    layer0_outputs(876) <= not((inputs(187)) or (inputs(152)));
    layer0_outputs(877) <= not((inputs(10)) or (inputs(176)));
    layer0_outputs(878) <= not(inputs(69)) or (inputs(116));
    layer0_outputs(879) <= inputs(193);
    layer0_outputs(880) <= (inputs(57)) and not (inputs(56));
    layer0_outputs(881) <= inputs(142);
    layer0_outputs(882) <= (inputs(132)) or (inputs(208));
    layer0_outputs(883) <= inputs(136);
    layer0_outputs(884) <= (inputs(188)) or (inputs(171));
    layer0_outputs(885) <= (inputs(167)) or (inputs(58));
    layer0_outputs(886) <= (inputs(5)) and not (inputs(159));
    layer0_outputs(887) <= not(inputs(85)) or (inputs(176));
    layer0_outputs(888) <= (inputs(95)) or (inputs(138));
    layer0_outputs(889) <= not(inputs(17));
    layer0_outputs(890) <= not(inputs(11)) or (inputs(25));
    layer0_outputs(891) <= not(inputs(104)) or (inputs(15));
    layer0_outputs(892) <= (inputs(182)) or (inputs(165));
    layer0_outputs(893) <= not(inputs(101)) or (inputs(2));
    layer0_outputs(894) <= (inputs(115)) and not (inputs(126));
    layer0_outputs(895) <= inputs(17);
    layer0_outputs(896) <= (inputs(101)) and not (inputs(207));
    layer0_outputs(897) <= (inputs(85)) and not (inputs(205));
    layer0_outputs(898) <= not(inputs(164)) or (inputs(98));
    layer0_outputs(899) <= not(inputs(104)) or (inputs(126));
    layer0_outputs(900) <= (inputs(31)) and (inputs(223));
    layer0_outputs(901) <= inputs(28);
    layer0_outputs(902) <= not(inputs(57)) or (inputs(8));
    layer0_outputs(903) <= (inputs(247)) and (inputs(164));
    layer0_outputs(904) <= inputs(101);
    layer0_outputs(905) <= (inputs(36)) and (inputs(25));
    layer0_outputs(906) <= inputs(179);
    layer0_outputs(907) <= inputs(171);
    layer0_outputs(908) <= not(inputs(125));
    layer0_outputs(909) <= inputs(50);
    layer0_outputs(910) <= (inputs(159)) or (inputs(72));
    layer0_outputs(911) <= (inputs(66)) and not (inputs(195));
    layer0_outputs(912) <= (inputs(159)) or (inputs(87));
    layer0_outputs(913) <= (inputs(132)) or (inputs(18));
    layer0_outputs(914) <= inputs(231);
    layer0_outputs(915) <= (inputs(112)) or (inputs(141));
    layer0_outputs(916) <= inputs(9);
    layer0_outputs(917) <= inputs(235);
    layer0_outputs(918) <= not((inputs(186)) or (inputs(47)));
    layer0_outputs(919) <= not(inputs(233));
    layer0_outputs(920) <= (inputs(132)) and not (inputs(48));
    layer0_outputs(921) <= inputs(116);
    layer0_outputs(922) <= not(inputs(183));
    layer0_outputs(923) <= inputs(117);
    layer0_outputs(924) <= (inputs(89)) and not (inputs(110));
    layer0_outputs(925) <= (inputs(171)) or (inputs(108));
    layer0_outputs(926) <= not((inputs(217)) or (inputs(250)));
    layer0_outputs(927) <= not((inputs(184)) and (inputs(202)));
    layer0_outputs(928) <= (inputs(82)) and not (inputs(132));
    layer0_outputs(929) <= inputs(71);
    layer0_outputs(930) <= inputs(228);
    layer0_outputs(931) <= (inputs(221)) or (inputs(120));
    layer0_outputs(932) <= not(inputs(8));
    layer0_outputs(933) <= (inputs(175)) xor (inputs(203));
    layer0_outputs(934) <= (inputs(253)) xor (inputs(85));
    layer0_outputs(935) <= not((inputs(195)) or (inputs(19)));
    layer0_outputs(936) <= (inputs(32)) or (inputs(138));
    layer0_outputs(937) <= not((inputs(74)) or (inputs(75)));
    layer0_outputs(938) <= (inputs(4)) and not (inputs(234));
    layer0_outputs(939) <= not((inputs(224)) or (inputs(212)));
    layer0_outputs(940) <= (inputs(124)) xor (inputs(34));
    layer0_outputs(941) <= not(inputs(167));
    layer0_outputs(942) <= inputs(239);
    layer0_outputs(943) <= not(inputs(206));
    layer0_outputs(944) <= not(inputs(153)) or (inputs(205));
    layer0_outputs(945) <= inputs(122);
    layer0_outputs(946) <= not(inputs(19));
    layer0_outputs(947) <= (inputs(97)) and not (inputs(63));
    layer0_outputs(948) <= (inputs(64)) or (inputs(196));
    layer0_outputs(949) <= not(inputs(199)) or (inputs(29));
    layer0_outputs(950) <= inputs(216);
    layer0_outputs(951) <= not((inputs(14)) and (inputs(77)));
    layer0_outputs(952) <= not((inputs(81)) xor (inputs(53)));
    layer0_outputs(953) <= inputs(158);
    layer0_outputs(954) <= not((inputs(127)) or (inputs(74)));
    layer0_outputs(955) <= (inputs(171)) and (inputs(89));
    layer0_outputs(956) <= not(inputs(228));
    layer0_outputs(957) <= '0';
    layer0_outputs(958) <= (inputs(161)) or (inputs(187));
    layer0_outputs(959) <= (inputs(136)) and not (inputs(205));
    layer0_outputs(960) <= not((inputs(122)) or (inputs(33)));
    layer0_outputs(961) <= (inputs(6)) and not (inputs(3));
    layer0_outputs(962) <= (inputs(171)) xor (inputs(90));
    layer0_outputs(963) <= not((inputs(154)) or (inputs(80)));
    layer0_outputs(964) <= not((inputs(133)) or (inputs(110)));
    layer0_outputs(965) <= not(inputs(167));
    layer0_outputs(966) <= (inputs(30)) or (inputs(217));
    layer0_outputs(967) <= not(inputs(153));
    layer0_outputs(968) <= not(inputs(195));
    layer0_outputs(969) <= not(inputs(229)) or (inputs(68));
    layer0_outputs(970) <= not(inputs(25));
    layer0_outputs(971) <= '1';
    layer0_outputs(972) <= not(inputs(253));
    layer0_outputs(973) <= (inputs(67)) and (inputs(67));
    layer0_outputs(974) <= (inputs(167)) and not (inputs(203));
    layer0_outputs(975) <= (inputs(167)) and not (inputs(225));
    layer0_outputs(976) <= (inputs(89)) and not (inputs(117));
    layer0_outputs(977) <= inputs(234);
    layer0_outputs(978) <= not((inputs(201)) or (inputs(222)));
    layer0_outputs(979) <= (inputs(33)) or (inputs(69));
    layer0_outputs(980) <= inputs(167);
    layer0_outputs(981) <= (inputs(5)) and not (inputs(185));
    layer0_outputs(982) <= not(inputs(69));
    layer0_outputs(983) <= (inputs(155)) xor (inputs(139));
    layer0_outputs(984) <= not((inputs(20)) or (inputs(164)));
    layer0_outputs(985) <= not(inputs(158)) or (inputs(113));
    layer0_outputs(986) <= (inputs(58)) xor (inputs(61));
    layer0_outputs(987) <= not(inputs(191));
    layer0_outputs(988) <= not((inputs(16)) or (inputs(19)));
    layer0_outputs(989) <= inputs(120);
    layer0_outputs(990) <= not((inputs(157)) xor (inputs(124)));
    layer0_outputs(991) <= not((inputs(157)) or (inputs(141)));
    layer0_outputs(992) <= inputs(183);
    layer0_outputs(993) <= not(inputs(217));
    layer0_outputs(994) <= not(inputs(151));
    layer0_outputs(995) <= inputs(97);
    layer0_outputs(996) <= inputs(112);
    layer0_outputs(997) <= (inputs(64)) xor (inputs(129));
    layer0_outputs(998) <= not(inputs(68)) or (inputs(191));
    layer0_outputs(999) <= not(inputs(247));
    layer0_outputs(1000) <= (inputs(199)) xor (inputs(254));
    layer0_outputs(1001) <= (inputs(79)) xor (inputs(172));
    layer0_outputs(1002) <= not((inputs(126)) or (inputs(196)));
    layer0_outputs(1003) <= (inputs(121)) and not (inputs(191));
    layer0_outputs(1004) <= (inputs(119)) and not (inputs(66));
    layer0_outputs(1005) <= inputs(150);
    layer0_outputs(1006) <= (inputs(251)) or (inputs(94));
    layer0_outputs(1007) <= not((inputs(219)) or (inputs(144)));
    layer0_outputs(1008) <= (inputs(183)) or (inputs(136));
    layer0_outputs(1009) <= not((inputs(65)) xor (inputs(93)));
    layer0_outputs(1010) <= inputs(118);
    layer0_outputs(1011) <= inputs(228);
    layer0_outputs(1012) <= (inputs(141)) and not (inputs(33));
    layer0_outputs(1013) <= (inputs(86)) or (inputs(205));
    layer0_outputs(1014) <= not(inputs(210));
    layer0_outputs(1015) <= not(inputs(190)) or (inputs(72));
    layer0_outputs(1016) <= inputs(100);
    layer0_outputs(1017) <= inputs(162);
    layer0_outputs(1018) <= inputs(145);
    layer0_outputs(1019) <= inputs(98);
    layer0_outputs(1020) <= not(inputs(236));
    layer0_outputs(1021) <= not(inputs(57)) or (inputs(145));
    layer0_outputs(1022) <= not((inputs(131)) or (inputs(159)));
    layer0_outputs(1023) <= inputs(111);
    layer0_outputs(1024) <= not(inputs(164));
    layer0_outputs(1025) <= inputs(221);
    layer0_outputs(1026) <= inputs(107);
    layer0_outputs(1027) <= not(inputs(81));
    layer0_outputs(1028) <= (inputs(196)) and not (inputs(112));
    layer0_outputs(1029) <= not((inputs(50)) or (inputs(67)));
    layer0_outputs(1030) <= (inputs(129)) or (inputs(113));
    layer0_outputs(1031) <= (inputs(62)) or (inputs(16));
    layer0_outputs(1032) <= inputs(231);
    layer0_outputs(1033) <= (inputs(102)) and not (inputs(49));
    layer0_outputs(1034) <= (inputs(207)) or (inputs(12));
    layer0_outputs(1035) <= (inputs(214)) or (inputs(15));
    layer0_outputs(1036) <= not((inputs(90)) or (inputs(17)));
    layer0_outputs(1037) <= (inputs(158)) or (inputs(172));
    layer0_outputs(1038) <= not(inputs(15));
    layer0_outputs(1039) <= (inputs(172)) xor (inputs(101));
    layer0_outputs(1040) <= not(inputs(39)) or (inputs(63));
    layer0_outputs(1041) <= inputs(137);
    layer0_outputs(1042) <= not(inputs(75));
    layer0_outputs(1043) <= (inputs(181)) xor (inputs(255));
    layer0_outputs(1044) <= inputs(213);
    layer0_outputs(1045) <= inputs(10);
    layer0_outputs(1046) <= not(inputs(199)) or (inputs(224));
    layer0_outputs(1047) <= inputs(68);
    layer0_outputs(1048) <= (inputs(83)) or (inputs(233));
    layer0_outputs(1049) <= not(inputs(25)) or (inputs(164));
    layer0_outputs(1050) <= not(inputs(168));
    layer0_outputs(1051) <= (inputs(85)) or (inputs(62));
    layer0_outputs(1052) <= inputs(23);
    layer0_outputs(1053) <= not((inputs(161)) or (inputs(203)));
    layer0_outputs(1054) <= (inputs(35)) or (inputs(17));
    layer0_outputs(1055) <= not(inputs(28));
    layer0_outputs(1056) <= (inputs(86)) xor (inputs(2));
    layer0_outputs(1057) <= not((inputs(100)) or (inputs(97)));
    layer0_outputs(1058) <= not(inputs(117)) or (inputs(155));
    layer0_outputs(1059) <= inputs(178);
    layer0_outputs(1060) <= not((inputs(148)) or (inputs(144)));
    layer0_outputs(1061) <= not(inputs(25));
    layer0_outputs(1062) <= (inputs(71)) and not (inputs(137));
    layer0_outputs(1063) <= (inputs(55)) and not (inputs(19));
    layer0_outputs(1064) <= (inputs(33)) and not (inputs(237));
    layer0_outputs(1065) <= not(inputs(46));
    layer0_outputs(1066) <= not((inputs(212)) or (inputs(70)));
    layer0_outputs(1067) <= (inputs(37)) and not (inputs(129));
    layer0_outputs(1068) <= not(inputs(190));
    layer0_outputs(1069) <= not(inputs(84)) or (inputs(163));
    layer0_outputs(1070) <= inputs(107);
    layer0_outputs(1071) <= not((inputs(16)) or (inputs(23)));
    layer0_outputs(1072) <= not((inputs(222)) or (inputs(103)));
    layer0_outputs(1073) <= inputs(245);
    layer0_outputs(1074) <= (inputs(4)) or (inputs(106));
    layer0_outputs(1075) <= inputs(32);
    layer0_outputs(1076) <= (inputs(236)) and not (inputs(39));
    layer0_outputs(1077) <= inputs(255);
    layer0_outputs(1078) <= inputs(116);
    layer0_outputs(1079) <= (inputs(56)) and not (inputs(6));
    layer0_outputs(1080) <= not(inputs(82));
    layer0_outputs(1081) <= inputs(86);
    layer0_outputs(1082) <= not(inputs(159));
    layer0_outputs(1083) <= not(inputs(69)) or (inputs(156));
    layer0_outputs(1084) <= (inputs(174)) xor (inputs(21));
    layer0_outputs(1085) <= not(inputs(135));
    layer0_outputs(1086) <= not(inputs(183));
    layer0_outputs(1087) <= (inputs(80)) or (inputs(181));
    layer0_outputs(1088) <= (inputs(165)) or (inputs(17));
    layer0_outputs(1089) <= (inputs(2)) or (inputs(168));
    layer0_outputs(1090) <= not(inputs(20));
    layer0_outputs(1091) <= not((inputs(74)) or (inputs(225)));
    layer0_outputs(1092) <= not(inputs(121));
    layer0_outputs(1093) <= (inputs(165)) xor (inputs(147));
    layer0_outputs(1094) <= not(inputs(99));
    layer0_outputs(1095) <= inputs(54);
    layer0_outputs(1096) <= inputs(23);
    layer0_outputs(1097) <= not(inputs(105));
    layer0_outputs(1098) <= inputs(244);
    layer0_outputs(1099) <= not((inputs(130)) or (inputs(161)));
    layer0_outputs(1100) <= not((inputs(230)) or (inputs(235)));
    layer0_outputs(1101) <= inputs(107);
    layer0_outputs(1102) <= (inputs(176)) or (inputs(75));
    layer0_outputs(1103) <= inputs(145);
    layer0_outputs(1104) <= not(inputs(144));
    layer0_outputs(1105) <= inputs(233);
    layer0_outputs(1106) <= inputs(151);
    layer0_outputs(1107) <= (inputs(116)) or (inputs(109));
    layer0_outputs(1108) <= not((inputs(128)) or (inputs(116)));
    layer0_outputs(1109) <= '1';
    layer0_outputs(1110) <= inputs(50);
    layer0_outputs(1111) <= (inputs(74)) xor (inputs(13));
    layer0_outputs(1112) <= not((inputs(66)) or (inputs(237)));
    layer0_outputs(1113) <= inputs(212);
    layer0_outputs(1114) <= '1';
    layer0_outputs(1115) <= not(inputs(247));
    layer0_outputs(1116) <= not(inputs(215));
    layer0_outputs(1117) <= not(inputs(205));
    layer0_outputs(1118) <= inputs(193);
    layer0_outputs(1119) <= (inputs(220)) and (inputs(215));
    layer0_outputs(1120) <= not(inputs(37));
    layer0_outputs(1121) <= (inputs(253)) and not (inputs(80));
    layer0_outputs(1122) <= not((inputs(167)) xor (inputs(100)));
    layer0_outputs(1123) <= inputs(179);
    layer0_outputs(1124) <= not(inputs(9)) or (inputs(169));
    layer0_outputs(1125) <= (inputs(101)) and not (inputs(251));
    layer0_outputs(1126) <= inputs(153);
    layer0_outputs(1127) <= not(inputs(122)) or (inputs(237));
    layer0_outputs(1128) <= not(inputs(232));
    layer0_outputs(1129) <= not(inputs(62));
    layer0_outputs(1130) <= (inputs(66)) and not (inputs(38));
    layer0_outputs(1131) <= inputs(6);
    layer0_outputs(1132) <= (inputs(246)) or (inputs(161));
    layer0_outputs(1133) <= not((inputs(79)) or (inputs(97)));
    layer0_outputs(1134) <= (inputs(58)) or (inputs(92));
    layer0_outputs(1135) <= (inputs(169)) xor (inputs(242));
    layer0_outputs(1136) <= inputs(40);
    layer0_outputs(1137) <= not((inputs(216)) and (inputs(244)));
    layer0_outputs(1138) <= (inputs(79)) or (inputs(156));
    layer0_outputs(1139) <= not(inputs(119)) or (inputs(83));
    layer0_outputs(1140) <= '0';
    layer0_outputs(1141) <= not(inputs(163));
    layer0_outputs(1142) <= inputs(100);
    layer0_outputs(1143) <= not(inputs(114));
    layer0_outputs(1144) <= not((inputs(210)) or (inputs(203)));
    layer0_outputs(1145) <= (inputs(96)) and not (inputs(1));
    layer0_outputs(1146) <= not(inputs(11)) or (inputs(240));
    layer0_outputs(1147) <= (inputs(108)) or (inputs(41));
    layer0_outputs(1148) <= (inputs(200)) or (inputs(3));
    layer0_outputs(1149) <= inputs(223);
    layer0_outputs(1150) <= not(inputs(68));
    layer0_outputs(1151) <= not(inputs(136));
    layer0_outputs(1152) <= not(inputs(114));
    layer0_outputs(1153) <= not((inputs(77)) or (inputs(18)));
    layer0_outputs(1154) <= not(inputs(65));
    layer0_outputs(1155) <= not(inputs(230));
    layer0_outputs(1156) <= (inputs(201)) or (inputs(48));
    layer0_outputs(1157) <= not((inputs(229)) or (inputs(32)));
    layer0_outputs(1158) <= inputs(167);
    layer0_outputs(1159) <= not(inputs(152));
    layer0_outputs(1160) <= inputs(8);
    layer0_outputs(1161) <= not(inputs(221)) or (inputs(82));
    layer0_outputs(1162) <= not(inputs(227));
    layer0_outputs(1163) <= not((inputs(220)) and (inputs(105)));
    layer0_outputs(1164) <= not(inputs(8));
    layer0_outputs(1165) <= inputs(46);
    layer0_outputs(1166) <= not((inputs(92)) or (inputs(177)));
    layer0_outputs(1167) <= not(inputs(38)) or (inputs(219));
    layer0_outputs(1168) <= not((inputs(19)) or (inputs(241)));
    layer0_outputs(1169) <= not(inputs(130));
    layer0_outputs(1170) <= (inputs(201)) or (inputs(192));
    layer0_outputs(1171) <= inputs(60);
    layer0_outputs(1172) <= (inputs(46)) or (inputs(13));
    layer0_outputs(1173) <= (inputs(70)) and not (inputs(79));
    layer0_outputs(1174) <= not(inputs(146));
    layer0_outputs(1175) <= (inputs(54)) and not (inputs(77));
    layer0_outputs(1176) <= not((inputs(98)) or (inputs(91)));
    layer0_outputs(1177) <= not(inputs(134)) or (inputs(159));
    layer0_outputs(1178) <= not((inputs(19)) or (inputs(211)));
    layer0_outputs(1179) <= not(inputs(105)) or (inputs(55));
    layer0_outputs(1180) <= not((inputs(87)) and (inputs(65)));
    layer0_outputs(1181) <= not(inputs(43));
    layer0_outputs(1182) <= not((inputs(193)) or (inputs(217)));
    layer0_outputs(1183) <= not(inputs(79)) or (inputs(244));
    layer0_outputs(1184) <= not((inputs(250)) xor (inputs(219)));
    layer0_outputs(1185) <= not(inputs(120));
    layer0_outputs(1186) <= (inputs(239)) or (inputs(137));
    layer0_outputs(1187) <= not((inputs(66)) and (inputs(218)));
    layer0_outputs(1188) <= not(inputs(55));
    layer0_outputs(1189) <= (inputs(245)) or (inputs(142));
    layer0_outputs(1190) <= (inputs(203)) and not (inputs(255));
    layer0_outputs(1191) <= (inputs(143)) or (inputs(190));
    layer0_outputs(1192) <= (inputs(57)) and not (inputs(18));
    layer0_outputs(1193) <= not((inputs(190)) or (inputs(6)));
    layer0_outputs(1194) <= (inputs(73)) and (inputs(40));
    layer0_outputs(1195) <= not(inputs(188));
    layer0_outputs(1196) <= inputs(161);
    layer0_outputs(1197) <= (inputs(73)) xor (inputs(61));
    layer0_outputs(1198) <= (inputs(74)) and not (inputs(34));
    layer0_outputs(1199) <= (inputs(148)) and not (inputs(191));
    layer0_outputs(1200) <= not(inputs(134)) or (inputs(207));
    layer0_outputs(1201) <= inputs(169);
    layer0_outputs(1202) <= not(inputs(73));
    layer0_outputs(1203) <= inputs(105);
    layer0_outputs(1204) <= (inputs(55)) or (inputs(142));
    layer0_outputs(1205) <= inputs(150);
    layer0_outputs(1206) <= not(inputs(169)) or (inputs(224));
    layer0_outputs(1207) <= (inputs(21)) or (inputs(127));
    layer0_outputs(1208) <= inputs(110);
    layer0_outputs(1209) <= not(inputs(237));
    layer0_outputs(1210) <= (inputs(21)) or (inputs(1));
    layer0_outputs(1211) <= not((inputs(46)) or (inputs(255)));
    layer0_outputs(1212) <= not((inputs(71)) xor (inputs(59)));
    layer0_outputs(1213) <= not((inputs(125)) or (inputs(126)));
    layer0_outputs(1214) <= inputs(18);
    layer0_outputs(1215) <= inputs(70);
    layer0_outputs(1216) <= not(inputs(174));
    layer0_outputs(1217) <= not(inputs(56));
    layer0_outputs(1218) <= (inputs(38)) and not (inputs(128));
    layer0_outputs(1219) <= not((inputs(58)) and (inputs(28)));
    layer0_outputs(1220) <= (inputs(93)) or (inputs(153));
    layer0_outputs(1221) <= inputs(173);
    layer0_outputs(1222) <= inputs(106);
    layer0_outputs(1223) <= not(inputs(145));
    layer0_outputs(1224) <= not((inputs(128)) or (inputs(80)));
    layer0_outputs(1225) <= not((inputs(84)) or (inputs(68)));
    layer0_outputs(1226) <= (inputs(24)) and not (inputs(160));
    layer0_outputs(1227) <= not(inputs(76)) or (inputs(31));
    layer0_outputs(1228) <= (inputs(190)) or (inputs(118));
    layer0_outputs(1229) <= not(inputs(175));
    layer0_outputs(1230) <= not(inputs(113));
    layer0_outputs(1231) <= inputs(231);
    layer0_outputs(1232) <= not(inputs(205));
    layer0_outputs(1233) <= not(inputs(233)) or (inputs(50));
    layer0_outputs(1234) <= not(inputs(43)) or (inputs(34));
    layer0_outputs(1235) <= inputs(168);
    layer0_outputs(1236) <= (inputs(201)) and not (inputs(86));
    layer0_outputs(1237) <= (inputs(192)) xor (inputs(178));
    layer0_outputs(1238) <= not((inputs(103)) or (inputs(68)));
    layer0_outputs(1239) <= inputs(102);
    layer0_outputs(1240) <= (inputs(149)) and (inputs(117));
    layer0_outputs(1241) <= (inputs(45)) and not (inputs(21));
    layer0_outputs(1242) <= (inputs(206)) or (inputs(39));
    layer0_outputs(1243) <= not(inputs(135));
    layer0_outputs(1244) <= not((inputs(188)) or (inputs(186)));
    layer0_outputs(1245) <= not(inputs(211));
    layer0_outputs(1246) <= (inputs(149)) and (inputs(196));
    layer0_outputs(1247) <= inputs(15);
    layer0_outputs(1248) <= not((inputs(195)) or (inputs(218)));
    layer0_outputs(1249) <= inputs(233);
    layer0_outputs(1250) <= not(inputs(210)) or (inputs(132));
    layer0_outputs(1251) <= not(inputs(25));
    layer0_outputs(1252) <= not(inputs(152));
    layer0_outputs(1253) <= (inputs(25)) and not (inputs(20));
    layer0_outputs(1254) <= (inputs(11)) and not (inputs(87));
    layer0_outputs(1255) <= not(inputs(38));
    layer0_outputs(1256) <= not(inputs(228));
    layer0_outputs(1257) <= (inputs(162)) xor (inputs(197));
    layer0_outputs(1258) <= not(inputs(73)) or (inputs(49));
    layer0_outputs(1259) <= inputs(90);
    layer0_outputs(1260) <= not(inputs(179));
    layer0_outputs(1261) <= not(inputs(77));
    layer0_outputs(1262) <= not((inputs(53)) or (inputs(174)));
    layer0_outputs(1263) <= not((inputs(161)) or (inputs(222)));
    layer0_outputs(1264) <= inputs(112);
    layer0_outputs(1265) <= (inputs(239)) xor (inputs(104));
    layer0_outputs(1266) <= inputs(225);
    layer0_outputs(1267) <= not(inputs(90)) or (inputs(112));
    layer0_outputs(1268) <= (inputs(137)) and not (inputs(55));
    layer0_outputs(1269) <= inputs(165);
    layer0_outputs(1270) <= inputs(162);
    layer0_outputs(1271) <= inputs(126);
    layer0_outputs(1272) <= (inputs(66)) and (inputs(20));
    layer0_outputs(1273) <= (inputs(115)) xor (inputs(113));
    layer0_outputs(1274) <= not((inputs(123)) or (inputs(145)));
    layer0_outputs(1275) <= (inputs(41)) or (inputs(160));
    layer0_outputs(1276) <= (inputs(115)) and not (inputs(209));
    layer0_outputs(1277) <= inputs(51);
    layer0_outputs(1278) <= (inputs(185)) or (inputs(127));
    layer0_outputs(1279) <= not((inputs(23)) xor (inputs(81)));
    layer0_outputs(1280) <= not(inputs(222));
    layer0_outputs(1281) <= not((inputs(140)) and (inputs(192)));
    layer0_outputs(1282) <= (inputs(96)) or (inputs(148));
    layer0_outputs(1283) <= not((inputs(238)) or (inputs(192)));
    layer0_outputs(1284) <= inputs(211);
    layer0_outputs(1285) <= not((inputs(46)) xor (inputs(244)));
    layer0_outputs(1286) <= inputs(141);
    layer0_outputs(1287) <= not(inputs(130));
    layer0_outputs(1288) <= (inputs(15)) or (inputs(37));
    layer0_outputs(1289) <= not(inputs(219)) or (inputs(93));
    layer0_outputs(1290) <= (inputs(120)) and not (inputs(220));
    layer0_outputs(1291) <= not(inputs(109)) or (inputs(252));
    layer0_outputs(1292) <= (inputs(215)) and not (inputs(4));
    layer0_outputs(1293) <= not(inputs(201)) or (inputs(159));
    layer0_outputs(1294) <= (inputs(106)) or (inputs(191));
    layer0_outputs(1295) <= not(inputs(133));
    layer0_outputs(1296) <= not(inputs(46));
    layer0_outputs(1297) <= not(inputs(178));
    layer0_outputs(1298) <= not(inputs(132));
    layer0_outputs(1299) <= not((inputs(71)) xor (inputs(97)));
    layer0_outputs(1300) <= (inputs(195)) xor (inputs(233));
    layer0_outputs(1301) <= not(inputs(22));
    layer0_outputs(1302) <= inputs(230);
    layer0_outputs(1303) <= not((inputs(119)) or (inputs(132)));
    layer0_outputs(1304) <= inputs(140);
    layer0_outputs(1305) <= not(inputs(52));
    layer0_outputs(1306) <= not((inputs(200)) or (inputs(143)));
    layer0_outputs(1307) <= (inputs(239)) and (inputs(78));
    layer0_outputs(1308) <= inputs(100);
    layer0_outputs(1309) <= not(inputs(185)) or (inputs(54));
    layer0_outputs(1310) <= (inputs(173)) or (inputs(93));
    layer0_outputs(1311) <= not(inputs(42));
    layer0_outputs(1312) <= not(inputs(93)) or (inputs(245));
    layer0_outputs(1313) <= not(inputs(220)) or (inputs(238));
    layer0_outputs(1314) <= inputs(139);
    layer0_outputs(1315) <= not(inputs(67)) or (inputs(224));
    layer0_outputs(1316) <= not((inputs(242)) or (inputs(11)));
    layer0_outputs(1317) <= (inputs(190)) or (inputs(197));
    layer0_outputs(1318) <= inputs(210);
    layer0_outputs(1319) <= (inputs(29)) and not (inputs(155));
    layer0_outputs(1320) <= not((inputs(125)) or (inputs(172)));
    layer0_outputs(1321) <= not((inputs(244)) or (inputs(234)));
    layer0_outputs(1322) <= not(inputs(232));
    layer0_outputs(1323) <= inputs(115);
    layer0_outputs(1324) <= inputs(22);
    layer0_outputs(1325) <= not(inputs(94)) or (inputs(176));
    layer0_outputs(1326) <= '0';
    layer0_outputs(1327) <= (inputs(51)) or (inputs(49));
    layer0_outputs(1328) <= (inputs(186)) or (inputs(204));
    layer0_outputs(1329) <= (inputs(206)) or (inputs(154));
    layer0_outputs(1330) <= not(inputs(217));
    layer0_outputs(1331) <= not(inputs(68));
    layer0_outputs(1332) <= not(inputs(171));
    layer0_outputs(1333) <= not(inputs(167));
    layer0_outputs(1334) <= (inputs(250)) and (inputs(220));
    layer0_outputs(1335) <= (inputs(59)) or (inputs(92));
    layer0_outputs(1336) <= (inputs(132)) or (inputs(27));
    layer0_outputs(1337) <= (inputs(197)) and not (inputs(50));
    layer0_outputs(1338) <= inputs(83);
    layer0_outputs(1339) <= (inputs(66)) or (inputs(54));
    layer0_outputs(1340) <= not(inputs(141));
    layer0_outputs(1341) <= inputs(190);
    layer0_outputs(1342) <= not((inputs(37)) or (inputs(94)));
    layer0_outputs(1343) <= not((inputs(23)) and (inputs(180)));
    layer0_outputs(1344) <= (inputs(143)) or (inputs(231));
    layer0_outputs(1345) <= not(inputs(90)) or (inputs(53));
    layer0_outputs(1346) <= not(inputs(105));
    layer0_outputs(1347) <= not(inputs(113));
    layer0_outputs(1348) <= not(inputs(74)) or (inputs(160));
    layer0_outputs(1349) <= not((inputs(115)) or (inputs(34)));
    layer0_outputs(1350) <= not(inputs(161));
    layer0_outputs(1351) <= inputs(132);
    layer0_outputs(1352) <= (inputs(127)) and (inputs(155));
    layer0_outputs(1353) <= not(inputs(243)) or (inputs(208));
    layer0_outputs(1354) <= (inputs(249)) or (inputs(160));
    layer0_outputs(1355) <= not(inputs(122)) or (inputs(111));
    layer0_outputs(1356) <= not(inputs(43));
    layer0_outputs(1357) <= (inputs(202)) or (inputs(72));
    layer0_outputs(1358) <= (inputs(135)) or (inputs(252));
    layer0_outputs(1359) <= not(inputs(102));
    layer0_outputs(1360) <= not(inputs(119));
    layer0_outputs(1361) <= (inputs(11)) and not (inputs(175));
    layer0_outputs(1362) <= (inputs(51)) and not (inputs(205));
    layer0_outputs(1363) <= (inputs(0)) xor (inputs(192));
    layer0_outputs(1364) <= not(inputs(193));
    layer0_outputs(1365) <= inputs(44);
    layer0_outputs(1366) <= not(inputs(228));
    layer0_outputs(1367) <= not(inputs(110));
    layer0_outputs(1368) <= (inputs(209)) or (inputs(54));
    layer0_outputs(1369) <= not((inputs(158)) or (inputs(202)));
    layer0_outputs(1370) <= inputs(106);
    layer0_outputs(1371) <= (inputs(42)) or (inputs(96));
    layer0_outputs(1372) <= (inputs(64)) or (inputs(186));
    layer0_outputs(1373) <= not((inputs(239)) or (inputs(103)));
    layer0_outputs(1374) <= inputs(46);
    layer0_outputs(1375) <= inputs(238);
    layer0_outputs(1376) <= (inputs(183)) and not (inputs(156));
    layer0_outputs(1377) <= (inputs(21)) or (inputs(198));
    layer0_outputs(1378) <= not((inputs(16)) or (inputs(146)));
    layer0_outputs(1379) <= (inputs(222)) or (inputs(134));
    layer0_outputs(1380) <= (inputs(67)) and (inputs(54));
    layer0_outputs(1381) <= (inputs(114)) or (inputs(69));
    layer0_outputs(1382) <= (inputs(49)) or (inputs(188));
    layer0_outputs(1383) <= not((inputs(215)) and (inputs(59)));
    layer0_outputs(1384) <= '0';
    layer0_outputs(1385) <= (inputs(16)) or (inputs(155));
    layer0_outputs(1386) <= (inputs(135)) and not (inputs(196));
    layer0_outputs(1387) <= inputs(245);
    layer0_outputs(1388) <= (inputs(30)) or (inputs(248));
    layer0_outputs(1389) <= not(inputs(212)) or (inputs(134));
    layer0_outputs(1390) <= inputs(18);
    layer0_outputs(1391) <= (inputs(214)) and not (inputs(225));
    layer0_outputs(1392) <= (inputs(165)) and not (inputs(48));
    layer0_outputs(1393) <= inputs(183);
    layer0_outputs(1394) <= not((inputs(140)) or (inputs(171)));
    layer0_outputs(1395) <= not(inputs(31));
    layer0_outputs(1396) <= inputs(166);
    layer0_outputs(1397) <= '0';
    layer0_outputs(1398) <= inputs(178);
    layer0_outputs(1399) <= (inputs(181)) and not (inputs(182));
    layer0_outputs(1400) <= inputs(91);
    layer0_outputs(1401) <= not((inputs(208)) or (inputs(191)));
    layer0_outputs(1402) <= not(inputs(165));
    layer0_outputs(1403) <= not((inputs(85)) and (inputs(60)));
    layer0_outputs(1404) <= inputs(91);
    layer0_outputs(1405) <= not(inputs(86));
    layer0_outputs(1406) <= inputs(195);
    layer0_outputs(1407) <= not(inputs(210)) or (inputs(219));
    layer0_outputs(1408) <= not(inputs(84)) or (inputs(143));
    layer0_outputs(1409) <= inputs(21);
    layer0_outputs(1410) <= (inputs(27)) or (inputs(225));
    layer0_outputs(1411) <= (inputs(171)) and not (inputs(6));
    layer0_outputs(1412) <= (inputs(246)) and not (inputs(252));
    layer0_outputs(1413) <= inputs(106);
    layer0_outputs(1414) <= not(inputs(190));
    layer0_outputs(1415) <= not((inputs(194)) or (inputs(36)));
    layer0_outputs(1416) <= not(inputs(165));
    layer0_outputs(1417) <= (inputs(48)) or (inputs(14));
    layer0_outputs(1418) <= not(inputs(228));
    layer0_outputs(1419) <= not((inputs(127)) or (inputs(186)));
    layer0_outputs(1420) <= not(inputs(94)) or (inputs(239));
    layer0_outputs(1421) <= inputs(131);
    layer0_outputs(1422) <= not((inputs(113)) or (inputs(192)));
    layer0_outputs(1423) <= inputs(164);
    layer0_outputs(1424) <= inputs(23);
    layer0_outputs(1425) <= (inputs(233)) or (inputs(175));
    layer0_outputs(1426) <= not((inputs(244)) or (inputs(255)));
    layer0_outputs(1427) <= (inputs(192)) and not (inputs(230));
    layer0_outputs(1428) <= not(inputs(26));
    layer0_outputs(1429) <= inputs(124);
    layer0_outputs(1430) <= not(inputs(133)) or (inputs(51));
    layer0_outputs(1431) <= (inputs(16)) or (inputs(153));
    layer0_outputs(1432) <= not((inputs(14)) or (inputs(232)));
    layer0_outputs(1433) <= (inputs(2)) or (inputs(159));
    layer0_outputs(1434) <= inputs(217);
    layer0_outputs(1435) <= not(inputs(44)) or (inputs(253));
    layer0_outputs(1436) <= (inputs(151)) and not (inputs(203));
    layer0_outputs(1437) <= not(inputs(76));
    layer0_outputs(1438) <= (inputs(70)) or (inputs(242));
    layer0_outputs(1439) <= not((inputs(78)) or (inputs(61)));
    layer0_outputs(1440) <= inputs(24);
    layer0_outputs(1441) <= not(inputs(99));
    layer0_outputs(1442) <= inputs(149);
    layer0_outputs(1443) <= (inputs(183)) or (inputs(168));
    layer0_outputs(1444) <= not(inputs(155)) or (inputs(222));
    layer0_outputs(1445) <= not((inputs(216)) or (inputs(219)));
    layer0_outputs(1446) <= not(inputs(33));
    layer0_outputs(1447) <= inputs(211);
    layer0_outputs(1448) <= inputs(248);
    layer0_outputs(1449) <= inputs(119);
    layer0_outputs(1450) <= not((inputs(90)) or (inputs(26)));
    layer0_outputs(1451) <= not((inputs(32)) or (inputs(232)));
    layer0_outputs(1452) <= (inputs(109)) and not (inputs(177));
    layer0_outputs(1453) <= not(inputs(151)) or (inputs(58));
    layer0_outputs(1454) <= (inputs(59)) and not (inputs(240));
    layer0_outputs(1455) <= inputs(175);
    layer0_outputs(1456) <= not(inputs(246)) or (inputs(144));
    layer0_outputs(1457) <= not(inputs(42)) or (inputs(31));
    layer0_outputs(1458) <= (inputs(92)) and (inputs(23));
    layer0_outputs(1459) <= not(inputs(227));
    layer0_outputs(1460) <= inputs(84);
    layer0_outputs(1461) <= not(inputs(70));
    layer0_outputs(1462) <= inputs(109);
    layer0_outputs(1463) <= not((inputs(188)) or (inputs(212)));
    layer0_outputs(1464) <= not(inputs(38)) or (inputs(208));
    layer0_outputs(1465) <= not(inputs(85));
    layer0_outputs(1466) <= not(inputs(180));
    layer0_outputs(1467) <= not((inputs(247)) or (inputs(212)));
    layer0_outputs(1468) <= not(inputs(253));
    layer0_outputs(1469) <= not(inputs(239));
    layer0_outputs(1470) <= (inputs(105)) and not (inputs(51));
    layer0_outputs(1471) <= not((inputs(73)) and (inputs(219)));
    layer0_outputs(1472) <= inputs(122);
    layer0_outputs(1473) <= not(inputs(173));
    layer0_outputs(1474) <= (inputs(249)) or (inputs(86));
    layer0_outputs(1475) <= (inputs(98)) or (inputs(87));
    layer0_outputs(1476) <= inputs(223);
    layer0_outputs(1477) <= not(inputs(213));
    layer0_outputs(1478) <= not(inputs(118)) or (inputs(124));
    layer0_outputs(1479) <= not((inputs(173)) and (inputs(182)));
    layer0_outputs(1480) <= not(inputs(43)) or (inputs(207));
    layer0_outputs(1481) <= not((inputs(146)) or (inputs(216)));
    layer0_outputs(1482) <= not(inputs(213)) or (inputs(68));
    layer0_outputs(1483) <= inputs(82);
    layer0_outputs(1484) <= inputs(118);
    layer0_outputs(1485) <= not(inputs(147));
    layer0_outputs(1486) <= (inputs(84)) and not (inputs(203));
    layer0_outputs(1487) <= not((inputs(53)) or (inputs(102)));
    layer0_outputs(1488) <= not((inputs(209)) or (inputs(23)));
    layer0_outputs(1489) <= (inputs(118)) and not (inputs(162));
    layer0_outputs(1490) <= not(inputs(24));
    layer0_outputs(1491) <= (inputs(215)) or (inputs(234));
    layer0_outputs(1492) <= not((inputs(68)) or (inputs(110)));
    layer0_outputs(1493) <= (inputs(217)) and (inputs(243));
    layer0_outputs(1494) <= inputs(195);
    layer0_outputs(1495) <= not(inputs(84));
    layer0_outputs(1496) <= inputs(34);
    layer0_outputs(1497) <= (inputs(106)) or (inputs(105));
    layer0_outputs(1498) <= inputs(73);
    layer0_outputs(1499) <= not((inputs(0)) xor (inputs(147)));
    layer0_outputs(1500) <= not(inputs(76));
    layer0_outputs(1501) <= not(inputs(197));
    layer0_outputs(1502) <= inputs(124);
    layer0_outputs(1503) <= not(inputs(79)) or (inputs(191));
    layer0_outputs(1504) <= (inputs(50)) or (inputs(31));
    layer0_outputs(1505) <= not((inputs(19)) or (inputs(124)));
    layer0_outputs(1506) <= (inputs(156)) or (inputs(165));
    layer0_outputs(1507) <= inputs(182);
    layer0_outputs(1508) <= not((inputs(98)) or (inputs(161)));
    layer0_outputs(1509) <= not(inputs(149));
    layer0_outputs(1510) <= (inputs(203)) and not (inputs(52));
    layer0_outputs(1511) <= (inputs(101)) and not (inputs(175));
    layer0_outputs(1512) <= not(inputs(26)) or (inputs(229));
    layer0_outputs(1513) <= not(inputs(107));
    layer0_outputs(1514) <= not(inputs(194));
    layer0_outputs(1515) <= (inputs(136)) and not (inputs(145));
    layer0_outputs(1516) <= (inputs(250)) and not (inputs(28));
    layer0_outputs(1517) <= not(inputs(151));
    layer0_outputs(1518) <= not(inputs(161)) or (inputs(34));
    layer0_outputs(1519) <= (inputs(68)) or (inputs(146));
    layer0_outputs(1520) <= (inputs(10)) or (inputs(6));
    layer0_outputs(1521) <= (inputs(205)) and not (inputs(189));
    layer0_outputs(1522) <= not((inputs(77)) or (inputs(90)));
    layer0_outputs(1523) <= (inputs(39)) or (inputs(239));
    layer0_outputs(1524) <= '0';
    layer0_outputs(1525) <= (inputs(167)) and not (inputs(114));
    layer0_outputs(1526) <= not(inputs(111));
    layer0_outputs(1527) <= (inputs(201)) xor (inputs(166));
    layer0_outputs(1528) <= inputs(228);
    layer0_outputs(1529) <= inputs(104);
    layer0_outputs(1530) <= (inputs(157)) or (inputs(4));
    layer0_outputs(1531) <= (inputs(60)) and not (inputs(87));
    layer0_outputs(1532) <= not((inputs(233)) or (inputs(65)));
    layer0_outputs(1533) <= inputs(98);
    layer0_outputs(1534) <= not(inputs(163)) or (inputs(169));
    layer0_outputs(1535) <= (inputs(131)) and not (inputs(238));
    layer0_outputs(1536) <= (inputs(59)) or (inputs(64));
    layer0_outputs(1537) <= (inputs(204)) or (inputs(157));
    layer0_outputs(1538) <= not(inputs(182));
    layer0_outputs(1539) <= not(inputs(242));
    layer0_outputs(1540) <= (inputs(95)) or (inputs(233));
    layer0_outputs(1541) <= not(inputs(98));
    layer0_outputs(1542) <= (inputs(20)) and not (inputs(254));
    layer0_outputs(1543) <= (inputs(62)) or (inputs(45));
    layer0_outputs(1544) <= (inputs(242)) or (inputs(127));
    layer0_outputs(1545) <= (inputs(248)) and (inputs(248));
    layer0_outputs(1546) <= inputs(254);
    layer0_outputs(1547) <= (inputs(209)) or (inputs(175));
    layer0_outputs(1548) <= not((inputs(245)) xor (inputs(178)));
    layer0_outputs(1549) <= inputs(205);
    layer0_outputs(1550) <= not(inputs(102));
    layer0_outputs(1551) <= not((inputs(65)) or (inputs(50)));
    layer0_outputs(1552) <= (inputs(129)) or (inputs(174));
    layer0_outputs(1553) <= inputs(133);
    layer0_outputs(1554) <= inputs(234);
    layer0_outputs(1555) <= (inputs(25)) and not (inputs(147));
    layer0_outputs(1556) <= (inputs(136)) and not (inputs(162));
    layer0_outputs(1557) <= (inputs(22)) or (inputs(81));
    layer0_outputs(1558) <= not(inputs(103));
    layer0_outputs(1559) <= not((inputs(222)) or (inputs(219)));
    layer0_outputs(1560) <= inputs(131);
    layer0_outputs(1561) <= inputs(85);
    layer0_outputs(1562) <= (inputs(147)) or (inputs(98));
    layer0_outputs(1563) <= inputs(228);
    layer0_outputs(1564) <= not(inputs(156)) or (inputs(46));
    layer0_outputs(1565) <= not(inputs(211)) or (inputs(111));
    layer0_outputs(1566) <= not((inputs(78)) xor (inputs(167)));
    layer0_outputs(1567) <= (inputs(227)) or (inputs(249));
    layer0_outputs(1568) <= (inputs(5)) and not (inputs(179));
    layer0_outputs(1569) <= inputs(200);
    layer0_outputs(1570) <= not(inputs(233)) or (inputs(70));
    layer0_outputs(1571) <= (inputs(241)) or (inputs(243));
    layer0_outputs(1572) <= not((inputs(54)) or (inputs(230)));
    layer0_outputs(1573) <= (inputs(88)) and not (inputs(34));
    layer0_outputs(1574) <= not(inputs(74));
    layer0_outputs(1575) <= not(inputs(82)) or (inputs(65));
    layer0_outputs(1576) <= (inputs(58)) and not (inputs(174));
    layer0_outputs(1577) <= (inputs(142)) or (inputs(207));
    layer0_outputs(1578) <= inputs(225);
    layer0_outputs(1579) <= (inputs(166)) or (inputs(185));
    layer0_outputs(1580) <= not(inputs(122)) or (inputs(178));
    layer0_outputs(1581) <= inputs(138);
    layer0_outputs(1582) <= inputs(99);
    layer0_outputs(1583) <= not(inputs(106)) or (inputs(242));
    layer0_outputs(1584) <= not(inputs(110));
    layer0_outputs(1585) <= not((inputs(35)) or (inputs(39)));
    layer0_outputs(1586) <= (inputs(104)) or (inputs(133));
    layer0_outputs(1587) <= not(inputs(156));
    layer0_outputs(1588) <= (inputs(212)) or (inputs(209));
    layer0_outputs(1589) <= not((inputs(81)) or (inputs(87)));
    layer0_outputs(1590) <= (inputs(194)) and not (inputs(55));
    layer0_outputs(1591) <= not(inputs(108)) or (inputs(135));
    layer0_outputs(1592) <= '1';
    layer0_outputs(1593) <= not(inputs(211));
    layer0_outputs(1594) <= not(inputs(57));
    layer0_outputs(1595) <= not(inputs(106));
    layer0_outputs(1596) <= not((inputs(241)) or (inputs(41)));
    layer0_outputs(1597) <= not(inputs(226));
    layer0_outputs(1598) <= (inputs(26)) and not (inputs(85));
    layer0_outputs(1599) <= inputs(100);
    layer0_outputs(1600) <= not((inputs(151)) or (inputs(251)));
    layer0_outputs(1601) <= (inputs(152)) and not (inputs(49));
    layer0_outputs(1602) <= inputs(102);
    layer0_outputs(1603) <= (inputs(165)) and not (inputs(47));
    layer0_outputs(1604) <= not((inputs(87)) and (inputs(65)));
    layer0_outputs(1605) <= not(inputs(168)) or (inputs(67));
    layer0_outputs(1606) <= '1';
    layer0_outputs(1607) <= not((inputs(19)) or (inputs(32)));
    layer0_outputs(1608) <= (inputs(51)) and not (inputs(123));
    layer0_outputs(1609) <= not((inputs(230)) and (inputs(153)));
    layer0_outputs(1610) <= (inputs(161)) xor (inputs(105));
    layer0_outputs(1611) <= (inputs(132)) and not (inputs(19));
    layer0_outputs(1612) <= not((inputs(92)) or (inputs(112)));
    layer0_outputs(1613) <= not((inputs(9)) or (inputs(99)));
    layer0_outputs(1614) <= not((inputs(89)) or (inputs(166)));
    layer0_outputs(1615) <= '1';
    layer0_outputs(1616) <= (inputs(8)) and not (inputs(177));
    layer0_outputs(1617) <= '0';
    layer0_outputs(1618) <= inputs(9);
    layer0_outputs(1619) <= not((inputs(174)) and (inputs(222)));
    layer0_outputs(1620) <= not(inputs(139)) or (inputs(153));
    layer0_outputs(1621) <= inputs(84);
    layer0_outputs(1622) <= not(inputs(240));
    layer0_outputs(1623) <= inputs(152);
    layer0_outputs(1624) <= inputs(114);
    layer0_outputs(1625) <= inputs(165);
    layer0_outputs(1626) <= not((inputs(233)) or (inputs(217)));
    layer0_outputs(1627) <= '1';
    layer0_outputs(1628) <= not(inputs(104)) or (inputs(12));
    layer0_outputs(1629) <= not(inputs(255)) or (inputs(98));
    layer0_outputs(1630) <= not(inputs(135)) or (inputs(164));
    layer0_outputs(1631) <= not((inputs(65)) or (inputs(238)));
    layer0_outputs(1632) <= inputs(232);
    layer0_outputs(1633) <= (inputs(45)) and not (inputs(239));
    layer0_outputs(1634) <= not((inputs(203)) or (inputs(103)));
    layer0_outputs(1635) <= (inputs(69)) or (inputs(84));
    layer0_outputs(1636) <= inputs(230);
    layer0_outputs(1637) <= inputs(12);
    layer0_outputs(1638) <= not((inputs(109)) or (inputs(175)));
    layer0_outputs(1639) <= not(inputs(43)) or (inputs(238));
    layer0_outputs(1640) <= inputs(248);
    layer0_outputs(1641) <= not(inputs(75));
    layer0_outputs(1642) <= (inputs(178)) or (inputs(235));
    layer0_outputs(1643) <= (inputs(105)) xor (inputs(175));
    layer0_outputs(1644) <= inputs(229);
    layer0_outputs(1645) <= (inputs(228)) and not (inputs(1));
    layer0_outputs(1646) <= inputs(4);
    layer0_outputs(1647) <= (inputs(7)) xor (inputs(217));
    layer0_outputs(1648) <= not(inputs(27));
    layer0_outputs(1649) <= not(inputs(188));
    layer0_outputs(1650) <= (inputs(233)) and (inputs(90));
    layer0_outputs(1651) <= (inputs(209)) or (inputs(15));
    layer0_outputs(1652) <= inputs(126);
    layer0_outputs(1653) <= not(inputs(180));
    layer0_outputs(1654) <= (inputs(172)) or (inputs(138));
    layer0_outputs(1655) <= not(inputs(178));
    layer0_outputs(1656) <= not(inputs(8));
    layer0_outputs(1657) <= (inputs(156)) xor (inputs(252));
    layer0_outputs(1658) <= inputs(78);
    layer0_outputs(1659) <= inputs(218);
    layer0_outputs(1660) <= inputs(33);
    layer0_outputs(1661) <= not((inputs(64)) or (inputs(254)));
    layer0_outputs(1662) <= (inputs(61)) and not (inputs(227));
    layer0_outputs(1663) <= not((inputs(156)) xor (inputs(253)));
    layer0_outputs(1664) <= (inputs(252)) xor (inputs(70));
    layer0_outputs(1665) <= not((inputs(170)) or (inputs(130)));
    layer0_outputs(1666) <= (inputs(109)) or (inputs(213));
    layer0_outputs(1667) <= inputs(131);
    layer0_outputs(1668) <= inputs(13);
    layer0_outputs(1669) <= inputs(70);
    layer0_outputs(1670) <= inputs(150);
    layer0_outputs(1671) <= inputs(78);
    layer0_outputs(1672) <= inputs(56);
    layer0_outputs(1673) <= not((inputs(218)) or (inputs(192)));
    layer0_outputs(1674) <= inputs(45);
    layer0_outputs(1675) <= not(inputs(230));
    layer0_outputs(1676) <= inputs(137);
    layer0_outputs(1677) <= (inputs(56)) or (inputs(7));
    layer0_outputs(1678) <= inputs(10);
    layer0_outputs(1679) <= (inputs(75)) or (inputs(5));
    layer0_outputs(1680) <= not(inputs(71));
    layer0_outputs(1681) <= not(inputs(102));
    layer0_outputs(1682) <= (inputs(156)) or (inputs(125));
    layer0_outputs(1683) <= not(inputs(213)) or (inputs(0));
    layer0_outputs(1684) <= inputs(141);
    layer0_outputs(1685) <= (inputs(87)) or (inputs(99));
    layer0_outputs(1686) <= not(inputs(42)) or (inputs(97));
    layer0_outputs(1687) <= not(inputs(231));
    layer0_outputs(1688) <= not((inputs(19)) xor (inputs(64)));
    layer0_outputs(1689) <= '1';
    layer0_outputs(1690) <= inputs(56);
    layer0_outputs(1691) <= not(inputs(229));
    layer0_outputs(1692) <= not(inputs(52)) or (inputs(252));
    layer0_outputs(1693) <= (inputs(39)) and not (inputs(248));
    layer0_outputs(1694) <= inputs(134);
    layer0_outputs(1695) <= not((inputs(32)) or (inputs(154)));
    layer0_outputs(1696) <= inputs(167);
    layer0_outputs(1697) <= inputs(218);
    layer0_outputs(1698) <= inputs(186);
    layer0_outputs(1699) <= not((inputs(80)) or (inputs(235)));
    layer0_outputs(1700) <= (inputs(88)) and not (inputs(202));
    layer0_outputs(1701) <= (inputs(182)) and not (inputs(127));
    layer0_outputs(1702) <= not(inputs(119));
    layer0_outputs(1703) <= (inputs(26)) or (inputs(192));
    layer0_outputs(1704) <= not(inputs(137)) or (inputs(215));
    layer0_outputs(1705) <= not(inputs(150));
    layer0_outputs(1706) <= (inputs(51)) and not (inputs(130));
    layer0_outputs(1707) <= not((inputs(18)) or (inputs(225)));
    layer0_outputs(1708) <= inputs(178);
    layer0_outputs(1709) <= not(inputs(217));
    layer0_outputs(1710) <= (inputs(152)) and not (inputs(112));
    layer0_outputs(1711) <= (inputs(156)) or (inputs(155));
    layer0_outputs(1712) <= not(inputs(69));
    layer0_outputs(1713) <= (inputs(218)) or (inputs(172));
    layer0_outputs(1714) <= not(inputs(79));
    layer0_outputs(1715) <= inputs(3);
    layer0_outputs(1716) <= not(inputs(137)) or (inputs(63));
    layer0_outputs(1717) <= inputs(91);
    layer0_outputs(1718) <= (inputs(197)) xor (inputs(12));
    layer0_outputs(1719) <= not(inputs(59));
    layer0_outputs(1720) <= (inputs(214)) and not (inputs(253));
    layer0_outputs(1721) <= not(inputs(156));
    layer0_outputs(1722) <= not((inputs(122)) or (inputs(90)));
    layer0_outputs(1723) <= not(inputs(228));
    layer0_outputs(1724) <= not(inputs(42)) or (inputs(128));
    layer0_outputs(1725) <= (inputs(226)) and not (inputs(113));
    layer0_outputs(1726) <= not(inputs(152));
    layer0_outputs(1727) <= not(inputs(179));
    layer0_outputs(1728) <= not(inputs(212)) or (inputs(26));
    layer0_outputs(1729) <= (inputs(208)) or (inputs(69));
    layer0_outputs(1730) <= inputs(49);
    layer0_outputs(1731) <= '0';
    layer0_outputs(1732) <= (inputs(139)) and not (inputs(14));
    layer0_outputs(1733) <= not(inputs(93)) or (inputs(97));
    layer0_outputs(1734) <= not(inputs(21));
    layer0_outputs(1735) <= (inputs(252)) xor (inputs(80));
    layer0_outputs(1736) <= not(inputs(211));
    layer0_outputs(1737) <= '1';
    layer0_outputs(1738) <= inputs(165);
    layer0_outputs(1739) <= not((inputs(208)) or (inputs(190)));
    layer0_outputs(1740) <= not((inputs(108)) or (inputs(8)));
    layer0_outputs(1741) <= (inputs(91)) or (inputs(182));
    layer0_outputs(1742) <= not((inputs(140)) or (inputs(187)));
    layer0_outputs(1743) <= not(inputs(38)) or (inputs(254));
    layer0_outputs(1744) <= not(inputs(209));
    layer0_outputs(1745) <= not((inputs(29)) or (inputs(78)));
    layer0_outputs(1746) <= (inputs(31)) xor (inputs(77));
    layer0_outputs(1747) <= not((inputs(72)) or (inputs(160)));
    layer0_outputs(1748) <= not(inputs(134));
    layer0_outputs(1749) <= inputs(223);
    layer0_outputs(1750) <= (inputs(173)) and not (inputs(64));
    layer0_outputs(1751) <= not(inputs(9));
    layer0_outputs(1752) <= not((inputs(255)) or (inputs(20)));
    layer0_outputs(1753) <= not(inputs(26));
    layer0_outputs(1754) <= inputs(218);
    layer0_outputs(1755) <= not((inputs(146)) or (inputs(119)));
    layer0_outputs(1756) <= not(inputs(98));
    layer0_outputs(1757) <= not(inputs(115)) or (inputs(77));
    layer0_outputs(1758) <= inputs(203);
    layer0_outputs(1759) <= (inputs(123)) or (inputs(176));
    layer0_outputs(1760) <= (inputs(235)) and not (inputs(134));
    layer0_outputs(1761) <= (inputs(76)) or (inputs(30));
    layer0_outputs(1762) <= inputs(69);
    layer0_outputs(1763) <= not((inputs(98)) or (inputs(158)));
    layer0_outputs(1764) <= not(inputs(41)) or (inputs(77));
    layer0_outputs(1765) <= (inputs(241)) xor (inputs(234));
    layer0_outputs(1766) <= not((inputs(113)) or (inputs(29)));
    layer0_outputs(1767) <= inputs(10);
    layer0_outputs(1768) <= (inputs(70)) and not (inputs(164));
    layer0_outputs(1769) <= not(inputs(176));
    layer0_outputs(1770) <= inputs(135);
    layer0_outputs(1771) <= (inputs(20)) or (inputs(111));
    layer0_outputs(1772) <= not(inputs(35));
    layer0_outputs(1773) <= (inputs(124)) and not (inputs(5));
    layer0_outputs(1774) <= inputs(232);
    layer0_outputs(1775) <= not(inputs(186));
    layer0_outputs(1776) <= not(inputs(247));
    layer0_outputs(1777) <= (inputs(229)) and not (inputs(15));
    layer0_outputs(1778) <= not((inputs(72)) or (inputs(56)));
    layer0_outputs(1779) <= (inputs(47)) and not (inputs(175));
    layer0_outputs(1780) <= not(inputs(42));
    layer0_outputs(1781) <= (inputs(119)) and not (inputs(142));
    layer0_outputs(1782) <= (inputs(76)) or (inputs(127));
    layer0_outputs(1783) <= not(inputs(247));
    layer0_outputs(1784) <= not((inputs(148)) or (inputs(224)));
    layer0_outputs(1785) <= inputs(34);
    layer0_outputs(1786) <= (inputs(22)) and not (inputs(99));
    layer0_outputs(1787) <= not((inputs(223)) or (inputs(102)));
    layer0_outputs(1788) <= inputs(209);
    layer0_outputs(1789) <= (inputs(169)) and (inputs(27));
    layer0_outputs(1790) <= not(inputs(36));
    layer0_outputs(1791) <= (inputs(107)) and (inputs(138));
    layer0_outputs(1792) <= not((inputs(161)) or (inputs(104)));
    layer0_outputs(1793) <= inputs(77);
    layer0_outputs(1794) <= not(inputs(212));
    layer0_outputs(1795) <= (inputs(108)) or (inputs(213));
    layer0_outputs(1796) <= (inputs(76)) or (inputs(217));
    layer0_outputs(1797) <= inputs(8);
    layer0_outputs(1798) <= '1';
    layer0_outputs(1799) <= not(inputs(189)) or (inputs(30));
    layer0_outputs(1800) <= inputs(62);
    layer0_outputs(1801) <= inputs(12);
    layer0_outputs(1802) <= inputs(145);
    layer0_outputs(1803) <= (inputs(115)) and not (inputs(79));
    layer0_outputs(1804) <= inputs(109);
    layer0_outputs(1805) <= inputs(200);
    layer0_outputs(1806) <= inputs(160);
    layer0_outputs(1807) <= inputs(52);
    layer0_outputs(1808) <= inputs(216);
    layer0_outputs(1809) <= '0';
    layer0_outputs(1810) <= not((inputs(55)) or (inputs(84)));
    layer0_outputs(1811) <= (inputs(35)) or (inputs(29));
    layer0_outputs(1812) <= (inputs(16)) or (inputs(245));
    layer0_outputs(1813) <= (inputs(156)) and not (inputs(35));
    layer0_outputs(1814) <= not(inputs(186)) or (inputs(143));
    layer0_outputs(1815) <= not((inputs(126)) or (inputs(14)));
    layer0_outputs(1816) <= not(inputs(19)) or (inputs(174));
    layer0_outputs(1817) <= not(inputs(22)) or (inputs(70));
    layer0_outputs(1818) <= '0';
    layer0_outputs(1819) <= inputs(212);
    layer0_outputs(1820) <= not((inputs(194)) or (inputs(146)));
    layer0_outputs(1821) <= not((inputs(236)) and (inputs(242)));
    layer0_outputs(1822) <= inputs(139);
    layer0_outputs(1823) <= inputs(60);
    layer0_outputs(1824) <= not(inputs(11));
    layer0_outputs(1825) <= inputs(232);
    layer0_outputs(1826) <= not((inputs(205)) or (inputs(173)));
    layer0_outputs(1827) <= inputs(121);
    layer0_outputs(1828) <= inputs(75);
    layer0_outputs(1829) <= (inputs(122)) or (inputs(202));
    layer0_outputs(1830) <= not(inputs(154));
    layer0_outputs(1831) <= inputs(129);
    layer0_outputs(1832) <= not(inputs(211));
    layer0_outputs(1833) <= (inputs(8)) or (inputs(210));
    layer0_outputs(1834) <= (inputs(20)) or (inputs(56));
    layer0_outputs(1835) <= (inputs(155)) and not (inputs(63));
    layer0_outputs(1836) <= (inputs(177)) or (inputs(131));
    layer0_outputs(1837) <= not(inputs(27));
    layer0_outputs(1838) <= (inputs(125)) and not (inputs(51));
    layer0_outputs(1839) <= not(inputs(142));
    layer0_outputs(1840) <= not((inputs(85)) or (inputs(114)));
    layer0_outputs(1841) <= not((inputs(168)) or (inputs(237)));
    layer0_outputs(1842) <= inputs(7);
    layer0_outputs(1843) <= (inputs(212)) and not (inputs(236));
    layer0_outputs(1844) <= not(inputs(83));
    layer0_outputs(1845) <= not(inputs(130));
    layer0_outputs(1846) <= inputs(90);
    layer0_outputs(1847) <= not((inputs(224)) and (inputs(204)));
    layer0_outputs(1848) <= (inputs(104)) and not (inputs(148));
    layer0_outputs(1849) <= not(inputs(53)) or (inputs(95));
    layer0_outputs(1850) <= (inputs(232)) and not (inputs(25));
    layer0_outputs(1851) <= inputs(226);
    layer0_outputs(1852) <= inputs(122);
    layer0_outputs(1853) <= not(inputs(53));
    layer0_outputs(1854) <= not(inputs(78));
    layer0_outputs(1855) <= not(inputs(96));
    layer0_outputs(1856) <= inputs(94);
    layer0_outputs(1857) <= '0';
    layer0_outputs(1858) <= (inputs(247)) or (inputs(133));
    layer0_outputs(1859) <= not((inputs(236)) or (inputs(191)));
    layer0_outputs(1860) <= not(inputs(23));
    layer0_outputs(1861) <= (inputs(47)) and not (inputs(224));
    layer0_outputs(1862) <= '0';
    layer0_outputs(1863) <= not(inputs(219)) or (inputs(93));
    layer0_outputs(1864) <= '1';
    layer0_outputs(1865) <= inputs(176);
    layer0_outputs(1866) <= not(inputs(119)) or (inputs(51));
    layer0_outputs(1867) <= not(inputs(140));
    layer0_outputs(1868) <= inputs(200);
    layer0_outputs(1869) <= not(inputs(232));
    layer0_outputs(1870) <= not(inputs(184)) or (inputs(111));
    layer0_outputs(1871) <= not((inputs(112)) xor (inputs(250)));
    layer0_outputs(1872) <= inputs(67);
    layer0_outputs(1873) <= (inputs(22)) and not (inputs(63));
    layer0_outputs(1874) <= not((inputs(53)) or (inputs(177)));
    layer0_outputs(1875) <= inputs(196);
    layer0_outputs(1876) <= not(inputs(163));
    layer0_outputs(1877) <= not((inputs(159)) or (inputs(86)));
    layer0_outputs(1878) <= (inputs(151)) and not (inputs(67));
    layer0_outputs(1879) <= '0';
    layer0_outputs(1880) <= inputs(145);
    layer0_outputs(1881) <= not(inputs(214)) or (inputs(92));
    layer0_outputs(1882) <= (inputs(195)) or (inputs(69));
    layer0_outputs(1883) <= (inputs(237)) and not (inputs(113));
    layer0_outputs(1884) <= (inputs(159)) and not (inputs(56));
    layer0_outputs(1885) <= (inputs(7)) or (inputs(9));
    layer0_outputs(1886) <= (inputs(239)) or (inputs(114));
    layer0_outputs(1887) <= inputs(164);
    layer0_outputs(1888) <= not(inputs(247)) or (inputs(145));
    layer0_outputs(1889) <= '1';
    layer0_outputs(1890) <= inputs(79);
    layer0_outputs(1891) <= not(inputs(43)) or (inputs(205));
    layer0_outputs(1892) <= not(inputs(23));
    layer0_outputs(1893) <= not(inputs(100));
    layer0_outputs(1894) <= not((inputs(104)) or (inputs(16)));
    layer0_outputs(1895) <= (inputs(246)) and not (inputs(163));
    layer0_outputs(1896) <= inputs(23);
    layer0_outputs(1897) <= not((inputs(237)) or (inputs(198)));
    layer0_outputs(1898) <= (inputs(110)) or (inputs(242));
    layer0_outputs(1899) <= not((inputs(28)) or (inputs(122)));
    layer0_outputs(1900) <= inputs(59);
    layer0_outputs(1901) <= not(inputs(84)) or (inputs(64));
    layer0_outputs(1902) <= not((inputs(27)) or (inputs(253)));
    layer0_outputs(1903) <= not(inputs(14));
    layer0_outputs(1904) <= inputs(226);
    layer0_outputs(1905) <= not(inputs(231));
    layer0_outputs(1906) <= inputs(248);
    layer0_outputs(1907) <= (inputs(166)) and not (inputs(77));
    layer0_outputs(1908) <= inputs(162);
    layer0_outputs(1909) <= (inputs(168)) and not (inputs(96));
    layer0_outputs(1910) <= (inputs(96)) and not (inputs(148));
    layer0_outputs(1911) <= not(inputs(206)) or (inputs(250));
    layer0_outputs(1912) <= (inputs(195)) or (inputs(77));
    layer0_outputs(1913) <= inputs(39);
    layer0_outputs(1914) <= (inputs(74)) and not (inputs(170));
    layer0_outputs(1915) <= inputs(126);
    layer0_outputs(1916) <= (inputs(166)) or (inputs(90));
    layer0_outputs(1917) <= not(inputs(243));
    layer0_outputs(1918) <= inputs(93);
    layer0_outputs(1919) <= not(inputs(172)) or (inputs(14));
    layer0_outputs(1920) <= (inputs(251)) or (inputs(189));
    layer0_outputs(1921) <= not((inputs(6)) or (inputs(61)));
    layer0_outputs(1922) <= '0';
    layer0_outputs(1923) <= inputs(231);
    layer0_outputs(1924) <= (inputs(59)) and not (inputs(45));
    layer0_outputs(1925) <= not(inputs(105));
    layer0_outputs(1926) <= not(inputs(18)) or (inputs(250));
    layer0_outputs(1927) <= not(inputs(153));
    layer0_outputs(1928) <= not(inputs(7)) or (inputs(25));
    layer0_outputs(1929) <= not(inputs(20)) or (inputs(255));
    layer0_outputs(1930) <= not(inputs(106)) or (inputs(161));
    layer0_outputs(1931) <= not((inputs(146)) or (inputs(188)));
    layer0_outputs(1932) <= inputs(139);
    layer0_outputs(1933) <= '1';
    layer0_outputs(1934) <= (inputs(48)) and not (inputs(243));
    layer0_outputs(1935) <= (inputs(36)) and not (inputs(128));
    layer0_outputs(1936) <= not(inputs(109)) or (inputs(65));
    layer0_outputs(1937) <= (inputs(190)) or (inputs(82));
    layer0_outputs(1938) <= (inputs(244)) or (inputs(16));
    layer0_outputs(1939) <= inputs(69);
    layer0_outputs(1940) <= (inputs(84)) xor (inputs(71));
    layer0_outputs(1941) <= inputs(140);
    layer0_outputs(1942) <= '1';
    layer0_outputs(1943) <= inputs(154);
    layer0_outputs(1944) <= not(inputs(50));
    layer0_outputs(1945) <= (inputs(116)) or (inputs(180));
    layer0_outputs(1946) <= not(inputs(168)) or (inputs(194));
    layer0_outputs(1947) <= (inputs(173)) or (inputs(7));
    layer0_outputs(1948) <= not(inputs(142));
    layer0_outputs(1949) <= (inputs(38)) and not (inputs(144));
    layer0_outputs(1950) <= not(inputs(116)) or (inputs(110));
    layer0_outputs(1951) <= inputs(101);
    layer0_outputs(1952) <= not(inputs(143)) or (inputs(34));
    layer0_outputs(1953) <= inputs(229);
    layer0_outputs(1954) <= (inputs(163)) or (inputs(207));
    layer0_outputs(1955) <= inputs(104);
    layer0_outputs(1956) <= not(inputs(93));
    layer0_outputs(1957) <= (inputs(193)) xor (inputs(101));
    layer0_outputs(1958) <= (inputs(93)) and not (inputs(48));
    layer0_outputs(1959) <= (inputs(200)) xor (inputs(241));
    layer0_outputs(1960) <= not((inputs(221)) or (inputs(226)));
    layer0_outputs(1961) <= not(inputs(17)) or (inputs(92));
    layer0_outputs(1962) <= not(inputs(18));
    layer0_outputs(1963) <= inputs(3);
    layer0_outputs(1964) <= not(inputs(85));
    layer0_outputs(1965) <= (inputs(99)) and not (inputs(50));
    layer0_outputs(1966) <= (inputs(60)) or (inputs(152));
    layer0_outputs(1967) <= inputs(108);
    layer0_outputs(1968) <= (inputs(40)) and (inputs(125));
    layer0_outputs(1969) <= not(inputs(6));
    layer0_outputs(1970) <= not(inputs(221));
    layer0_outputs(1971) <= (inputs(115)) and not (inputs(154));
    layer0_outputs(1972) <= not((inputs(239)) or (inputs(38)));
    layer0_outputs(1973) <= not(inputs(221));
    layer0_outputs(1974) <= inputs(28);
    layer0_outputs(1975) <= not(inputs(36));
    layer0_outputs(1976) <= not(inputs(148));
    layer0_outputs(1977) <= not(inputs(232));
    layer0_outputs(1978) <= inputs(126);
    layer0_outputs(1979) <= inputs(223);
    layer0_outputs(1980) <= not(inputs(198)) or (inputs(143));
    layer0_outputs(1981) <= not(inputs(140));
    layer0_outputs(1982) <= (inputs(187)) and (inputs(184));
    layer0_outputs(1983) <= not(inputs(89)) or (inputs(210));
    layer0_outputs(1984) <= (inputs(113)) or (inputs(187));
    layer0_outputs(1985) <= not((inputs(171)) or (inputs(98)));
    layer0_outputs(1986) <= (inputs(65)) or (inputs(180));
    layer0_outputs(1987) <= not(inputs(3));
    layer0_outputs(1988) <= (inputs(220)) and not (inputs(13));
    layer0_outputs(1989) <= (inputs(179)) and not (inputs(145));
    layer0_outputs(1990) <= not(inputs(150));
    layer0_outputs(1991) <= not((inputs(162)) or (inputs(17)));
    layer0_outputs(1992) <= inputs(107);
    layer0_outputs(1993) <= not((inputs(66)) or (inputs(129)));
    layer0_outputs(1994) <= not(inputs(117));
    layer0_outputs(1995) <= inputs(48);
    layer0_outputs(1996) <= not(inputs(163));
    layer0_outputs(1997) <= not(inputs(36));
    layer0_outputs(1998) <= (inputs(145)) and not (inputs(254));
    layer0_outputs(1999) <= not(inputs(156));
    layer0_outputs(2000) <= inputs(93);
    layer0_outputs(2001) <= not(inputs(132)) or (inputs(16));
    layer0_outputs(2002) <= inputs(174);
    layer0_outputs(2003) <= not(inputs(160)) or (inputs(30));
    layer0_outputs(2004) <= not((inputs(107)) or (inputs(103)));
    layer0_outputs(2005) <= inputs(246);
    layer0_outputs(2006) <= inputs(231);
    layer0_outputs(2007) <= not(inputs(26)) or (inputs(164));
    layer0_outputs(2008) <= not((inputs(187)) or (inputs(124)));
    layer0_outputs(2009) <= (inputs(54)) xor (inputs(23));
    layer0_outputs(2010) <= inputs(134);
    layer0_outputs(2011) <= (inputs(104)) and not (inputs(112));
    layer0_outputs(2012) <= inputs(173);
    layer0_outputs(2013) <= not(inputs(69)) or (inputs(221));
    layer0_outputs(2014) <= inputs(14);
    layer0_outputs(2015) <= not(inputs(228));
    layer0_outputs(2016) <= inputs(83);
    layer0_outputs(2017) <= not((inputs(123)) or (inputs(238)));
    layer0_outputs(2018) <= not((inputs(242)) or (inputs(208)));
    layer0_outputs(2019) <= (inputs(46)) or (inputs(245));
    layer0_outputs(2020) <= not(inputs(116));
    layer0_outputs(2021) <= not((inputs(180)) or (inputs(248)));
    layer0_outputs(2022) <= not((inputs(102)) or (inputs(178)));
    layer0_outputs(2023) <= not(inputs(128));
    layer0_outputs(2024) <= inputs(36);
    layer0_outputs(2025) <= (inputs(24)) or (inputs(11));
    layer0_outputs(2026) <= not(inputs(151));
    layer0_outputs(2027) <= not(inputs(212)) or (inputs(247));
    layer0_outputs(2028) <= (inputs(107)) and not (inputs(205));
    layer0_outputs(2029) <= not(inputs(225)) or (inputs(2));
    layer0_outputs(2030) <= not(inputs(63)) or (inputs(245));
    layer0_outputs(2031) <= not((inputs(21)) xor (inputs(72)));
    layer0_outputs(2032) <= (inputs(183)) and not (inputs(116));
    layer0_outputs(2033) <= not((inputs(101)) or (inputs(127)));
    layer0_outputs(2034) <= not(inputs(169));
    layer0_outputs(2035) <= not(inputs(150)) or (inputs(247));
    layer0_outputs(2036) <= not((inputs(99)) or (inputs(145)));
    layer0_outputs(2037) <= not(inputs(85));
    layer0_outputs(2038) <= (inputs(4)) and not (inputs(79));
    layer0_outputs(2039) <= not(inputs(219));
    layer0_outputs(2040) <= '1';
    layer0_outputs(2041) <= not((inputs(231)) or (inputs(215)));
    layer0_outputs(2042) <= not(inputs(108)) or (inputs(144));
    layer0_outputs(2043) <= not((inputs(204)) or (inputs(207)));
    layer0_outputs(2044) <= '0';
    layer0_outputs(2045) <= not((inputs(58)) or (inputs(79)));
    layer0_outputs(2046) <= (inputs(194)) and (inputs(194));
    layer0_outputs(2047) <= not(inputs(7));
    layer0_outputs(2048) <= (inputs(184)) xor (inputs(167));
    layer0_outputs(2049) <= (inputs(245)) or (inputs(130));
    layer0_outputs(2050) <= not(inputs(135)) or (inputs(24));
    layer0_outputs(2051) <= not((inputs(234)) or (inputs(61)));
    layer0_outputs(2052) <= not((inputs(179)) or (inputs(209)));
    layer0_outputs(2053) <= not(inputs(247)) or (inputs(107));
    layer0_outputs(2054) <= inputs(58);
    layer0_outputs(2055) <= inputs(144);
    layer0_outputs(2056) <= not((inputs(110)) and (inputs(29)));
    layer0_outputs(2057) <= inputs(148);
    layer0_outputs(2058) <= inputs(86);
    layer0_outputs(2059) <= not((inputs(47)) or (inputs(62)));
    layer0_outputs(2060) <= '1';
    layer0_outputs(2061) <= not(inputs(99));
    layer0_outputs(2062) <= (inputs(217)) or (inputs(213));
    layer0_outputs(2063) <= (inputs(169)) and not (inputs(184));
    layer0_outputs(2064) <= inputs(145);
    layer0_outputs(2065) <= (inputs(70)) and not (inputs(32));
    layer0_outputs(2066) <= not(inputs(67));
    layer0_outputs(2067) <= (inputs(122)) and not (inputs(223));
    layer0_outputs(2068) <= (inputs(214)) and not (inputs(79));
    layer0_outputs(2069) <= not(inputs(230)) or (inputs(182));
    layer0_outputs(2070) <= (inputs(95)) xor (inputs(45));
    layer0_outputs(2071) <= not((inputs(76)) or (inputs(110)));
    layer0_outputs(2072) <= not((inputs(3)) or (inputs(13)));
    layer0_outputs(2073) <= not(inputs(0));
    layer0_outputs(2074) <= not((inputs(207)) or (inputs(192)));
    layer0_outputs(2075) <= inputs(118);
    layer0_outputs(2076) <= not((inputs(114)) xor (inputs(117)));
    layer0_outputs(2077) <= '1';
    layer0_outputs(2078) <= inputs(226);
    layer0_outputs(2079) <= not(inputs(39)) or (inputs(187));
    layer0_outputs(2080) <= inputs(27);
    layer0_outputs(2081) <= (inputs(188)) or (inputs(229));
    layer0_outputs(2082) <= inputs(190);
    layer0_outputs(2083) <= not(inputs(27));
    layer0_outputs(2084) <= (inputs(223)) or (inputs(117));
    layer0_outputs(2085) <= not(inputs(126));
    layer0_outputs(2086) <= inputs(174);
    layer0_outputs(2087) <= not(inputs(248)) or (inputs(0));
    layer0_outputs(2088) <= not((inputs(0)) or (inputs(30)));
    layer0_outputs(2089) <= inputs(178);
    layer0_outputs(2090) <= (inputs(215)) or (inputs(2));
    layer0_outputs(2091) <= not(inputs(176));
    layer0_outputs(2092) <= inputs(77);
    layer0_outputs(2093) <= (inputs(101)) and not (inputs(75));
    layer0_outputs(2094) <= (inputs(55)) and not (inputs(137));
    layer0_outputs(2095) <= (inputs(50)) and (inputs(51));
    layer0_outputs(2096) <= inputs(98);
    layer0_outputs(2097) <= not((inputs(207)) and (inputs(160)));
    layer0_outputs(2098) <= not((inputs(73)) and (inputs(202)));
    layer0_outputs(2099) <= not(inputs(199)) or (inputs(93));
    layer0_outputs(2100) <= not(inputs(177)) or (inputs(126));
    layer0_outputs(2101) <= (inputs(53)) and not (inputs(227));
    layer0_outputs(2102) <= inputs(73);
    layer0_outputs(2103) <= not((inputs(3)) or (inputs(93)));
    layer0_outputs(2104) <= (inputs(144)) or (inputs(210));
    layer0_outputs(2105) <= not(inputs(190));
    layer0_outputs(2106) <= (inputs(222)) and not (inputs(142));
    layer0_outputs(2107) <= not(inputs(149));
    layer0_outputs(2108) <= (inputs(133)) and not (inputs(64));
    layer0_outputs(2109) <= (inputs(249)) and not (inputs(61));
    layer0_outputs(2110) <= not(inputs(218));
    layer0_outputs(2111) <= not((inputs(121)) and (inputs(28)));
    layer0_outputs(2112) <= (inputs(214)) and not (inputs(83));
    layer0_outputs(2113) <= '0';
    layer0_outputs(2114) <= not(inputs(154)) or (inputs(184));
    layer0_outputs(2115) <= inputs(115);
    layer0_outputs(2116) <= (inputs(57)) and not (inputs(107));
    layer0_outputs(2117) <= (inputs(191)) or (inputs(182));
    layer0_outputs(2118) <= not((inputs(37)) or (inputs(81)));
    layer0_outputs(2119) <= inputs(146);
    layer0_outputs(2120) <= (inputs(187)) and not (inputs(20));
    layer0_outputs(2121) <= inputs(130);
    layer0_outputs(2122) <= (inputs(222)) and not (inputs(40));
    layer0_outputs(2123) <= not(inputs(119)) or (inputs(74));
    layer0_outputs(2124) <= (inputs(159)) and not (inputs(109));
    layer0_outputs(2125) <= inputs(10);
    layer0_outputs(2126) <= not(inputs(56)) or (inputs(254));
    layer0_outputs(2127) <= (inputs(51)) or (inputs(162));
    layer0_outputs(2128) <= not((inputs(101)) or (inputs(5)));
    layer0_outputs(2129) <= inputs(232);
    layer0_outputs(2130) <= inputs(131);
    layer0_outputs(2131) <= not(inputs(25));
    layer0_outputs(2132) <= (inputs(8)) and not (inputs(229));
    layer0_outputs(2133) <= inputs(61);
    layer0_outputs(2134) <= (inputs(162)) or (inputs(32));
    layer0_outputs(2135) <= not(inputs(133));
    layer0_outputs(2136) <= inputs(172);
    layer0_outputs(2137) <= not(inputs(144));
    layer0_outputs(2138) <= '0';
    layer0_outputs(2139) <= (inputs(46)) or (inputs(107));
    layer0_outputs(2140) <= (inputs(33)) or (inputs(38));
    layer0_outputs(2141) <= inputs(165);
    layer0_outputs(2142) <= not(inputs(153));
    layer0_outputs(2143) <= '1';
    layer0_outputs(2144) <= inputs(122);
    layer0_outputs(2145) <= not(inputs(253));
    layer0_outputs(2146) <= (inputs(221)) and not (inputs(248));
    layer0_outputs(2147) <= not((inputs(22)) or (inputs(32)));
    layer0_outputs(2148) <= (inputs(230)) and not (inputs(74));
    layer0_outputs(2149) <= '0';
    layer0_outputs(2150) <= not(inputs(177)) or (inputs(61));
    layer0_outputs(2151) <= not((inputs(90)) and (inputs(246)));
    layer0_outputs(2152) <= not(inputs(155)) or (inputs(208));
    layer0_outputs(2153) <= not((inputs(188)) or (inputs(80)));
    layer0_outputs(2154) <= (inputs(86)) and not (inputs(110));
    layer0_outputs(2155) <= not(inputs(53)) or (inputs(255));
    layer0_outputs(2156) <= not(inputs(89));
    layer0_outputs(2157) <= not((inputs(213)) or (inputs(165)));
    layer0_outputs(2158) <= (inputs(96)) or (inputs(82));
    layer0_outputs(2159) <= (inputs(39)) and not (inputs(223));
    layer0_outputs(2160) <= (inputs(194)) or (inputs(65));
    layer0_outputs(2161) <= (inputs(120)) or (inputs(87));
    layer0_outputs(2162) <= not((inputs(252)) or (inputs(251)));
    layer0_outputs(2163) <= not(inputs(33));
    layer0_outputs(2164) <= (inputs(197)) or (inputs(255));
    layer0_outputs(2165) <= not((inputs(188)) or (inputs(148)));
    layer0_outputs(2166) <= not((inputs(64)) and (inputs(1)));
    layer0_outputs(2167) <= (inputs(14)) and not (inputs(249));
    layer0_outputs(2168) <= inputs(143);
    layer0_outputs(2169) <= inputs(148);
    layer0_outputs(2170) <= not((inputs(131)) or (inputs(180)));
    layer0_outputs(2171) <= not((inputs(228)) or (inputs(64)));
    layer0_outputs(2172) <= not(inputs(125));
    layer0_outputs(2173) <= (inputs(188)) or (inputs(72));
    layer0_outputs(2174) <= (inputs(222)) and (inputs(36));
    layer0_outputs(2175) <= (inputs(14)) or (inputs(193));
    layer0_outputs(2176) <= not(inputs(6));
    layer0_outputs(2177) <= inputs(70);
    layer0_outputs(2178) <= not((inputs(35)) or (inputs(247)));
    layer0_outputs(2179) <= (inputs(112)) or (inputs(231));
    layer0_outputs(2180) <= (inputs(49)) or (inputs(239));
    layer0_outputs(2181) <= (inputs(127)) or (inputs(198));
    layer0_outputs(2182) <= inputs(34);
    layer0_outputs(2183) <= not(inputs(134));
    layer0_outputs(2184) <= (inputs(184)) xor (inputs(0));
    layer0_outputs(2185) <= not((inputs(30)) or (inputs(146)));
    layer0_outputs(2186) <= not(inputs(166));
    layer0_outputs(2187) <= inputs(26);
    layer0_outputs(2188) <= not(inputs(39));
    layer0_outputs(2189) <= not(inputs(181));
    layer0_outputs(2190) <= (inputs(35)) or (inputs(3));
    layer0_outputs(2191) <= not(inputs(217)) or (inputs(224));
    layer0_outputs(2192) <= (inputs(92)) and (inputs(43));
    layer0_outputs(2193) <= not((inputs(128)) and (inputs(118)));
    layer0_outputs(2194) <= (inputs(89)) and not (inputs(150));
    layer0_outputs(2195) <= inputs(109);
    layer0_outputs(2196) <= '0';
    layer0_outputs(2197) <= not(inputs(195)) or (inputs(108));
    layer0_outputs(2198) <= (inputs(116)) or (inputs(252));
    layer0_outputs(2199) <= not(inputs(176)) or (inputs(255));
    layer0_outputs(2200) <= (inputs(108)) and not (inputs(234));
    layer0_outputs(2201) <= not(inputs(149)) or (inputs(46));
    layer0_outputs(2202) <= not(inputs(147));
    layer0_outputs(2203) <= (inputs(94)) or (inputs(147));
    layer0_outputs(2204) <= not((inputs(159)) or (inputs(163)));
    layer0_outputs(2205) <= (inputs(198)) and not (inputs(223));
    layer0_outputs(2206) <= not(inputs(27));
    layer0_outputs(2207) <= (inputs(6)) or (inputs(52));
    layer0_outputs(2208) <= not(inputs(231)) or (inputs(184));
    layer0_outputs(2209) <= inputs(181);
    layer0_outputs(2210) <= not(inputs(245));
    layer0_outputs(2211) <= (inputs(244)) or (inputs(181));
    layer0_outputs(2212) <= (inputs(227)) and not (inputs(105));
    layer0_outputs(2213) <= (inputs(180)) or (inputs(52));
    layer0_outputs(2214) <= not(inputs(188));
    layer0_outputs(2215) <= (inputs(29)) or (inputs(20));
    layer0_outputs(2216) <= (inputs(129)) xor (inputs(126));
    layer0_outputs(2217) <= inputs(66);
    layer0_outputs(2218) <= inputs(181);
    layer0_outputs(2219) <= (inputs(36)) and not (inputs(120));
    layer0_outputs(2220) <= inputs(116);
    layer0_outputs(2221) <= not(inputs(104));
    layer0_outputs(2222) <= (inputs(115)) or (inputs(52));
    layer0_outputs(2223) <= not(inputs(229));
    layer0_outputs(2224) <= inputs(178);
    layer0_outputs(2225) <= not((inputs(16)) and (inputs(244)));
    layer0_outputs(2226) <= not(inputs(131)) or (inputs(193));
    layer0_outputs(2227) <= not(inputs(37));
    layer0_outputs(2228) <= inputs(172);
    layer0_outputs(2229) <= (inputs(42)) and not (inputs(128));
    layer0_outputs(2230) <= inputs(162);
    layer0_outputs(2231) <= not(inputs(23)) or (inputs(146));
    layer0_outputs(2232) <= '0';
    layer0_outputs(2233) <= not(inputs(220));
    layer0_outputs(2234) <= not(inputs(248));
    layer0_outputs(2235) <= not(inputs(122));
    layer0_outputs(2236) <= (inputs(2)) xor (inputs(128));
    layer0_outputs(2237) <= inputs(244);
    layer0_outputs(2238) <= not(inputs(219));
    layer0_outputs(2239) <= not(inputs(65));
    layer0_outputs(2240) <= inputs(197);
    layer0_outputs(2241) <= not(inputs(119)) or (inputs(160));
    layer0_outputs(2242) <= inputs(32);
    layer0_outputs(2243) <= not((inputs(4)) or (inputs(155)));
    layer0_outputs(2244) <= not(inputs(110));
    layer0_outputs(2245) <= inputs(105);
    layer0_outputs(2246) <= inputs(199);
    layer0_outputs(2247) <= not(inputs(24));
    layer0_outputs(2248) <= not((inputs(86)) or (inputs(69)));
    layer0_outputs(2249) <= (inputs(123)) or (inputs(211));
    layer0_outputs(2250) <= not((inputs(18)) or (inputs(243)));
    layer0_outputs(2251) <= not((inputs(112)) or (inputs(176)));
    layer0_outputs(2252) <= (inputs(22)) or (inputs(125));
    layer0_outputs(2253) <= (inputs(75)) and not (inputs(252));
    layer0_outputs(2254) <= (inputs(113)) or (inputs(115));
    layer0_outputs(2255) <= not((inputs(55)) or (inputs(155)));
    layer0_outputs(2256) <= not(inputs(183)) or (inputs(156));
    layer0_outputs(2257) <= (inputs(28)) and not (inputs(10));
    layer0_outputs(2258) <= not((inputs(54)) xor (inputs(132)));
    layer0_outputs(2259) <= not(inputs(146));
    layer0_outputs(2260) <= (inputs(250)) or (inputs(49));
    layer0_outputs(2261) <= inputs(25);
    layer0_outputs(2262) <= inputs(104);
    layer0_outputs(2263) <= inputs(117);
    layer0_outputs(2264) <= inputs(151);
    layer0_outputs(2265) <= not(inputs(228));
    layer0_outputs(2266) <= (inputs(8)) or (inputs(143));
    layer0_outputs(2267) <= (inputs(23)) and not (inputs(238));
    layer0_outputs(2268) <= '1';
    layer0_outputs(2269) <= (inputs(227)) or (inputs(208));
    layer0_outputs(2270) <= not(inputs(176));
    layer0_outputs(2271) <= (inputs(153)) or (inputs(126));
    layer0_outputs(2272) <= (inputs(189)) or (inputs(209));
    layer0_outputs(2273) <= (inputs(241)) or (inputs(121));
    layer0_outputs(2274) <= (inputs(233)) or (inputs(114));
    layer0_outputs(2275) <= inputs(44);
    layer0_outputs(2276) <= not(inputs(76));
    layer0_outputs(2277) <= not(inputs(65)) or (inputs(31));
    layer0_outputs(2278) <= not(inputs(170));
    layer0_outputs(2279) <= '1';
    layer0_outputs(2280) <= (inputs(44)) and not (inputs(175));
    layer0_outputs(2281) <= not((inputs(41)) or (inputs(15)));
    layer0_outputs(2282) <= not(inputs(97));
    layer0_outputs(2283) <= not((inputs(183)) or (inputs(198)));
    layer0_outputs(2284) <= (inputs(194)) or (inputs(6));
    layer0_outputs(2285) <= (inputs(226)) or (inputs(128));
    layer0_outputs(2286) <= not(inputs(132));
    layer0_outputs(2287) <= not((inputs(54)) or (inputs(129)));
    layer0_outputs(2288) <= not(inputs(83));
    layer0_outputs(2289) <= inputs(2);
    layer0_outputs(2290) <= not((inputs(186)) or (inputs(215)));
    layer0_outputs(2291) <= inputs(218);
    layer0_outputs(2292) <= not((inputs(88)) xor (inputs(41)));
    layer0_outputs(2293) <= (inputs(136)) and not (inputs(52));
    layer0_outputs(2294) <= not((inputs(99)) or (inputs(170)));
    layer0_outputs(2295) <= not((inputs(244)) or (inputs(11)));
    layer0_outputs(2296) <= not((inputs(157)) or (inputs(43)));
    layer0_outputs(2297) <= not((inputs(222)) or (inputs(218)));
    layer0_outputs(2298) <= (inputs(92)) and not (inputs(1));
    layer0_outputs(2299) <= inputs(224);
    layer0_outputs(2300) <= not((inputs(8)) or (inputs(10)));
    layer0_outputs(2301) <= not(inputs(44)) or (inputs(254));
    layer0_outputs(2302) <= not((inputs(241)) or (inputs(95)));
    layer0_outputs(2303) <= inputs(125);
    layer0_outputs(2304) <= not((inputs(202)) or (inputs(122)));
    layer0_outputs(2305) <= not((inputs(197)) xor (inputs(60)));
    layer0_outputs(2306) <= not((inputs(130)) or (inputs(67)));
    layer0_outputs(2307) <= (inputs(100)) xor (inputs(129));
    layer0_outputs(2308) <= (inputs(53)) or (inputs(51));
    layer0_outputs(2309) <= (inputs(5)) xor (inputs(78));
    layer0_outputs(2310) <= inputs(101);
    layer0_outputs(2311) <= inputs(180);
    layer0_outputs(2312) <= inputs(124);
    layer0_outputs(2313) <= not(inputs(8));
    layer0_outputs(2314) <= (inputs(152)) and not (inputs(113));
    layer0_outputs(2315) <= (inputs(87)) and not (inputs(255));
    layer0_outputs(2316) <= not(inputs(29));
    layer0_outputs(2317) <= not(inputs(148));
    layer0_outputs(2318) <= not(inputs(245));
    layer0_outputs(2319) <= not(inputs(244)) or (inputs(144));
    layer0_outputs(2320) <= not((inputs(88)) or (inputs(177)));
    layer0_outputs(2321) <= not(inputs(157));
    layer0_outputs(2322) <= inputs(48);
    layer0_outputs(2323) <= '0';
    layer0_outputs(2324) <= not(inputs(217));
    layer0_outputs(2325) <= inputs(229);
    layer0_outputs(2326) <= (inputs(134)) and not (inputs(2));
    layer0_outputs(2327) <= not(inputs(75));
    layer0_outputs(2328) <= inputs(130);
    layer0_outputs(2329) <= (inputs(235)) or (inputs(131));
    layer0_outputs(2330) <= not(inputs(246)) or (inputs(206));
    layer0_outputs(2331) <= not(inputs(163)) or (inputs(175));
    layer0_outputs(2332) <= not(inputs(57)) or (inputs(19));
    layer0_outputs(2333) <= (inputs(7)) and not (inputs(128));
    layer0_outputs(2334) <= not(inputs(73));
    layer0_outputs(2335) <= (inputs(235)) and not (inputs(10));
    layer0_outputs(2336) <= (inputs(196)) or (inputs(140));
    layer0_outputs(2337) <= not(inputs(120));
    layer0_outputs(2338) <= inputs(82);
    layer0_outputs(2339) <= (inputs(18)) or (inputs(58));
    layer0_outputs(2340) <= (inputs(233)) and not (inputs(199));
    layer0_outputs(2341) <= inputs(75);
    layer0_outputs(2342) <= not((inputs(210)) or (inputs(0)));
    layer0_outputs(2343) <= (inputs(248)) or (inputs(128));
    layer0_outputs(2344) <= not(inputs(15));
    layer0_outputs(2345) <= (inputs(89)) or (inputs(181));
    layer0_outputs(2346) <= inputs(160);
    layer0_outputs(2347) <= not(inputs(231));
    layer0_outputs(2348) <= not((inputs(99)) or (inputs(116)));
    layer0_outputs(2349) <= not(inputs(200));
    layer0_outputs(2350) <= (inputs(204)) and not (inputs(1));
    layer0_outputs(2351) <= inputs(181);
    layer0_outputs(2352) <= not(inputs(75));
    layer0_outputs(2353) <= (inputs(129)) or (inputs(130));
    layer0_outputs(2354) <= not(inputs(111));
    layer0_outputs(2355) <= not(inputs(136)) or (inputs(207));
    layer0_outputs(2356) <= not(inputs(25));
    layer0_outputs(2357) <= (inputs(150)) or (inputs(98));
    layer0_outputs(2358) <= not(inputs(22)) or (inputs(245));
    layer0_outputs(2359) <= inputs(223);
    layer0_outputs(2360) <= (inputs(187)) or (inputs(175));
    layer0_outputs(2361) <= (inputs(133)) or (inputs(208));
    layer0_outputs(2362) <= inputs(137);
    layer0_outputs(2363) <= not(inputs(136));
    layer0_outputs(2364) <= not((inputs(179)) or (inputs(95)));
    layer0_outputs(2365) <= inputs(149);
    layer0_outputs(2366) <= not(inputs(140));
    layer0_outputs(2367) <= (inputs(113)) or (inputs(5));
    layer0_outputs(2368) <= inputs(9);
    layer0_outputs(2369) <= not((inputs(176)) or (inputs(132)));
    layer0_outputs(2370) <= inputs(210);
    layer0_outputs(2371) <= not(inputs(120));
    layer0_outputs(2372) <= not(inputs(92));
    layer0_outputs(2373) <= not(inputs(215));
    layer0_outputs(2374) <= not(inputs(182));
    layer0_outputs(2375) <= inputs(179);
    layer0_outputs(2376) <= not(inputs(72)) or (inputs(117));
    layer0_outputs(2377) <= not(inputs(212));
    layer0_outputs(2378) <= not((inputs(47)) or (inputs(233)));
    layer0_outputs(2379) <= (inputs(89)) and not (inputs(14));
    layer0_outputs(2380) <= (inputs(88)) and not (inputs(145));
    layer0_outputs(2381) <= inputs(149);
    layer0_outputs(2382) <= not((inputs(215)) or (inputs(198)));
    layer0_outputs(2383) <= inputs(209);
    layer0_outputs(2384) <= (inputs(47)) or (inputs(218));
    layer0_outputs(2385) <= not(inputs(22)) or (inputs(150));
    layer0_outputs(2386) <= not((inputs(192)) xor (inputs(207)));
    layer0_outputs(2387) <= (inputs(164)) or (inputs(210));
    layer0_outputs(2388) <= not(inputs(251)) or (inputs(206));
    layer0_outputs(2389) <= (inputs(5)) or (inputs(90));
    layer0_outputs(2390) <= not((inputs(197)) xor (inputs(212)));
    layer0_outputs(2391) <= not((inputs(82)) or (inputs(160)));
    layer0_outputs(2392) <= not(inputs(196));
    layer0_outputs(2393) <= not(inputs(185)) or (inputs(89));
    layer0_outputs(2394) <= not(inputs(146));
    layer0_outputs(2395) <= not(inputs(6)) or (inputs(1));
    layer0_outputs(2396) <= (inputs(202)) and not (inputs(127));
    layer0_outputs(2397) <= inputs(104);
    layer0_outputs(2398) <= not((inputs(8)) xor (inputs(1)));
    layer0_outputs(2399) <= not((inputs(77)) or (inputs(106)));
    layer0_outputs(2400) <= not(inputs(138));
    layer0_outputs(2401) <= not((inputs(74)) or (inputs(78)));
    layer0_outputs(2402) <= not(inputs(254));
    layer0_outputs(2403) <= not((inputs(227)) or (inputs(224)));
    layer0_outputs(2404) <= (inputs(76)) or (inputs(45));
    layer0_outputs(2405) <= not((inputs(3)) or (inputs(221)));
    layer0_outputs(2406) <= inputs(1);
    layer0_outputs(2407) <= inputs(139);
    layer0_outputs(2408) <= not((inputs(145)) or (inputs(172)));
    layer0_outputs(2409) <= not(inputs(228));
    layer0_outputs(2410) <= (inputs(47)) and not (inputs(111));
    layer0_outputs(2411) <= not(inputs(133)) or (inputs(196));
    layer0_outputs(2412) <= inputs(193);
    layer0_outputs(2413) <= not(inputs(71));
    layer0_outputs(2414) <= not((inputs(69)) or (inputs(21)));
    layer0_outputs(2415) <= (inputs(9)) xor (inputs(11));
    layer0_outputs(2416) <= not((inputs(213)) or (inputs(62)));
    layer0_outputs(2417) <= (inputs(237)) xor (inputs(173));
    layer0_outputs(2418) <= not((inputs(236)) or (inputs(136)));
    layer0_outputs(2419) <= not(inputs(85));
    layer0_outputs(2420) <= inputs(116);
    layer0_outputs(2421) <= inputs(163);
    layer0_outputs(2422) <= not(inputs(163));
    layer0_outputs(2423) <= not(inputs(154)) or (inputs(6));
    layer0_outputs(2424) <= not(inputs(94)) or (inputs(94));
    layer0_outputs(2425) <= not(inputs(40)) or (inputs(202));
    layer0_outputs(2426) <= (inputs(7)) and not (inputs(158));
    layer0_outputs(2427) <= not((inputs(224)) or (inputs(150)));
    layer0_outputs(2428) <= inputs(91);
    layer0_outputs(2429) <= (inputs(194)) or (inputs(20));
    layer0_outputs(2430) <= inputs(214);
    layer0_outputs(2431) <= not((inputs(54)) or (inputs(197)));
    layer0_outputs(2432) <= not(inputs(234)) or (inputs(77));
    layer0_outputs(2433) <= not(inputs(219));
    layer0_outputs(2434) <= not(inputs(24));
    layer0_outputs(2435) <= not(inputs(90));
    layer0_outputs(2436) <= (inputs(237)) or (inputs(56));
    layer0_outputs(2437) <= (inputs(4)) or (inputs(211));
    layer0_outputs(2438) <= not(inputs(99)) or (inputs(241));
    layer0_outputs(2439) <= inputs(249);
    layer0_outputs(2440) <= (inputs(66)) or (inputs(29));
    layer0_outputs(2441) <= (inputs(199)) and not (inputs(59));
    layer0_outputs(2442) <= (inputs(0)) or (inputs(125));
    layer0_outputs(2443) <= '0';
    layer0_outputs(2444) <= inputs(106);
    layer0_outputs(2445) <= (inputs(221)) and not (inputs(49));
    layer0_outputs(2446) <= (inputs(107)) or (inputs(95));
    layer0_outputs(2447) <= not(inputs(230));
    layer0_outputs(2448) <= '0';
    layer0_outputs(2449) <= (inputs(93)) or (inputs(145));
    layer0_outputs(2450) <= not(inputs(201)) or (inputs(49));
    layer0_outputs(2451) <= '1';
    layer0_outputs(2452) <= inputs(119);
    layer0_outputs(2453) <= '0';
    layer0_outputs(2454) <= (inputs(110)) or (inputs(142));
    layer0_outputs(2455) <= not((inputs(200)) or (inputs(161)));
    layer0_outputs(2456) <= inputs(165);
    layer0_outputs(2457) <= inputs(18);
    layer0_outputs(2458) <= not((inputs(1)) or (inputs(3)));
    layer0_outputs(2459) <= (inputs(23)) and not (inputs(229));
    layer0_outputs(2460) <= inputs(144);
    layer0_outputs(2461) <= (inputs(125)) xor (inputs(140));
    layer0_outputs(2462) <= (inputs(238)) or (inputs(109));
    layer0_outputs(2463) <= inputs(86);
    layer0_outputs(2464) <= (inputs(47)) xor (inputs(48));
    layer0_outputs(2465) <= (inputs(58)) and (inputs(143));
    layer0_outputs(2466) <= not((inputs(252)) xor (inputs(203)));
    layer0_outputs(2467) <= (inputs(162)) and not (inputs(153));
    layer0_outputs(2468) <= '1';
    layer0_outputs(2469) <= (inputs(38)) or (inputs(181));
    layer0_outputs(2470) <= inputs(92);
    layer0_outputs(2471) <= (inputs(220)) or (inputs(181));
    layer0_outputs(2472) <= not(inputs(149));
    layer0_outputs(2473) <= not(inputs(172));
    layer0_outputs(2474) <= not((inputs(0)) and (inputs(40)));
    layer0_outputs(2475) <= not(inputs(43)) or (inputs(251));
    layer0_outputs(2476) <= not(inputs(247));
    layer0_outputs(2477) <= (inputs(231)) and not (inputs(206));
    layer0_outputs(2478) <= not((inputs(6)) or (inputs(28)));
    layer0_outputs(2479) <= inputs(108);
    layer0_outputs(2480) <= (inputs(252)) or (inputs(93));
    layer0_outputs(2481) <= inputs(219);
    layer0_outputs(2482) <= not(inputs(226)) or (inputs(175));
    layer0_outputs(2483) <= (inputs(57)) or (inputs(184));
    layer0_outputs(2484) <= (inputs(128)) or (inputs(252));
    layer0_outputs(2485) <= inputs(92);
    layer0_outputs(2486) <= (inputs(134)) and not (inputs(2));
    layer0_outputs(2487) <= (inputs(96)) or (inputs(237));
    layer0_outputs(2488) <= inputs(178);
    layer0_outputs(2489) <= (inputs(60)) or (inputs(114));
    layer0_outputs(2490) <= inputs(164);
    layer0_outputs(2491) <= '0';
    layer0_outputs(2492) <= not(inputs(40));
    layer0_outputs(2493) <= not(inputs(189)) or (inputs(12));
    layer0_outputs(2494) <= inputs(173);
    layer0_outputs(2495) <= not((inputs(138)) xor (inputs(200)));
    layer0_outputs(2496) <= inputs(212);
    layer0_outputs(2497) <= inputs(151);
    layer0_outputs(2498) <= inputs(103);
    layer0_outputs(2499) <= (inputs(181)) or (inputs(208));
    layer0_outputs(2500) <= (inputs(17)) or (inputs(52));
    layer0_outputs(2501) <= inputs(126);
    layer0_outputs(2502) <= inputs(186);
    layer0_outputs(2503) <= not((inputs(185)) or (inputs(132)));
    layer0_outputs(2504) <= inputs(178);
    layer0_outputs(2505) <= (inputs(165)) or (inputs(221));
    layer0_outputs(2506) <= (inputs(210)) or (inputs(129));
    layer0_outputs(2507) <= not(inputs(16));
    layer0_outputs(2508) <= (inputs(234)) or (inputs(144));
    layer0_outputs(2509) <= not((inputs(83)) or (inputs(131)));
    layer0_outputs(2510) <= not((inputs(117)) or (inputs(178)));
    layer0_outputs(2511) <= not(inputs(214));
    layer0_outputs(2512) <= not(inputs(182)) or (inputs(128));
    layer0_outputs(2513) <= not((inputs(17)) and (inputs(236)));
    layer0_outputs(2514) <= not((inputs(211)) or (inputs(193)));
    layer0_outputs(2515) <= (inputs(223)) or (inputs(120));
    layer0_outputs(2516) <= not(inputs(210)) or (inputs(144));
    layer0_outputs(2517) <= (inputs(209)) or (inputs(50));
    layer0_outputs(2518) <= not((inputs(212)) or (inputs(211)));
    layer0_outputs(2519) <= inputs(166);
    layer0_outputs(2520) <= not(inputs(181));
    layer0_outputs(2521) <= not(inputs(30));
    layer0_outputs(2522) <= inputs(42);
    layer0_outputs(2523) <= not(inputs(25));
    layer0_outputs(2524) <= not((inputs(225)) or (inputs(64)));
    layer0_outputs(2525) <= not(inputs(25));
    layer0_outputs(2526) <= inputs(67);
    layer0_outputs(2527) <= not(inputs(38));
    layer0_outputs(2528) <= not(inputs(38)) or (inputs(204));
    layer0_outputs(2529) <= not(inputs(9));
    layer0_outputs(2530) <= (inputs(22)) or (inputs(225));
    layer0_outputs(2531) <= not((inputs(135)) or (inputs(49)));
    layer0_outputs(2532) <= (inputs(118)) and not (inputs(254));
    layer0_outputs(2533) <= '0';
    layer0_outputs(2534) <= not((inputs(154)) or (inputs(131)));
    layer0_outputs(2535) <= not(inputs(129)) or (inputs(236));
    layer0_outputs(2536) <= not(inputs(223)) or (inputs(157));
    layer0_outputs(2537) <= (inputs(102)) and (inputs(45));
    layer0_outputs(2538) <= inputs(244);
    layer0_outputs(2539) <= not(inputs(179));
    layer0_outputs(2540) <= not(inputs(136));
    layer0_outputs(2541) <= (inputs(34)) or (inputs(227));
    layer0_outputs(2542) <= not((inputs(226)) or (inputs(13)));
    layer0_outputs(2543) <= (inputs(164)) and not (inputs(0));
    layer0_outputs(2544) <= (inputs(61)) and not (inputs(237));
    layer0_outputs(2545) <= not(inputs(169));
    layer0_outputs(2546) <= (inputs(109)) or (inputs(20));
    layer0_outputs(2547) <= (inputs(146)) or (inputs(54));
    layer0_outputs(2548) <= inputs(112);
    layer0_outputs(2549) <= not((inputs(3)) and (inputs(87)));
    layer0_outputs(2550) <= '1';
    layer0_outputs(2551) <= not(inputs(134)) or (inputs(166));
    layer0_outputs(2552) <= (inputs(167)) or (inputs(164));
    layer0_outputs(2553) <= (inputs(19)) or (inputs(238));
    layer0_outputs(2554) <= (inputs(208)) and not (inputs(61));
    layer0_outputs(2555) <= inputs(204);
    layer0_outputs(2556) <= not(inputs(56)) or (inputs(222));
    layer0_outputs(2557) <= (inputs(188)) and not (inputs(79));
    layer0_outputs(2558) <= not(inputs(95)) or (inputs(0));
    layer0_outputs(2559) <= (inputs(150)) or (inputs(252));
    outputs(0) <= layer0_outputs(2034);
    outputs(1) <= not(layer0_outputs(2075));
    outputs(2) <= not((layer0_outputs(2242)) or (layer0_outputs(892)));
    outputs(3) <= layer0_outputs(1808);
    outputs(4) <= not(layer0_outputs(144)) or (layer0_outputs(1062));
    outputs(5) <= not((layer0_outputs(1879)) xor (layer0_outputs(585)));
    outputs(6) <= not(layer0_outputs(2515));
    outputs(7) <= not((layer0_outputs(2071)) or (layer0_outputs(507)));
    outputs(8) <= not(layer0_outputs(1174));
    outputs(9) <= (layer0_outputs(1192)) or (layer0_outputs(476));
    outputs(10) <= (layer0_outputs(201)) and not (layer0_outputs(2095));
    outputs(11) <= layer0_outputs(2298);
    outputs(12) <= not((layer0_outputs(1290)) or (layer0_outputs(364)));
    outputs(13) <= not((layer0_outputs(1351)) xor (layer0_outputs(1508)));
    outputs(14) <= layer0_outputs(2130);
    outputs(15) <= not(layer0_outputs(355));
    outputs(16) <= layer0_outputs(1429);
    outputs(17) <= layer0_outputs(1658);
    outputs(18) <= (layer0_outputs(1402)) and not (layer0_outputs(173));
    outputs(19) <= not(layer0_outputs(2332));
    outputs(20) <= layer0_outputs(915);
    outputs(21) <= not(layer0_outputs(1099));
    outputs(22) <= (layer0_outputs(582)) and not (layer0_outputs(157));
    outputs(23) <= (layer0_outputs(1196)) and not (layer0_outputs(2138));
    outputs(24) <= not(layer0_outputs(286));
    outputs(25) <= layer0_outputs(1357);
    outputs(26) <= (layer0_outputs(394)) xor (layer0_outputs(864));
    outputs(27) <= layer0_outputs(941);
    outputs(28) <= not(layer0_outputs(504)) or (layer0_outputs(1971));
    outputs(29) <= (layer0_outputs(281)) xor (layer0_outputs(1657));
    outputs(30) <= not(layer0_outputs(273));
    outputs(31) <= layer0_outputs(1204);
    outputs(32) <= (layer0_outputs(1151)) and (layer0_outputs(1275));
    outputs(33) <= not((layer0_outputs(1756)) and (layer0_outputs(1435)));
    outputs(34) <= (layer0_outputs(68)) and (layer0_outputs(632));
    outputs(35) <= layer0_outputs(1711);
    outputs(36) <= layer0_outputs(1782);
    outputs(37) <= (layer0_outputs(2388)) and (layer0_outputs(1185));
    outputs(38) <= not(layer0_outputs(21));
    outputs(39) <= (layer0_outputs(1469)) and not (layer0_outputs(847));
    outputs(40) <= layer0_outputs(581);
    outputs(41) <= not(layer0_outputs(82));
    outputs(42) <= not((layer0_outputs(26)) and (layer0_outputs(1534)));
    outputs(43) <= (layer0_outputs(2254)) and not (layer0_outputs(2122));
    outputs(44) <= (layer0_outputs(401)) and (layer0_outputs(486));
    outputs(45) <= not(layer0_outputs(3)) or (layer0_outputs(2298));
    outputs(46) <= (layer0_outputs(1395)) and (layer0_outputs(2449));
    outputs(47) <= not(layer0_outputs(538));
    outputs(48) <= layer0_outputs(605);
    outputs(49) <= layer0_outputs(661);
    outputs(50) <= (layer0_outputs(253)) and (layer0_outputs(1038));
    outputs(51) <= layer0_outputs(87);
    outputs(52) <= layer0_outputs(1880);
    outputs(53) <= layer0_outputs(329);
    outputs(54) <= layer0_outputs(1318);
    outputs(55) <= (layer0_outputs(1608)) or (layer0_outputs(1118));
    outputs(56) <= not((layer0_outputs(1199)) xor (layer0_outputs(2277)));
    outputs(57) <= not((layer0_outputs(1358)) or (layer0_outputs(911)));
    outputs(58) <= (layer0_outputs(499)) xor (layer0_outputs(2344));
    outputs(59) <= (layer0_outputs(2006)) and (layer0_outputs(275));
    outputs(60) <= layer0_outputs(299);
    outputs(61) <= not((layer0_outputs(1626)) or (layer0_outputs(493)));
    outputs(62) <= (layer0_outputs(965)) and not (layer0_outputs(200));
    outputs(63) <= (layer0_outputs(706)) and not (layer0_outputs(1676));
    outputs(64) <= not(layer0_outputs(808));
    outputs(65) <= (layer0_outputs(126)) and not (layer0_outputs(81));
    outputs(66) <= layer0_outputs(1600);
    outputs(67) <= not(layer0_outputs(1876));
    outputs(68) <= layer0_outputs(834);
    outputs(69) <= layer0_outputs(1609);
    outputs(70) <= not(layer0_outputs(116));
    outputs(71) <= (layer0_outputs(1955)) xor (layer0_outputs(469));
    outputs(72) <= (layer0_outputs(647)) xor (layer0_outputs(2148));
    outputs(73) <= layer0_outputs(243);
    outputs(74) <= (layer0_outputs(1659)) or (layer0_outputs(617));
    outputs(75) <= not(layer0_outputs(1005));
    outputs(76) <= not((layer0_outputs(217)) and (layer0_outputs(1420)));
    outputs(77) <= (layer0_outputs(45)) or (layer0_outputs(2168));
    outputs(78) <= layer0_outputs(1990);
    outputs(79) <= (layer0_outputs(1908)) or (layer0_outputs(2346));
    outputs(80) <= not(layer0_outputs(2265));
    outputs(81) <= not(layer0_outputs(534));
    outputs(82) <= layer0_outputs(2496);
    outputs(83) <= layer0_outputs(1614);
    outputs(84) <= layer0_outputs(1671);
    outputs(85) <= (layer0_outputs(483)) and not (layer0_outputs(1668));
    outputs(86) <= not((layer0_outputs(1326)) xor (layer0_outputs(1186)));
    outputs(87) <= layer0_outputs(1125);
    outputs(88) <= layer0_outputs(1915);
    outputs(89) <= layer0_outputs(391);
    outputs(90) <= layer0_outputs(1180);
    outputs(91) <= not(layer0_outputs(2248));
    outputs(92) <= not(layer0_outputs(2386)) or (layer0_outputs(2086));
    outputs(93) <= (layer0_outputs(1973)) and (layer0_outputs(1595));
    outputs(94) <= layer0_outputs(2325);
    outputs(95) <= layer0_outputs(791);
    outputs(96) <= layer0_outputs(1918);
    outputs(97) <= layer0_outputs(2212);
    outputs(98) <= not((layer0_outputs(1948)) and (layer0_outputs(872)));
    outputs(99) <= (layer0_outputs(1373)) and not (layer0_outputs(182));
    outputs(100) <= not(layer0_outputs(980));
    outputs(101) <= (layer0_outputs(235)) or (layer0_outputs(1998));
    outputs(102) <= layer0_outputs(2195);
    outputs(103) <= not(layer0_outputs(117)) or (layer0_outputs(863));
    outputs(104) <= not(layer0_outputs(1499));
    outputs(105) <= not((layer0_outputs(1714)) and (layer0_outputs(59)));
    outputs(106) <= not(layer0_outputs(705)) or (layer0_outputs(1813));
    outputs(107) <= not(layer0_outputs(751));
    outputs(108) <= (layer0_outputs(2035)) and not (layer0_outputs(1227));
    outputs(109) <= (layer0_outputs(2531)) and not (layer0_outputs(1457));
    outputs(110) <= (layer0_outputs(135)) or (layer0_outputs(518));
    outputs(111) <= (layer0_outputs(2374)) and (layer0_outputs(1339));
    outputs(112) <= layer0_outputs(2522);
    outputs(113) <= not(layer0_outputs(454));
    outputs(114) <= layer0_outputs(1189);
    outputs(115) <= layer0_outputs(586);
    outputs(116) <= not((layer0_outputs(422)) or (layer0_outputs(2015)));
    outputs(117) <= layer0_outputs(1836);
    outputs(118) <= not(layer0_outputs(1306)) or (layer0_outputs(408));
    outputs(119) <= not(layer0_outputs(624));
    outputs(120) <= not(layer0_outputs(1820));
    outputs(121) <= not(layer0_outputs(2085));
    outputs(122) <= (layer0_outputs(1446)) and not (layer0_outputs(742));
    outputs(123) <= not((layer0_outputs(756)) and (layer0_outputs(59)));
    outputs(124) <= not(layer0_outputs(285));
    outputs(125) <= not(layer0_outputs(813)) or (layer0_outputs(255));
    outputs(126) <= (layer0_outputs(533)) and (layer0_outputs(788));
    outputs(127) <= not((layer0_outputs(2146)) or (layer0_outputs(742)));
    outputs(128) <= layer0_outputs(2130);
    outputs(129) <= not(layer0_outputs(2085)) or (layer0_outputs(24));
    outputs(130) <= not((layer0_outputs(1909)) or (layer0_outputs(1166)));
    outputs(131) <= not((layer0_outputs(2023)) and (layer0_outputs(1727)));
    outputs(132) <= (layer0_outputs(940)) or (layer0_outputs(288));
    outputs(133) <= layer0_outputs(1252);
    outputs(134) <= not(layer0_outputs(503));
    outputs(135) <= (layer0_outputs(2418)) and not (layer0_outputs(376));
    outputs(136) <= layer0_outputs(63);
    outputs(137) <= (layer0_outputs(764)) or (layer0_outputs(1208));
    outputs(138) <= not(layer0_outputs(1594));
    outputs(139) <= not((layer0_outputs(2199)) and (layer0_outputs(2204)));
    outputs(140) <= (layer0_outputs(1462)) or (layer0_outputs(635));
    outputs(141) <= (layer0_outputs(1702)) and not (layer0_outputs(895));
    outputs(142) <= not(layer0_outputs(1403)) or (layer0_outputs(1897));
    outputs(143) <= (layer0_outputs(833)) or (layer0_outputs(1608));
    outputs(144) <= not(layer0_outputs(1389));
    outputs(145) <= not((layer0_outputs(128)) or (layer0_outputs(1149)));
    outputs(146) <= not(layer0_outputs(1840));
    outputs(147) <= not(layer0_outputs(300));
    outputs(148) <= layer0_outputs(391);
    outputs(149) <= layer0_outputs(1215);
    outputs(150) <= (layer0_outputs(540)) and not (layer0_outputs(1245));
    outputs(151) <= (layer0_outputs(2008)) xor (layer0_outputs(1015));
    outputs(152) <= layer0_outputs(1804);
    outputs(153) <= layer0_outputs(1978);
    outputs(154) <= not(layer0_outputs(1133));
    outputs(155) <= not((layer0_outputs(130)) and (layer0_outputs(2330)));
    outputs(156) <= not(layer0_outputs(1104));
    outputs(157) <= (layer0_outputs(240)) and not (layer0_outputs(223));
    outputs(158) <= not(layer0_outputs(2015));
    outputs(159) <= not(layer0_outputs(358));
    outputs(160) <= not((layer0_outputs(367)) and (layer0_outputs(65)));
    outputs(161) <= not((layer0_outputs(2362)) or (layer0_outputs(1418)));
    outputs(162) <= not(layer0_outputs(1343)) or (layer0_outputs(69));
    outputs(163) <= layer0_outputs(1843);
    outputs(164) <= (layer0_outputs(802)) or (layer0_outputs(1774));
    outputs(165) <= not(layer0_outputs(2345));
    outputs(166) <= not(layer0_outputs(727)) or (layer0_outputs(947));
    outputs(167) <= layer0_outputs(515);
    outputs(168) <= not((layer0_outputs(2459)) or (layer0_outputs(2365)));
    outputs(169) <= not(layer0_outputs(1008));
    outputs(170) <= layer0_outputs(717);
    outputs(171) <= (layer0_outputs(2488)) or (layer0_outputs(2055));
    outputs(172) <= not(layer0_outputs(2372));
    outputs(173) <= (layer0_outputs(1092)) and not (layer0_outputs(2322));
    outputs(174) <= layer0_outputs(1802);
    outputs(175) <= not(layer0_outputs(1827));
    outputs(176) <= not(layer0_outputs(1557)) or (layer0_outputs(1019));
    outputs(177) <= layer0_outputs(2547);
    outputs(178) <= layer0_outputs(275);
    outputs(179) <= not(layer0_outputs(618));
    outputs(180) <= layer0_outputs(834);
    outputs(181) <= not((layer0_outputs(440)) or (layer0_outputs(115)));
    outputs(182) <= not(layer0_outputs(1152));
    outputs(183) <= not(layer0_outputs(726));
    outputs(184) <= not(layer0_outputs(215));
    outputs(185) <= layer0_outputs(2540);
    outputs(186) <= (layer0_outputs(234)) and not (layer0_outputs(2475));
    outputs(187) <= layer0_outputs(1446);
    outputs(188) <= (layer0_outputs(2142)) and (layer0_outputs(674));
    outputs(189) <= not(layer0_outputs(1439)) or (layer0_outputs(1910));
    outputs(190) <= not(layer0_outputs(1262)) or (layer0_outputs(688));
    outputs(191) <= (layer0_outputs(909)) xor (layer0_outputs(907));
    outputs(192) <= (layer0_outputs(1257)) or (layer0_outputs(1831));
    outputs(193) <= not(layer0_outputs(704));
    outputs(194) <= (layer0_outputs(972)) and not (layer0_outputs(3));
    outputs(195) <= not(layer0_outputs(74)) or (layer0_outputs(2267));
    outputs(196) <= layer0_outputs(2253);
    outputs(197) <= not(layer0_outputs(1364)) or (layer0_outputs(2316));
    outputs(198) <= not(layer0_outputs(989));
    outputs(199) <= not(layer0_outputs(1956));
    outputs(200) <= layer0_outputs(1344);
    outputs(201) <= layer0_outputs(536);
    outputs(202) <= not(layer0_outputs(703)) or (layer0_outputs(451));
    outputs(203) <= not(layer0_outputs(918)) or (layer0_outputs(1558));
    outputs(204) <= layer0_outputs(1535);
    outputs(205) <= not(layer0_outputs(273));
    outputs(206) <= not(layer0_outputs(587));
    outputs(207) <= not((layer0_outputs(792)) or (layer0_outputs(1089)));
    outputs(208) <= (layer0_outputs(1360)) and not (layer0_outputs(2014));
    outputs(209) <= layer0_outputs(2545);
    outputs(210) <= not((layer0_outputs(924)) or (layer0_outputs(2182)));
    outputs(211) <= (layer0_outputs(1170)) or (layer0_outputs(745));
    outputs(212) <= layer0_outputs(1984);
    outputs(213) <= (layer0_outputs(54)) xor (layer0_outputs(233));
    outputs(214) <= not(layer0_outputs(2137)) or (layer0_outputs(1856));
    outputs(215) <= not(layer0_outputs(1322)) or (layer0_outputs(1103));
    outputs(216) <= not(layer0_outputs(346));
    outputs(217) <= layer0_outputs(111);
    outputs(218) <= not(layer0_outputs(1586));
    outputs(219) <= layer0_outputs(1762);
    outputs(220) <= layer0_outputs(1894);
    outputs(221) <= not((layer0_outputs(206)) and (layer0_outputs(458)));
    outputs(222) <= (layer0_outputs(1984)) and not (layer0_outputs(992));
    outputs(223) <= (layer0_outputs(1580)) and (layer0_outputs(1271));
    outputs(224) <= not(layer0_outputs(785));
    outputs(225) <= (layer0_outputs(2004)) and not (layer0_outputs(1670));
    outputs(226) <= (layer0_outputs(105)) or (layer0_outputs(1561));
    outputs(227) <= not((layer0_outputs(1521)) or (layer0_outputs(1003)));
    outputs(228) <= not(layer0_outputs(1492));
    outputs(229) <= not(layer0_outputs(162)) or (layer0_outputs(1524));
    outputs(230) <= (layer0_outputs(252)) and not (layer0_outputs(2289));
    outputs(231) <= layer0_outputs(403);
    outputs(232) <= not(layer0_outputs(1694));
    outputs(233) <= not(layer0_outputs(1443));
    outputs(234) <= (layer0_outputs(775)) or (layer0_outputs(2449));
    outputs(235) <= (layer0_outputs(2266)) and not (layer0_outputs(1932));
    outputs(236) <= layer0_outputs(1012);
    outputs(237) <= layer0_outputs(372);
    outputs(238) <= layer0_outputs(2221);
    outputs(239) <= layer0_outputs(1666);
    outputs(240) <= layer0_outputs(1050);
    outputs(241) <= (layer0_outputs(1416)) and not (layer0_outputs(756));
    outputs(242) <= not(layer0_outputs(2273));
    outputs(243) <= not(layer0_outputs(908)) or (layer0_outputs(1371));
    outputs(244) <= (layer0_outputs(771)) and not (layer0_outputs(1377));
    outputs(245) <= layer0_outputs(412);
    outputs(246) <= (layer0_outputs(1198)) or (layer0_outputs(1695));
    outputs(247) <= not(layer0_outputs(1415)) or (layer0_outputs(143));
    outputs(248) <= not(layer0_outputs(1437));
    outputs(249) <= layer0_outputs(2340);
    outputs(250) <= layer0_outputs(259);
    outputs(251) <= not((layer0_outputs(1665)) or (layer0_outputs(1696)));
    outputs(252) <= not(layer0_outputs(1964));
    outputs(253) <= not(layer0_outputs(2332)) or (layer0_outputs(2496));
    outputs(254) <= not(layer0_outputs(830));
    outputs(255) <= (layer0_outputs(2142)) and not (layer0_outputs(1555));
    outputs(256) <= '0';
    outputs(257) <= (layer0_outputs(1619)) and not (layer0_outputs(2557));
    outputs(258) <= (layer0_outputs(1559)) and (layer0_outputs(654));
    outputs(259) <= layer0_outputs(1470);
    outputs(260) <= (layer0_outputs(1757)) and not (layer0_outputs(2353));
    outputs(261) <= (layer0_outputs(1090)) and not (layer0_outputs(715));
    outputs(262) <= (layer0_outputs(2521)) and (layer0_outputs(261));
    outputs(263) <= (layer0_outputs(1874)) and not (layer0_outputs(1833));
    outputs(264) <= (layer0_outputs(2011)) and not (layer0_outputs(2081));
    outputs(265) <= (layer0_outputs(1623)) and not (layer0_outputs(2000));
    outputs(266) <= not((layer0_outputs(1812)) or (layer0_outputs(615)));
    outputs(267) <= (layer0_outputs(641)) and (layer0_outputs(383));
    outputs(268) <= (layer0_outputs(1663)) and (layer0_outputs(2155));
    outputs(269) <= (layer0_outputs(1770)) and (layer0_outputs(1394));
    outputs(270) <= not((layer0_outputs(108)) or (layer0_outputs(76)));
    outputs(271) <= (layer0_outputs(138)) and not (layer0_outputs(882));
    outputs(272) <= (layer0_outputs(1720)) and not (layer0_outputs(805));
    outputs(273) <= (layer0_outputs(1347)) and not (layer0_outputs(1920));
    outputs(274) <= layer0_outputs(1740);
    outputs(275) <= not((layer0_outputs(824)) or (layer0_outputs(466)));
    outputs(276) <= (layer0_outputs(1470)) and (layer0_outputs(2));
    outputs(277) <= (layer0_outputs(641)) and (layer0_outputs(1572));
    outputs(278) <= (layer0_outputs(1899)) and not (layer0_outputs(2024));
    outputs(279) <= (layer0_outputs(668)) and not (layer0_outputs(10));
    outputs(280) <= not((layer0_outputs(949)) or (layer0_outputs(191)));
    outputs(281) <= (layer0_outputs(1775)) and not (layer0_outputs(250));
    outputs(282) <= '0';
    outputs(283) <= (layer0_outputs(1242)) xor (layer0_outputs(1589));
    outputs(284) <= (layer0_outputs(964)) and not (layer0_outputs(1664));
    outputs(285) <= (layer0_outputs(2184)) and (layer0_outputs(1601));
    outputs(286) <= (layer0_outputs(698)) and not (layer0_outputs(1379));
    outputs(287) <= (layer0_outputs(1556)) and not (layer0_outputs(559));
    outputs(288) <= not((layer0_outputs(1715)) or (layer0_outputs(415)));
    outputs(289) <= (layer0_outputs(622)) and (layer0_outputs(1178));
    outputs(290) <= (layer0_outputs(1183)) and not (layer0_outputs(958));
    outputs(291) <= not(layer0_outputs(2361));
    outputs(292) <= not((layer0_outputs(2464)) or (layer0_outputs(2221)));
    outputs(293) <= (layer0_outputs(1784)) and not (layer0_outputs(1310));
    outputs(294) <= (layer0_outputs(319)) and not (layer0_outputs(1599));
    outputs(295) <= (layer0_outputs(1009)) and (layer0_outputs(1349));
    outputs(296) <= (layer0_outputs(1320)) and (layer0_outputs(2091));
    outputs(297) <= layer0_outputs(203);
    outputs(298) <= layer0_outputs(2497);
    outputs(299) <= (layer0_outputs(7)) and not (layer0_outputs(1749));
    outputs(300) <= not((layer0_outputs(1201)) or (layer0_outputs(1842)));
    outputs(301) <= (layer0_outputs(2441)) and not (layer0_outputs(550));
    outputs(302) <= (layer0_outputs(1991)) and not (layer0_outputs(192));
    outputs(303) <= not((layer0_outputs(2190)) or (layer0_outputs(2093)));
    outputs(304) <= not((layer0_outputs(772)) or (layer0_outputs(47)));
    outputs(305) <= (layer0_outputs(1827)) and not (layer0_outputs(525));
    outputs(306) <= (layer0_outputs(2135)) and not (layer0_outputs(1560));
    outputs(307) <= not(layer0_outputs(2355));
    outputs(308) <= (layer0_outputs(729)) and (layer0_outputs(2510));
    outputs(309) <= (layer0_outputs(982)) and (layer0_outputs(2036));
    outputs(310) <= (layer0_outputs(655)) and (layer0_outputs(574));
    outputs(311) <= (layer0_outputs(2483)) and not (layer0_outputs(1228));
    outputs(312) <= (layer0_outputs(133)) and not (layer0_outputs(1605));
    outputs(313) <= not((layer0_outputs(743)) or (layer0_outputs(1968)));
    outputs(314) <= (layer0_outputs(1004)) and not (layer0_outputs(2119));
    outputs(315) <= (layer0_outputs(2379)) and (layer0_outputs(2415));
    outputs(316) <= not((layer0_outputs(211)) or (layer0_outputs(1427)));
    outputs(317) <= not((layer0_outputs(588)) or (layer0_outputs(1013)));
    outputs(318) <= (layer0_outputs(898)) and not (layer0_outputs(185));
    outputs(319) <= (layer0_outputs(1500)) and not (layer0_outputs(1898));
    outputs(320) <= (layer0_outputs(12)) and (layer0_outputs(456));
    outputs(321) <= (layer0_outputs(623)) and not (layer0_outputs(1833));
    outputs(322) <= (layer0_outputs(2233)) and not (layer0_outputs(2261));
    outputs(323) <= not(layer0_outputs(330));
    outputs(324) <= not((layer0_outputs(977)) or (layer0_outputs(553)));
    outputs(325) <= layer0_outputs(1878);
    outputs(326) <= (layer0_outputs(1976)) and (layer0_outputs(1473));
    outputs(327) <= (layer0_outputs(1456)) and not (layer0_outputs(1698));
    outputs(328) <= (layer0_outputs(2074)) and not (layer0_outputs(2489));
    outputs(329) <= not((layer0_outputs(1517)) or (layer0_outputs(2490)));
    outputs(330) <= (layer0_outputs(2210)) and (layer0_outputs(2103));
    outputs(331) <= (layer0_outputs(2181)) and not (layer0_outputs(1327));
    outputs(332) <= (layer0_outputs(195)) and not (layer0_outputs(1795));
    outputs(333) <= not((layer0_outputs(2312)) or (layer0_outputs(379)));
    outputs(334) <= (layer0_outputs(428)) and not (layer0_outputs(916));
    outputs(335) <= (layer0_outputs(93)) and (layer0_outputs(2473));
    outputs(336) <= not((layer0_outputs(1056)) or (layer0_outputs(223)));
    outputs(337) <= (layer0_outputs(984)) and not (layer0_outputs(1986));
    outputs(338) <= not(layer0_outputs(890));
    outputs(339) <= not((layer0_outputs(740)) or (layer0_outputs(1726)));
    outputs(340) <= (layer0_outputs(823)) and (layer0_outputs(946));
    outputs(341) <= (layer0_outputs(731)) and not (layer0_outputs(2429));
    outputs(342) <= not((layer0_outputs(1861)) or (layer0_outputs(408)));
    outputs(343) <= not((layer0_outputs(2322)) or (layer0_outputs(1021)));
    outputs(344) <= (layer0_outputs(684)) and not (layer0_outputs(293));
    outputs(345) <= not((layer0_outputs(933)) or (layer0_outputs(2256)));
    outputs(346) <= (layer0_outputs(2206)) and not (layer0_outputs(1718));
    outputs(347) <= not((layer0_outputs(2236)) or (layer0_outputs(979)));
    outputs(348) <= (layer0_outputs(564)) and (layer0_outputs(2248));
    outputs(349) <= (layer0_outputs(103)) and not (layer0_outputs(1630));
    outputs(350) <= (layer0_outputs(2400)) and (layer0_outputs(1534));
    outputs(351) <= (layer0_outputs(586)) and not (layer0_outputs(852));
    outputs(352) <= (layer0_outputs(1527)) and not (layer0_outputs(2222));
    outputs(353) <= (layer0_outputs(2400)) and not (layer0_outputs(1382));
    outputs(354) <= (layer0_outputs(1340)) and not (layer0_outputs(665));
    outputs(355) <= layer0_outputs(84);
    outputs(356) <= not((layer0_outputs(1294)) or (layer0_outputs(1865)));
    outputs(357) <= (layer0_outputs(2394)) and not (layer0_outputs(913));
    outputs(358) <= (layer0_outputs(44)) and not (layer0_outputs(16));
    outputs(359) <= (layer0_outputs(355)) and not (layer0_outputs(2084));
    outputs(360) <= '0';
    outputs(361) <= '0';
    outputs(362) <= (layer0_outputs(267)) and not (layer0_outputs(1365));
    outputs(363) <= (layer0_outputs(2251)) and (layer0_outputs(931));
    outputs(364) <= (layer0_outputs(990)) and (layer0_outputs(2243));
    outputs(365) <= (layer0_outputs(203)) and not (layer0_outputs(888));
    outputs(366) <= (layer0_outputs(453)) and not (layer0_outputs(2156));
    outputs(367) <= layer0_outputs(1907);
    outputs(368) <= (layer0_outputs(860)) and (layer0_outputs(436));
    outputs(369) <= not((layer0_outputs(2055)) or (layer0_outputs(416)));
    outputs(370) <= (layer0_outputs(280)) and not (layer0_outputs(1171));
    outputs(371) <= not((layer0_outputs(799)) or (layer0_outputs(429)));
    outputs(372) <= not((layer0_outputs(1304)) or (layer0_outputs(1111)));
    outputs(373) <= (layer0_outputs(1383)) and (layer0_outputs(2534));
    outputs(374) <= not((layer0_outputs(1666)) xor (layer0_outputs(2255)));
    outputs(375) <= (layer0_outputs(292)) and not (layer0_outputs(598));
    outputs(376) <= (layer0_outputs(1931)) and not (layer0_outputs(1025));
    outputs(377) <= (layer0_outputs(1699)) and not (layer0_outputs(1765));
    outputs(378) <= not((layer0_outputs(515)) or (layer0_outputs(1047)));
    outputs(379) <= (layer0_outputs(269)) and not (layer0_outputs(1054));
    outputs(380) <= not(layer0_outputs(330));
    outputs(381) <= not((layer0_outputs(2336)) or (layer0_outputs(1237)));
    outputs(382) <= (layer0_outputs(1859)) and (layer0_outputs(642));
    outputs(383) <= (layer0_outputs(1312)) and not (layer0_outputs(1336));
    outputs(384) <= not((layer0_outputs(2260)) or (layer0_outputs(489)));
    outputs(385) <= layer0_outputs(1722);
    outputs(386) <= not(layer0_outputs(1210)) or (layer0_outputs(64));
    outputs(387) <= (layer0_outputs(2293)) and not (layer0_outputs(945));
    outputs(388) <= (layer0_outputs(596)) and not (layer0_outputs(2087));
    outputs(389) <= layer0_outputs(116);
    outputs(390) <= (layer0_outputs(1244)) and not (layer0_outputs(340));
    outputs(391) <= '0';
    outputs(392) <= (layer0_outputs(1790)) and not (layer0_outputs(1566));
    outputs(393) <= not((layer0_outputs(214)) or (layer0_outputs(492)));
    outputs(394) <= (layer0_outputs(1029)) and not (layer0_outputs(1789));
    outputs(395) <= '0';
    outputs(396) <= not((layer0_outputs(266)) or (layer0_outputs(1797)));
    outputs(397) <= not((layer0_outputs(2224)) or (layer0_outputs(2127)));
    outputs(398) <= layer0_outputs(1225);
    outputs(399) <= not((layer0_outputs(288)) or (layer0_outputs(1543)));
    outputs(400) <= (layer0_outputs(2153)) and not (layer0_outputs(829));
    outputs(401) <= (layer0_outputs(1815)) and (layer0_outputs(1712));
    outputs(402) <= not((layer0_outputs(1138)) or (layer0_outputs(95)));
    outputs(403) <= (layer0_outputs(1700)) and (layer0_outputs(2391));
    outputs(404) <= not((layer0_outputs(1372)) or (layer0_outputs(179)));
    outputs(405) <= not(layer0_outputs(1039));
    outputs(406) <= (layer0_outputs(274)) and not (layer0_outputs(831));
    outputs(407) <= (layer0_outputs(2518)) and not (layer0_outputs(627));
    outputs(408) <= (layer0_outputs(2354)) and not (layer0_outputs(714));
    outputs(409) <= not((layer0_outputs(997)) or (layer0_outputs(2424)));
    outputs(410) <= '0';
    outputs(411) <= (layer0_outputs(1166)) and not (layer0_outputs(2412));
    outputs(412) <= (layer0_outputs(569)) and not (layer0_outputs(1732));
    outputs(413) <= (layer0_outputs(1211)) and not (layer0_outputs(644));
    outputs(414) <= not((layer0_outputs(1156)) or (layer0_outputs(1382)));
    outputs(415) <= not((layer0_outputs(2343)) or (layer0_outputs(902)));
    outputs(416) <= (layer0_outputs(2294)) and not (layer0_outputs(772));
    outputs(417) <= not((layer0_outputs(1811)) or (layer0_outputs(351)));
    outputs(418) <= not((layer0_outputs(677)) or (layer0_outputs(1442)));
    outputs(419) <= (layer0_outputs(35)) and (layer0_outputs(1944));
    outputs(420) <= not(layer0_outputs(1351));
    outputs(421) <= (layer0_outputs(2399)) and (layer0_outputs(1468));
    outputs(422) <= (layer0_outputs(736)) and not (layer0_outputs(646));
    outputs(423) <= not((layer0_outputs(740)) or (layer0_outputs(2479)));
    outputs(424) <= not((layer0_outputs(2338)) or (layer0_outputs(1703)));
    outputs(425) <= (layer0_outputs(1060)) and not (layer0_outputs(1729));
    outputs(426) <= (layer0_outputs(1585)) and (layer0_outputs(1859));
    outputs(427) <= not((layer0_outputs(2303)) or (layer0_outputs(1937)));
    outputs(428) <= (layer0_outputs(1993)) and not (layer0_outputs(155));
    outputs(429) <= not((layer0_outputs(681)) or (layer0_outputs(819)));
    outputs(430) <= (layer0_outputs(2503)) and not (layer0_outputs(1932));
    outputs(431) <= not((layer0_outputs(2547)) or (layer0_outputs(413)));
    outputs(432) <= not(layer0_outputs(71)) or (layer0_outputs(974));
    outputs(433) <= (layer0_outputs(443)) and not (layer0_outputs(1946));
    outputs(434) <= not((layer0_outputs(1954)) or (layer0_outputs(1363)));
    outputs(435) <= (layer0_outputs(11)) and not (layer0_outputs(1476));
    outputs(436) <= (layer0_outputs(592)) and not (layer0_outputs(799));
    outputs(437) <= (layer0_outputs(110)) and (layer0_outputs(1295));
    outputs(438) <= not((layer0_outputs(1829)) or (layer0_outputs(2500)));
    outputs(439) <= (layer0_outputs(851)) xor (layer0_outputs(2521));
    outputs(440) <= (layer0_outputs(2551)) and (layer0_outputs(338));
    outputs(441) <= (layer0_outputs(1251)) and not (layer0_outputs(152));
    outputs(442) <= layer0_outputs(1487);
    outputs(443) <= (layer0_outputs(2107)) and (layer0_outputs(1690));
    outputs(444) <= not(layer0_outputs(2256));
    outputs(445) <= layer0_outputs(2503);
    outputs(446) <= not(layer0_outputs(1453)) or (layer0_outputs(1279));
    outputs(447) <= (layer0_outputs(1100)) and not (layer0_outputs(372));
    outputs(448) <= not((layer0_outputs(858)) or (layer0_outputs(1317)));
    outputs(449) <= (layer0_outputs(1369)) and (layer0_outputs(346));
    outputs(450) <= (layer0_outputs(244)) and not (layer0_outputs(780));
    outputs(451) <= (layer0_outputs(1985)) and (layer0_outputs(1826));
    outputs(452) <= (layer0_outputs(172)) and not (layer0_outputs(602));
    outputs(453) <= (layer0_outputs(2128)) and not (layer0_outputs(445));
    outputs(454) <= (layer0_outputs(509)) and (layer0_outputs(1000));
    outputs(455) <= (layer0_outputs(1069)) and not (layer0_outputs(747));
    outputs(456) <= not((layer0_outputs(1645)) or (layer0_outputs(2260)));
    outputs(457) <= (layer0_outputs(735)) and (layer0_outputs(228));
    outputs(458) <= (layer0_outputs(2433)) and not (layer0_outputs(2546));
    outputs(459) <= (layer0_outputs(1153)) and not (layer0_outputs(1980));
    outputs(460) <= (layer0_outputs(463)) and (layer0_outputs(1959));
    outputs(461) <= not((layer0_outputs(1431)) or (layer0_outputs(316)));
    outputs(462) <= (layer0_outputs(1649)) and not (layer0_outputs(367));
    outputs(463) <= (layer0_outputs(1830)) and not (layer0_outputs(23));
    outputs(464) <= (layer0_outputs(165)) and (layer0_outputs(654));
    outputs(465) <= (layer0_outputs(376)) and (layer0_outputs(1661));
    outputs(466) <= layer0_outputs(1450);
    outputs(467) <= (layer0_outputs(2558)) and not (layer0_outputs(1754));
    outputs(468) <= not((layer0_outputs(2271)) or (layer0_outputs(839)));
    outputs(469) <= (layer0_outputs(220)) and not (layer0_outputs(2553));
    outputs(470) <= (layer0_outputs(555)) and (layer0_outputs(78));
    outputs(471) <= not((layer0_outputs(1170)) or (layer0_outputs(863)));
    outputs(472) <= not((layer0_outputs(2089)) or (layer0_outputs(1873)));
    outputs(473) <= (layer0_outputs(2304)) and not (layer0_outputs(2249));
    outputs(474) <= (layer0_outputs(1960)) and (layer0_outputs(2199));
    outputs(475) <= (layer0_outputs(1487)) and not (layer0_outputs(1654));
    outputs(476) <= (layer0_outputs(1551)) and not (layer0_outputs(1870));
    outputs(477) <= (layer0_outputs(411)) and (layer0_outputs(678));
    outputs(478) <= (layer0_outputs(1734)) and (layer0_outputs(56));
    outputs(479) <= not((layer0_outputs(558)) or (layer0_outputs(1678)));
    outputs(480) <= not(layer0_outputs(899));
    outputs(481) <= not(layer0_outputs(884));
    outputs(482) <= not((layer0_outputs(1557)) or (layer0_outputs(605)));
    outputs(483) <= (layer0_outputs(731)) and not (layer0_outputs(2546));
    outputs(484) <= (layer0_outputs(2386)) and not (layer0_outputs(1951));
    outputs(485) <= (layer0_outputs(69)) and not (layer0_outputs(2410));
    outputs(486) <= not((layer0_outputs(1102)) or (layer0_outputs(182)));
    outputs(487) <= (layer0_outputs(690)) and not (layer0_outputs(1107));
    outputs(488) <= not((layer0_outputs(247)) xor (layer0_outputs(2111)));
    outputs(489) <= not((layer0_outputs(1957)) or (layer0_outputs(966)));
    outputs(490) <= (layer0_outputs(883)) and not (layer0_outputs(2016));
    outputs(491) <= not((layer0_outputs(1385)) or (layer0_outputs(1013)));
    outputs(492) <= (layer0_outputs(844)) and not (layer0_outputs(30));
    outputs(493) <= (layer0_outputs(1415)) and not (layer0_outputs(1243));
    outputs(494) <= (layer0_outputs(2527)) and (layer0_outputs(1830));
    outputs(495) <= not(layer0_outputs(2367));
    outputs(496) <= not(layer0_outputs(2308));
    outputs(497) <= not((layer0_outputs(2136)) or (layer0_outputs(1236)));
    outputs(498) <= (layer0_outputs(1062)) and not (layer0_outputs(1278));
    outputs(499) <= not(layer0_outputs(1758));
    outputs(500) <= not((layer0_outputs(925)) or (layer0_outputs(1410)));
    outputs(501) <= (layer0_outputs(840)) and not (layer0_outputs(1324));
    outputs(502) <= (layer0_outputs(2414)) and not (layer0_outputs(936));
    outputs(503) <= (layer0_outputs(766)) and not (layer0_outputs(2454));
    outputs(504) <= (layer0_outputs(1525)) and not (layer0_outputs(850));
    outputs(505) <= (layer0_outputs(2559)) and not (layer0_outputs(1311));
    outputs(506) <= layer0_outputs(750);
    outputs(507) <= (layer0_outputs(1612)) and not (layer0_outputs(317));
    outputs(508) <= (layer0_outputs(984)) and not (layer0_outputs(865));
    outputs(509) <= (layer0_outputs(620)) and not (layer0_outputs(1947));
    outputs(510) <= (layer0_outputs(968)) and not (layer0_outputs(1679));
    outputs(511) <= (layer0_outputs(15)) and (layer0_outputs(763));
    outputs(512) <= (layer0_outputs(1005)) and not (layer0_outputs(1386));
    outputs(513) <= layer0_outputs(603);
    outputs(514) <= not(layer0_outputs(2290));
    outputs(515) <= not(layer0_outputs(1286)) or (layer0_outputs(554));
    outputs(516) <= not(layer0_outputs(612)) or (layer0_outputs(992));
    outputs(517) <= not((layer0_outputs(1694)) and (layer0_outputs(2153)));
    outputs(518) <= (layer0_outputs(382)) or (layer0_outputs(92));
    outputs(519) <= not(layer0_outputs(357));
    outputs(520) <= not(layer0_outputs(326)) or (layer0_outputs(1642));
    outputs(521) <= layer0_outputs(2517);
    outputs(522) <= not((layer0_outputs(797)) or (layer0_outputs(1448)));
    outputs(523) <= not((layer0_outputs(2236)) xor (layer0_outputs(656)));
    outputs(524) <= not(layer0_outputs(2440)) or (layer0_outputs(2396));
    outputs(525) <= not(layer0_outputs(1068)) or (layer0_outputs(2436));
    outputs(526) <= layer0_outputs(1866);
    outputs(527) <= not(layer0_outputs(1980));
    outputs(528) <= (layer0_outputs(1432)) or (layer0_outputs(1084));
    outputs(529) <= layer0_outputs(2504);
    outputs(530) <= (layer0_outputs(267)) and not (layer0_outputs(923));
    outputs(531) <= not(layer0_outputs(1484));
    outputs(532) <= not(layer0_outputs(510)) or (layer0_outputs(1697));
    outputs(533) <= (layer0_outputs(184)) and not (layer0_outputs(1802));
    outputs(534) <= not(layer0_outputs(40));
    outputs(535) <= not((layer0_outputs(227)) and (layer0_outputs(91)));
    outputs(536) <= (layer0_outputs(2000)) xor (layer0_outputs(1771));
    outputs(537) <= not(layer0_outputs(1539));
    outputs(538) <= not(layer0_outputs(687));
    outputs(539) <= (layer0_outputs(181)) xor (layer0_outputs(1774));
    outputs(540) <= not(layer0_outputs(2292));
    outputs(541) <= not(layer0_outputs(1602));
    outputs(542) <= (layer0_outputs(1824)) and not (layer0_outputs(1221));
    outputs(543) <= not(layer0_outputs(922)) or (layer0_outputs(327));
    outputs(544) <= not((layer0_outputs(1319)) or (layer0_outputs(1078)));
    outputs(545) <= layer0_outputs(1084);
    outputs(546) <= (layer0_outputs(1873)) or (layer0_outputs(492));
    outputs(547) <= not(layer0_outputs(511)) or (layer0_outputs(639));
    outputs(548) <= (layer0_outputs(2296)) or (layer0_outputs(1601));
    outputs(549) <= not(layer0_outputs(521));
    outputs(550) <= (layer0_outputs(854)) xor (layer0_outputs(449));
    outputs(551) <= not((layer0_outputs(2136)) xor (layer0_outputs(2039)));
    outputs(552) <= layer0_outputs(1284);
    outputs(553) <= not(layer0_outputs(1604)) or (layer0_outputs(869));
    outputs(554) <= layer0_outputs(1148);
    outputs(555) <= (layer0_outputs(2286)) and not (layer0_outputs(956));
    outputs(556) <= not((layer0_outputs(209)) and (layer0_outputs(1068)));
    outputs(557) <= not((layer0_outputs(969)) xor (layer0_outputs(762)));
    outputs(558) <= not((layer0_outputs(1501)) and (layer0_outputs(2422)));
    outputs(559) <= not(layer0_outputs(1140)) or (layer0_outputs(61));
    outputs(560) <= not(layer0_outputs(1917));
    outputs(561) <= layer0_outputs(1447);
    outputs(562) <= (layer0_outputs(1619)) and not (layer0_outputs(474));
    outputs(563) <= (layer0_outputs(1725)) and (layer0_outputs(0));
    outputs(564) <= not(layer0_outputs(532)) or (layer0_outputs(2230));
    outputs(565) <= not((layer0_outputs(1669)) xor (layer0_outputs(2308)));
    outputs(566) <= (layer0_outputs(1840)) and not (layer0_outputs(995));
    outputs(567) <= layer0_outputs(2033);
    outputs(568) <= not(layer0_outputs(1264));
    outputs(569) <= (layer0_outputs(306)) and (layer0_outputs(311));
    outputs(570) <= not(layer0_outputs(927)) or (layer0_outputs(1989));
    outputs(571) <= not(layer0_outputs(2516));
    outputs(572) <= not((layer0_outputs(1638)) xor (layer0_outputs(1074)));
    outputs(573) <= not(layer0_outputs(1707));
    outputs(574) <= (layer0_outputs(819)) xor (layer0_outputs(1197));
    outputs(575) <= layer0_outputs(134);
    outputs(576) <= (layer0_outputs(2411)) and not (layer0_outputs(486));
    outputs(577) <= layer0_outputs(1179);
    outputs(578) <= not(layer0_outputs(1009));
    outputs(579) <= not(layer0_outputs(1739));
    outputs(580) <= not(layer0_outputs(250));
    outputs(581) <= not((layer0_outputs(426)) and (layer0_outputs(2274)));
    outputs(582) <= not(layer0_outputs(1667));
    outputs(583) <= (layer0_outputs(1988)) or (layer0_outputs(148));
    outputs(584) <= not(layer0_outputs(263)) or (layer0_outputs(1979));
    outputs(585) <= not(layer0_outputs(2377));
    outputs(586) <= layer0_outputs(347);
    outputs(587) <= (layer0_outputs(707)) and (layer0_outputs(842));
    outputs(588) <= layer0_outputs(1901);
    outputs(589) <= layer0_outputs(2037);
    outputs(590) <= layer0_outputs(793);
    outputs(591) <= (layer0_outputs(954)) or (layer0_outputs(2327));
    outputs(592) <= not(layer0_outputs(1814));
    outputs(593) <= not((layer0_outputs(1425)) xor (layer0_outputs(1134)));
    outputs(594) <= not(layer0_outputs(1142));
    outputs(595) <= not(layer0_outputs(51));
    outputs(596) <= not(layer0_outputs(2244)) or (layer0_outputs(757));
    outputs(597) <= not(layer0_outputs(613)) or (layer0_outputs(2078));
    outputs(598) <= (layer0_outputs(13)) xor (layer0_outputs(1290));
    outputs(599) <= (layer0_outputs(1795)) or (layer0_outputs(1834));
    outputs(600) <= layer0_outputs(286);
    outputs(601) <= not(layer0_outputs(1463));
    outputs(602) <= layer0_outputs(430);
    outputs(603) <= not(layer0_outputs(1469)) or (layer0_outputs(1735));
    outputs(604) <= not(layer0_outputs(1637));
    outputs(605) <= layer0_outputs(1236);
    outputs(606) <= layer0_outputs(776);
    outputs(607) <= layer0_outputs(446);
    outputs(608) <= (layer0_outputs(395)) xor (layer0_outputs(1380));
    outputs(609) <= layer0_outputs(2218);
    outputs(610) <= not(layer0_outputs(1280));
    outputs(611) <= not(layer0_outputs(434));
    outputs(612) <= not(layer0_outputs(352));
    outputs(613) <= not(layer0_outputs(1414)) or (layer0_outputs(373));
    outputs(614) <= not(layer0_outputs(1974)) or (layer0_outputs(2531));
    outputs(615) <= layer0_outputs(2185);
    outputs(616) <= not(layer0_outputs(1685));
    outputs(617) <= (layer0_outputs(144)) xor (layer0_outputs(2163));
    outputs(618) <= not(layer0_outputs(2035));
    outputs(619) <= not(layer0_outputs(791));
    outputs(620) <= (layer0_outputs(562)) and (layer0_outputs(413));
    outputs(621) <= (layer0_outputs(1752)) xor (layer0_outputs(1500));
    outputs(622) <= not((layer0_outputs(1981)) xor (layer0_outputs(1435)));
    outputs(623) <= layer0_outputs(1025);
    outputs(624) <= layer0_outputs(1783);
    outputs(625) <= (layer0_outputs(1766)) and not (layer0_outputs(151));
    outputs(626) <= not(layer0_outputs(2466));
    outputs(627) <= (layer0_outputs(725)) and not (layer0_outputs(2328));
    outputs(628) <= not((layer0_outputs(1924)) xor (layer0_outputs(1371)));
    outputs(629) <= (layer0_outputs(2050)) and (layer0_outputs(368));
    outputs(630) <= (layer0_outputs(1148)) and not (layer0_outputs(995));
    outputs(631) <= (layer0_outputs(2321)) and not (layer0_outputs(1051));
    outputs(632) <= not(layer0_outputs(1573));
    outputs(633) <= (layer0_outputs(1359)) and not (layer0_outputs(640));
    outputs(634) <= (layer0_outputs(457)) and (layer0_outputs(893));
    outputs(635) <= not(layer0_outputs(1293)) or (layer0_outputs(2242));
    outputs(636) <= not(layer0_outputs(544)) or (layer0_outputs(1546));
    outputs(637) <= not((layer0_outputs(1631)) and (layer0_outputs(1714)));
    outputs(638) <= (layer0_outputs(713)) or (layer0_outputs(2351));
    outputs(639) <= not(layer0_outputs(1250));
    outputs(640) <= not(layer0_outputs(1112));
    outputs(641) <= (layer0_outputs(306)) and (layer0_outputs(1027));
    outputs(642) <= (layer0_outputs(1708)) or (layer0_outputs(906));
    outputs(643) <= not(layer0_outputs(1911));
    outputs(644) <= not(layer0_outputs(1161));
    outputs(645) <= layer0_outputs(1113);
    outputs(646) <= (layer0_outputs(1028)) and not (layer0_outputs(1030));
    outputs(647) <= not(layer0_outputs(337));
    outputs(648) <= not(layer0_outputs(2096));
    outputs(649) <= not((layer0_outputs(88)) or (layer0_outputs(2161)));
    outputs(650) <= layer0_outputs(893);
    outputs(651) <= layer0_outputs(2519);
    outputs(652) <= (layer0_outputs(1085)) xor (layer0_outputs(1196));
    outputs(653) <= (layer0_outputs(2087)) and (layer0_outputs(777));
    outputs(654) <= layer0_outputs(1022);
    outputs(655) <= layer0_outputs(109);
    outputs(656) <= not(layer0_outputs(668));
    outputs(657) <= (layer0_outputs(295)) and not (layer0_outputs(535));
    outputs(658) <= (layer0_outputs(34)) and not (layer0_outputs(2121));
    outputs(659) <= layer0_outputs(2033);
    outputs(660) <= (layer0_outputs(724)) and (layer0_outputs(657));
    outputs(661) <= layer0_outputs(971);
    outputs(662) <= not((layer0_outputs(1667)) and (layer0_outputs(987)));
    outputs(663) <= layer0_outputs(1480);
    outputs(664) <= not((layer0_outputs(2096)) or (layer0_outputs(434)));
    outputs(665) <= not(layer0_outputs(353));
    outputs(666) <= (layer0_outputs(1146)) and (layer0_outputs(2301));
    outputs(667) <= not(layer0_outputs(278));
    outputs(668) <= (layer0_outputs(2141)) or (layer0_outputs(335));
    outputs(669) <= layer0_outputs(1805);
    outputs(670) <= (layer0_outputs(673)) and not (layer0_outputs(1841));
    outputs(671) <= not(layer0_outputs(474));
    outputs(672) <= not((layer0_outputs(409)) or (layer0_outputs(626)));
    outputs(673) <= not(layer0_outputs(7));
    outputs(674) <= (layer0_outputs(693)) xor (layer0_outputs(148));
    outputs(675) <= layer0_outputs(2456);
    outputs(676) <= not(layer0_outputs(2027));
    outputs(677) <= (layer0_outputs(370)) xor (layer0_outputs(1229));
    outputs(678) <= layer0_outputs(1507);
    outputs(679) <= (layer0_outputs(1210)) or (layer0_outputs(2240));
    outputs(680) <= (layer0_outputs(33)) or (layer0_outputs(839));
    outputs(681) <= (layer0_outputs(2246)) or (layer0_outputs(1899));
    outputs(682) <= not((layer0_outputs(2105)) xor (layer0_outputs(552)));
    outputs(683) <= (layer0_outputs(589)) or (layer0_outputs(1428));
    outputs(684) <= (layer0_outputs(1131)) and not (layer0_outputs(196));
    outputs(685) <= not((layer0_outputs(1141)) and (layer0_outputs(1775)));
    outputs(686) <= layer0_outputs(2146);
    outputs(687) <= not(layer0_outputs(440));
    outputs(688) <= not(layer0_outputs(2150)) or (layer0_outputs(1583));
    outputs(689) <= not(layer0_outputs(1338));
    outputs(690) <= (layer0_outputs(1151)) and (layer0_outputs(669));
    outputs(691) <= (layer0_outputs(1219)) and not (layer0_outputs(773));
    outputs(692) <= not(layer0_outputs(1137)) or (layer0_outputs(1935));
    outputs(693) <= not(layer0_outputs(160));
    outputs(694) <= (layer0_outputs(433)) and not (layer0_outputs(1272));
    outputs(695) <= (layer0_outputs(2117)) and not (layer0_outputs(1635));
    outputs(696) <= not(layer0_outputs(2186));
    outputs(697) <= not(layer0_outputs(96));
    outputs(698) <= not((layer0_outputs(1728)) and (layer0_outputs(103)));
    outputs(699) <= (layer0_outputs(1230)) and (layer0_outputs(128));
    outputs(700) <= layer0_outputs(1710);
    outputs(701) <= not((layer0_outputs(585)) xor (layer0_outputs(1871)));
    outputs(702) <= layer0_outputs(202);
    outputs(703) <= not(layer0_outputs(2275)) or (layer0_outputs(917));
    outputs(704) <= layer0_outputs(2505);
    outputs(705) <= not((layer0_outputs(1816)) and (layer0_outputs(994)));
    outputs(706) <= not(layer0_outputs(305));
    outputs(707) <= (layer0_outputs(356)) or (layer0_outputs(2314));
    outputs(708) <= not(layer0_outputs(2403)) or (layer0_outputs(281));
    outputs(709) <= (layer0_outputs(2438)) and not (layer0_outputs(2220));
    outputs(710) <= not(layer0_outputs(838));
    outputs(711) <= layer0_outputs(1269);
    outputs(712) <= not(layer0_outputs(343)) or (layer0_outputs(2399));
    outputs(713) <= not(layer0_outputs(1232));
    outputs(714) <= (layer0_outputs(1054)) or (layer0_outputs(827));
    outputs(715) <= layer0_outputs(1408);
    outputs(716) <= not((layer0_outputs(477)) xor (layer0_outputs(2129)));
    outputs(717) <= layer0_outputs(1741);
    outputs(718) <= (layer0_outputs(1329)) and not (layer0_outputs(1130));
    outputs(719) <= not((layer0_outputs(2393)) and (layer0_outputs(736)));
    outputs(720) <= not((layer0_outputs(809)) or (layer0_outputs(1459)));
    outputs(721) <= layer0_outputs(1954);
    outputs(722) <= (layer0_outputs(2214)) xor (layer0_outputs(2238));
    outputs(723) <= layer0_outputs(1851);
    outputs(724) <= (layer0_outputs(1875)) or (layer0_outputs(1883));
    outputs(725) <= not(layer0_outputs(1483));
    outputs(726) <= not(layer0_outputs(503));
    outputs(727) <= (layer0_outputs(1660)) or (layer0_outputs(2502));
    outputs(728) <= not(layer0_outputs(2343));
    outputs(729) <= not(layer0_outputs(576));
    outputs(730) <= not(layer0_outputs(653));
    outputs(731) <= layer0_outputs(2383);
    outputs(732) <= layer0_outputs(90);
    outputs(733) <= (layer0_outputs(1315)) and not (layer0_outputs(390));
    outputs(734) <= not((layer0_outputs(640)) or (layer0_outputs(939)));
    outputs(735) <= not((layer0_outputs(2179)) and (layer0_outputs(463)));
    outputs(736) <= layer0_outputs(2112);
    outputs(737) <= layer0_outputs(1893);
    outputs(738) <= layer0_outputs(1620);
    outputs(739) <= not(layer0_outputs(432));
    outputs(740) <= (layer0_outputs(395)) and not (layer0_outputs(218));
    outputs(741) <= not((layer0_outputs(2512)) and (layer0_outputs(142)));
    outputs(742) <= (layer0_outputs(451)) and not (layer0_outputs(1474));
    outputs(743) <= (layer0_outputs(865)) and not (layer0_outputs(619));
    outputs(744) <= (layer0_outputs(1427)) or (layer0_outputs(378));
    outputs(745) <= not(layer0_outputs(1182));
    outputs(746) <= layer0_outputs(1156);
    outputs(747) <= (layer0_outputs(146)) xor (layer0_outputs(2465));
    outputs(748) <= (layer0_outputs(2089)) and not (layer0_outputs(121));
    outputs(749) <= layer0_outputs(1875);
    outputs(750) <= not(layer0_outputs(2150)) or (layer0_outputs(874));
    outputs(751) <= layer0_outputs(1447);
    outputs(752) <= not(layer0_outputs(2461));
    outputs(753) <= layer0_outputs(821);
    outputs(754) <= not((layer0_outputs(2262)) and (layer0_outputs(1154)));
    outputs(755) <= (layer0_outputs(1730)) or (layer0_outputs(2106));
    outputs(756) <= not((layer0_outputs(960)) xor (layer0_outputs(1036)));
    outputs(757) <= not((layer0_outputs(2524)) and (layer0_outputs(1906)));
    outputs(758) <= (layer0_outputs(1058)) and not (layer0_outputs(466));
    outputs(759) <= not((layer0_outputs(1801)) or (layer0_outputs(1483)));
    outputs(760) <= not((layer0_outputs(89)) and (layer0_outputs(212)));
    outputs(761) <= not(layer0_outputs(341));
    outputs(762) <= (layer0_outputs(993)) xor (layer0_outputs(2408));
    outputs(763) <= not(layer0_outputs(737)) or (layer0_outputs(1555));
    outputs(764) <= (layer0_outputs(1658)) xor (layer0_outputs(695));
    outputs(765) <= (layer0_outputs(823)) and not (layer0_outputs(1972));
    outputs(766) <= not(layer0_outputs(666));
    outputs(767) <= layer0_outputs(739);
    outputs(768) <= not(layer0_outputs(1129)) or (layer0_outputs(761));
    outputs(769) <= (layer0_outputs(2539)) and not (layer0_outputs(625));
    outputs(770) <= not(layer0_outputs(1579));
    outputs(771) <= not((layer0_outputs(1673)) or (layer0_outputs(1836)));
    outputs(772) <= not((layer0_outputs(229)) or (layer0_outputs(1634)));
    outputs(773) <= not((layer0_outputs(1261)) xor (layer0_outputs(1568)));
    outputs(774) <= (layer0_outputs(2282)) and not (layer0_outputs(564));
    outputs(775) <= layer0_outputs(981);
    outputs(776) <= not(layer0_outputs(1355));
    outputs(777) <= layer0_outputs(502);
    outputs(778) <= not(layer0_outputs(345));
    outputs(779) <= not(layer0_outputs(631));
    outputs(780) <= not(layer0_outputs(849)) or (layer0_outputs(2502));
    outputs(781) <= not(layer0_outputs(393));
    outputs(782) <= (layer0_outputs(1600)) and not (layer0_outputs(1244));
    outputs(783) <= not(layer0_outputs(2098)) or (layer0_outputs(289));
    outputs(784) <= not((layer0_outputs(1494)) or (layer0_outputs(1436)));
    outputs(785) <= not(layer0_outputs(604));
    outputs(786) <= layer0_outputs(2013);
    outputs(787) <= not(layer0_outputs(2319));
    outputs(788) <= not(layer0_outputs(1233));
    outputs(789) <= not(layer0_outputs(985));
    outputs(790) <= not(layer0_outputs(1281)) or (layer0_outputs(2530));
    outputs(791) <= not(layer0_outputs(1216));
    outputs(792) <= not(layer0_outputs(1635));
    outputs(793) <= (layer0_outputs(880)) or (layer0_outputs(238));
    outputs(794) <= (layer0_outputs(2173)) and (layer0_outputs(1542));
    outputs(795) <= not(layer0_outputs(1471));
    outputs(796) <= not((layer0_outputs(1389)) and (layer0_outputs(1418)));
    outputs(797) <= (layer0_outputs(199)) and not (layer0_outputs(1742));
    outputs(798) <= layer0_outputs(732);
    outputs(799) <= layer0_outputs(1472);
    outputs(800) <= (layer0_outputs(1143)) and not (layer0_outputs(596));
    outputs(801) <= not(layer0_outputs(646));
    outputs(802) <= not(layer0_outputs(62)) or (layer0_outputs(2002));
    outputs(803) <= (layer0_outputs(2129)) and (layer0_outputs(1584));
    outputs(804) <= not((layer0_outputs(1049)) or (layer0_outputs(1675)));
    outputs(805) <= (layer0_outputs(1094)) and (layer0_outputs(965));
    outputs(806) <= not(layer0_outputs(1565)) or (layer0_outputs(1312));
    outputs(807) <= not(layer0_outputs(855));
    outputs(808) <= (layer0_outputs(594)) and (layer0_outputs(1206));
    outputs(809) <= layer0_outputs(1822);
    outputs(810) <= (layer0_outputs(636)) and not (layer0_outputs(1831));
    outputs(811) <= (layer0_outputs(1331)) and (layer0_outputs(1174));
    outputs(812) <= not((layer0_outputs(1282)) or (layer0_outputs(2222)));
    outputs(813) <= layer0_outputs(2067);
    outputs(814) <= not((layer0_outputs(2319)) or (layer0_outputs(64)));
    outputs(815) <= layer0_outputs(1844);
    outputs(816) <= layer0_outputs(1633);
    outputs(817) <= not(layer0_outputs(855));
    outputs(818) <= not((layer0_outputs(2177)) or (layer0_outputs(764)));
    outputs(819) <= (layer0_outputs(1631)) and (layer0_outputs(1040));
    outputs(820) <= not((layer0_outputs(2513)) xor (layer0_outputs(2464)));
    outputs(821) <= not(layer0_outputs(2313));
    outputs(822) <= layer0_outputs(847);
    outputs(823) <= not(layer0_outputs(1322));
    outputs(824) <= not((layer0_outputs(2110)) and (layer0_outputs(2395)));
    outputs(825) <= not((layer0_outputs(276)) xor (layer0_outputs(2152)));
    outputs(826) <= not((layer0_outputs(1460)) or (layer0_outputs(2337)));
    outputs(827) <= not((layer0_outputs(398)) and (layer0_outputs(437)));
    outputs(828) <= (layer0_outputs(2124)) or (layer0_outputs(2534));
    outputs(829) <= not(layer0_outputs(1289));
    outputs(830) <= not(layer0_outputs(2007));
    outputs(831) <= (layer0_outputs(2402)) and not (layer0_outputs(2324));
    outputs(832) <= layer0_outputs(828);
    outputs(833) <= (layer0_outputs(1228)) and not (layer0_outputs(2127));
    outputs(834) <= layer0_outputs(982);
    outputs(835) <= not(layer0_outputs(21)) or (layer0_outputs(648));
    outputs(836) <= (layer0_outputs(313)) and not (layer0_outputs(5));
    outputs(837) <= layer0_outputs(1037);
    outputs(838) <= layer0_outputs(410);
    outputs(839) <= not(layer0_outputs(604));
    outputs(840) <= layer0_outputs(1050);
    outputs(841) <= not(layer0_outputs(1624));
    outputs(842) <= layer0_outputs(1086);
    outputs(843) <= layer0_outputs(1231);
    outputs(844) <= not(layer0_outputs(2500));
    outputs(845) <= layer0_outputs(801);
    outputs(846) <= (layer0_outputs(1515)) and not (layer0_outputs(2324));
    outputs(847) <= (layer0_outputs(245)) and (layer0_outputs(754));
    outputs(848) <= not(layer0_outputs(282));
    outputs(849) <= (layer0_outputs(310)) and (layer0_outputs(2288));
    outputs(850) <= layer0_outputs(1413);
    outputs(851) <= (layer0_outputs(99)) or (layer0_outputs(160));
    outputs(852) <= layer0_outputs(2306);
    outputs(853) <= not(layer0_outputs(1277));
    outputs(854) <= not((layer0_outputs(219)) or (layer0_outputs(1738)));
    outputs(855) <= layer0_outputs(2194);
    outputs(856) <= layer0_outputs(1650);
    outputs(857) <= layer0_outputs(1080);
    outputs(858) <= (layer0_outputs(91)) xor (layer0_outputs(939));
    outputs(859) <= layer0_outputs(158);
    outputs(860) <= (layer0_outputs(2309)) or (layer0_outputs(1160));
    outputs(861) <= (layer0_outputs(1529)) and not (layer0_outputs(1710));
    outputs(862) <= layer0_outputs(2431);
    outputs(863) <= not(layer0_outputs(987)) or (layer0_outputs(1424));
    outputs(864) <= (layer0_outputs(166)) and not (layer0_outputs(1986));
    outputs(865) <= (layer0_outputs(1224)) and (layer0_outputs(1260));
    outputs(866) <= layer0_outputs(595);
    outputs(867) <= (layer0_outputs(1842)) and (layer0_outputs(566));
    outputs(868) <= not(layer0_outputs(2466));
    outputs(869) <= layer0_outputs(2011);
    outputs(870) <= not(layer0_outputs(1721)) or (layer0_outputs(983));
    outputs(871) <= layer0_outputs(265);
    outputs(872) <= layer0_outputs(1876);
    outputs(873) <= not(layer0_outputs(1258)) or (layer0_outputs(1800));
    outputs(874) <= layer0_outputs(163);
    outputs(875) <= not(layer0_outputs(671));
    outputs(876) <= not((layer0_outputs(2257)) or (layer0_outputs(2366)));
    outputs(877) <= not(layer0_outputs(2210));
    outputs(878) <= not(layer0_outputs(1507));
    outputs(879) <= (layer0_outputs(922)) and (layer0_outputs(727));
    outputs(880) <= layer0_outputs(950);
    outputs(881) <= not(layer0_outputs(1925));
    outputs(882) <= layer0_outputs(2391);
    outputs(883) <= layer0_outputs(936);
    outputs(884) <= layer0_outputs(2031);
    outputs(885) <= not(layer0_outputs(584)) or (layer0_outputs(2369));
    outputs(886) <= layer0_outputs(1041);
    outputs(887) <= (layer0_outputs(1405)) and not (layer0_outputs(1016));
    outputs(888) <= layer0_outputs(1885);
    outputs(889) <= not(layer0_outputs(513));
    outputs(890) <= not(layer0_outputs(937));
    outputs(891) <= not(layer0_outputs(817)) or (layer0_outputs(1862));
    outputs(892) <= (layer0_outputs(630)) and (layer0_outputs(765));
    outputs(893) <= layer0_outputs(868);
    outputs(894) <= (layer0_outputs(2380)) and not (layer0_outputs(2257));
    outputs(895) <= not(layer0_outputs(846));
    outputs(896) <= (layer0_outputs(1101)) or (layer0_outputs(1715));
    outputs(897) <= not((layer0_outputs(1201)) or (layer0_outputs(904)));
    outputs(898) <= not(layer0_outputs(1092));
    outputs(899) <= not((layer0_outputs(1863)) and (layer0_outputs(1321)));
    outputs(900) <= layer0_outputs(875);
    outputs(901) <= (layer0_outputs(2485)) xor (layer0_outputs(475));
    outputs(902) <= not((layer0_outputs(25)) or (layer0_outputs(225)));
    outputs(903) <= layer0_outputs(1852);
    outputs(904) <= not(layer0_outputs(2433)) or (layer0_outputs(1493));
    outputs(905) <= (layer0_outputs(1786)) and not (layer0_outputs(659));
    outputs(906) <= layer0_outputs(660);
    outputs(907) <= not(layer0_outputs(2549)) or (layer0_outputs(210));
    outputs(908) <= not(layer0_outputs(2151));
    outputs(909) <= not((layer0_outputs(1320)) and (layer0_outputs(2114)));
    outputs(910) <= (layer0_outputs(1996)) and not (layer0_outputs(1103));
    outputs(911) <= (layer0_outputs(1855)) and (layer0_outputs(512));
    outputs(912) <= (layer0_outputs(1964)) and (layer0_outputs(617));
    outputs(913) <= not((layer0_outputs(1945)) or (layer0_outputs(1806)));
    outputs(914) <= not((layer0_outputs(2224)) or (layer0_outputs(969)));
    outputs(915) <= not((layer0_outputs(477)) xor (layer0_outputs(1648)));
    outputs(916) <= not((layer0_outputs(589)) xor (layer0_outputs(1346)));
    outputs(917) <= (layer0_outputs(2082)) or (layer0_outputs(2410));
    outputs(918) <= not((layer0_outputs(1144)) or (layer0_outputs(683)));
    outputs(919) <= layer0_outputs(523);
    outputs(920) <= (layer0_outputs(2331)) and (layer0_outputs(1846));
    outputs(921) <= (layer0_outputs(2061)) and not (layer0_outputs(942));
    outputs(922) <= not(layer0_outputs(709));
    outputs(923) <= layer0_outputs(1197);
    outputs(924) <= not(layer0_outputs(378));
    outputs(925) <= not((layer0_outputs(2115)) or (layer0_outputs(2069)));
    outputs(926) <= not((layer0_outputs(820)) or (layer0_outputs(1030)));
    outputs(927) <= not(layer0_outputs(1235));
    outputs(928) <= layer0_outputs(1203);
    outputs(929) <= (layer0_outputs(1726)) or (layer0_outputs(1237));
    outputs(930) <= layer0_outputs(1150);
    outputs(931) <= not(layer0_outputs(339));
    outputs(932) <= not(layer0_outputs(461)) or (layer0_outputs(2465));
    outputs(933) <= layer0_outputs(2189);
    outputs(934) <= not(layer0_outputs(2476));
    outputs(935) <= not(layer0_outputs(1817)) or (layer0_outputs(1577));
    outputs(936) <= not(layer0_outputs(1195)) or (layer0_outputs(881));
    outputs(937) <= (layer0_outputs(77)) xor (layer0_outputs(1925));
    outputs(938) <= not(layer0_outputs(1625));
    outputs(939) <= not(layer0_outputs(2526));
    outputs(940) <= not((layer0_outputs(1356)) xor (layer0_outputs(1672)));
    outputs(941) <= layer0_outputs(40);
    outputs(942) <= not(layer0_outputs(825));
    outputs(943) <= not(layer0_outputs(1872));
    outputs(944) <= (layer0_outputs(2003)) and not (layer0_outputs(615));
    outputs(945) <= not((layer0_outputs(1973)) and (layer0_outputs(2373)));
    outputs(946) <= not(layer0_outputs(381)) or (layer0_outputs(17));
    outputs(947) <= (layer0_outputs(1712)) or (layer0_outputs(1433));
    outputs(948) <= (layer0_outputs(1122)) and not (layer0_outputs(1087));
    outputs(949) <= layer0_outputs(1567);
    outputs(950) <= (layer0_outputs(2494)) and not (layer0_outputs(2501));
    outputs(951) <= (layer0_outputs(159)) and not (layer0_outputs(1175));
    outputs(952) <= (layer0_outputs(1509)) and not (layer0_outputs(1071));
    outputs(953) <= not(layer0_outputs(1345)) or (layer0_outputs(1549));
    outputs(954) <= (layer0_outputs(1404)) and (layer0_outputs(1793));
    outputs(955) <= layer0_outputs(2237);
    outputs(956) <= (layer0_outputs(826)) and not (layer0_outputs(2213));
    outputs(957) <= (layer0_outputs(290)) and not (layer0_outputs(1940));
    outputs(958) <= (layer0_outputs(1425)) and not (layer0_outputs(2499));
    outputs(959) <= not(layer0_outputs(437)) or (layer0_outputs(2192));
    outputs(960) <= not(layer0_outputs(300));
    outputs(961) <= layer0_outputs(1222);
    outputs(962) <= layer0_outputs(2228);
    outputs(963) <= (layer0_outputs(733)) and not (layer0_outputs(1780));
    outputs(964) <= layer0_outputs(1029);
    outputs(965) <= (layer0_outputs(163)) and not (layer0_outputs(1533));
    outputs(966) <= not(layer0_outputs(1267)) or (layer0_outputs(1075));
    outputs(967) <= not(layer0_outputs(862)) or (layer0_outputs(224));
    outputs(968) <= (layer0_outputs(1209)) and not (layer0_outputs(2356));
    outputs(969) <= (layer0_outputs(1122)) and (layer0_outputs(1798));
    outputs(970) <= (layer0_outputs(1655)) and (layer0_outputs(2339));
    outputs(971) <= (layer0_outputs(1541)) and not (layer0_outputs(1570));
    outputs(972) <= (layer0_outputs(326)) and not (layer0_outputs(1279));
    outputs(973) <= not(layer0_outputs(2487));
    outputs(974) <= (layer0_outputs(1485)) and not (layer0_outputs(431));
    outputs(975) <= not((layer0_outputs(1869)) or (layer0_outputs(178)));
    outputs(976) <= not((layer0_outputs(2434)) or (layer0_outputs(371)));
    outputs(977) <= not(layer0_outputs(2493));
    outputs(978) <= not((layer0_outputs(257)) or (layer0_outputs(1270)));
    outputs(979) <= (layer0_outputs(2066)) and not (layer0_outputs(2094));
    outputs(980) <= not((layer0_outputs(387)) and (layer0_outputs(377)));
    outputs(981) <= (layer0_outputs(1461)) and not (layer0_outputs(2043));
    outputs(982) <= layer0_outputs(386);
    outputs(983) <= (layer0_outputs(697)) and (layer0_outputs(1581));
    outputs(984) <= layer0_outputs(2509);
    outputs(985) <= not(layer0_outputs(2371));
    outputs(986) <= not((layer0_outputs(1939)) or (layer0_outputs(1366)));
    outputs(987) <= layer0_outputs(1024);
    outputs(988) <= (layer0_outputs(1825)) and (layer0_outputs(2287));
    outputs(989) <= not((layer0_outputs(331)) or (layer0_outputs(1735)));
    outputs(990) <= not((layer0_outputs(2233)) and (layer0_outputs(852)));
    outputs(991) <= (layer0_outputs(645)) and not (layer0_outputs(343));
    outputs(992) <= (layer0_outputs(539)) and (layer0_outputs(1526));
    outputs(993) <= (layer0_outputs(1304)) or (layer0_outputs(881));
    outputs(994) <= layer0_outputs(1895);
    outputs(995) <= layer0_outputs(1328);
    outputs(996) <= (layer0_outputs(2145)) and not (layer0_outputs(2484));
    outputs(997) <= not(layer0_outputs(2313));
    outputs(998) <= layer0_outputs(174);
    outputs(999) <= not((layer0_outputs(175)) or (layer0_outputs(127)));
    outputs(1000) <= not(layer0_outputs(1270));
    outputs(1001) <= layer0_outputs(2509);
    outputs(1002) <= layer0_outputs(439);
    outputs(1003) <= layer0_outputs(611);
    outputs(1004) <= layer0_outputs(810);
    outputs(1005) <= not(layer0_outputs(1393));
    outputs(1006) <= layer0_outputs(156);
    outputs(1007) <= layer0_outputs(1226);
    outputs(1008) <= layer0_outputs(1765);
    outputs(1009) <= not(layer0_outputs(738));
    outputs(1010) <= not(layer0_outputs(1459)) or (layer0_outputs(134));
    outputs(1011) <= not(layer0_outputs(2421));
    outputs(1012) <= not((layer0_outputs(2198)) or (layer0_outputs(2353)));
    outputs(1013) <= not(layer0_outputs(2176));
    outputs(1014) <= (layer0_outputs(870)) and (layer0_outputs(2333));
    outputs(1015) <= (layer0_outputs(1370)) and not (layer0_outputs(2378));
    outputs(1016) <= layer0_outputs(1510);
    outputs(1017) <= (layer0_outputs(310)) or (layer0_outputs(1387));
    outputs(1018) <= not(layer0_outputs(2469));
    outputs(1019) <= (layer0_outputs(1223)) and not (layer0_outputs(249));
    outputs(1020) <= not(layer0_outputs(2385));
    outputs(1021) <= not(layer0_outputs(1135));
    outputs(1022) <= layer0_outputs(1655);
    outputs(1023) <= (layer0_outputs(149)) and (layer0_outputs(2515));
    outputs(1024) <= layer0_outputs(1482);
    outputs(1025) <= (layer0_outputs(529)) and not (layer0_outputs(662));
    outputs(1026) <= layer0_outputs(1778);
    outputs(1027) <= (layer0_outputs(1773)) or (layer0_outputs(1941));
    outputs(1028) <= (layer0_outputs(2478)) or (layer0_outputs(556));
    outputs(1029) <= (layer0_outputs(655)) and not (layer0_outputs(967));
    outputs(1030) <= (layer0_outputs(1643)) and not (layer0_outputs(2082));
    outputs(1031) <= layer0_outputs(1245);
    outputs(1032) <= not(layer0_outputs(1225));
    outputs(1033) <= layer0_outputs(851);
    outputs(1034) <= (layer0_outputs(889)) and not (layer0_outputs(2417));
    outputs(1035) <= (layer0_outputs(1514)) and not (layer0_outputs(741));
    outputs(1036) <= layer0_outputs(417);
    outputs(1037) <= not(layer0_outputs(636));
    outputs(1038) <= (layer0_outputs(1597)) and not (layer0_outputs(232));
    outputs(1039) <= not(layer0_outputs(405));
    outputs(1040) <= (layer0_outputs(959)) and not (layer0_outputs(1150));
    outputs(1041) <= not(layer0_outputs(1845));
    outputs(1042) <= layer0_outputs(1157);
    outputs(1043) <= layer0_outputs(1477);
    outputs(1044) <= layer0_outputs(1905);
    outputs(1045) <= (layer0_outputs(2100)) and not (layer0_outputs(916));
    outputs(1046) <= (layer0_outputs(2302)) and not (layer0_outputs(769));
    outputs(1047) <= not(layer0_outputs(944));
    outputs(1048) <= (layer0_outputs(1368)) xor (layer0_outputs(971));
    outputs(1049) <= (layer0_outputs(1803)) and not (layer0_outputs(1455));
    outputs(1050) <= (layer0_outputs(488)) and (layer0_outputs(1737));
    outputs(1051) <= not(layer0_outputs(2202));
    outputs(1052) <= layer0_outputs(1203);
    outputs(1053) <= not(layer0_outputs(705));
    outputs(1054) <= not(layer0_outputs(1127));
    outputs(1055) <= not((layer0_outputs(39)) or (layer0_outputs(2481)));
    outputs(1056) <= (layer0_outputs(2432)) and (layer0_outputs(949));
    outputs(1057) <= not((layer0_outputs(293)) or (layer0_outputs(1640)));
    outputs(1058) <= layer0_outputs(2365);
    outputs(1059) <= layer0_outputs(1753);
    outputs(1060) <= layer0_outputs(1255);
    outputs(1061) <= (layer0_outputs(1451)) and not (layer0_outputs(1191));
    outputs(1062) <= layer0_outputs(877);
    outputs(1063) <= not(layer0_outputs(1060));
    outputs(1064) <= (layer0_outputs(363)) and not (layer0_outputs(1190));
    outputs(1065) <= not((layer0_outputs(94)) xor (layer0_outputs(1832)));
    outputs(1066) <= not(layer0_outputs(2411));
    outputs(1067) <= not(layer0_outputs(1896));
    outputs(1068) <= not(layer0_outputs(1994));
    outputs(1069) <= not((layer0_outputs(1152)) or (layer0_outputs(2109)));
    outputs(1070) <= (layer0_outputs(1124)) and (layer0_outputs(1490));
    outputs(1071) <= layer0_outputs(2514);
    outputs(1072) <= layer0_outputs(2188);
    outputs(1073) <= layer0_outputs(50);
    outputs(1074) <= (layer0_outputs(1531)) or (layer0_outputs(2455));
    outputs(1075) <= (layer0_outputs(2420)) and not (layer0_outputs(213));
    outputs(1076) <= not((layer0_outputs(685)) or (layer0_outputs(2229)));
    outputs(1077) <= (layer0_outputs(112)) and (layer0_outputs(1562));
    outputs(1078) <= layer0_outputs(1268);
    outputs(1079) <= not(layer0_outputs(132));
    outputs(1080) <= layer0_outputs(135);
    outputs(1081) <= (layer0_outputs(2405)) and not (layer0_outputs(1571));
    outputs(1082) <= not((layer0_outputs(753)) xor (layer0_outputs(506)));
    outputs(1083) <= (layer0_outputs(2559)) or (layer0_outputs(900));
    outputs(1084) <= not(layer0_outputs(1440));
    outputs(1085) <= (layer0_outputs(1607)) and not (layer0_outputs(929));
    outputs(1086) <= not((layer0_outputs(438)) or (layer0_outputs(2006)));
    outputs(1087) <= (layer0_outputs(576)) and not (layer0_outputs(1176));
    outputs(1088) <= (layer0_outputs(2198)) and not (layer0_outputs(423));
    outputs(1089) <= (layer0_outputs(353)) and (layer0_outputs(1407));
    outputs(1090) <= (layer0_outputs(627)) and not (layer0_outputs(2315));
    outputs(1091) <= not((layer0_outputs(406)) or (layer0_outputs(1521)));
    outputs(1092) <= (layer0_outputs(2208)) and not (layer0_outputs(1064));
    outputs(1093) <= layer0_outputs(970);
    outputs(1094) <= (layer0_outputs(1969)) and (layer0_outputs(563));
    outputs(1095) <= not((layer0_outputs(697)) or (layer0_outputs(521)));
    outputs(1096) <= not(layer0_outputs(1377));
    outputs(1097) <= layer0_outputs(258);
    outputs(1098) <= layer0_outputs(1049);
    outputs(1099) <= (layer0_outputs(1596)) and not (layer0_outputs(732));
    outputs(1100) <= not((layer0_outputs(2095)) or (layer0_outputs(1746)));
    outputs(1101) <= not(layer0_outputs(1309));
    outputs(1102) <= (layer0_outputs(1128)) and not (layer0_outputs(906));
    outputs(1103) <= (layer0_outputs(1917)) and not (layer0_outputs(841));
    outputs(1104) <= not(layer0_outputs(1913));
    outputs(1105) <= layer0_outputs(1532);
    outputs(1106) <= not(layer0_outputs(2211));
    outputs(1107) <= not(layer0_outputs(967));
    outputs(1108) <= layer0_outputs(555);
    outputs(1109) <= (layer0_outputs(1180)) and (layer0_outputs(172));
    outputs(1110) <= not((layer0_outputs(1001)) or (layer0_outputs(2360)));
    outputs(1111) <= (layer0_outputs(1116)) and not (layer0_outputs(289));
    outputs(1112) <= not(layer0_outputs(800));
    outputs(1113) <= not((layer0_outputs(264)) and (layer0_outputs(1704)));
    outputs(1114) <= not(layer0_outputs(1441));
    outputs(1115) <= not(layer0_outputs(1520));
    outputs(1116) <= (layer0_outputs(1115)) and (layer0_outputs(2425));
    outputs(1117) <= layer0_outputs(303);
    outputs(1118) <= not((layer0_outputs(2412)) or (layer0_outputs(1444)));
    outputs(1119) <= not(layer0_outputs(1678));
    outputs(1120) <= not((layer0_outputs(2182)) or (layer0_outputs(1938)));
    outputs(1121) <= layer0_outputs(601);
    outputs(1122) <= not(layer0_outputs(392));
    outputs(1123) <= not(layer0_outputs(1588));
    outputs(1124) <= (layer0_outputs(514)) and not (layer0_outputs(752));
    outputs(1125) <= layer0_outputs(462);
    outputs(1126) <= layer0_outputs(2057);
    outputs(1127) <= (layer0_outputs(283)) and not (layer0_outputs(862));
    outputs(1128) <= layer0_outputs(1533);
    outputs(1129) <= (layer0_outputs(599)) and not (layer0_outputs(757));
    outputs(1130) <= not(layer0_outputs(802));
    outputs(1131) <= (layer0_outputs(1680)) and not (layer0_outputs(671));
    outputs(1132) <= (layer0_outputs(808)) and not (layer0_outputs(1672));
    outputs(1133) <= (layer0_outputs(1436)) and not (layer0_outputs(694));
    outputs(1134) <= (layer0_outputs(696)) xor (layer0_outputs(2462));
    outputs(1135) <= not(layer0_outputs(20));
    outputs(1136) <= (layer0_outputs(2382)) and not (layer0_outputs(99));
    outputs(1137) <= layer0_outputs(608);
    outputs(1138) <= (layer0_outputs(419)) xor (layer0_outputs(1864));
    outputs(1139) <= (layer0_outputs(1597)) and not (layer0_outputs(1075));
    outputs(1140) <= layer0_outputs(897);
    outputs(1141) <= layer0_outputs(2171);
    outputs(1142) <= (layer0_outputs(1764)) and not (layer0_outputs(1458));
    outputs(1143) <= (layer0_outputs(1239)) or (layer0_outputs(973));
    outputs(1144) <= not(layer0_outputs(126)) or (layer0_outputs(131));
    outputs(1145) <= layer0_outputs(1101);
    outputs(1146) <= (layer0_outputs(872)) and (layer0_outputs(1146));
    outputs(1147) <= (layer0_outputs(2083)) and not (layer0_outputs(80));
    outputs(1148) <= not((layer0_outputs(34)) xor (layer0_outputs(2154)));
    outputs(1149) <= (layer0_outputs(2069)) and (layer0_outputs(943));
    outputs(1150) <= (layer0_outputs(125)) and (layer0_outputs(2543));
    outputs(1151) <= layer0_outputs(1519);
    outputs(1152) <= (layer0_outputs(1157)) and not (layer0_outputs(1851));
    outputs(1153) <= not((layer0_outputs(867)) or (layer0_outputs(2345)));
    outputs(1154) <= layer0_outputs(1158);
    outputs(1155) <= (layer0_outputs(248)) and not (layer0_outputs(1524));
    outputs(1156) <= not(layer0_outputs(347));
    outputs(1157) <= (layer0_outputs(795)) and not (layer0_outputs(439));
    outputs(1158) <= layer0_outputs(664);
    outputs(1159) <= (layer0_outputs(970)) and (layer0_outputs(550));
    outputs(1160) <= not(layer0_outputs(1755));
    outputs(1161) <= (layer0_outputs(2529)) and not (layer0_outputs(2429));
    outputs(1162) <= not(layer0_outputs(610)) or (layer0_outputs(1519));
    outputs(1163) <= not(layer0_outputs(2036));
    outputs(1164) <= layer0_outputs(1560);
    outputs(1165) <= (layer0_outputs(734)) and (layer0_outputs(112));
    outputs(1166) <= not(layer0_outputs(1207));
    outputs(1167) <= (layer0_outputs(356)) xor (layer0_outputs(360));
    outputs(1168) <= (layer0_outputs(2513)) and not (layer0_outputs(2125));
    outputs(1169) <= (layer0_outputs(2271)) and not (layer0_outputs(1671));
    outputs(1170) <= layer0_outputs(1193);
    outputs(1171) <= (layer0_outputs(607)) xor (layer0_outputs(1677));
    outputs(1172) <= layer0_outputs(1276);
    outputs(1173) <= not(layer0_outputs(1885));
    outputs(1174) <= layer0_outputs(1943);
    outputs(1175) <= layer0_outputs(748);
    outputs(1176) <= (layer0_outputs(816)) and not (layer0_outputs(2192));
    outputs(1177) <= not((layer0_outputs(1583)) and (layer0_outputs(1287)));
    outputs(1178) <= not(layer0_outputs(735));
    outputs(1179) <= not(layer0_outputs(805)) or (layer0_outputs(938));
    outputs(1180) <= (layer0_outputs(1021)) and not (layer0_outputs(146));
    outputs(1181) <= not(layer0_outputs(2140)) or (layer0_outputs(68));
    outputs(1182) <= (layer0_outputs(445)) or (layer0_outputs(241));
    outputs(1183) <= (layer0_outputs(458)) and not (layer0_outputs(543));
    outputs(1184) <= layer0_outputs(1488);
    outputs(1185) <= (layer0_outputs(849)) and not (layer0_outputs(2164));
    outputs(1186) <= not(layer0_outputs(2072)) or (layer0_outputs(1838));
    outputs(1187) <= not((layer0_outputs(1525)) or (layer0_outputs(2109)));
    outputs(1188) <= layer0_outputs(1217);
    outputs(1189) <= (layer0_outputs(609)) and (layer0_outputs(397));
    outputs(1190) <= (layer0_outputs(843)) and not (layer0_outputs(361));
    outputs(1191) <= not(layer0_outputs(1767));
    outputs(1192) <= not((layer0_outputs(592)) and (layer0_outputs(679)));
    outputs(1193) <= (layer0_outputs(1456)) and (layer0_outputs(1829));
    outputs(1194) <= layer0_outputs(1014);
    outputs(1195) <= (layer0_outputs(514)) and not (layer0_outputs(2187));
    outputs(1196) <= not((layer0_outputs(24)) or (layer0_outputs(452)));
    outputs(1197) <= layer0_outputs(2357);
    outputs(1198) <= (layer0_outputs(42)) and not (layer0_outputs(588));
    outputs(1199) <= (layer0_outputs(140)) and (layer0_outputs(2389));
    outputs(1200) <= layer0_outputs(2041);
    outputs(1201) <= (layer0_outputs(560)) and not (layer0_outputs(1200));
    outputs(1202) <= (layer0_outputs(2537)) or (layer0_outputs(1878));
    outputs(1203) <= not(layer0_outputs(1179));
    outputs(1204) <= not(layer0_outputs(2202)) or (layer0_outputs(1586));
    outputs(1205) <= not(layer0_outputs(656));
    outputs(1206) <= layer0_outputs(58);
    outputs(1207) <= not((layer0_outputs(208)) xor (layer0_outputs(2553)));
    outputs(1208) <= not(layer0_outputs(455));
    outputs(1209) <= (layer0_outputs(2536)) and not (layer0_outputs(1409));
    outputs(1210) <= not(layer0_outputs(444));
    outputs(1211) <= (layer0_outputs(1003)) and not (layer0_outputs(2554));
    outputs(1212) <= not((layer0_outputs(1177)) xor (layer0_outputs(1396)));
    outputs(1213) <= (layer0_outputs(1975)) and (layer0_outputs(1987));
    outputs(1214) <= not(layer0_outputs(807));
    outputs(1215) <= layer0_outputs(1582);
    outputs(1216) <= (layer0_outputs(1688)) and (layer0_outputs(978));
    outputs(1217) <= not((layer0_outputs(1982)) or (layer0_outputs(1708)));
    outputs(1218) <= (layer0_outputs(472)) and not (layer0_outputs(1716));
    outputs(1219) <= not((layer0_outputs(2299)) or (layer0_outputs(2457)));
    outputs(1220) <= layer0_outputs(98);
    outputs(1221) <= not(layer0_outputs(1324));
    outputs(1222) <= layer0_outputs(1593);
    outputs(1223) <= layer0_outputs(462);
    outputs(1224) <= (layer0_outputs(1329)) and (layer0_outputs(1977));
    outputs(1225) <= not(layer0_outputs(204));
    outputs(1226) <= not((layer0_outputs(1495)) or (layer0_outputs(804)));
    outputs(1227) <= not(layer0_outputs(2370));
    outputs(1228) <= (layer0_outputs(2492)) and not (layer0_outputs(976));
    outputs(1229) <= layer0_outputs(1639);
    outputs(1230) <= (layer0_outputs(1527)) or (layer0_outputs(2537));
    outputs(1231) <= not((layer0_outputs(2436)) or (layer0_outputs(1785)));
    outputs(1232) <= (layer0_outputs(11)) and (layer0_outputs(2));
    outputs(1233) <= layer0_outputs(896);
    outputs(1234) <= not((layer0_outputs(1419)) and (layer0_outputs(1903)));
    outputs(1235) <= not((layer0_outputs(2545)) or (layer0_outputs(728)));
    outputs(1236) <= not(layer0_outputs(2418));
    outputs(1237) <= not((layer0_outputs(73)) or (layer0_outputs(1376)));
    outputs(1238) <= not((layer0_outputs(1946)) or (layer0_outputs(1098)));
    outputs(1239) <= not(layer0_outputs(1825));
    outputs(1240) <= layer0_outputs(784);
    outputs(1241) <= not(layer0_outputs(400)) or (layer0_outputs(1916));
    outputs(1242) <= layer0_outputs(31);
    outputs(1243) <= not(layer0_outputs(1567));
    outputs(1244) <= not(layer0_outputs(120));
    outputs(1245) <= (layer0_outputs(2455)) and not (layer0_outputs(866));
    outputs(1246) <= not(layer0_outputs(2423));
    outputs(1247) <= layer0_outputs(2413);
    outputs(1248) <= (layer0_outputs(606)) and (layer0_outputs(1977));
    outputs(1249) <= (layer0_outputs(424)) and (layer0_outputs(1314));
    outputs(1250) <= not(layer0_outputs(389));
    outputs(1251) <= not((layer0_outputs(2282)) and (layer0_outputs(663)));
    outputs(1252) <= (layer0_outputs(1117)) and (layer0_outputs(1259));
    outputs(1253) <= not(layer0_outputs(1509));
    outputs(1254) <= not(layer0_outputs(670));
    outputs(1255) <= (layer0_outputs(782)) and not (layer0_outputs(2174));
    outputs(1256) <= layer0_outputs(1623);
    outputs(1257) <= not(layer0_outputs(1159));
    outputs(1258) <= not(layer0_outputs(1032));
    outputs(1259) <= not(layer0_outputs(2402)) or (layer0_outputs(644));
    outputs(1260) <= layer0_outputs(717);
    outputs(1261) <= not(layer0_outputs(2185)) or (layer0_outputs(2532));
    outputs(1262) <= layer0_outputs(2018);
    outputs(1263) <= layer0_outputs(2223);
    outputs(1264) <= (layer0_outputs(921)) and (layer0_outputs(638));
    outputs(1265) <= layer0_outputs(1561);
    outputs(1266) <= not((layer0_outputs(364)) xor (layer0_outputs(94)));
    outputs(1267) <= (layer0_outputs(2003)) and (layer0_outputs(803));
    outputs(1268) <= (layer0_outputs(243)) and (layer0_outputs(321));
    outputs(1269) <= (layer0_outputs(584)) and not (layer0_outputs(1045));
    outputs(1270) <= not((layer0_outputs(44)) or (layer0_outputs(1118)));
    outputs(1271) <= not((layer0_outputs(1493)) or (layer0_outputs(2472)));
    outputs(1272) <= layer0_outputs(188);
    outputs(1273) <= not(layer0_outputs(2172)) or (layer0_outputs(480));
    outputs(1274) <= layer0_outputs(1502);
    outputs(1275) <= not(layer0_outputs(2226));
    outputs(1276) <= not(layer0_outputs(400));
    outputs(1277) <= not(layer0_outputs(2259));
    outputs(1278) <= layer0_outputs(1316);
    outputs(1279) <= not((layer0_outputs(1410)) and (layer0_outputs(610)));
    outputs(1280) <= (layer0_outputs(1378)) and not (layer0_outputs(1764));
    outputs(1281) <= not(layer0_outputs(1687)) or (layer0_outputs(2358));
    outputs(1282) <= layer0_outputs(1599);
    outputs(1283) <= not((layer0_outputs(2348)) or (layer0_outputs(1006)));
    outputs(1284) <= not(layer0_outputs(2264));
    outputs(1285) <= not(layer0_outputs(925)) or (layer0_outputs(1388));
    outputs(1286) <= (layer0_outputs(1605)) and not (layer0_outputs(1238));
    outputs(1287) <= not((layer0_outputs(2444)) and (layer0_outputs(580)));
    outputs(1288) <= layer0_outputs(1727);
    outputs(1289) <= (layer0_outputs(1466)) and (layer0_outputs(846));
    outputs(1290) <= not(layer0_outputs(195)) or (layer0_outputs(1033));
    outputs(1291) <= layer0_outputs(2398);
    outputs(1292) <= not(layer0_outputs(1717));
    outputs(1293) <= not((layer0_outputs(2004)) xor (layer0_outputs(1999)));
    outputs(1294) <= (layer0_outputs(1231)) and (layer0_outputs(597));
    outputs(1295) <= (layer0_outputs(1002)) and not (layer0_outputs(888));
    outputs(1296) <= (layer0_outputs(1976)) and (layer0_outputs(1125));
    outputs(1297) <= not(layer0_outputs(322));
    outputs(1298) <= (layer0_outputs(712)) and not (layer0_outputs(2359));
    outputs(1299) <= layer0_outputs(2276);
    outputs(1300) <= layer0_outputs(1638);
    outputs(1301) <= layer0_outputs(2305);
    outputs(1302) <= not((layer0_outputs(1692)) or (layer0_outputs(1838)));
    outputs(1303) <= not(layer0_outputs(1246));
    outputs(1304) <= (layer0_outputs(760)) and not (layer0_outputs(1465));
    outputs(1305) <= (layer0_outputs(192)) and not (layer0_outputs(1400));
    outputs(1306) <= not(layer0_outputs(1191)) or (layer0_outputs(2487));
    outputs(1307) <= not((layer0_outputs(1043)) xor (layer0_outputs(412)));
    outputs(1308) <= not(layer0_outputs(1310));
    outputs(1309) <= not(layer0_outputs(1028)) or (layer0_outputs(561));
    outputs(1310) <= (layer0_outputs(2529)) xor (layer0_outputs(2431));
    outputs(1311) <= layer0_outputs(1308);
    outputs(1312) <= not(layer0_outputs(924));
    outputs(1313) <= not(layer0_outputs(1916));
    outputs(1314) <= layer0_outputs(167);
    outputs(1315) <= not(layer0_outputs(145));
    outputs(1316) <= not(layer0_outputs(1006));
    outputs(1317) <= (layer0_outputs(937)) and (layer0_outputs(484));
    outputs(1318) <= not(layer0_outputs(1757));
    outputs(1319) <= (layer0_outputs(2041)) xor (layer0_outputs(388));
    outputs(1320) <= layer0_outputs(344);
    outputs(1321) <= (layer0_outputs(1682)) xor (layer0_outputs(339));
    outputs(1322) <= not((layer0_outputs(859)) xor (layer0_outputs(1490)));
    outputs(1323) <= not((layer0_outputs(678)) and (layer0_outputs(27)));
    outputs(1324) <= (layer0_outputs(1032)) xor (layer0_outputs(1450));
    outputs(1325) <= not(layer0_outputs(566)) or (layer0_outputs(1768));
    outputs(1326) <= not(layer0_outputs(23));
    outputs(1327) <= not(layer0_outputs(2030));
    outputs(1328) <= layer0_outputs(773);
    outputs(1329) <= (layer0_outputs(1046)) and not (layer0_outputs(150));
    outputs(1330) <= not(layer0_outputs(1285));
    outputs(1331) <= not((layer0_outputs(759)) or (layer0_outputs(2501)));
    outputs(1332) <= layer0_outputs(1142);
    outputs(1333) <= not((layer0_outputs(2359)) or (layer0_outputs(1853)));
    outputs(1334) <= (layer0_outputs(28)) and not (layer0_outputs(70));
    outputs(1335) <= not(layer0_outputs(2369)) or (layer0_outputs(1547));
    outputs(1336) <= not((layer0_outputs(189)) or (layer0_outputs(723)));
    outputs(1337) <= not((layer0_outputs(579)) or (layer0_outputs(2119)));
    outputs(1338) <= not((layer0_outputs(1023)) or (layer0_outputs(1572)));
    outputs(1339) <= layer0_outputs(305);
    outputs(1340) <= not(layer0_outputs(1950));
    outputs(1341) <= not((layer0_outputs(739)) or (layer0_outputs(680)));
    outputs(1342) <= not(layer0_outputs(184));
    outputs(1343) <= (layer0_outputs(1949)) or (layer0_outputs(1241));
    outputs(1344) <= not(layer0_outputs(1643)) or (layer0_outputs(1272));
    outputs(1345) <= layer0_outputs(854);
    outputs(1346) <= not((layer0_outputs(2490)) or (layer0_outputs(2480)));
    outputs(1347) <= not((layer0_outputs(676)) xor (layer0_outputs(1595)));
    outputs(1348) <= (layer0_outputs(1460)) and not (layer0_outputs(2442));
    outputs(1349) <= (layer0_outputs(890)) and not (layer0_outputs(2027));
    outputs(1350) <= not((layer0_outputs(2235)) xor (layer0_outputs(1867)));
    outputs(1351) <= not(layer0_outputs(294)) or (layer0_outputs(43));
    outputs(1352) <= not((layer0_outputs(512)) or (layer0_outputs(2122)));
    outputs(1353) <= not((layer0_outputs(150)) or (layer0_outputs(1458)));
    outputs(1354) <= not((layer0_outputs(65)) and (layer0_outputs(599)));
    outputs(1355) <= not(layer0_outputs(1205));
    outputs(1356) <= (layer0_outputs(1879)) xor (layer0_outputs(2307));
    outputs(1357) <= layer0_outputs(864);
    outputs(1358) <= not(layer0_outputs(1069));
    outputs(1359) <= (layer0_outputs(205)) and (layer0_outputs(342));
    outputs(1360) <= not((layer0_outputs(974)) or (layer0_outputs(384)));
    outputs(1361) <= layer0_outputs(194);
    outputs(1362) <= (layer0_outputs(429)) and (layer0_outputs(397));
    outputs(1363) <= not(layer0_outputs(1462));
    outputs(1364) <= (layer0_outputs(1353)) and not (layer0_outputs(2252));
    outputs(1365) <= layer0_outputs(990);
    outputs(1366) <= not(layer0_outputs(1497));
    outputs(1367) <= (layer0_outputs(2374)) and not (layer0_outputs(1366));
    outputs(1368) <= not(layer0_outputs(1099)) or (layer0_outputs(318));
    outputs(1369) <= (layer0_outputs(1042)) and not (layer0_outputs(1810));
    outputs(1370) <= not(layer0_outputs(527));
    outputs(1371) <= (layer0_outputs(643)) and (layer0_outputs(1926));
    outputs(1372) <= (layer0_outputs(363)) xor (layer0_outputs(672));
    outputs(1373) <= (layer0_outputs(520)) and (layer0_outputs(682));
    outputs(1374) <= not(layer0_outputs(1548));
    outputs(1375) <= not(layer0_outputs(580));
    outputs(1376) <= (layer0_outputs(1779)) or (layer0_outputs(2334));
    outputs(1377) <= layer0_outputs(573);
    outputs(1378) <= not((layer0_outputs(2117)) and (layer0_outputs(667)));
    outputs(1379) <= (layer0_outputs(522)) or (layer0_outputs(1867));
    outputs(1380) <= (layer0_outputs(95)) xor (layer0_outputs(392));
    outputs(1381) <= (layer0_outputs(1779)) or (layer0_outputs(320));
    outputs(1382) <= not((layer0_outputs(2100)) or (layer0_outputs(850)));
    outputs(1383) <= (layer0_outputs(452)) and not (layer0_outputs(2230));
    outputs(1384) <= layer0_outputs(525);
    outputs(1385) <= not((layer0_outputs(1906)) xor (layer0_outputs(1537)));
    outputs(1386) <= layer0_outputs(374);
    outputs(1387) <= (layer0_outputs(1045)) xor (layer0_outputs(2046));
    outputs(1388) <= not((layer0_outputs(394)) xor (layer0_outputs(2416)));
    outputs(1389) <= layer0_outputs(2317);
    outputs(1390) <= layer0_outputs(130);
    outputs(1391) <= not(layer0_outputs(386));
    outputs(1392) <= not(layer0_outputs(1887));
    outputs(1393) <= layer0_outputs(1274);
    outputs(1394) <= not(layer0_outputs(2482));
    outputs(1395) <= not(layer0_outputs(2544)) or (layer0_outputs(2290));
    outputs(1396) <= (layer0_outputs(572)) and (layer0_outputs(1213));
    outputs(1397) <= layer0_outputs(2305);
    outputs(1398) <= (layer0_outputs(1718)) or (layer0_outputs(97));
    outputs(1399) <= (layer0_outputs(1928)) and not (layer0_outputs(129));
    outputs(1400) <= layer0_outputs(75);
    outputs(1401) <= (layer0_outputs(291)) and (layer0_outputs(520));
    outputs(1402) <= not((layer0_outputs(377)) or (layer0_outputs(1995)));
    outputs(1403) <= not(layer0_outputs(465));
    outputs(1404) <= not(layer0_outputs(1679));
    outputs(1405) <= not(layer0_outputs(2114)) or (layer0_outputs(798));
    outputs(1406) <= (layer0_outputs(2539)) and not (layer0_outputs(2341));
    outputs(1407) <= layer0_outputs(2058);
    outputs(1408) <= not(layer0_outputs(1550));
    outputs(1409) <= not(layer0_outputs(1));
    outputs(1410) <= layer0_outputs(1566);
    outputs(1411) <= not((layer0_outputs(446)) or (layer0_outputs(1066)));
    outputs(1412) <= not(layer0_outputs(1670));
    outputs(1413) <= not((layer0_outputs(86)) xor (layer0_outputs(696)));
    outputs(1414) <= layer0_outputs(414);
    outputs(1415) <= (layer0_outputs(6)) and not (layer0_outputs(1797));
    outputs(1416) <= not((layer0_outputs(471)) xor (layer0_outputs(913)));
    outputs(1417) <= not(layer0_outputs(1610));
    outputs(1418) <= not(layer0_outputs(537));
    outputs(1419) <= not(layer0_outputs(1027)) or (layer0_outputs(214));
    outputs(1420) <= not(layer0_outputs(48));
    outputs(1421) <= not(layer0_outputs(1837));
    outputs(1422) <= not((layer0_outputs(416)) xor (layer0_outputs(1632)));
    outputs(1423) <= layer0_outputs(701);
    outputs(1424) <= layer0_outputs(896);
    outputs(1425) <= layer0_outputs(2520);
    outputs(1426) <= layer0_outputs(2325);
    outputs(1427) <= layer0_outputs(340);
    outputs(1428) <= (layer0_outputs(22)) and not (layer0_outputs(2207));
    outputs(1429) <= layer0_outputs(2300);
    outputs(1430) <= not((layer0_outputs(1077)) or (layer0_outputs(482)));
    outputs(1431) <= not(layer0_outputs(1220));
    outputs(1432) <= (layer0_outputs(1079)) and not (layer0_outputs(1988));
    outputs(1433) <= layer0_outputs(22);
    outputs(1434) <= not((layer0_outputs(980)) and (layer0_outputs(1756)));
    outputs(1435) <= not((layer0_outputs(2239)) xor (layer0_outputs(379)));
    outputs(1436) <= not(layer0_outputs(524));
    outputs(1437) <= not((layer0_outputs(844)) or (layer0_outputs(942)));
    outputs(1438) <= not(layer0_outputs(1187)) or (layer0_outputs(177));
    outputs(1439) <= (layer0_outputs(876)) or (layer0_outputs(1363));
    outputs(1440) <= (layer0_outputs(2278)) xor (layer0_outputs(218));
    outputs(1441) <= not(layer0_outputs(1408));
    outputs(1442) <= (layer0_outputs(1328)) xor (layer0_outputs(33));
    outputs(1443) <= (layer0_outputs(2548)) xor (layer0_outputs(1665));
    outputs(1444) <= (layer0_outputs(1284)) and not (layer0_outputs(1064));
    outputs(1445) <= (layer0_outputs(2178)) xor (layer0_outputs(101));
    outputs(1446) <= layer0_outputs(1740);
    outputs(1447) <= not(layer0_outputs(2551));
    outputs(1448) <= not((layer0_outputs(2138)) or (layer0_outputs(41)));
    outputs(1449) <= layer0_outputs(960);
    outputs(1450) <= not(layer0_outputs(173));
    outputs(1451) <= (layer0_outputs(1333)) and not (layer0_outputs(1498));
    outputs(1452) <= not(layer0_outputs(875));
    outputs(1453) <= not(layer0_outputs(2203));
    outputs(1454) <= layer0_outputs(894);
    outputs(1455) <= (layer0_outputs(2244)) and not (layer0_outputs(2552));
    outputs(1456) <= (layer0_outputs(1518)) xor (layer0_outputs(2131));
    outputs(1457) <= layer0_outputs(622);
    outputs(1458) <= layer0_outputs(221);
    outputs(1459) <= (layer0_outputs(1046)) or (layer0_outputs(920));
    outputs(1460) <= (layer0_outputs(529)) xor (layer0_outputs(1565));
    outputs(1461) <= (layer0_outputs(2493)) and not (layer0_outputs(155));
    outputs(1462) <= (layer0_outputs(1937)) and (layer0_outputs(1302));
    outputs(1463) <= layer0_outputs(749);
    outputs(1464) <= (layer0_outputs(1731)) or (layer0_outputs(825));
    outputs(1465) <= (layer0_outputs(442)) xor (layer0_outputs(1467));
    outputs(1466) <= not((layer0_outputs(533)) xor (layer0_outputs(2430)));
    outputs(1467) <= (layer0_outputs(2364)) and not (layer0_outputs(2200));
    outputs(1468) <= (layer0_outputs(689)) and not (layer0_outputs(224));
    outputs(1469) <= not((layer0_outputs(1181)) xor (layer0_outputs(2349)));
    outputs(1470) <= not(layer0_outputs(39)) or (layer0_outputs(1861));
    outputs(1471) <= layer0_outputs(194);
    outputs(1472) <= not(layer0_outputs(2347)) or (layer0_outputs(1085));
    outputs(1473) <= not((layer0_outputs(2181)) or (layer0_outputs(371)));
    outputs(1474) <= (layer0_outputs(1627)) xor (layer0_outputs(543));
    outputs(1475) <= layer0_outputs(447);
    outputs(1476) <= not(layer0_outputs(1732));
    outputs(1477) <= (layer0_outputs(2162)) and not (layer0_outputs(1026));
    outputs(1478) <= not(layer0_outputs(2375)) or (layer0_outputs(2165));
    outputs(1479) <= not((layer0_outputs(478)) xor (layer0_outputs(1912)));
    outputs(1480) <= (layer0_outputs(1716)) and not (layer0_outputs(2195));
    outputs(1481) <= (layer0_outputs(1792)) and (layer0_outputs(689));
    outputs(1482) <= layer0_outputs(1522);
    outputs(1483) <= not(layer0_outputs(1520)) or (layer0_outputs(1574));
    outputs(1484) <= not((layer0_outputs(873)) xor (layer0_outputs(53)));
    outputs(1485) <= not(layer0_outputs(1057));
    outputs(1486) <= not(layer0_outputs(2020));
    outputs(1487) <= (layer0_outputs(287)) or (layer0_outputs(1475));
    outputs(1488) <= not(layer0_outputs(789));
    outputs(1489) <= (layer0_outputs(2071)) and not (layer0_outputs(986));
    outputs(1490) <= not(layer0_outputs(884));
    outputs(1491) <= not(layer0_outputs(1844));
    outputs(1492) <= (layer0_outputs(1378)) and not (layer0_outputs(48));
    outputs(1493) <= (layer0_outputs(2372)) and not (layer0_outputs(2032));
    outputs(1494) <= layer0_outputs(934);
    outputs(1495) <= (layer0_outputs(666)) and (layer0_outputs(1479));
    outputs(1496) <= layer0_outputs(43);
    outputs(1497) <= not((layer0_outputs(1370)) or (layer0_outputs(45)));
    outputs(1498) <= layer0_outputs(1212);
    outputs(1499) <= not((layer0_outputs(812)) and (layer0_outputs(1794)));
    outputs(1500) <= (layer0_outputs(1438)) and (layer0_outputs(1340));
    outputs(1501) <= not((layer0_outputs(1696)) xor (layer0_outputs(2094)));
    outputs(1502) <= (layer0_outputs(726)) and not (layer0_outputs(2306));
    outputs(1503) <= layer0_outputs(268);
    outputs(1504) <= layer0_outputs(1628);
    outputs(1505) <= layer0_outputs(545);
    outputs(1506) <= not(layer0_outputs(975));
    outputs(1507) <= (layer0_outputs(2333)) xor (layer0_outputs(1192));
    outputs(1508) <= layer0_outputs(2463);
    outputs(1509) <= layer0_outputs(1457);
    outputs(1510) <= not(layer0_outputs(226));
    outputs(1511) <= (layer0_outputs(506)) and not (layer0_outputs(14));
    outputs(1512) <= not(layer0_outputs(261)) or (layer0_outputs(996));
    outputs(1513) <= layer0_outputs(2422);
    outputs(1514) <= layer0_outputs(1499);
    outputs(1515) <= layer0_outputs(611);
    outputs(1516) <= (layer0_outputs(1582)) and not (layer0_outputs(2470));
    outputs(1517) <= (layer0_outputs(2070)) and not (layer0_outputs(470));
    outputs(1518) <= layer0_outputs(1644);
    outputs(1519) <= layer0_outputs(921);
    outputs(1520) <= (layer0_outputs(1759)) xor (layer0_outputs(1514));
    outputs(1521) <= (layer0_outputs(813)) and not (layer0_outputs(118));
    outputs(1522) <= not((layer0_outputs(1909)) or (layer0_outputs(359)));
    outputs(1523) <= layer0_outputs(1768);
    outputs(1524) <= not(layer0_outputs(885));
    outputs(1525) <= (layer0_outputs(294)) xor (layer0_outputs(1723));
    outputs(1526) <= not((layer0_outputs(2049)) xor (layer0_outputs(2270)));
    outputs(1527) <= not(layer0_outputs(2542));
    outputs(1528) <= not((layer0_outputs(257)) xor (layer0_outputs(2178)));
    outputs(1529) <= (layer0_outputs(324)) and not (layer0_outputs(1924));
    outputs(1530) <= not(layer0_outputs(1947));
    outputs(1531) <= (layer0_outputs(1882)) and (layer0_outputs(771));
    outputs(1532) <= not((layer0_outputs(1531)) or (layer0_outputs(2417)));
    outputs(1533) <= layer0_outputs(1489);
    outputs(1534) <= layer0_outputs(1621);
    outputs(1535) <= (layer0_outputs(549)) or (layer0_outputs(567));
    outputs(1536) <= (layer0_outputs(1065)) and not (layer0_outputs(119));
    outputs(1537) <= layer0_outputs(1505);
    outputs(1538) <= not(layer0_outputs(2426));
    outputs(1539) <= not((layer0_outputs(467)) and (layer0_outputs(212)));
    outputs(1540) <= layer0_outputs(977);
    outputs(1541) <= layer0_outputs(2120);
    outputs(1542) <= layer0_outputs(1391);
    outputs(1543) <= not((layer0_outputs(1298)) or (layer0_outputs(244)));
    outputs(1544) <= not((layer0_outputs(2009)) or (layer0_outputs(1380)));
    outputs(1545) <= (layer0_outputs(790)) and not (layer0_outputs(1365));
    outputs(1546) <= (layer0_outputs(602)) xor (layer0_outputs(1489));
    outputs(1547) <= not((layer0_outputs(2516)) xor (layer0_outputs(1901)));
    outputs(1548) <= (layer0_outputs(767)) and (layer0_outputs(1594));
    outputs(1549) <= not((layer0_outputs(1676)) and (layer0_outputs(207)));
    outputs(1550) <= layer0_outputs(2301);
    outputs(1551) <= (layer0_outputs(1962)) and (layer0_outputs(37));
    outputs(1552) <= (layer0_outputs(1503)) and (layer0_outputs(297));
    outputs(1553) <= not((layer0_outputs(1453)) and (layer0_outputs(783)));
    outputs(1554) <= not((layer0_outputs(1763)) xor (layer0_outputs(2108)));
    outputs(1555) <= (layer0_outputs(591)) and not (layer0_outputs(380));
    outputs(1556) <= (layer0_outputs(498)) and not (layer0_outputs(1504));
    outputs(1557) <= (layer0_outputs(2446)) xor (layer0_outputs(181));
    outputs(1558) <= (layer0_outputs(354)) and not (layer0_outputs(266));
    outputs(1559) <= layer0_outputs(498);
    outputs(1560) <= not(layer0_outputs(2009));
    outputs(1561) <= layer0_outputs(2478);
    outputs(1562) <= layer0_outputs(1411);
    outputs(1563) <= (layer0_outputs(840)) and not (layer0_outputs(782));
    outputs(1564) <= not(layer0_outputs(781));
    outputs(1565) <= (layer0_outputs(2376)) and not (layer0_outputs(691));
    outputs(1566) <= not((layer0_outputs(1995)) or (layer0_outputs(621)));
    outputs(1567) <= layer0_outputs(164);
    outputs(1568) <= layer0_outputs(2188);
    outputs(1569) <= (layer0_outputs(52)) and not (layer0_outputs(1031));
    outputs(1570) <= (layer0_outputs(469)) and not (layer0_outputs(577));
    outputs(1571) <= not(layer0_outputs(2201));
    outputs(1572) <= not(layer0_outputs(475));
    outputs(1573) <= (layer0_outputs(2381)) or (layer0_outputs(2012));
    outputs(1574) <= not(layer0_outputs(919));
    outputs(1575) <= (layer0_outputs(1387)) and (layer0_outputs(1745));
    outputs(1576) <= layer0_outputs(2068);
    outputs(1577) <= not(layer0_outputs(2266));
    outputs(1578) <= not(layer0_outputs(1761));
    outputs(1579) <= not(layer0_outputs(2520));
    outputs(1580) <= layer0_outputs(1356);
    outputs(1581) <= not((layer0_outputs(1051)) or (layer0_outputs(422)));
    outputs(1582) <= (layer0_outputs(1132)) and not (layer0_outputs(1218));
    outputs(1583) <= (layer0_outputs(1301)) and (layer0_outputs(1283));
    outputs(1584) <= (layer0_outputs(167)) xor (layer0_outputs(1056));
    outputs(1585) <= not(layer0_outputs(526));
    outputs(1586) <= (layer0_outputs(441)) and not (layer0_outputs(2452));
    outputs(1587) <= not((layer0_outputs(236)) and (layer0_outputs(2226)));
    outputs(1588) <= (layer0_outputs(442)) xor (layer0_outputs(79));
    outputs(1589) <= (layer0_outputs(528)) and not (layer0_outputs(1823));
    outputs(1590) <= (layer0_outputs(418)) and (layer0_outputs(1097));
    outputs(1591) <= (layer0_outputs(2205)) and not (layer0_outputs(1375));
    outputs(1592) <= (layer0_outputs(892)) and (layer0_outputs(1604));
    outputs(1593) <= (layer0_outputs(2059)) and not (layer0_outputs(100));
    outputs(1594) <= layer0_outputs(2148);
    outputs(1595) <= not(layer0_outputs(1700));
    outputs(1596) <= not(layer0_outputs(234));
    outputs(1597) <= (layer0_outputs(1311)) and (layer0_outputs(1202));
    outputs(1598) <= not((layer0_outputs(2157)) or (layer0_outputs(120)));
    outputs(1599) <= layer0_outputs(2005);
    outputs(1600) <= not(layer0_outputs(2110));
    outputs(1601) <= (layer0_outputs(1733)) and not (layer0_outputs(651));
    outputs(1602) <= not(layer0_outputs(886));
    outputs(1603) <= not(layer0_outputs(2349));
    outputs(1604) <= layer0_outputs(190);
    outputs(1605) <= (layer0_outputs(1824)) and not (layer0_outputs(425));
    outputs(1606) <= layer0_outputs(1923);
    outputs(1607) <= not(layer0_outputs(523));
    outputs(1608) <= layer0_outputs(147);
    outputs(1609) <= (layer0_outputs(842)) or (layer0_outputs(2335));
    outputs(1610) <= not(layer0_outputs(2054));
    outputs(1611) <= not(layer0_outputs(2284)) or (layer0_outputs(1421));
    outputs(1612) <= not((layer0_outputs(1374)) or (layer0_outputs(1823)));
    outputs(1613) <= (layer0_outputs(129)) or (layer0_outputs(920));
    outputs(1614) <= not(layer0_outputs(999));
    outputs(1615) <= (layer0_outputs(1734)) and not (layer0_outputs(1900));
    outputs(1616) <= not(layer0_outputs(20));
    outputs(1617) <= (layer0_outputs(766)) xor (layer0_outputs(390));
    outputs(1618) <= not((layer0_outputs(259)) xor (layer0_outputs(714)));
    outputs(1619) <= (layer0_outputs(619)) and not (layer0_outputs(2133));
    outputs(1620) <= (layer0_outputs(199)) and (layer0_outputs(575));
    outputs(1621) <= (layer0_outputs(1713)) and (layer0_outputs(1620));
    outputs(1622) <= not(layer0_outputs(1593)) or (layer0_outputs(2311));
    outputs(1623) <= not(layer0_outputs(49));
    outputs(1624) <= layer0_outputs(2018);
    outputs(1625) <= not(layer0_outputs(2140));
    outputs(1626) <= not((layer0_outputs(2479)) or (layer0_outputs(1440)));
    outputs(1627) <= (layer0_outputs(170)) and not (layer0_outputs(633));
    outputs(1628) <= layer0_outputs(1923);
    outputs(1629) <= (layer0_outputs(724)) and (layer0_outputs(1395));
    outputs(1630) <= (layer0_outputs(1037)) and (layer0_outputs(497));
    outputs(1631) <= not(layer0_outputs(374)) or (layer0_outputs(2445));
    outputs(1632) <= layer0_outputs(1113);
    outputs(1633) <= (layer0_outputs(52)) and not (layer0_outputs(2215));
    outputs(1634) <= layer0_outputs(903);
    outputs(1635) <= layer0_outputs(1819);
    outputs(1636) <= not(layer0_outputs(2234));
    outputs(1637) <= layer0_outputs(1611);
    outputs(1638) <= (layer0_outputs(1391)) and not (layer0_outputs(156));
    outputs(1639) <= not(layer0_outputs(1856));
    outputs(1640) <= not(layer0_outputs(1609));
    outputs(1641) <= layer0_outputs(405);
    outputs(1642) <= not(layer0_outputs(785)) or (layer0_outputs(1860));
    outputs(1643) <= not(layer0_outputs(2092));
    outputs(1644) <= not(layer0_outputs(1430));
    outputs(1645) <= not(layer0_outputs(2283));
    outputs(1646) <= (layer0_outputs(1628)) and (layer0_outputs(2505));
    outputs(1647) <= layer0_outputs(479);
    outputs(1648) <= not(layer0_outputs(302));
    outputs(1649) <= (layer0_outputs(1011)) and (layer0_outputs(958));
    outputs(1650) <= not(layer0_outputs(1828));
    outputs(1651) <= not(layer0_outputs(829));
    outputs(1652) <= (layer0_outputs(1105)) and not (layer0_outputs(568));
    outputs(1653) <= (layer0_outputs(183)) and not (layer0_outputs(976));
    outputs(1654) <= (layer0_outputs(1097)) and not (layer0_outputs(940));
    outputs(1655) <= not(layer0_outputs(1165));
    outputs(1656) <= (layer0_outputs(1822)) and (layer0_outputs(2302));
    outputs(1657) <= not((layer0_outputs(2133)) or (layer0_outputs(538)));
    outputs(1658) <= (layer0_outputs(1484)) xor (layer0_outputs(535));
    outputs(1659) <= not(layer0_outputs(510));
    outputs(1660) <= not(layer0_outputs(110));
    outputs(1661) <= (layer0_outputs(1987)) and (layer0_outputs(1997));
    outputs(1662) <= layer0_outputs(1437);
    outputs(1663) <= not(layer0_outputs(1783));
    outputs(1664) <= (layer0_outputs(1816)) and not (layer0_outputs(1313));
    outputs(1665) <= (layer0_outputs(53)) and (layer0_outputs(1713));
    outputs(1666) <= (layer0_outputs(1008)) and not (layer0_outputs(1781));
    outputs(1667) <= (layer0_outputs(2354)) and not (layer0_outputs(369));
    outputs(1668) <= (layer0_outputs(107)) and not (layer0_outputs(1674));
    outputs(1669) <= layer0_outputs(1123);
    outputs(1670) <= (layer0_outputs(2093)) and (layer0_outputs(358));
    outputs(1671) <= layer0_outputs(2527);
    outputs(1672) <= not((layer0_outputs(1368)) and (layer0_outputs(2286)));
    outputs(1673) <= not((layer0_outputs(1759)) or (layer0_outputs(2217)));
    outputs(1674) <= not(layer0_outputs(2197));
    outputs(1675) <= (layer0_outputs(1407)) and (layer0_outputs(930));
    outputs(1676) <= layer0_outputs(2421);
    outputs(1677) <= layer0_outputs(2557);
    outputs(1678) <= not((layer0_outputs(1626)) or (layer0_outputs(1544)));
    outputs(1679) <= (layer0_outputs(1091)) and not (layer0_outputs(816));
    outputs(1680) <= (layer0_outputs(2535)) xor (layer0_outputs(2144));
    outputs(1681) <= not((layer0_outputs(1497)) or (layer0_outputs(639)));
    outputs(1682) <= (layer0_outputs(1302)) and (layer0_outputs(1337));
    outputs(1683) <= layer0_outputs(598);
    outputs(1684) <= not(layer0_outputs(1564));
    outputs(1685) <= (layer0_outputs(1506)) and (layer0_outputs(61));
    outputs(1686) <= not(layer0_outputs(1015)) or (layer0_outputs(1342));
    outputs(1687) <= not(layer0_outputs(2076));
    outputs(1688) <= (layer0_outputs(2507)) and not (layer0_outputs(594));
    outputs(1689) <= (layer0_outputs(295)) and (layer0_outputs(2316));
    outputs(1690) <= layer0_outputs(1850);
    outputs(1691) <= (layer0_outputs(1629)) and (layer0_outputs(1044));
    outputs(1692) <= not(layer0_outputs(1536));
    outputs(1693) <= not(layer0_outputs(1653));
    outputs(1694) <= not(layer0_outputs(2392));
    outputs(1695) <= (layer0_outputs(860)) xor (layer0_outputs(2149));
    outputs(1696) <= layer0_outputs(2281);
    outputs(1697) <= (layer0_outputs(424)) and not (layer0_outputs(2180));
    outputs(1698) <= (layer0_outputs(235)) and (layer0_outputs(2274));
    outputs(1699) <= (layer0_outputs(1448)) and (layer0_outputs(1367));
    outputs(1700) <= layer0_outputs(2241);
    outputs(1701) <= not(layer0_outputs(2397)) or (layer0_outputs(470));
    outputs(1702) <= (layer0_outputs(1580)) and not (layer0_outputs(905));
    outputs(1703) <= (layer0_outputs(2458)) and not (layer0_outputs(1881));
    outputs(1704) <= (layer0_outputs(779)) xor (layer0_outputs(712));
    outputs(1705) <= not(layer0_outputs(342));
    outputs(1706) <= (layer0_outputs(1961)) and (layer0_outputs(247));
    outputs(1707) <= not(layer0_outputs(1445));
    outputs(1708) <= not(layer0_outputs(2191));
    outputs(1709) <= layer0_outputs(1273);
    outputs(1710) <= not(layer0_outputs(2511));
    outputs(1711) <= (layer0_outputs(490)) and not (layer0_outputs(230));
    outputs(1712) <= (layer0_outputs(1392)) and not (layer0_outputs(728));
    outputs(1713) <= not((layer0_outputs(495)) and (layer0_outputs(1350)));
    outputs(1714) <= (layer0_outputs(1961)) and not (layer0_outputs(1782));
    outputs(1715) <= not((layer0_outputs(200)) or (layer0_outputs(869)));
    outputs(1716) <= (layer0_outputs(2471)) and (layer0_outputs(271));
    outputs(1717) <= layer0_outputs(2045);
    outputs(1718) <= (layer0_outputs(2013)) and (layer0_outputs(1661));
    outputs(1719) <= not((layer0_outputs(941)) or (layer0_outputs(2167)));
    outputs(1720) <= not(layer0_outputs(1082)) or (layer0_outputs(542));
    outputs(1721) <= not(layer0_outputs(312));
    outputs(1722) <= (layer0_outputs(1636)) and not (layer0_outputs(548));
    outputs(1723) <= not(layer0_outputs(380));
    outputs(1724) <= not((layer0_outputs(1288)) and (layer0_outputs(1663)));
    outputs(1725) <= not(layer0_outputs(1266));
    outputs(1726) <= not((layer0_outputs(1299)) or (layer0_outputs(500)));
    outputs(1727) <= not(layer0_outputs(1333));
    outputs(1728) <= not((layer0_outputs(431)) xor (layer0_outputs(1931)));
    outputs(1729) <= (layer0_outputs(1641)) and not (layer0_outputs(188));
    outputs(1730) <= not(layer0_outputs(1233));
    outputs(1731) <= (layer0_outputs(18)) and (layer0_outputs(1442));
    outputs(1732) <= not((layer0_outputs(485)) or (layer0_outputs(711)));
    outputs(1733) <= (layer0_outputs(215)) and not (layer0_outputs(1066));
    outputs(1734) <= (layer0_outputs(2270)) and (layer0_outputs(37));
    outputs(1735) <= (layer0_outputs(972)) and not (layer0_outputs(388));
    outputs(1736) <= not(layer0_outputs(291));
    outputs(1737) <= not(layer0_outputs(1007));
    outputs(1738) <= not(layer0_outputs(491));
    outputs(1739) <= layer0_outputs(1261);
    outputs(1740) <= (layer0_outputs(878)) and not (layer0_outputs(1706));
    outputs(1741) <= layer0_outputs(309);
    outputs(1742) <= (layer0_outputs(497)) or (layer0_outputs(1334));
    outputs(1743) <= (layer0_outputs(706)) and not (layer0_outputs(1968));
    outputs(1744) <= not((layer0_outputs(1289)) or (layer0_outputs(168)));
    outputs(1745) <= (layer0_outputs(1792)) and not (layer0_outputs(2001));
    outputs(1746) <= (layer0_outputs(1772)) and not (layer0_outputs(650));
    outputs(1747) <= not(layer0_outputs(2152)) or (layer0_outputs(1273));
    outputs(1748) <= (layer0_outputs(838)) xor (layer0_outputs(912));
    outputs(1749) <= (layer0_outputs(404)) and not (layer0_outputs(1905));
    outputs(1750) <= layer0_outputs(2147);
    outputs(1751) <= (layer0_outputs(285)) and not (layer0_outputs(1523));
    outputs(1752) <= not((layer0_outputs(2404)) or (layer0_outputs(2309)));
    outputs(1753) <= layer0_outputs(2156);
    outputs(1754) <= not((layer0_outputs(1814)) or (layer0_outputs(2132)));
    outputs(1755) <= not(layer0_outputs(747)) or (layer0_outputs(2356));
    outputs(1756) <= not((layer0_outputs(1330)) or (layer0_outputs(1266)));
    outputs(1757) <= layer0_outputs(2042);
    outputs(1758) <= (layer0_outputs(1510)) or (layer0_outputs(928));
    outputs(1759) <= not(layer0_outputs(1479)) or (layer0_outputs(240));
    outputs(1760) <= not(layer0_outputs(1002)) or (layer0_outputs(1908));
    outputs(1761) <= (layer0_outputs(1036)) and (layer0_outputs(1342));
    outputs(1762) <= not(layer0_outputs(351));
    outputs(1763) <= layer0_outputs(2327);
    outputs(1764) <= (layer0_outputs(333)) and (layer0_outputs(2088));
    outputs(1765) <= not(layer0_outputs(2070));
    outputs(1766) <= not((layer0_outputs(352)) xor (layer0_outputs(1033)));
    outputs(1767) <= layer0_outputs(760);
    outputs(1768) <= (layer0_outputs(1858)) and (layer0_outputs(1719));
    outputs(1769) <= not(layer0_outputs(2321)) or (layer0_outputs(1603));
    outputs(1770) <= (layer0_outputs(398)) and not (layer0_outputs(1896));
    outputs(1771) <= layer0_outputs(1808);
    outputs(1772) <= layer0_outputs(1434);
    outputs(1773) <= layer0_outputs(2231);
    outputs(1774) <= (layer0_outputs(878)) and not (layer0_outputs(1794));
    outputs(1775) <= not(layer0_outputs(316));
    outputs(1776) <= not(layer0_outputs(2444));
    outputs(1777) <= not(layer0_outputs(1501)) or (layer0_outputs(176));
    outputs(1778) <= (layer0_outputs(190)) and (layer0_outputs(1584));
    outputs(1779) <= layer0_outputs(1902);
    outputs(1780) <= not((layer0_outputs(1771)) xor (layer0_outputs(1145)));
    outputs(1781) <= not(layer0_outputs(926)) or (layer0_outputs(1249));
    outputs(1782) <= layer0_outputs(565);
    outputs(1783) <= not(layer0_outputs(1223)) or (layer0_outputs(137));
    outputs(1784) <= (layer0_outputs(2158)) xor (layer0_outputs(638));
    outputs(1785) <= not(layer0_outputs(1846));
    outputs(1786) <= not(layer0_outputs(1869));
    outputs(1787) <= not((layer0_outputs(1252)) or (layer0_outputs(485)));
    outputs(1788) <= (layer0_outputs(2371)) and not (layer0_outputs(1472));
    outputs(1789) <= layer0_outputs(328);
    outputs(1790) <= layer0_outputs(1642);
    outputs(1791) <= (layer0_outputs(1211)) and not (layer0_outputs(335));
    outputs(1792) <= layer0_outputs(1785);
    outputs(1793) <= (layer0_outputs(1007)) and (layer0_outputs(142));
    outputs(1794) <= (layer0_outputs(820)) and (layer0_outputs(832));
    outputs(1795) <= (layer0_outputs(1728)) and not (layer0_outputs(2057));
    outputs(1796) <= not((layer0_outputs(260)) or (layer0_outputs(628)));
    outputs(1797) <= (layer0_outputs(1256)) and not (layer0_outputs(741));
    outputs(1798) <= (layer0_outputs(1776)) and (layer0_outputs(1136));
    outputs(1799) <= layer0_outputs(1761);
    outputs(1800) <= layer0_outputs(1598);
    outputs(1801) <= (layer0_outputs(1417)) or (layer0_outputs(1576));
    outputs(1802) <= (layer0_outputs(1155)) and not (layer0_outputs(25));
    outputs(1803) <= layer0_outputs(517);
    outputs(1804) <= not((layer0_outputs(1591)) and (layer0_outputs(2508)));
    outputs(1805) <= not((layer0_outputs(532)) and (layer0_outputs(2550)));
    outputs(1806) <= not(layer0_outputs(660));
    outputs(1807) <= (layer0_outputs(1135)) and (layer0_outputs(794));
    outputs(1808) <= (layer0_outputs(1575)) and not (layer0_outputs(1305));
    outputs(1809) <= not((layer0_outputs(213)) or (layer0_outputs(1087)));
    outputs(1810) <= layer0_outputs(1755);
    outputs(1811) <= not(layer0_outputs(304));
    outputs(1812) <= layer0_outputs(496);
    outputs(1813) <= (layer0_outputs(1589)) and not (layer0_outputs(2177));
    outputs(1814) <= layer0_outputs(2223);
    outputs(1815) <= layer0_outputs(421);
    outputs(1816) <= (layer0_outputs(780)) and not (layer0_outputs(2486));
    outputs(1817) <= not(layer0_outputs(2081));
    outputs(1818) <= (layer0_outputs(763)) and (layer0_outputs(157));
    outputs(1819) <= not((layer0_outputs(2460)) or (layer0_outputs(2499)));
    outputs(1820) <= not(layer0_outputs(1858));
    outputs(1821) <= not((layer0_outputs(1090)) or (layer0_outputs(1516)));
    outputs(1822) <= '0';
    outputs(1823) <= not(layer0_outputs(1835));
    outputs(1824) <= (layer0_outputs(1810)) and not (layer0_outputs(1149));
    outputs(1825) <= layer0_outputs(1662);
    outputs(1826) <= (layer0_outputs(278)) and (layer0_outputs(1072));
    outputs(1827) <= layer0_outputs(1481);
    outputs(1828) <= not(layer0_outputs(2220));
    outputs(1829) <= not(layer0_outputs(401));
    outputs(1830) <= (layer0_outputs(2067)) and not (layer0_outputs(931));
    outputs(1831) <= not(layer0_outputs(1048));
    outputs(1832) <= (layer0_outputs(46)) and not (layer0_outputs(191));
    outputs(1833) <= layer0_outputs(2022);
    outputs(1834) <= not(layer0_outputs(296));
    outputs(1835) <= (layer0_outputs(1550)) and (layer0_outputs(2514));
    outputs(1836) <= not(layer0_outputs(1554));
    outputs(1837) <= (layer0_outputs(1169)) and (layer0_outputs(2197));
    outputs(1838) <= not((layer0_outputs(125)) and (layer0_outputs(308)));
    outputs(1839) <= not((layer0_outputs(1010)) or (layer0_outputs(30)));
    outputs(1840) <= not((layer0_outputs(2461)) or (layer0_outputs(2064)));
    outputs(1841) <= (layer0_outputs(1108)) and (layer0_outputs(2394));
    outputs(1842) <= (layer0_outputs(2207)) and (layer0_outputs(1263));
    outputs(1843) <= layer0_outputs(1207);
    outputs(1844) <= not((layer0_outputs(797)) or (layer0_outputs(2396)));
    outputs(1845) <= (layer0_outputs(1362)) and not (layer0_outputs(2012));
    outputs(1846) <= not(layer0_outputs(1398));
    outputs(1847) <= not((layer0_outputs(1017)) or (layer0_outputs(634)));
    outputs(1848) <= layer0_outputs(119);
    outputs(1849) <= not(layer0_outputs(31));
    outputs(1850) <= layer0_outputs(1226);
    outputs(1851) <= not((layer0_outputs(2086)) or (layer0_outputs(36)));
    outputs(1852) <= (layer0_outputs(2472)) and not (layer0_outputs(75));
    outputs(1853) <= layer0_outputs(1298);
    outputs(1854) <= (layer0_outputs(725)) and not (layer0_outputs(2141));
    outputs(1855) <= not((layer0_outputs(2329)) or (layer0_outputs(448)));
    outputs(1856) <= (layer0_outputs(624)) and not (layer0_outputs(626));
    outputs(1857) <= not((layer0_outputs(815)) or (layer0_outputs(2307)));
    outputs(1858) <= not((layer0_outputs(1185)) xor (layer0_outputs(2157)));
    outputs(1859) <= layer0_outputs(2080);
    outputs(1860) <= not(layer0_outputs(154)) or (layer0_outputs(63));
    outputs(1861) <= not(layer0_outputs(29)) or (layer0_outputs(597));
    outputs(1862) <= (layer0_outputs(1736)) and not (layer0_outputs(1215));
    outputs(1863) <= not((layer0_outputs(385)) and (layer0_outputs(2425)));
    outputs(1864) <= '0';
    outputs(1865) <= not((layer0_outputs(14)) or (layer0_outputs(2237)));
    outputs(1866) <= (layer0_outputs(1784)) and not (layer0_outputs(109));
    outputs(1867) <= (layer0_outputs(1646)) or (layer0_outputs(2280));
    outputs(1868) <= not((layer0_outputs(2160)) or (layer0_outputs(709)));
    outputs(1869) <= layer0_outputs(702);
    outputs(1870) <= layer0_outputs(338);
    outputs(1871) <= not(layer0_outputs(1127));
    outputs(1872) <= not(layer0_outputs(744));
    outputs(1873) <= not(layer0_outputs(583));
    outputs(1874) <= (layer0_outputs(494)) and not (layer0_outputs(1724));
    outputs(1875) <= not(layer0_outputs(246));
    outputs(1876) <= (layer0_outputs(382)) and not (layer0_outputs(435));
    outputs(1877) <= not((layer0_outputs(2311)) or (layer0_outputs(561)));
    outputs(1878) <= not(layer0_outputs(2269));
    outputs(1879) <= (layer0_outputs(487)) and (layer0_outputs(1303));
    outputs(1880) <= (layer0_outputs(986)) and not (layer0_outputs(955));
    outputs(1881) <= not(layer0_outputs(856)) or (layer0_outputs(1390));
    outputs(1882) <= not((layer0_outputs(298)) or (layer0_outputs(1940)));
    outputs(1883) <= (layer0_outputs(1967)) and not (layer0_outputs(1904));
    outputs(1884) <= (layer0_outputs(459)) and not (layer0_outputs(175));
    outputs(1885) <= not(layer0_outputs(41));
    outputs(1886) <= not((layer0_outputs(1183)) and (layer0_outputs(902)));
    outputs(1887) <= not(layer0_outputs(433));
    outputs(1888) <= (layer0_outputs(1751)) xor (layer0_outputs(9));
    outputs(1889) <= not(layer0_outputs(1423));
    outputs(1890) <= not(layer0_outputs(254)) or (layer0_outputs(2190));
    outputs(1891) <= not((layer0_outputs(1055)) or (layer0_outputs(950)));
    outputs(1892) <= layer0_outputs(1361);
    outputs(1893) <= (layer0_outputs(1541)) and not (layer0_outputs(1292));
    outputs(1894) <= not(layer0_outputs(161)) or (layer0_outputs(2406));
    outputs(1895) <= (layer0_outputs(2037)) and (layer0_outputs(2137));
    outputs(1896) <= (layer0_outputs(1769)) and (layer0_outputs(601));
    outputs(1897) <= layer0_outputs(556);
    outputs(1898) <= not((layer0_outputs(1645)) or (layer0_outputs(770)));
    outputs(1899) <= (layer0_outputs(1243)) and not (layer0_outputs(1018));
    outputs(1900) <= not(layer0_outputs(2506));
    outputs(1901) <= layer0_outputs(1960);
    outputs(1902) <= not(layer0_outputs(1464));
    outputs(1903) <= not((layer0_outputs(1886)) or (layer0_outputs(1001)));
    outputs(1904) <= not(layer0_outputs(571)) or (layer0_outputs(425));
    outputs(1905) <= (layer0_outputs(2029)) and not (layer0_outputs(464));
    outputs(1906) <= not(layer0_outputs(1686));
    outputs(1907) <= (layer0_outputs(1070)) and not (layer0_outputs(1399));
    outputs(1908) <= not((layer0_outputs(189)) xor (layer0_outputs(2239)));
    outputs(1909) <= (layer0_outputs(2053)) and not (layer0_outputs(542));
    outputs(1910) <= not((layer0_outputs(1341)) or (layer0_outputs(1379)));
    outputs(1911) <= layer0_outputs(1287);
    outputs(1912) <= not((layer0_outputs(2216)) xor (layer0_outputs(1271)));
    outputs(1913) <= layer0_outputs(631);
    outputs(1914) <= (layer0_outputs(547)) and not (layer0_outputs(784));
    outputs(1915) <= (layer0_outputs(968)) and not (layer0_outputs(1860));
    outputs(1916) <= (layer0_outputs(720)) and not (layer0_outputs(1891));
    outputs(1917) <= (layer0_outputs(919)) and not (layer0_outputs(105));
    outputs(1918) <= (layer0_outputs(2470)) and (layer0_outputs(1229));
    outputs(1919) <= not((layer0_outputs(1189)) or (layer0_outputs(2295)));
    outputs(1920) <= not((layer0_outputs(1749)) or (layer0_outputs(1817)));
    outputs(1921) <= not(layer0_outputs(1607));
    outputs(1922) <= layer0_outputs(1405);
    outputs(1923) <= (layer0_outputs(2170)) and not (layer0_outputs(2350));
    outputs(1924) <= (layer0_outputs(1683)) and not (layer0_outputs(923));
    outputs(1925) <= (layer0_outputs(1163)) and not (layer0_outputs(107));
    outputs(1926) <= not(layer0_outputs(1120));
    outputs(1927) <= not(layer0_outputs(1921)) or (layer0_outputs(1730));
    outputs(1928) <= (layer0_outputs(1871)) and not (layer0_outputs(1563));
    outputs(1929) <= not((layer0_outputs(1614)) xor (layer0_outputs(19)));
    outputs(1930) <= not(layer0_outputs(381)) or (layer0_outputs(2303));
    outputs(1931) <= layer0_outputs(1832);
    outputs(1932) <= layer0_outputs(1297);
    outputs(1933) <= (layer0_outputs(547)) and (layer0_outputs(1184));
    outputs(1934) <= not(layer0_outputs(1016));
    outputs(1935) <= (layer0_outputs(2277)) and (layer0_outputs(2389));
    outputs(1936) <= not((layer0_outputs(216)) or (layer0_outputs(2385)));
    outputs(1937) <= not(layer0_outputs(1929));
    outputs(1938) <= (layer0_outputs(674)) and (layer0_outputs(1634));
    outputs(1939) <= layer0_outputs(830);
    outputs(1940) <= not((layer0_outputs(2212)) or (layer0_outputs(1743)));
    outputs(1941) <= (layer0_outputs(1877)) and (layer0_outputs(1297));
    outputs(1942) <= (layer0_outputs(2524)) and (layer0_outputs(1820));
    outputs(1943) <= not((layer0_outputs(1529)) or (layer0_outputs(143)));
    outputs(1944) <= (layer0_outputs(2285)) xor (layer0_outputs(2363));
    outputs(1945) <= not(layer0_outputs(1109)) or (layer0_outputs(1504));
    outputs(1946) <= (layer0_outputs(698)) and not (layer0_outputs(444));
    outputs(1947) <= not((layer0_outputs(1956)) and (layer0_outputs(2475)));
    outputs(1948) <= (layer0_outputs(2364)) and (layer0_outputs(2495));
    outputs(1949) <= not(layer0_outputs(930));
    outputs(1950) <= (layer0_outputs(2123)) and not (layer0_outputs(201));
    outputs(1951) <= layer0_outputs(1637);
    outputs(1952) <= not((layer0_outputs(334)) and (layer0_outputs(1790)));
    outputs(1953) <= (layer0_outputs(899)) and not (layer0_outputs(1123));
    outputs(1954) <= not((layer0_outputs(693)) or (layer0_outputs(2384)));
    outputs(1955) <= not(layer0_outputs(1120));
    outputs(1956) <= (layer0_outputs(2348)) and not (layer0_outputs(2346));
    outputs(1957) <= not((layer0_outputs(2065)) or (layer0_outputs(57)));
    outputs(1958) <= (layer0_outputs(676)) and not (layer0_outputs(1975));
    outputs(1959) <= layer0_outputs(1067);
    outputs(1960) <= (layer0_outputs(1116)) and not (layer0_outputs(328));
    outputs(1961) <= not((layer0_outputs(98)) or (layer0_outputs(2504)));
    outputs(1962) <= not((layer0_outputs(2494)) or (layer0_outputs(1772)));
    outputs(1963) <= (layer0_outputs(2139)) and not (layer0_outputs(688));
    outputs(1964) <= layer0_outputs(1913);
    outputs(1965) <= (layer0_outputs(2135)) and (layer0_outputs(1258));
    outputs(1966) <= (layer0_outputs(722)) and not (layer0_outputs(149));
    outputs(1967) <= (layer0_outputs(1426)) and not (layer0_outputs(973));
    outputs(1968) <= not(layer0_outputs(833));
    outputs(1969) <= layer0_outputs(1799);
    outputs(1970) <= (layer0_outputs(1067)) and (layer0_outputs(370));
    outputs(1971) <= layer0_outputs(2043);
    outputs(1972) <= not(layer0_outputs(193)) or (layer0_outputs(229));
    outputs(1973) <= not((layer0_outputs(1406)) xor (layer0_outputs(2078)));
    outputs(1974) <= not((layer0_outputs(1449)) or (layer0_outputs(603)));
    outputs(1975) <= (layer0_outputs(2026)) and not (layer0_outputs(1513));
    outputs(1976) <= not(layer0_outputs(1545));
    outputs(1977) <= (layer0_outputs(2320)) and (layer0_outputs(1748));
    outputs(1978) <= (layer0_outputs(1996)) and not (layer0_outputs(1439));
    outputs(1979) <= not((layer0_outputs(692)) xor (layer0_outputs(1927)));
    outputs(1980) <= (layer0_outputs(62)) and (layer0_outputs(1147));
    outputs(1981) <= (layer0_outputs(2183)) and (layer0_outputs(2427));
    outputs(1982) <= not(layer0_outputs(2163)) or (layer0_outputs(2048));
    outputs(1983) <= not((layer0_outputs(1547)) or (layer0_outputs(1205)));
    outputs(1984) <= not(layer0_outputs(60));
    outputs(1985) <= (layer0_outputs(1020)) and not (layer0_outputs(2508));
    outputs(1986) <= not((layer0_outputs(1552)) or (layer0_outputs(307)));
    outputs(1987) <= (layer0_outputs(1364)) and not (layer0_outputs(2397));
    outputs(1988) <= (layer0_outputs(145)) and not (layer0_outputs(456));
    outputs(1989) <= (layer0_outputs(1581)) and not (layer0_outputs(841));
    outputs(1990) <= (layer0_outputs(652)) and not (layer0_outputs(1168));
    outputs(1991) <= not((layer0_outputs(2414)) or (layer0_outputs(1884)));
    outputs(1992) <= not((layer0_outputs(843)) or (layer0_outputs(1545)));
    outputs(1993) <= (layer0_outputs(1900)) and not (layer0_outputs(441));
    outputs(1994) <= not((layer0_outputs(1325)) or (layer0_outputs(2164)));
    outputs(1995) <= not(layer0_outputs(4)) or (layer0_outputs(1110));
    outputs(1996) <= layer0_outputs(901);
    outputs(1997) <= (layer0_outputs(245)) and (layer0_outputs(1014));
    outputs(1998) <= (layer0_outputs(2469)) and not (layer0_outputs(1249));
    outputs(1999) <= not(layer0_outputs(354));
    outputs(2000) <= not(layer0_outputs(1955));
    outputs(2001) <= not(layer0_outputs(642));
    outputs(2002) <= (layer0_outputs(1169)) and (layer0_outputs(2536));
    outputs(2003) <= not(layer0_outputs(399)) or (layer0_outputs(1935));
    outputs(2004) <= (layer0_outputs(858)) or (layer0_outputs(1914));
    outputs(2005) <= not(layer0_outputs(1733));
    outputs(2006) <= not((layer0_outputs(744)) or (layer0_outputs(540)));
    outputs(2007) <= not(layer0_outputs(1381));
    outputs(2008) <= layer0_outputs(557);
    outputs(2009) <= not(layer0_outputs(396));
    outputs(2010) <= not((layer0_outputs(1173)) or (layer0_outputs(1657)));
    outputs(2011) <= not((layer0_outputs(2506)) or (layer0_outputs(770)));
    outputs(2012) <= (layer0_outputs(1022)) and (layer0_outputs(1687));
    outputs(2013) <= layer0_outputs(2544);
    outputs(2014) <= not((layer0_outputs(856)) or (layer0_outputs(1904)));
    outputs(2015) <= not(layer0_outputs(2272));
    outputs(2016) <= layer0_outputs(681);
    outputs(2017) <= not((layer0_outputs(1476)) or (layer0_outputs(637)));
    outputs(2018) <= layer0_outputs(1893);
    outputs(2019) <= not((layer0_outputs(778)) and (layer0_outputs(2172)));
    outputs(2020) <= layer0_outputs(743);
    outputs(2021) <= layer0_outputs(74);
    outputs(2022) <= not((layer0_outputs(567)) or (layer0_outputs(331)));
    outputs(2023) <= (layer0_outputs(1082)) and not (layer0_outputs(637));
    outputs(2024) <= not(layer0_outputs(1296));
    outputs(2025) <= not((layer0_outputs(67)) and (layer0_outputs(1055)));
    outputs(2026) <= layer0_outputs(1254);
    outputs(2027) <= not((layer0_outputs(270)) or (layer0_outputs(2104)));
    outputs(2028) <= (layer0_outputs(1172)) and not (layer0_outputs(303));
    outputs(2029) <= not(layer0_outputs(350));
    outputs(2030) <= layer0_outputs(1452);
    outputs(2031) <= (layer0_outputs(70)) xor (layer0_outputs(877));
    outputs(2032) <= not(layer0_outputs(2492));
    outputs(2033) <= (layer0_outputs(938)) or (layer0_outputs(1949));
    outputs(2034) <= (layer0_outputs(962)) and not (layer0_outputs(1398));
    outputs(2035) <= not((layer0_outputs(1883)) or (layer0_outputs(1648)));
    outputs(2036) <= not(layer0_outputs(2016));
    outputs(2037) <= (layer0_outputs(1347)) and (layer0_outputs(209));
    outputs(2038) <= (layer0_outputs(2170)) and not (layer0_outputs(186));
    outputs(2039) <= not(layer0_outputs(139));
    outputs(2040) <= (layer0_outputs(1134)) or (layer0_outputs(1660));
    outputs(2041) <= not(layer0_outputs(632));
    outputs(2042) <= not(layer0_outputs(1059));
    outputs(2043) <= layer0_outputs(2318);
    outputs(2044) <= (layer0_outputs(832)) and (layer0_outputs(793));
    outputs(2045) <= not((layer0_outputs(287)) or (layer0_outputs(1004)));
    outputs(2046) <= not((layer0_outputs(1722)) or (layer0_outputs(2291)));
    outputs(2047) <= not((layer0_outputs(634)) xor (layer0_outputs(911)));
    outputs(2048) <= (layer0_outputs(1327)) and not (layer0_outputs(476));
    outputs(2049) <= layer0_outputs(904);
    outputs(2050) <= layer0_outputs(633);
    outputs(2051) <= (layer0_outputs(774)) and (layer0_outputs(1821));
    outputs(2052) <= not(layer0_outputs(1492));
    outputs(2053) <= (layer0_outputs(1332)) and not (layer0_outputs(811));
    outputs(2054) <= layer0_outputs(1777);
    outputs(2055) <= not(layer0_outputs(581)) or (layer0_outputs(1553));
    outputs(2056) <= (layer0_outputs(1970)) xor (layer0_outputs(947));
    outputs(2057) <= layer0_outputs(2452);
    outputs(2058) <= not(layer0_outputs(2189)) or (layer0_outputs(1494));
    outputs(2059) <= not(layer0_outputs(1187)) or (layer0_outputs(1419));
    outputs(2060) <= not(layer0_outputs(1286));
    outputs(2061) <= not((layer0_outputs(578)) or (layer0_outputs(473)));
    outputs(2062) <= layer0_outputs(2498);
    outputs(2063) <= not(layer0_outputs(1558));
    outputs(2064) <= layer0_outputs(1358);
    outputs(2065) <= not(layer0_outputs(2525));
    outputs(2066) <= layer0_outputs(2532);
    outputs(2067) <= not(layer0_outputs(2318)) or (layer0_outputs(1644));
    outputs(2068) <= layer0_outputs(2326);
    outputs(2069) <= layer0_outputs(323);
    outputs(2070) <= layer0_outputs(2456);
    outputs(2071) <= layer0_outputs(745);
    outputs(2072) <= (layer0_outputs(1647)) xor (layer0_outputs(1796));
    outputs(2073) <= not((layer0_outputs(1821)) xor (layer0_outputs(1911)));
    outputs(2074) <= layer0_outputs(2538);
    outputs(2075) <= not(layer0_outputs(1684));
    outputs(2076) <= not((layer0_outputs(612)) and (layer0_outputs(290)));
    outputs(2077) <= not(layer0_outputs(2523));
    outputs(2078) <= (layer0_outputs(1625)) xor (layer0_outputs(1862));
    outputs(2079) <= not(layer0_outputs(108));
    outputs(2080) <= layer0_outputs(1936);
    outputs(2081) <= layer0_outputs(1239);
    outputs(2082) <= layer0_outputs(751);
    outputs(2083) <= (layer0_outputs(1132)) xor (layer0_outputs(2350));
    outputs(2084) <= not(layer0_outputs(2254));
    outputs(2085) <= not((layer0_outputs(1121)) or (layer0_outputs(546)));
    outputs(2086) <= not((layer0_outputs(824)) xor (layer0_outputs(1452)));
    outputs(2087) <= not(layer0_outputs(127));
    outputs(2088) <= not((layer0_outputs(1711)) xor (layer0_outputs(917)));
    outputs(2089) <= not(layer0_outputs(848));
    outputs(2090) <= not((layer0_outputs(222)) xor (layer0_outputs(675)));
    outputs(2091) <= layer0_outputs(301);
    outputs(2092) <= not(layer0_outputs(1488));
    outputs(2093) <= (layer0_outputs(1412)) or (layer0_outputs(409));
    outputs(2094) <= (layer0_outputs(1796)) and not (layer0_outputs(2329));
    outputs(2095) <= not(layer0_outputs(1024));
    outputs(2096) <= not((layer0_outputs(749)) and (layer0_outputs(2079)));
    outputs(2097) <= (layer0_outputs(1777)) and not (layer0_outputs(1167));
    outputs(2098) <= (layer0_outputs(1540)) xor (layer0_outputs(268));
    outputs(2099) <= layer0_outputs(750);
    outputs(2100) <= not((layer0_outputs(524)) or (layer0_outputs(1535)));
    outputs(2101) <= not(layer0_outputs(1141));
    outputs(2102) <= not(layer0_outputs(114));
    outputs(2103) <= not(layer0_outputs(1465));
    outputs(2104) <= layer0_outputs(2543);
    outputs(2105) <= not(layer0_outputs(1420)) or (layer0_outputs(314));
    outputs(2106) <= (layer0_outputs(1815)) and not (layer0_outputs(2038));
    outputs(2107) <= not((layer0_outputs(2116)) or (layer0_outputs(625)));
    outputs(2108) <= not(layer0_outputs(758));
    outputs(2109) <= (layer0_outputs(152)) or (layer0_outputs(645));
    outputs(2110) <= not(layer0_outputs(1315)) or (layer0_outputs(909));
    outputs(2111) <= (layer0_outputs(1629)) and not (layer0_outputs(183));
    outputs(2112) <= (layer0_outputs(817)) and (layer0_outputs(1966));
    outputs(2113) <= layer0_outputs(517);
    outputs(2114) <= layer0_outputs(2010);
    outputs(2115) <= not(layer0_outputs(593));
    outputs(2116) <= not(layer0_outputs(1941));
    outputs(2117) <= (layer0_outputs(758)) xor (layer0_outputs(1109));
    outputs(2118) <= (layer0_outputs(1807)) xor (layer0_outputs(1095));
    outputs(2119) <= not(layer0_outputs(1854)) or (layer0_outputs(2310));
    outputs(2120) <= not(layer0_outputs(501)) or (layer0_outputs(686));
    outputs(2121) <= (layer0_outputs(1548)) xor (layer0_outputs(682));
    outputs(2122) <= not(layer0_outputs(1748));
    outputs(2123) <= layer0_outputs(1826);
    outputs(2124) <= (layer0_outputs(1847)) and not (layer0_outputs(541));
    outputs(2125) <= not((layer0_outputs(815)) or (layer0_outputs(2554)));
    outputs(2126) <= (layer0_outputs(948)) or (layer0_outputs(1706));
    outputs(2127) <= layer0_outputs(1396);
    outputs(2128) <= layer0_outputs(1300);
    outputs(2129) <= not(layer0_outputs(38));
    outputs(2130) <= layer0_outputs(2477);
    outputs(2131) <= not(layer0_outputs(205));
    outputs(2132) <= not(layer0_outputs(1058));
    outputs(2133) <= not(layer0_outputs(132)) or (layer0_outputs(2458));
    outputs(2134) <= layer0_outputs(2517);
    outputs(2135) <= layer0_outputs(302);
    outputs(2136) <= not(layer0_outputs(493));
    outputs(2137) <= (layer0_outputs(222)) xor (layer0_outputs(1646));
    outputs(2138) <= layer0_outputs(230);
    outputs(2139) <= layer0_outputs(323);
    outputs(2140) <= (layer0_outputs(1306)) and not (layer0_outputs(298));
    outputs(2141) <= not((layer0_outputs(2445)) and (layer0_outputs(1133)));
    outputs(2142) <= layer0_outputs(704);
    outputs(2143) <= not(layer0_outputs(491)) or (layer0_outputs(2211));
    outputs(2144) <= (layer0_outputs(2097)) xor (layer0_outputs(670));
    outputs(2145) <= not((layer0_outputs(1079)) or (layer0_outputs(260)));
    outputs(2146) <= not(layer0_outputs(1517));
    outputs(2147) <= not(layer0_outputs(1705));
    outputs(2148) <= layer0_outputs(701);
    outputs(2149) <= (layer0_outputs(2555)) xor (layer0_outputs(1073));
    outputs(2150) <= (layer0_outputs(2304)) and (layer0_outputs(1404));
    outputs(2151) <= not(layer0_outputs(1892));
    outputs(2152) <= layer0_outputs(1650);
    outputs(2153) <= not((layer0_outputs(786)) and (layer0_outputs(952)));
    outputs(2154) <= (layer0_outputs(1374)) or (layer0_outputs(539));
    outputs(2155) <= not(layer0_outputs(1994));
    outputs(2156) <= not(layer0_outputs(2147));
    outputs(2157) <= (layer0_outputs(263)) and (layer0_outputs(1491));
    outputs(2158) <= (layer0_outputs(1703)) and (layer0_outputs(1043));
    outputs(2159) <= not(layer0_outputs(2390));
    outputs(2160) <= not(layer0_outputs(1813));
    outputs(2161) <= layer0_outputs(1685);
    outputs(2162) <= (layer0_outputs(2259)) and (layer0_outputs(2552));
    outputs(2163) <= layer0_outputs(242);
    outputs(2164) <= not((layer0_outputs(2097)) xor (layer0_outputs(2530)));
    outputs(2165) <= (layer0_outputs(2507)) and not (layer0_outputs(1888));
    outputs(2166) <= (layer0_outputs(460)) and (layer0_outputs(708));
    outputs(2167) <= not(layer0_outputs(2052)) or (layer0_outputs(961));
    outputs(2168) <= (layer0_outputs(207)) and not (layer0_outputs(836));
    outputs(2169) <= not((layer0_outputs(2200)) or (layer0_outputs(796)));
    outputs(2170) <= layer0_outputs(1081);
    outputs(2171) <= not(layer0_outputs(455));
    outputs(2172) <= layer0_outputs(1257);
    outputs(2173) <= layer0_outputs(1738);
    outputs(2174) <= (layer0_outputs(1701)) and not (layer0_outputs(1776));
    outputs(2175) <= not(layer0_outputs(1128));
    outputs(2176) <= not((layer0_outputs(1162)) xor (layer0_outputs(1632)));
    outputs(2177) <= layer0_outputs(775);
    outputs(2178) <= (layer0_outputs(1209)) and not (layer0_outputs(720));
    outputs(2179) <= (layer0_outputs(1939)) xor (layer0_outputs(1323));
    outputs(2180) <= layer0_outputs(124);
    outputs(2181) <= layer0_outputs(755);
    outputs(2182) <= not(layer0_outputs(593));
    outputs(2183) <= (layer0_outputs(1441)) and (layer0_outputs(1195));
    outputs(2184) <= (layer0_outputs(537)) xor (layer0_outputs(2008));
    outputs(2185) <= (layer0_outputs(1361)) or (layer0_outputs(1863));
    outputs(2186) <= not(layer0_outputs(270));
    outputs(2187) <= not(layer0_outputs(1478));
    outputs(2188) <= not((layer0_outputs(528)) xor (layer0_outputs(2526)));
    outputs(2189) <= not(layer0_outputs(1061));
    outputs(2190) <= (layer0_outputs(765)) xor (layer0_outputs(1538));
    outputs(2191) <= layer0_outputs(1989);
    outputs(2192) <= (layer0_outputs(613)) and not (layer0_outputs(141));
    outputs(2193) <= not(layer0_outputs(910));
    outputs(2194) <= not(layer0_outputs(402));
    outputs(2195) <= (layer0_outputs(663)) and not (layer0_outputs(1522));
    outputs(2196) <= layer0_outputs(2245);
    outputs(2197) <= layer0_outputs(2314);
    outputs(2198) <= (layer0_outputs(185)) xor (layer0_outputs(781));
    outputs(2199) <= not(layer0_outputs(1888));
    outputs(2200) <= (layer0_outputs(2467)) or (layer0_outputs(1729));
    outputs(2201) <= not(layer0_outputs(337)) or (layer0_outputs(2416));
    outputs(2202) <= layer0_outputs(2024);
    outputs(2203) <= (layer0_outputs(2017)) or (layer0_outputs(1590));
    outputs(2204) <= (layer0_outputs(1839)) and not (layer0_outputs(2228));
    outputs(2205) <= (layer0_outputs(1083)) xor (layer0_outputs(1855));
    outputs(2206) <= layer0_outputs(1882);
    outputs(2207) <= (layer0_outputs(1588)) and not (layer0_outputs(1806));
    outputs(2208) <= (layer0_outputs(417)) and not (layer0_outputs(1965));
    outputs(2209) <= layer0_outputs(554);
    outputs(2210) <= (layer0_outputs(1184)) and not (layer0_outputs(1251));
    outputs(2211) <= (layer0_outputs(1543)) or (layer0_outputs(2404));
    outputs(2212) <= not(layer0_outputs(707)) or (layer0_outputs(2092));
    outputs(2213) <= (layer0_outputs(1473)) and not (layer0_outputs(658));
    outputs(2214) <= layer0_outputs(410);
    outputs(2215) <= (layer0_outputs(1690)) xor (layer0_outputs(71));
    outputs(2216) <= not(layer0_outputs(2312));
    outputs(2217) <= (layer0_outputs(9)) and (layer0_outputs(2160));
    outputs(2218) <= layer0_outputs(1131);
    outputs(2219) <= layer0_outputs(2217);
    outputs(2220) <= not(layer0_outputs(262));
    outputs(2221) <= not((layer0_outputs(66)) or (layer0_outputs(2128)));
    outputs(2222) <= layer0_outputs(718);
    outputs(2223) <= (layer0_outputs(1354)) and (layer0_outputs(2251));
    outputs(2224) <= not((layer0_outputs(2447)) or (layer0_outputs(1963)));
    outputs(2225) <= layer0_outputs(241);
    outputs(2226) <= layer0_outputs(2263);
    outputs(2227) <= not((layer0_outputs(478)) or (layer0_outputs(1208)));
    outputs(2228) <= (layer0_outputs(2437)) xor (layer0_outputs(2235));
    outputs(2229) <= not(layer0_outputs(2523));
    outputs(2230) <= not((layer0_outputs(806)) xor (layer0_outputs(956)));
    outputs(2231) <= not(layer0_outputs(220));
    outputs(2232) <= (layer0_outputs(2368)) and (layer0_outputs(1952));
    outputs(2233) <= (layer0_outputs(489)) and (layer0_outputs(1269));
    outputs(2234) <= (layer0_outputs(1445)) xor (layer0_outputs(1673));
    outputs(2235) <= (layer0_outputs(1770)) and not (layer0_outputs(1577));
    outputs(2236) <= (layer0_outputs(722)) and (layer0_outputs(187));
    outputs(2237) <= not((layer0_outputs(2419)) and (layer0_outputs(334)));
    outputs(2238) <= (layer0_outputs(1669)) and (layer0_outputs(1742));
    outputs(2239) <= not(layer0_outputs(6));
    outputs(2240) <= layer0_outputs(1424);
    outputs(2241) <= (layer0_outputs(1653)) xor (layer0_outputs(28));
    outputs(2242) <= (layer0_outputs(1786)) or (layer0_outputs(1870));
    outputs(2243) <= layer0_outputs(2262);
    outputs(2244) <= not(layer0_outputs(853)) or (layer0_outputs(978));
    outputs(2245) <= (layer0_outputs(1332)) and not (layer0_outputs(835));
    outputs(2246) <= not(layer0_outputs(35));
    outputs(2247) <= (layer0_outputs(1482)) or (layer0_outputs(1130));
    outputs(2248) <= (layer0_outputs(430)) and (layer0_outputs(985));
    outputs(2249) <= not((layer0_outputs(530)) or (layer0_outputs(176)));
    outputs(2250) <= not(layer0_outputs(1552)) or (layer0_outputs(1076));
    outputs(2251) <= not(layer0_outputs(1853));
    outputs(2252) <= layer0_outputs(2415);
    outputs(2253) <= not(layer0_outputs(1537));
    outputs(2254) <= layer0_outputs(667);
    outputs(2255) <= not((layer0_outputs(473)) or (layer0_outputs(1910)));
    outputs(2256) <= not((layer0_outputs(2231)) and (layer0_outputs(2171)));
    outputs(2257) <= (layer0_outputs(450)) and not (layer0_outputs(699));
    outputs(2258) <= not(layer0_outputs(2330));
    outputs(2259) <= (layer0_outputs(2118)) xor (layer0_outputs(1688));
    outputs(2260) <= (layer0_outputs(2074)) xor (layer0_outputs(1260));
    outputs(2261) <= not((layer0_outputs(2549)) xor (layer0_outputs(2125)));
    outputs(2262) <= (layer0_outputs(139)) and (layer0_outputs(1847));
    outputs(2263) <= (layer0_outputs(1622)) and (layer0_outputs(360));
    outputs(2264) <= layer0_outputs(1265);
    outputs(2265) <= (layer0_outputs(1999)) and (layer0_outputs(1912));
    outputs(2266) <= not(layer0_outputs(1416));
    outputs(2267) <= (layer0_outputs(315)) and not (layer0_outputs(1803));
    outputs(2268) <= not((layer0_outputs(623)) xor (layer0_outputs(1868)));
    outputs(2269) <= not(layer0_outputs(2183));
    outputs(2270) <= not((layer0_outputs(664)) or (layer0_outputs(448)));
    outputs(2271) <= (layer0_outputs(789)) and (layer0_outputs(1250));
    outputs(2272) <= layer0_outputs(1274);
    outputs(2273) <= not((layer0_outputs(1865)) or (layer0_outputs(1194)));
    outputs(2274) <= not(layer0_outputs(1750));
    outputs(2275) <= not((layer0_outputs(2234)) xor (layer0_outputs(1898)));
    outputs(2276) <= not(layer0_outputs(471));
    outputs(2277) <= not(layer0_outputs(2247)) or (layer0_outputs(2159));
    outputs(2278) <= not(layer0_outputs(887));
    outputs(2279) <= (layer0_outputs(575)) and (layer0_outputs(2209));
    outputs(2280) <= layer0_outputs(1966);
    outputs(2281) <= not(layer0_outputs(1295));
    outputs(2282) <= not(layer0_outputs(1841)) or (layer0_outputs(2046));
    outputs(2283) <= not(layer0_outputs(887)) or (layer0_outputs(1474));
    outputs(2284) <= not(layer0_outputs(2026));
    outputs(2285) <= (layer0_outputs(1143)) and not (layer0_outputs(2347));
    outputs(2286) <= not((layer0_outputs(894)) or (layer0_outputs(516)));
    outputs(2287) <= layer0_outputs(1160);
    outputs(2288) <= (layer0_outputs(1563)) and (layer0_outputs(680));
    outputs(2289) <= not((layer0_outputs(721)) or (layer0_outputs(2398)));
    outputs(2290) <= not(layer0_outputs(2021));
    outputs(2291) <= (layer0_outputs(2477)) or (layer0_outputs(1386));
    outputs(2292) <= not(layer0_outputs(1598)) or (layer0_outputs(1059));
    outputs(2293) <= not(layer0_outputs(1681)) or (layer0_outputs(1240));
    outputs(2294) <= (layer0_outputs(1491)) xor (layer0_outputs(284));
    outputs(2295) <= layer0_outputs(2519);
    outputs(2296) <= not(layer0_outputs(2107));
    outputs(2297) <= not((layer0_outputs(699)) or (layer0_outputs(19)));
    outputs(2298) <= layer0_outputs(1202);
    outputs(2299) <= layer0_outputs(151);
    outputs(2300) <= (layer0_outputs(1890)) or (layer0_outputs(2498));
    outputs(2301) <= not(layer0_outputs(2151));
    outputs(2302) <= (layer0_outputs(1811)) and not (layer0_outputs(141));
    outputs(2303) <= not(layer0_outputs(792));
    outputs(2304) <= not(layer0_outputs(348));
    outputs(2305) <= not(layer0_outputs(57));
    outputs(2306) <= not(layer0_outputs(2090));
    outputs(2307) <= not(layer0_outputs(1164)) or (layer0_outputs(1767));
    outputs(2308) <= (layer0_outputs(2214)) xor (layer0_outputs(713));
    outputs(2309) <= not(layer0_outputs(2384));
    outputs(2310) <= layer0_outputs(1096);
    outputs(2311) <= layer0_outputs(1958);
    outputs(2312) <= (layer0_outputs(927)) and not (layer0_outputs(499));
    outputs(2313) <= not((layer0_outputs(1392)) or (layer0_outputs(1651)));
    outputs(2314) <= (layer0_outputs(159)) and not (layer0_outputs(464));
    outputs(2315) <= (layer0_outputs(1538)) and not (layer0_outputs(531));
    outputs(2316) <= (layer0_outputs(511)) and (layer0_outputs(436));
    outputs(2317) <= layer0_outputs(1413);
    outputs(2318) <= layer0_outputs(2342);
    outputs(2319) <= layer0_outputs(822);
    outputs(2320) <= (layer0_outputs(2075)) and not (layer0_outputs(1018));
    outputs(2321) <= layer0_outputs(1741);
    outputs(2322) <= (layer0_outputs(590)) and (layer0_outputs(1336));
    outputs(2323) <= (layer0_outputs(1222)) and (layer0_outputs(861));
    outputs(2324) <= not((layer0_outputs(1167)) or (layer0_outputs(1668)));
    outputs(2325) <= not(layer0_outputs(2175));
    outputs(2326) <= (layer0_outputs(1957)) and (layer0_outputs(943));
    outputs(2327) <= layer0_outputs(2459);
    outputs(2328) <= (layer0_outputs(58)) or (layer0_outputs(1186));
    outputs(2329) <= not(layer0_outputs(733)) or (layer0_outputs(2031));
    outputs(2330) <= not(layer0_outputs(2434));
    outputs(2331) <= not((layer0_outputs(88)) or (layer0_outputs(90)));
    outputs(2332) <= not((layer0_outputs(161)) or (layer0_outputs(1571)));
    outputs(2333) <= (layer0_outputs(652)) and (layer0_outputs(897));
    outputs(2334) <= (layer0_outputs(1745)) and (layer0_outputs(101));
    outputs(2335) <= not((layer0_outputs(15)) or (layer0_outputs(635)));
    outputs(2336) <= not(layer0_outputs(432));
    outputs(2337) <= (layer0_outputs(1881)) and not (layer0_outputs(277));
    outputs(2338) <= (layer0_outputs(708)) and (layer0_outputs(609));
    outputs(2339) <= layer0_outputs(1691);
    outputs(2340) <= (layer0_outputs(369)) and (layer0_outputs(2408));
    outputs(2341) <= (layer0_outputs(562)) and (layer0_outputs(122));
    outputs(2342) <= (layer0_outputs(2084)) and (layer0_outputs(2091));
    outputs(2343) <= layer0_outputs(27);
    outputs(2344) <= (layer0_outputs(662)) and not (layer0_outputs(1496));
    outputs(2345) <= layer0_outputs(1967);
    outputs(2346) <= (layer0_outputs(271)) and not (layer0_outputs(2439));
    outputs(2347) <= (layer0_outputs(996)) or (layer0_outputs(600));
    outputs(2348) <= layer0_outputs(1618);
    outputs(2349) <= layer0_outputs(2342);
    outputs(2350) <= not((layer0_outputs(2296)) or (layer0_outputs(1760)));
    outputs(2351) <= not((layer0_outputs(1929)) xor (layer0_outputs(1526)));
    outputs(2352) <= not(layer0_outputs(1464));
    outputs(2353) <= (layer0_outputs(198)) and not (layer0_outputs(2219));
    outputs(2354) <= (layer0_outputs(653)) and (layer0_outputs(2413));
    outputs(2355) <= layer0_outputs(2261);
    outputs(2356) <= layer0_outputs(1744);
    outputs(2357) <= (layer0_outputs(675)) and (layer0_outputs(861));
    outputs(2358) <= not(layer0_outputs(2272));
    outputs(2359) <= not((layer0_outputs(279)) or (layer0_outputs(46)));
    outputs(2360) <= layer0_outputs(835);
    outputs(2361) <= layer0_outputs(1253);
    outputs(2362) <= (layer0_outputs(748)) or (layer0_outputs(1486));
    outputs(2363) <= (layer0_outputs(1622)) and not (layer0_outputs(186));
    outputs(2364) <= (layer0_outputs(1313)) and not (layer0_outputs(1093));
    outputs(2365) <= not((layer0_outputs(516)) or (layer0_outputs(1214)));
    outputs(2366) <= not(layer0_outputs(2352));
    outputs(2367) <= not(layer0_outputs(669));
    outputs(2368) <= not(layer0_outputs(730));
    outputs(2369) <= (layer0_outputs(1198)) and (layer0_outputs(2208));
    outputs(2370) <= not((layer0_outputs(1455)) or (layer0_outputs(2169)));
    outputs(2371) <= layer0_outputs(468);
    outputs(2372) <= not(layer0_outputs(1061));
    outputs(2373) <= not((layer0_outputs(755)) or (layer0_outputs(553)));
    outputs(2374) <= not(layer0_outputs(649));
    outputs(2375) <= layer0_outputs(122);
    outputs(2376) <= layer0_outputs(926);
    outputs(2377) <= layer0_outputs(1256);
    outputs(2378) <= not((layer0_outputs(719)) or (layer0_outputs(1318)));
    outputs(2379) <= not((layer0_outputs(1921)) or (layer0_outputs(2184)));
    outputs(2380) <= layer0_outputs(1330);
    outputs(2381) <= (layer0_outputs(2255)) and not (layer0_outputs(301));
    outputs(2382) <= (layer0_outputs(508)) and (layer0_outputs(505));
    outputs(2383) <= layer0_outputs(988);
    outputs(2384) <= not(layer0_outputs(1230)) or (layer0_outputs(630));
    outputs(2385) <= layer0_outputs(647);
    outputs(2386) <= not(layer0_outputs(2047));
    outputs(2387) <= not(layer0_outputs(2437));
    outputs(2388) <= not(layer0_outputs(914));
    outputs(2389) <= (layer0_outputs(239)) and (layer0_outputs(1793));
    outputs(2390) <= not((layer0_outputs(1341)) or (layer0_outputs(366)));
    outputs(2391) <= (layer0_outputs(449)) and not (layer0_outputs(879));
    outputs(2392) <= (layer0_outputs(1683)) and not (layer0_outputs(895));
    outputs(2393) <= (layer0_outputs(1762)) and not (layer0_outputs(746));
    outputs(2394) <= layer0_outputs(468);
    outputs(2395) <= not(layer0_outputs(1751));
    outputs(2396) <= not(layer0_outputs(2388));
    outputs(2397) <= not(layer0_outputs(804));
    outputs(2398) <= (layer0_outputs(1971)) or (layer0_outputs(2144));
    outputs(2399) <= not((layer0_outputs(2497)) and (layer0_outputs(531)));
    outputs(2400) <= (layer0_outputs(898)) and not (layer0_outputs(1317));
    outputs(2401) <= (layer0_outputs(219)) and (layer0_outputs(2029));
    outputs(2402) <= not(layer0_outputs(810));
    outputs(2403) <= (layer0_outputs(2265)) and not (layer0_outputs(92));
    outputs(2404) <= layer0_outputs(1039);
    outputs(2405) <= layer0_outputs(2101);
    outputs(2406) <= layer0_outputs(484);
    outputs(2407) <= not((layer0_outputs(541)) xor (layer0_outputs(2169)));
    outputs(2408) <= not((layer0_outputs(1248)) xor (layer0_outputs(1864)));
    outputs(2409) <= not(layer0_outputs(438));
    outputs(2410) <= (layer0_outputs(587)) and not (layer0_outputs(1554));
    outputs(2411) <= (layer0_outputs(1766)) and not (layer0_outputs(546));
    outputs(2412) <= (layer0_outputs(1467)) and not (layer0_outputs(1613));
    outputs(2413) <= (layer0_outputs(1052)) and (layer0_outputs(2432));
    outputs(2414) <= (layer0_outputs(716)) and not (layer0_outputs(1569));
    outputs(2415) <= (layer0_outputs(1188)) and not (layer0_outputs(1035));
    outputs(2416) <= layer0_outputs(1602);
    outputs(2417) <= (layer0_outputs(1401)) and not (layer0_outputs(1542));
    outputs(2418) <= not((layer0_outputs(818)) or (layer0_outputs(1682)));
    outputs(2419) <= (layer0_outputs(2317)) and (layer0_outputs(2366));
    outputs(2420) <= not((layer0_outputs(1247)) or (layer0_outputs(2241)));
    outputs(2421) <= not(layer0_outputs(616)) or (layer0_outputs(692));
    outputs(2422) <= (layer0_outputs(113)) and not (layer0_outputs(700));
    outputs(2423) <= layer0_outputs(1253);
    outputs(2424) <= (layer0_outputs(193)) and not (layer0_outputs(1636));
    outputs(2425) <= layer0_outputs(1481);
    outputs(2426) <= (layer0_outputs(113)) and (layer0_outputs(1052));
    outputs(2427) <= (layer0_outputs(687)) and (layer0_outputs(1263));
    outputs(2428) <= not((layer0_outputs(1017)) or (layer0_outputs(1800)));
    outputs(2429) <= (layer0_outputs(115)) and not (layer0_outputs(404));
    outputs(2430) <= not(layer0_outputs(1512));
    outputs(2431) <= (layer0_outputs(1335)) and not (layer0_outputs(1438));
    outputs(2432) <= (layer0_outputs(1662)) or (layer0_outputs(1848));
    outputs(2433) <= layer0_outputs(945);
    outputs(2434) <= (layer0_outputs(1992)) and not (layer0_outputs(1982));
    outputs(2435) <= not((layer0_outputs(1750)) or (layer0_outputs(1930)));
    outputs(2436) <= not(layer0_outputs(551));
    outputs(2437) <= (layer0_outputs(2073)) and (layer0_outputs(1962));
    outputs(2438) <= (layer0_outputs(2102)) or (layer0_outputs(104));
    outputs(2439) <= (layer0_outputs(208)) xor (layer0_outputs(2048));
    outputs(2440) <= (layer0_outputs(42)) and not (layer0_outputs(1578));
    outputs(2441) <= layer0_outputs(1616);
    outputs(2442) <= layer0_outputs(312);
    outputs(2443) <= not((layer0_outputs(2180)) xor (layer0_outputs(1834)));
    outputs(2444) <= not((layer0_outputs(2439)) or (layer0_outputs(233)));
    outputs(2445) <= not(layer0_outputs(2179));
    outputs(2446) <= (layer0_outputs(1990)) and not (layer0_outputs(368));
    outputs(2447) <= not(layer0_outputs(929));
    outputs(2448) <= (layer0_outputs(1570)) and (layer0_outputs(1747));
    outputs(2449) <= not(layer0_outputs(513));
    outputs(2450) <= layer0_outputs(2377);
    outputs(2451) <= not((layer0_outputs(2442)) or (layer0_outputs(2351)));
    outputs(2452) <= not(layer0_outputs(1983));
    outputs(2453) <= not((layer0_outputs(2118)) and (layer0_outputs(2079)));
    outputs(2454) <= not(layer0_outputs(1758));
    outputs(2455) <= (layer0_outputs(774)) and (layer0_outputs(494));
    outputs(2456) <= (layer0_outputs(544)) and (layer0_outputs(1511));
    outputs(2457) <= (layer0_outputs(2556)) and (layer0_outputs(710));
    outputs(2458) <= (layer0_outputs(786)) and not (layer0_outputs(2528));
    outputs(2459) <= layer0_outputs(1265);
    outputs(2460) <= not(layer0_outputs(1512));
    outputs(2461) <= (layer0_outputs(1178)) and (layer0_outputs(1649));
    outputs(2462) <= not(layer0_outputs(2358));
    outputs(2463) <= layer0_outputs(866);
    outputs(2464) <= not(layer0_outputs(2387));
    outputs(2465) <= not(layer0_outputs(1972));
    outputs(2466) <= not((layer0_outputs(1088)) or (layer0_outputs(2387)));
    outputs(2467) <= not((layer0_outputs(1354)) or (layer0_outputs(1406)));
    outputs(2468) <= (layer0_outputs(1137)) and not (layer0_outputs(519));
    outputs(2469) <= not((layer0_outputs(1433)) or (layer0_outputs(2430)));
    outputs(2470) <= not(layer0_outputs(1042));
    outputs(2471) <= not(layer0_outputs(730));
    outputs(2472) <= layer0_outputs(621);
    outputs(2473) <= (layer0_outputs(508)) and (layer0_outputs(918));
    outputs(2474) <= layer0_outputs(79);
    outputs(2475) <= not((layer0_outputs(1485)) xor (layer0_outputs(29)));
    outputs(2476) <= (layer0_outputs(333)) and not (layer0_outputs(246));
    outputs(2477) <= (layer0_outputs(935)) and not (layer0_outputs(1963));
    outputs(2478) <= not(layer0_outputs(2007));
    outputs(2479) <= (layer0_outputs(325)) and not (layer0_outputs(1907));
    outputs(2480) <= (layer0_outputs(2194)) and not (layer0_outputs(136));
    outputs(2481) <= not(layer0_outputs(1468));
    outputs(2482) <= layer0_outputs(1992);
    outputs(2483) <= layer0_outputs(2368);
    outputs(2484) <= (layer0_outputs(415)) and (layer0_outputs(502));
    outputs(2485) <= (layer0_outputs(2323)) xor (layer0_outputs(1752));
    outputs(2486) <= not(layer0_outputs(1388));
    outputs(2487) <= (layer0_outputs(123)) and not (layer0_outputs(672));
    outputs(2488) <= (layer0_outputs(2072)) and not (layer0_outputs(2218));
    outputs(2489) <= not(layer0_outputs(1953));
    outputs(2490) <= not((layer0_outputs(953)) or (layer0_outputs(871)));
    outputs(2491) <= (layer0_outputs(1691)) and not (layer0_outputs(2541));
    outputs(2492) <= (layer0_outputs(1486)) and not (layer0_outputs(1652));
    outputs(2493) <= (layer0_outputs(396)) and not (layer0_outputs(685));
    outputs(2494) <= (layer0_outputs(1849)) xor (layer0_outputs(1154));
    outputs(2495) <= not((layer0_outputs(1417)) or (layer0_outputs(2049)));
    outputs(2496) <= not(layer0_outputs(2227));
    outputs(2497) <= (layer0_outputs(1107)) and not (layer0_outputs(2019));
    outputs(2498) <= not(layer0_outputs(1530));
    outputs(2499) <= layer0_outputs(1402);
    outputs(2500) <= layer0_outputs(988);
    outputs(2501) <= layer0_outputs(822);
    outputs(2502) <= layer0_outputs(552);
    outputs(2503) <= (layer0_outputs(1451)) and (layer0_outputs(1952));
    outputs(2504) <= not((layer0_outputs(1953)) or (layer0_outputs(932)));
    outputs(2505) <= not((layer0_outputs(2460)) or (layer0_outputs(2300)));
    outputs(2506) <= not(layer0_outputs(2131));
    outputs(2507) <= (layer0_outputs(2447)) and not (layer0_outputs(2090));
    outputs(2508) <= (layer0_outputs(1254)) or (layer0_outputs(357));
    outputs(2509) <= not((layer0_outputs(2375)) or (layer0_outputs(1902)));
    outputs(2510) <= layer0_outputs(665);
    outputs(2511) <= layer0_outputs(1918);
    outputs(2512) <= (layer0_outputs(2393)) and (layer0_outputs(768));
    outputs(2513) <= not((layer0_outputs(2283)) xor (layer0_outputs(18)));
    outputs(2514) <= not(layer0_outputs(673)) or (layer0_outputs(2115));
    outputs(2515) <= not((layer0_outputs(2315)) xor (layer0_outputs(264)));
    outputs(2516) <= (layer0_outputs(138)) and not (layer0_outputs(573));
    outputs(2517) <= (layer0_outputs(1053)) and (layer0_outputs(1394));
    outputs(2518) <= (layer0_outputs(2028)) and not (layer0_outputs(1979));
    outputs(2519) <= (layer0_outputs(2331)) and not (layer0_outputs(1495));
    outputs(2520) <= (layer0_outputs(1213)) and not (layer0_outputs(1513));
    outputs(2521) <= (layer0_outputs(1839)) and (layer0_outputs(1161));
    outputs(2522) <= (layer0_outputs(428)) and (layer0_outputs(1852));
    outputs(2523) <= (layer0_outputs(2052)) and not (layer0_outputs(879));
    outputs(2524) <= (layer0_outputs(1375)) xor (layer0_outputs(1393));
    outputs(2525) <= not(layer0_outputs(2435));
    outputs(2526) <= (layer0_outputs(807)) or (layer0_outputs(934));
    outputs(2527) <= (layer0_outputs(231)) and (layer0_outputs(718));
    outputs(2528) <= (layer0_outputs(1475)) and not (layer0_outputs(2173));
    outputs(2529) <= not(layer0_outputs(1355));
    outputs(2530) <= not((layer0_outputs(2216)) or (layer0_outputs(526)));
    outputs(2531) <= (layer0_outputs(12)) and not (layer0_outputs(265));
    outputs(2532) <= (layer0_outputs(329)) and (layer0_outputs(1414));
    outputs(2533) <= layer0_outputs(1338);
    outputs(2534) <= layer0_outputs(2446);
    outputs(2535) <= (layer0_outputs(716)) and not (layer0_outputs(848));
    outputs(2536) <= not((layer0_outputs(953)) or (layer0_outputs(1112)));
    outputs(2537) <= (layer0_outputs(1546)) or (layer0_outputs(1515));
    outputs(2538) <= not(layer0_outputs(252));
    outputs(2539) <= not(layer0_outputs(1412));
    outputs(2540) <= (layer0_outputs(857)) and not (layer0_outputs(1544));
    outputs(2541) <= not(layer0_outputs(998));
    outputs(2542) <= layer0_outputs(2132);
    outputs(2543) <= (layer0_outputs(2297)) and not (layer0_outputs(2336));
    outputs(2544) <= (layer0_outputs(460)) and not (layer0_outputs(2454));
    outputs(2545) <= not(layer0_outputs(1656));
    outputs(2546) <= (layer0_outputs(1096)) xor (layer0_outputs(2323));
    outputs(2547) <= layer0_outputs(447);
    outputs(2548) <= (layer0_outputs(2378)) and not (layer0_outputs(262));
    outputs(2549) <= (layer0_outputs(299)) and (layer0_outputs(2023));
    outputs(2550) <= (layer0_outputs(795)) and not (layer0_outputs(423));
    outputs(2551) <= layer0_outputs(935);
    outputs(2552) <= not((layer0_outputs(1788)) or (layer0_outputs(2134)));
    outputs(2553) <= layer0_outputs(557);
    outputs(2554) <= (layer0_outputs(577)) and not (layer0_outputs(891));
    outputs(2555) <= (layer0_outputs(481)) and not (layer0_outputs(1612));
    outputs(2556) <= layer0_outputs(1168);
    outputs(2557) <= (layer0_outputs(1945)) and not (layer0_outputs(1887));
    outputs(2558) <= (layer0_outputs(703)) and (layer0_outputs(414));
    outputs(2559) <= layer0_outputs(1621);

end Behavioral;
