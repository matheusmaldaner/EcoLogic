library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logic_network is
    port (
        inputs : in std_logic_vector(255 downto 0);
        outputs : out std_logic_vector(5119 downto 0)
    );
end logic_network;

architecture Behavioral of logic_network is
    signal layer0_outputs : std_logic_vector(5119 downto 0);

begin

    layer0_outputs(0) <= not(inputs(233)) or (inputs(111));
    layer0_outputs(1) <= not(inputs(54));
    layer0_outputs(2) <= not(inputs(122));
    layer0_outputs(3) <= inputs(120);
    layer0_outputs(4) <= inputs(216);
    layer0_outputs(5) <= (inputs(182)) and (inputs(4));
    layer0_outputs(6) <= (inputs(54)) or (inputs(177));
    layer0_outputs(7) <= not(inputs(207));
    layer0_outputs(8) <= '1';
    layer0_outputs(9) <= not(inputs(141));
    layer0_outputs(10) <= (inputs(106)) xor (inputs(158));
    layer0_outputs(11) <= not(inputs(101));
    layer0_outputs(12) <= not((inputs(2)) xor (inputs(77)));
    layer0_outputs(13) <= not(inputs(205));
    layer0_outputs(14) <= not((inputs(73)) or (inputs(57)));
    layer0_outputs(15) <= not(inputs(227));
    layer0_outputs(16) <= inputs(148);
    layer0_outputs(17) <= not(inputs(85));
    layer0_outputs(18) <= not(inputs(234));
    layer0_outputs(19) <= not(inputs(33));
    layer0_outputs(20) <= not(inputs(71)) or (inputs(125));
    layer0_outputs(21) <= (inputs(53)) xor (inputs(20));
    layer0_outputs(22) <= (inputs(71)) xor (inputs(96));
    layer0_outputs(23) <= not((inputs(13)) or (inputs(109)));
    layer0_outputs(24) <= not((inputs(158)) and (inputs(127)));
    layer0_outputs(25) <= not(inputs(7)) or (inputs(126));
    layer0_outputs(26) <= not((inputs(188)) and (inputs(171)));
    layer0_outputs(27) <= not(inputs(84));
    layer0_outputs(28) <= (inputs(222)) or (inputs(89));
    layer0_outputs(29) <= (inputs(127)) or (inputs(163));
    layer0_outputs(30) <= inputs(105);
    layer0_outputs(31) <= not((inputs(95)) or (inputs(179)));
    layer0_outputs(32) <= not((inputs(92)) xor (inputs(139)));
    layer0_outputs(33) <= (inputs(182)) and not (inputs(80));
    layer0_outputs(34) <= inputs(119);
    layer0_outputs(35) <= not(inputs(60));
    layer0_outputs(36) <= inputs(167);
    layer0_outputs(37) <= not(inputs(30));
    layer0_outputs(38) <= not((inputs(121)) or (inputs(153)));
    layer0_outputs(39) <= not((inputs(33)) or (inputs(58)));
    layer0_outputs(40) <= not(inputs(64)) or (inputs(128));
    layer0_outputs(41) <= not(inputs(145));
    layer0_outputs(42) <= not(inputs(23)) or (inputs(249));
    layer0_outputs(43) <= not((inputs(240)) or (inputs(197)));
    layer0_outputs(44) <= not((inputs(128)) or (inputs(146)));
    layer0_outputs(45) <= inputs(181);
    layer0_outputs(46) <= '1';
    layer0_outputs(47) <= not((inputs(128)) or (inputs(226)));
    layer0_outputs(48) <= not(inputs(228));
    layer0_outputs(49) <= inputs(70);
    layer0_outputs(50) <= (inputs(58)) xor (inputs(216));
    layer0_outputs(51) <= (inputs(211)) and not (inputs(86));
    layer0_outputs(52) <= (inputs(218)) and not (inputs(43));
    layer0_outputs(53) <= '1';
    layer0_outputs(54) <= (inputs(133)) and not (inputs(6));
    layer0_outputs(55) <= (inputs(54)) and not (inputs(127));
    layer0_outputs(56) <= not((inputs(185)) or (inputs(207)));
    layer0_outputs(57) <= inputs(147);
    layer0_outputs(58) <= not((inputs(109)) xor (inputs(103)));
    layer0_outputs(59) <= not(inputs(140));
    layer0_outputs(60) <= not((inputs(68)) or (inputs(6)));
    layer0_outputs(61) <= inputs(10);
    layer0_outputs(62) <= not(inputs(249)) or (inputs(51));
    layer0_outputs(63) <= not(inputs(40));
    layer0_outputs(64) <= not(inputs(181)) or (inputs(113));
    layer0_outputs(65) <= not((inputs(236)) xor (inputs(166)));
    layer0_outputs(66) <= (inputs(204)) or (inputs(225));
    layer0_outputs(67) <= not((inputs(62)) xor (inputs(34)));
    layer0_outputs(68) <= inputs(230);
    layer0_outputs(69) <= not(inputs(78));
    layer0_outputs(70) <= not((inputs(189)) or (inputs(216)));
    layer0_outputs(71) <= inputs(149);
    layer0_outputs(72) <= not(inputs(148));
    layer0_outputs(73) <= inputs(133);
    layer0_outputs(74) <= not(inputs(190));
    layer0_outputs(75) <= inputs(174);
    layer0_outputs(76) <= (inputs(143)) or (inputs(188));
    layer0_outputs(77) <= (inputs(27)) and not (inputs(190));
    layer0_outputs(78) <= not((inputs(222)) or (inputs(24)));
    layer0_outputs(79) <= (inputs(209)) or (inputs(188));
    layer0_outputs(80) <= not(inputs(146));
    layer0_outputs(81) <= (inputs(113)) or (inputs(160));
    layer0_outputs(82) <= inputs(10);
    layer0_outputs(83) <= (inputs(219)) or (inputs(203));
    layer0_outputs(84) <= inputs(248);
    layer0_outputs(85) <= not(inputs(109));
    layer0_outputs(86) <= (inputs(189)) and not (inputs(12));
    layer0_outputs(87) <= not((inputs(175)) or (inputs(192)));
    layer0_outputs(88) <= (inputs(34)) xor (inputs(20));
    layer0_outputs(89) <= (inputs(7)) or (inputs(222));
    layer0_outputs(90) <= (inputs(161)) or (inputs(189));
    layer0_outputs(91) <= (inputs(107)) and not (inputs(163));
    layer0_outputs(92) <= (inputs(87)) or (inputs(103));
    layer0_outputs(93) <= not(inputs(44));
    layer0_outputs(94) <= not((inputs(99)) or (inputs(144)));
    layer0_outputs(95) <= (inputs(125)) and not (inputs(64));
    layer0_outputs(96) <= inputs(38);
    layer0_outputs(97) <= not((inputs(197)) or (inputs(161)));
    layer0_outputs(98) <= not(inputs(122)) or (inputs(210));
    layer0_outputs(99) <= (inputs(187)) xor (inputs(80));
    layer0_outputs(100) <= (inputs(209)) or (inputs(24));
    layer0_outputs(101) <= (inputs(173)) xor (inputs(104));
    layer0_outputs(102) <= (inputs(211)) or (inputs(64));
    layer0_outputs(103) <= not(inputs(152)) or (inputs(223));
    layer0_outputs(104) <= not(inputs(245)) or (inputs(182));
    layer0_outputs(105) <= not(inputs(181));
    layer0_outputs(106) <= inputs(159);
    layer0_outputs(107) <= (inputs(254)) xor (inputs(96));
    layer0_outputs(108) <= not(inputs(87));
    layer0_outputs(109) <= not(inputs(27));
    layer0_outputs(110) <= not(inputs(124));
    layer0_outputs(111) <= not(inputs(117));
    layer0_outputs(112) <= not(inputs(243)) or (inputs(65));
    layer0_outputs(113) <= (inputs(22)) and not (inputs(102));
    layer0_outputs(114) <= not((inputs(27)) and (inputs(51)));
    layer0_outputs(115) <= (inputs(118)) or (inputs(235));
    layer0_outputs(116) <= inputs(138);
    layer0_outputs(117) <= not((inputs(19)) or (inputs(23)));
    layer0_outputs(118) <= (inputs(52)) or (inputs(31));
    layer0_outputs(119) <= (inputs(212)) xor (inputs(137));
    layer0_outputs(120) <= not(inputs(195));
    layer0_outputs(121) <= not(inputs(13)) or (inputs(192));
    layer0_outputs(122) <= inputs(133);
    layer0_outputs(123) <= not(inputs(26));
    layer0_outputs(124) <= not(inputs(114));
    layer0_outputs(125) <= inputs(66);
    layer0_outputs(126) <= '0';
    layer0_outputs(127) <= inputs(136);
    layer0_outputs(128) <= not(inputs(126));
    layer0_outputs(129) <= (inputs(84)) and not (inputs(73));
    layer0_outputs(130) <= (inputs(241)) and not (inputs(11));
    layer0_outputs(131) <= '1';
    layer0_outputs(132) <= (inputs(59)) and not (inputs(250));
    layer0_outputs(133) <= not((inputs(45)) and (inputs(58)));
    layer0_outputs(134) <= not((inputs(93)) or (inputs(162)));
    layer0_outputs(135) <= (inputs(232)) xor (inputs(160));
    layer0_outputs(136) <= not((inputs(42)) xor (inputs(45)));
    layer0_outputs(137) <= not((inputs(78)) xor (inputs(188)));
    layer0_outputs(138) <= not(inputs(103));
    layer0_outputs(139) <= (inputs(63)) and (inputs(59));
    layer0_outputs(140) <= inputs(4);
    layer0_outputs(141) <= not((inputs(180)) xor (inputs(79)));
    layer0_outputs(142) <= not((inputs(33)) xor (inputs(230)));
    layer0_outputs(143) <= not(inputs(228));
    layer0_outputs(144) <= inputs(116);
    layer0_outputs(145) <= (inputs(187)) or (inputs(213));
    layer0_outputs(146) <= not(inputs(106)) or (inputs(224));
    layer0_outputs(147) <= (inputs(206)) and not (inputs(110));
    layer0_outputs(148) <= not(inputs(116));
    layer0_outputs(149) <= not(inputs(99));
    layer0_outputs(150) <= not(inputs(99));
    layer0_outputs(151) <= (inputs(67)) or (inputs(7));
    layer0_outputs(152) <= not((inputs(0)) or (inputs(201)));
    layer0_outputs(153) <= (inputs(253)) or (inputs(184));
    layer0_outputs(154) <= inputs(24);
    layer0_outputs(155) <= not((inputs(80)) or (inputs(36)));
    layer0_outputs(156) <= not((inputs(200)) or (inputs(253)));
    layer0_outputs(157) <= not((inputs(73)) or (inputs(89)));
    layer0_outputs(158) <= not(inputs(38));
    layer0_outputs(159) <= not(inputs(212)) or (inputs(35));
    layer0_outputs(160) <= (inputs(99)) and not (inputs(191));
    layer0_outputs(161) <= (inputs(104)) or (inputs(9));
    layer0_outputs(162) <= inputs(10);
    layer0_outputs(163) <= (inputs(15)) or (inputs(53));
    layer0_outputs(164) <= (inputs(128)) xor (inputs(255));
    layer0_outputs(165) <= (inputs(117)) or (inputs(29));
    layer0_outputs(166) <= not(inputs(180));
    layer0_outputs(167) <= (inputs(236)) or (inputs(129));
    layer0_outputs(168) <= (inputs(205)) or (inputs(161));
    layer0_outputs(169) <= '0';
    layer0_outputs(170) <= inputs(114);
    layer0_outputs(171) <= not(inputs(102));
    layer0_outputs(172) <= not(inputs(34));
    layer0_outputs(173) <= inputs(121);
    layer0_outputs(174) <= (inputs(240)) or (inputs(200));
    layer0_outputs(175) <= inputs(112);
    layer0_outputs(176) <= not(inputs(190)) or (inputs(58));
    layer0_outputs(177) <= not((inputs(134)) or (inputs(101)));
    layer0_outputs(178) <= not(inputs(101)) or (inputs(255));
    layer0_outputs(179) <= not((inputs(243)) or (inputs(135)));
    layer0_outputs(180) <= (inputs(112)) xor (inputs(23));
    layer0_outputs(181) <= not((inputs(181)) or (inputs(13)));
    layer0_outputs(182) <= (inputs(89)) or (inputs(253));
    layer0_outputs(183) <= not((inputs(159)) or (inputs(191)));
    layer0_outputs(184) <= not((inputs(224)) or (inputs(248)));
    layer0_outputs(185) <= inputs(191);
    layer0_outputs(186) <= not((inputs(211)) xor (inputs(207)));
    layer0_outputs(187) <= (inputs(102)) and not (inputs(228));
    layer0_outputs(188) <= not((inputs(24)) or (inputs(38)));
    layer0_outputs(189) <= (inputs(222)) xor (inputs(10));
    layer0_outputs(190) <= not(inputs(158));
    layer0_outputs(191) <= inputs(163);
    layer0_outputs(192) <= (inputs(3)) xor (inputs(169));
    layer0_outputs(193) <= not(inputs(148)) or (inputs(191));
    layer0_outputs(194) <= not(inputs(156));
    layer0_outputs(195) <= inputs(74);
    layer0_outputs(196) <= inputs(232);
    layer0_outputs(197) <= (inputs(207)) or (inputs(80));
    layer0_outputs(198) <= not((inputs(189)) or (inputs(138)));
    layer0_outputs(199) <= '0';
    layer0_outputs(200) <= (inputs(243)) and not (inputs(164));
    layer0_outputs(201) <= not(inputs(102));
    layer0_outputs(202) <= not((inputs(114)) or (inputs(213)));
    layer0_outputs(203) <= not(inputs(98));
    layer0_outputs(204) <= not(inputs(151));
    layer0_outputs(205) <= (inputs(233)) and not (inputs(240));
    layer0_outputs(206) <= (inputs(208)) or (inputs(204));
    layer0_outputs(207) <= (inputs(114)) and (inputs(16));
    layer0_outputs(208) <= not(inputs(50));
    layer0_outputs(209) <= not((inputs(172)) xor (inputs(70)));
    layer0_outputs(210) <= (inputs(121)) and not (inputs(180));
    layer0_outputs(211) <= inputs(131);
    layer0_outputs(212) <= (inputs(4)) or (inputs(193));
    layer0_outputs(213) <= not(inputs(179)) or (inputs(158));
    layer0_outputs(214) <= not(inputs(213));
    layer0_outputs(215) <= inputs(193);
    layer0_outputs(216) <= inputs(27);
    layer0_outputs(217) <= inputs(148);
    layer0_outputs(218) <= not(inputs(250)) or (inputs(155));
    layer0_outputs(219) <= not(inputs(88)) or (inputs(117));
    layer0_outputs(220) <= not(inputs(88));
    layer0_outputs(221) <= not(inputs(201)) or (inputs(30));
    layer0_outputs(222) <= inputs(105);
    layer0_outputs(223) <= '0';
    layer0_outputs(224) <= not(inputs(13)) or (inputs(241));
    layer0_outputs(225) <= (inputs(244)) xor (inputs(223));
    layer0_outputs(226) <= not(inputs(166));
    layer0_outputs(227) <= not(inputs(40));
    layer0_outputs(228) <= not(inputs(77));
    layer0_outputs(229) <= inputs(116);
    layer0_outputs(230) <= (inputs(40)) and not (inputs(170));
    layer0_outputs(231) <= not(inputs(130));
    layer0_outputs(232) <= not(inputs(107));
    layer0_outputs(233) <= not(inputs(118)) or (inputs(17));
    layer0_outputs(234) <= not(inputs(182)) or (inputs(96));
    layer0_outputs(235) <= inputs(124);
    layer0_outputs(236) <= not(inputs(24)) or (inputs(254));
    layer0_outputs(237) <= (inputs(91)) and not (inputs(161));
    layer0_outputs(238) <= (inputs(60)) and not (inputs(36));
    layer0_outputs(239) <= not((inputs(199)) or (inputs(174)));
    layer0_outputs(240) <= not(inputs(181)) or (inputs(66));
    layer0_outputs(241) <= inputs(134);
    layer0_outputs(242) <= (inputs(70)) or (inputs(128));
    layer0_outputs(243) <= inputs(85);
    layer0_outputs(244) <= inputs(116);
    layer0_outputs(245) <= (inputs(129)) xor (inputs(204));
    layer0_outputs(246) <= inputs(14);
    layer0_outputs(247) <= inputs(81);
    layer0_outputs(248) <= (inputs(31)) xor (inputs(6));
    layer0_outputs(249) <= not(inputs(82));
    layer0_outputs(250) <= (inputs(205)) or (inputs(243));
    layer0_outputs(251) <= not(inputs(10));
    layer0_outputs(252) <= inputs(87);
    layer0_outputs(253) <= not(inputs(108));
    layer0_outputs(254) <= (inputs(169)) or (inputs(205));
    layer0_outputs(255) <= (inputs(81)) and not (inputs(105));
    layer0_outputs(256) <= inputs(163);
    layer0_outputs(257) <= not(inputs(101));
    layer0_outputs(258) <= (inputs(21)) xor (inputs(160));
    layer0_outputs(259) <= (inputs(245)) and not (inputs(35));
    layer0_outputs(260) <= (inputs(99)) and not (inputs(178));
    layer0_outputs(261) <= not(inputs(24));
    layer0_outputs(262) <= inputs(180);
    layer0_outputs(263) <= (inputs(141)) and not (inputs(66));
    layer0_outputs(264) <= inputs(103);
    layer0_outputs(265) <= not((inputs(43)) or (inputs(124)));
    layer0_outputs(266) <= not(inputs(190)) or (inputs(96));
    layer0_outputs(267) <= not(inputs(93));
    layer0_outputs(268) <= not((inputs(159)) or (inputs(91)));
    layer0_outputs(269) <= (inputs(121)) and not (inputs(84));
    layer0_outputs(270) <= not(inputs(178));
    layer0_outputs(271) <= (inputs(66)) or (inputs(147));
    layer0_outputs(272) <= (inputs(245)) and not (inputs(255));
    layer0_outputs(273) <= (inputs(11)) and not (inputs(238));
    layer0_outputs(274) <= not(inputs(99));
    layer0_outputs(275) <= not((inputs(140)) or (inputs(109)));
    layer0_outputs(276) <= not((inputs(101)) or (inputs(195)));
    layer0_outputs(277) <= not((inputs(47)) or (inputs(249)));
    layer0_outputs(278) <= not((inputs(223)) xor (inputs(171)));
    layer0_outputs(279) <= (inputs(212)) and not (inputs(129));
    layer0_outputs(280) <= inputs(111);
    layer0_outputs(281) <= not((inputs(209)) or (inputs(16)));
    layer0_outputs(282) <= (inputs(71)) and not (inputs(238));
    layer0_outputs(283) <= inputs(220);
    layer0_outputs(284) <= (inputs(83)) or (inputs(95));
    layer0_outputs(285) <= inputs(168);
    layer0_outputs(286) <= (inputs(4)) or (inputs(153));
    layer0_outputs(287) <= (inputs(188)) or (inputs(169));
    layer0_outputs(288) <= not((inputs(133)) or (inputs(6)));
    layer0_outputs(289) <= not(inputs(198)) or (inputs(202));
    layer0_outputs(290) <= '1';
    layer0_outputs(291) <= (inputs(65)) or (inputs(191));
    layer0_outputs(292) <= not(inputs(191)) or (inputs(65));
    layer0_outputs(293) <= '0';
    layer0_outputs(294) <= not(inputs(200));
    layer0_outputs(295) <= inputs(103);
    layer0_outputs(296) <= (inputs(230)) xor (inputs(79));
    layer0_outputs(297) <= not(inputs(184)) or (inputs(210));
    layer0_outputs(298) <= (inputs(219)) and not (inputs(149));
    layer0_outputs(299) <= inputs(236);
    layer0_outputs(300) <= not(inputs(94));
    layer0_outputs(301) <= not(inputs(104)) or (inputs(236));
    layer0_outputs(302) <= (inputs(195)) or (inputs(8));
    layer0_outputs(303) <= (inputs(219)) or (inputs(193));
    layer0_outputs(304) <= not(inputs(142));
    layer0_outputs(305) <= not(inputs(192));
    layer0_outputs(306) <= not(inputs(113));
    layer0_outputs(307) <= not(inputs(73));
    layer0_outputs(308) <= '0';
    layer0_outputs(309) <= not(inputs(6)) or (inputs(110));
    layer0_outputs(310) <= (inputs(83)) or (inputs(62));
    layer0_outputs(311) <= not(inputs(193)) or (inputs(156));
    layer0_outputs(312) <= not(inputs(208)) or (inputs(190));
    layer0_outputs(313) <= not(inputs(5));
    layer0_outputs(314) <= not((inputs(32)) xor (inputs(138)));
    layer0_outputs(315) <= not(inputs(52));
    layer0_outputs(316) <= not(inputs(165));
    layer0_outputs(317) <= not((inputs(190)) xor (inputs(253)));
    layer0_outputs(318) <= not(inputs(41));
    layer0_outputs(319) <= (inputs(6)) and not (inputs(127));
    layer0_outputs(320) <= not(inputs(101)) or (inputs(209));
    layer0_outputs(321) <= (inputs(156)) and (inputs(110));
    layer0_outputs(322) <= (inputs(30)) and (inputs(60));
    layer0_outputs(323) <= (inputs(25)) and not (inputs(103));
    layer0_outputs(324) <= not(inputs(17));
    layer0_outputs(325) <= not(inputs(236));
    layer0_outputs(326) <= not((inputs(212)) or (inputs(146)));
    layer0_outputs(327) <= not(inputs(57));
    layer0_outputs(328) <= (inputs(251)) and not (inputs(0));
    layer0_outputs(329) <= not(inputs(93)) or (inputs(239));
    layer0_outputs(330) <= not((inputs(45)) xor (inputs(131)));
    layer0_outputs(331) <= (inputs(188)) or (inputs(174));
    layer0_outputs(332) <= (inputs(182)) and not (inputs(139));
    layer0_outputs(333) <= (inputs(132)) and not (inputs(61));
    layer0_outputs(334) <= not(inputs(27));
    layer0_outputs(335) <= inputs(187);
    layer0_outputs(336) <= (inputs(221)) or (inputs(139));
    layer0_outputs(337) <= (inputs(234)) and not (inputs(100));
    layer0_outputs(338) <= (inputs(82)) or (inputs(70));
    layer0_outputs(339) <= not((inputs(170)) or (inputs(216)));
    layer0_outputs(340) <= not(inputs(84)) or (inputs(191));
    layer0_outputs(341) <= not(inputs(48)) or (inputs(12));
    layer0_outputs(342) <= (inputs(196)) xor (inputs(152));
    layer0_outputs(343) <= not(inputs(13));
    layer0_outputs(344) <= (inputs(206)) or (inputs(247));
    layer0_outputs(345) <= not(inputs(114)) or (inputs(140));
    layer0_outputs(346) <= inputs(166);
    layer0_outputs(347) <= (inputs(106)) or (inputs(34));
    layer0_outputs(348) <= inputs(119);
    layer0_outputs(349) <= not(inputs(156)) or (inputs(66));
    layer0_outputs(350) <= inputs(147);
    layer0_outputs(351) <= (inputs(10)) or (inputs(77));
    layer0_outputs(352) <= (inputs(104)) and not (inputs(236));
    layer0_outputs(353) <= not(inputs(134));
    layer0_outputs(354) <= not((inputs(93)) and (inputs(136)));
    layer0_outputs(355) <= (inputs(175)) xor (inputs(76));
    layer0_outputs(356) <= not((inputs(219)) or (inputs(203)));
    layer0_outputs(357) <= not(inputs(119));
    layer0_outputs(358) <= not(inputs(27));
    layer0_outputs(359) <= inputs(114);
    layer0_outputs(360) <= inputs(13);
    layer0_outputs(361) <= not(inputs(232));
    layer0_outputs(362) <= (inputs(161)) or (inputs(54));
    layer0_outputs(363) <= not(inputs(180)) or (inputs(31));
    layer0_outputs(364) <= not(inputs(41)) or (inputs(47));
    layer0_outputs(365) <= (inputs(62)) or (inputs(191));
    layer0_outputs(366) <= not(inputs(84)) or (inputs(164));
    layer0_outputs(367) <= inputs(144);
    layer0_outputs(368) <= not((inputs(64)) and (inputs(67)));
    layer0_outputs(369) <= (inputs(37)) or (inputs(95));
    layer0_outputs(370) <= inputs(101);
    layer0_outputs(371) <= inputs(94);
    layer0_outputs(372) <= inputs(78);
    layer0_outputs(373) <= not(inputs(209));
    layer0_outputs(374) <= not((inputs(159)) or (inputs(76)));
    layer0_outputs(375) <= inputs(243);
    layer0_outputs(376) <= (inputs(249)) and not (inputs(15));
    layer0_outputs(377) <= not((inputs(65)) or (inputs(149)));
    layer0_outputs(378) <= inputs(113);
    layer0_outputs(379) <= (inputs(101)) or (inputs(163));
    layer0_outputs(380) <= (inputs(235)) or (inputs(236));
    layer0_outputs(381) <= not(inputs(187));
    layer0_outputs(382) <= not(inputs(29)) or (inputs(26));
    layer0_outputs(383) <= not(inputs(198));
    layer0_outputs(384) <= not(inputs(90));
    layer0_outputs(385) <= (inputs(148)) or (inputs(196));
    layer0_outputs(386) <= (inputs(114)) and not (inputs(71));
    layer0_outputs(387) <= inputs(151);
    layer0_outputs(388) <= '1';
    layer0_outputs(389) <= not(inputs(59));
    layer0_outputs(390) <= not(inputs(152)) or (inputs(86));
    layer0_outputs(391) <= inputs(27);
    layer0_outputs(392) <= (inputs(3)) or (inputs(124));
    layer0_outputs(393) <= not(inputs(124)) or (inputs(81));
    layer0_outputs(394) <= not(inputs(164));
    layer0_outputs(395) <= not((inputs(215)) or (inputs(191)));
    layer0_outputs(396) <= (inputs(43)) and not (inputs(30));
    layer0_outputs(397) <= not(inputs(221)) or (inputs(112));
    layer0_outputs(398) <= not(inputs(122)) or (inputs(20));
    layer0_outputs(399) <= (inputs(185)) and not (inputs(72));
    layer0_outputs(400) <= not((inputs(161)) or (inputs(227)));
    layer0_outputs(401) <= not((inputs(18)) or (inputs(164)));
    layer0_outputs(402) <= not(inputs(8));
    layer0_outputs(403) <= not(inputs(185));
    layer0_outputs(404) <= not(inputs(1)) or (inputs(97));
    layer0_outputs(405) <= not(inputs(182)) or (inputs(194));
    layer0_outputs(406) <= not((inputs(175)) xor (inputs(21)));
    layer0_outputs(407) <= (inputs(182)) xor (inputs(196));
    layer0_outputs(408) <= not((inputs(218)) and (inputs(103)));
    layer0_outputs(409) <= not((inputs(94)) or (inputs(57)));
    layer0_outputs(410) <= inputs(108);
    layer0_outputs(411) <= not(inputs(177));
    layer0_outputs(412) <= not(inputs(230));
    layer0_outputs(413) <= not((inputs(189)) xor (inputs(4)));
    layer0_outputs(414) <= (inputs(186)) and not (inputs(255));
    layer0_outputs(415) <= not(inputs(183)) or (inputs(235));
    layer0_outputs(416) <= not(inputs(227)) or (inputs(254));
    layer0_outputs(417) <= (inputs(10)) xor (inputs(17));
    layer0_outputs(418) <= (inputs(246)) and not (inputs(89));
    layer0_outputs(419) <= '0';
    layer0_outputs(420) <= not(inputs(252));
    layer0_outputs(421) <= (inputs(245)) and not (inputs(7));
    layer0_outputs(422) <= (inputs(175)) and (inputs(72));
    layer0_outputs(423) <= inputs(133);
    layer0_outputs(424) <= inputs(132);
    layer0_outputs(425) <= not(inputs(97));
    layer0_outputs(426) <= not(inputs(68));
    layer0_outputs(427) <= (inputs(205)) and not (inputs(118));
    layer0_outputs(428) <= not((inputs(0)) or (inputs(8)));
    layer0_outputs(429) <= not(inputs(241)) or (inputs(97));
    layer0_outputs(430) <= inputs(131);
    layer0_outputs(431) <= not((inputs(236)) xor (inputs(164)));
    layer0_outputs(432) <= (inputs(22)) and not (inputs(173));
    layer0_outputs(433) <= not(inputs(214));
    layer0_outputs(434) <= (inputs(60)) xor (inputs(91));
    layer0_outputs(435) <= inputs(18);
    layer0_outputs(436) <= not((inputs(226)) or (inputs(198)));
    layer0_outputs(437) <= not((inputs(62)) or (inputs(139)));
    layer0_outputs(438) <= inputs(226);
    layer0_outputs(439) <= not(inputs(118));
    layer0_outputs(440) <= (inputs(172)) xor (inputs(252));
    layer0_outputs(441) <= (inputs(145)) and not (inputs(138));
    layer0_outputs(442) <= (inputs(153)) and (inputs(107));
    layer0_outputs(443) <= not((inputs(143)) or (inputs(248)));
    layer0_outputs(444) <= not((inputs(119)) xor (inputs(88)));
    layer0_outputs(445) <= not((inputs(223)) or (inputs(238)));
    layer0_outputs(446) <= (inputs(117)) or (inputs(31));
    layer0_outputs(447) <= inputs(168);
    layer0_outputs(448) <= inputs(178);
    layer0_outputs(449) <= not(inputs(211)) or (inputs(123));
    layer0_outputs(450) <= (inputs(64)) and not (inputs(236));
    layer0_outputs(451) <= not(inputs(13));
    layer0_outputs(452) <= inputs(233);
    layer0_outputs(453) <= (inputs(22)) or (inputs(14));
    layer0_outputs(454) <= not((inputs(32)) and (inputs(211)));
    layer0_outputs(455) <= not(inputs(57));
    layer0_outputs(456) <= (inputs(115)) and not (inputs(185));
    layer0_outputs(457) <= not(inputs(249));
    layer0_outputs(458) <= not((inputs(220)) or (inputs(0)));
    layer0_outputs(459) <= not((inputs(133)) or (inputs(117)));
    layer0_outputs(460) <= not(inputs(106)) or (inputs(24));
    layer0_outputs(461) <= not(inputs(145));
    layer0_outputs(462) <= not(inputs(160));
    layer0_outputs(463) <= (inputs(152)) and (inputs(136));
    layer0_outputs(464) <= '1';
    layer0_outputs(465) <= (inputs(64)) xor (inputs(59));
    layer0_outputs(466) <= (inputs(152)) and not (inputs(42));
    layer0_outputs(467) <= (inputs(90)) or (inputs(254));
    layer0_outputs(468) <= inputs(181);
    layer0_outputs(469) <= not(inputs(210));
    layer0_outputs(470) <= (inputs(241)) or (inputs(60));
    layer0_outputs(471) <= not((inputs(85)) or (inputs(86)));
    layer0_outputs(472) <= not(inputs(76));
    layer0_outputs(473) <= (inputs(73)) or (inputs(90));
    layer0_outputs(474) <= inputs(138);
    layer0_outputs(475) <= not(inputs(187));
    layer0_outputs(476) <= not(inputs(0));
    layer0_outputs(477) <= not(inputs(61));
    layer0_outputs(478) <= (inputs(99)) and not (inputs(232));
    layer0_outputs(479) <= not(inputs(197));
    layer0_outputs(480) <= '0';
    layer0_outputs(481) <= not((inputs(252)) or (inputs(223)));
    layer0_outputs(482) <= not(inputs(29)) or (inputs(192));
    layer0_outputs(483) <= (inputs(111)) or (inputs(71));
    layer0_outputs(484) <= (inputs(169)) or (inputs(185));
    layer0_outputs(485) <= inputs(149);
    layer0_outputs(486) <= not(inputs(13)) or (inputs(237));
    layer0_outputs(487) <= (inputs(151)) xor (inputs(252));
    layer0_outputs(488) <= not(inputs(104)) or (inputs(203));
    layer0_outputs(489) <= not(inputs(201));
    layer0_outputs(490) <= (inputs(83)) and not (inputs(175));
    layer0_outputs(491) <= (inputs(21)) or (inputs(175));
    layer0_outputs(492) <= not(inputs(151)) or (inputs(54));
    layer0_outputs(493) <= '0';
    layer0_outputs(494) <= not((inputs(172)) xor (inputs(128)));
    layer0_outputs(495) <= (inputs(8)) and not (inputs(124));
    layer0_outputs(496) <= inputs(178);
    layer0_outputs(497) <= not(inputs(174));
    layer0_outputs(498) <= inputs(145);
    layer0_outputs(499) <= (inputs(5)) and not (inputs(117));
    layer0_outputs(500) <= (inputs(30)) and (inputs(1));
    layer0_outputs(501) <= (inputs(24)) or (inputs(240));
    layer0_outputs(502) <= not(inputs(135)) or (inputs(18));
    layer0_outputs(503) <= (inputs(85)) xor (inputs(113));
    layer0_outputs(504) <= (inputs(230)) or (inputs(224));
    layer0_outputs(505) <= not(inputs(31)) or (inputs(84));
    layer0_outputs(506) <= inputs(100);
    layer0_outputs(507) <= not(inputs(57)) or (inputs(18));
    layer0_outputs(508) <= not(inputs(39)) or (inputs(250));
    layer0_outputs(509) <= (inputs(215)) and (inputs(228));
    layer0_outputs(510) <= inputs(229);
    layer0_outputs(511) <= (inputs(163)) or (inputs(237));
    layer0_outputs(512) <= not(inputs(189)) or (inputs(167));
    layer0_outputs(513) <= inputs(46);
    layer0_outputs(514) <= inputs(39);
    layer0_outputs(515) <= not((inputs(156)) xor (inputs(107)));
    layer0_outputs(516) <= (inputs(117)) and not (inputs(211));
    layer0_outputs(517) <= not((inputs(253)) or (inputs(96)));
    layer0_outputs(518) <= (inputs(76)) or (inputs(189));
    layer0_outputs(519) <= (inputs(51)) and not (inputs(33));
    layer0_outputs(520) <= not((inputs(46)) xor (inputs(88)));
    layer0_outputs(521) <= (inputs(195)) and not (inputs(16));
    layer0_outputs(522) <= (inputs(211)) or (inputs(172));
    layer0_outputs(523) <= not(inputs(221));
    layer0_outputs(524) <= not((inputs(87)) xor (inputs(133)));
    layer0_outputs(525) <= inputs(192);
    layer0_outputs(526) <= not(inputs(212));
    layer0_outputs(527) <= not((inputs(220)) xor (inputs(172)));
    layer0_outputs(528) <= (inputs(248)) or (inputs(180));
    layer0_outputs(529) <= (inputs(126)) or (inputs(149));
    layer0_outputs(530) <= not(inputs(199));
    layer0_outputs(531) <= (inputs(40)) xor (inputs(18));
    layer0_outputs(532) <= not(inputs(56));
    layer0_outputs(533) <= (inputs(33)) or (inputs(44));
    layer0_outputs(534) <= not(inputs(235));
    layer0_outputs(535) <= not((inputs(5)) or (inputs(63)));
    layer0_outputs(536) <= (inputs(102)) or (inputs(83));
    layer0_outputs(537) <= inputs(147);
    layer0_outputs(538) <= (inputs(113)) or (inputs(183));
    layer0_outputs(539) <= not(inputs(217)) or (inputs(107));
    layer0_outputs(540) <= not((inputs(186)) xor (inputs(90)));
    layer0_outputs(541) <= (inputs(163)) or (inputs(52));
    layer0_outputs(542) <= not(inputs(167));
    layer0_outputs(543) <= inputs(141);
    layer0_outputs(544) <= not(inputs(211)) or (inputs(114));
    layer0_outputs(545) <= not(inputs(229)) or (inputs(15));
    layer0_outputs(546) <= (inputs(17)) and not (inputs(206));
    layer0_outputs(547) <= not((inputs(226)) or (inputs(33)));
    layer0_outputs(548) <= not(inputs(239));
    layer0_outputs(549) <= (inputs(53)) and not (inputs(142));
    layer0_outputs(550) <= (inputs(22)) and not (inputs(15));
    layer0_outputs(551) <= not(inputs(57));
    layer0_outputs(552) <= not(inputs(74)) or (inputs(157));
    layer0_outputs(553) <= not((inputs(85)) or (inputs(162)));
    layer0_outputs(554) <= (inputs(196)) xor (inputs(232));
    layer0_outputs(555) <= not(inputs(187));
    layer0_outputs(556) <= not(inputs(94));
    layer0_outputs(557) <= (inputs(157)) and not (inputs(49));
    layer0_outputs(558) <= not(inputs(230));
    layer0_outputs(559) <= not((inputs(174)) and (inputs(188)));
    layer0_outputs(560) <= not((inputs(34)) or (inputs(244)));
    layer0_outputs(561) <= not(inputs(154));
    layer0_outputs(562) <= not((inputs(40)) or (inputs(248)));
    layer0_outputs(563) <= not((inputs(18)) xor (inputs(146)));
    layer0_outputs(564) <= (inputs(186)) and not (inputs(140));
    layer0_outputs(565) <= not((inputs(20)) or (inputs(142)));
    layer0_outputs(566) <= not((inputs(237)) or (inputs(238)));
    layer0_outputs(567) <= not(inputs(21)) or (inputs(127));
    layer0_outputs(568) <= not(inputs(233));
    layer0_outputs(569) <= not((inputs(124)) or (inputs(109)));
    layer0_outputs(570) <= (inputs(223)) xor (inputs(204));
    layer0_outputs(571) <= (inputs(87)) or (inputs(79));
    layer0_outputs(572) <= not((inputs(152)) and (inputs(248)));
    layer0_outputs(573) <= inputs(35);
    layer0_outputs(574) <= inputs(199);
    layer0_outputs(575) <= not(inputs(168));
    layer0_outputs(576) <= (inputs(94)) or (inputs(65));
    layer0_outputs(577) <= (inputs(89)) xor (inputs(80));
    layer0_outputs(578) <= '0';
    layer0_outputs(579) <= (inputs(164)) and not (inputs(97));
    layer0_outputs(580) <= not(inputs(115));
    layer0_outputs(581) <= not(inputs(194));
    layer0_outputs(582) <= not(inputs(123)) or (inputs(214));
    layer0_outputs(583) <= inputs(163);
    layer0_outputs(584) <= not(inputs(211));
    layer0_outputs(585) <= not((inputs(29)) or (inputs(140)));
    layer0_outputs(586) <= not(inputs(11)) or (inputs(44));
    layer0_outputs(587) <= not((inputs(158)) xor (inputs(100)));
    layer0_outputs(588) <= (inputs(124)) xor (inputs(0));
    layer0_outputs(589) <= (inputs(46)) or (inputs(17));
    layer0_outputs(590) <= (inputs(107)) xor (inputs(120));
    layer0_outputs(591) <= (inputs(215)) and not (inputs(13));
    layer0_outputs(592) <= not((inputs(218)) or (inputs(62)));
    layer0_outputs(593) <= (inputs(74)) xor (inputs(24));
    layer0_outputs(594) <= not(inputs(83));
    layer0_outputs(595) <= inputs(116);
    layer0_outputs(596) <= inputs(154);
    layer0_outputs(597) <= (inputs(130)) or (inputs(180));
    layer0_outputs(598) <= (inputs(123)) and not (inputs(98));
    layer0_outputs(599) <= not(inputs(120));
    layer0_outputs(600) <= not(inputs(31));
    layer0_outputs(601) <= not((inputs(37)) and (inputs(37)));
    layer0_outputs(602) <= (inputs(225)) xor (inputs(209));
    layer0_outputs(603) <= not((inputs(199)) and (inputs(7)));
    layer0_outputs(604) <= not((inputs(231)) xor (inputs(60)));
    layer0_outputs(605) <= not(inputs(105)) or (inputs(145));
    layer0_outputs(606) <= not(inputs(133));
    layer0_outputs(607) <= '0';
    layer0_outputs(608) <= not(inputs(102));
    layer0_outputs(609) <= (inputs(88)) and not (inputs(47));
    layer0_outputs(610) <= not((inputs(139)) and (inputs(52)));
    layer0_outputs(611) <= inputs(195);
    layer0_outputs(612) <= not(inputs(132));
    layer0_outputs(613) <= not(inputs(41));
    layer0_outputs(614) <= (inputs(198)) and not (inputs(66));
    layer0_outputs(615) <= not(inputs(121)) or (inputs(64));
    layer0_outputs(616) <= inputs(161);
    layer0_outputs(617) <= not((inputs(23)) or (inputs(157)));
    layer0_outputs(618) <= not((inputs(144)) xor (inputs(211)));
    layer0_outputs(619) <= (inputs(196)) and not (inputs(158));
    layer0_outputs(620) <= (inputs(250)) and not (inputs(70));
    layer0_outputs(621) <= not(inputs(216));
    layer0_outputs(622) <= inputs(176);
    layer0_outputs(623) <= inputs(118);
    layer0_outputs(624) <= not(inputs(145));
    layer0_outputs(625) <= not(inputs(89));
    layer0_outputs(626) <= inputs(137);
    layer0_outputs(627) <= not(inputs(212)) or (inputs(145));
    layer0_outputs(628) <= not(inputs(171));
    layer0_outputs(629) <= (inputs(232)) and not (inputs(111));
    layer0_outputs(630) <= (inputs(15)) or (inputs(117));
    layer0_outputs(631) <= (inputs(46)) and not (inputs(170));
    layer0_outputs(632) <= inputs(177);
    layer0_outputs(633) <= not((inputs(94)) xor (inputs(122)));
    layer0_outputs(634) <= (inputs(219)) and not (inputs(44));
    layer0_outputs(635) <= inputs(144);
    layer0_outputs(636) <= not(inputs(132));
    layer0_outputs(637) <= not(inputs(196));
    layer0_outputs(638) <= (inputs(74)) and not (inputs(70));
    layer0_outputs(639) <= (inputs(77)) and not (inputs(89));
    layer0_outputs(640) <= not((inputs(135)) or (inputs(86)));
    layer0_outputs(641) <= (inputs(118)) or (inputs(164));
    layer0_outputs(642) <= not(inputs(181)) or (inputs(73));
    layer0_outputs(643) <= (inputs(74)) or (inputs(3));
    layer0_outputs(644) <= (inputs(42)) and not (inputs(158));
    layer0_outputs(645) <= inputs(75);
    layer0_outputs(646) <= inputs(152);
    layer0_outputs(647) <= inputs(71);
    layer0_outputs(648) <= not((inputs(253)) or (inputs(121)));
    layer0_outputs(649) <= (inputs(83)) or (inputs(66));
    layer0_outputs(650) <= inputs(19);
    layer0_outputs(651) <= not(inputs(145));
    layer0_outputs(652) <= not(inputs(93));
    layer0_outputs(653) <= (inputs(142)) and not (inputs(14));
    layer0_outputs(654) <= '1';
    layer0_outputs(655) <= not((inputs(174)) or (inputs(218)));
    layer0_outputs(656) <= not(inputs(78)) or (inputs(239));
    layer0_outputs(657) <= not(inputs(122));
    layer0_outputs(658) <= (inputs(68)) and not (inputs(111));
    layer0_outputs(659) <= (inputs(147)) or (inputs(121));
    layer0_outputs(660) <= not(inputs(147));
    layer0_outputs(661) <= not((inputs(19)) or (inputs(240)));
    layer0_outputs(662) <= not((inputs(251)) and (inputs(235)));
    layer0_outputs(663) <= '0';
    layer0_outputs(664) <= not((inputs(132)) xor (inputs(66)));
    layer0_outputs(665) <= not(inputs(40));
    layer0_outputs(666) <= '0';
    layer0_outputs(667) <= inputs(69);
    layer0_outputs(668) <= not((inputs(239)) or (inputs(6)));
    layer0_outputs(669) <= (inputs(76)) or (inputs(201));
    layer0_outputs(670) <= (inputs(37)) xor (inputs(73));
    layer0_outputs(671) <= not(inputs(113));
    layer0_outputs(672) <= not((inputs(237)) or (inputs(253)));
    layer0_outputs(673) <= inputs(163);
    layer0_outputs(674) <= not((inputs(92)) and (inputs(51)));
    layer0_outputs(675) <= (inputs(223)) xor (inputs(106));
    layer0_outputs(676) <= inputs(93);
    layer0_outputs(677) <= (inputs(101)) or (inputs(82));
    layer0_outputs(678) <= (inputs(35)) or (inputs(48));
    layer0_outputs(679) <= not(inputs(99)) or (inputs(170));
    layer0_outputs(680) <= not(inputs(235)) or (inputs(128));
    layer0_outputs(681) <= not(inputs(131));
    layer0_outputs(682) <= not(inputs(168)) or (inputs(168));
    layer0_outputs(683) <= not((inputs(174)) or (inputs(224)));
    layer0_outputs(684) <= not(inputs(124)) or (inputs(35));
    layer0_outputs(685) <= not(inputs(109));
    layer0_outputs(686) <= not(inputs(128));
    layer0_outputs(687) <= (inputs(36)) and not (inputs(70));
    layer0_outputs(688) <= inputs(152);
    layer0_outputs(689) <= '0';
    layer0_outputs(690) <= (inputs(243)) xor (inputs(211));
    layer0_outputs(691) <= not((inputs(222)) xor (inputs(8)));
    layer0_outputs(692) <= (inputs(142)) and not (inputs(58));
    layer0_outputs(693) <= (inputs(179)) and not (inputs(93));
    layer0_outputs(694) <= (inputs(203)) xor (inputs(219));
    layer0_outputs(695) <= not(inputs(159)) or (inputs(47));
    layer0_outputs(696) <= not((inputs(229)) or (inputs(208)));
    layer0_outputs(697) <= (inputs(4)) or (inputs(21));
    layer0_outputs(698) <= not(inputs(161)) or (inputs(165));
    layer0_outputs(699) <= not(inputs(101)) or (inputs(44));
    layer0_outputs(700) <= not(inputs(151));
    layer0_outputs(701) <= (inputs(212)) and not (inputs(24));
    layer0_outputs(702) <= '0';
    layer0_outputs(703) <= not((inputs(10)) or (inputs(132)));
    layer0_outputs(704) <= (inputs(62)) xor (inputs(11));
    layer0_outputs(705) <= not(inputs(47));
    layer0_outputs(706) <= inputs(91);
    layer0_outputs(707) <= not(inputs(217)) or (inputs(81));
    layer0_outputs(708) <= not(inputs(86));
    layer0_outputs(709) <= not(inputs(86));
    layer0_outputs(710) <= not(inputs(181)) or (inputs(12));
    layer0_outputs(711) <= not((inputs(179)) xor (inputs(87)));
    layer0_outputs(712) <= (inputs(212)) and not (inputs(5));
    layer0_outputs(713) <= not((inputs(180)) or (inputs(239)));
    layer0_outputs(714) <= (inputs(154)) and not (inputs(45));
    layer0_outputs(715) <= (inputs(68)) and not (inputs(91));
    layer0_outputs(716) <= (inputs(89)) and not (inputs(64));
    layer0_outputs(717) <= inputs(83);
    layer0_outputs(718) <= not((inputs(17)) or (inputs(32)));
    layer0_outputs(719) <= not(inputs(152)) or (inputs(65));
    layer0_outputs(720) <= inputs(197);
    layer0_outputs(721) <= (inputs(121)) and not (inputs(144));
    layer0_outputs(722) <= inputs(141);
    layer0_outputs(723) <= not((inputs(27)) xor (inputs(72)));
    layer0_outputs(724) <= not((inputs(20)) or (inputs(120)));
    layer0_outputs(725) <= inputs(130);
    layer0_outputs(726) <= not(inputs(11));
    layer0_outputs(727) <= inputs(229);
    layer0_outputs(728) <= (inputs(103)) and not (inputs(35));
    layer0_outputs(729) <= inputs(127);
    layer0_outputs(730) <= (inputs(112)) and not (inputs(240));
    layer0_outputs(731) <= inputs(90);
    layer0_outputs(732) <= not(inputs(197)) or (inputs(171));
    layer0_outputs(733) <= inputs(151);
    layer0_outputs(734) <= (inputs(135)) and not (inputs(13));
    layer0_outputs(735) <= inputs(158);
    layer0_outputs(736) <= not(inputs(173));
    layer0_outputs(737) <= (inputs(216)) and not (inputs(107));
    layer0_outputs(738) <= (inputs(154)) and not (inputs(254));
    layer0_outputs(739) <= not(inputs(83)) or (inputs(76));
    layer0_outputs(740) <= not(inputs(119));
    layer0_outputs(741) <= not(inputs(87));
    layer0_outputs(742) <= inputs(106);
    layer0_outputs(743) <= (inputs(10)) and not (inputs(218));
    layer0_outputs(744) <= not(inputs(104)) or (inputs(209));
    layer0_outputs(745) <= not((inputs(6)) xor (inputs(54)));
    layer0_outputs(746) <= inputs(151);
    layer0_outputs(747) <= inputs(141);
    layer0_outputs(748) <= inputs(44);
    layer0_outputs(749) <= not(inputs(28)) or (inputs(159));
    layer0_outputs(750) <= not(inputs(228));
    layer0_outputs(751) <= (inputs(82)) and (inputs(210));
    layer0_outputs(752) <= inputs(211);
    layer0_outputs(753) <= inputs(92);
    layer0_outputs(754) <= not((inputs(126)) or (inputs(139)));
    layer0_outputs(755) <= not((inputs(36)) xor (inputs(193)));
    layer0_outputs(756) <= not(inputs(183));
    layer0_outputs(757) <= not(inputs(214)) or (inputs(172));
    layer0_outputs(758) <= (inputs(157)) or (inputs(122));
    layer0_outputs(759) <= not((inputs(241)) or (inputs(9)));
    layer0_outputs(760) <= not(inputs(10));
    layer0_outputs(761) <= (inputs(12)) and not (inputs(162));
    layer0_outputs(762) <= (inputs(117)) or (inputs(4));
    layer0_outputs(763) <= (inputs(234)) and not (inputs(88));
    layer0_outputs(764) <= not((inputs(237)) or (inputs(11)));
    layer0_outputs(765) <= not(inputs(227));
    layer0_outputs(766) <= '0';
    layer0_outputs(767) <= (inputs(185)) and not (inputs(40));
    layer0_outputs(768) <= not(inputs(24));
    layer0_outputs(769) <= (inputs(79)) or (inputs(84));
    layer0_outputs(770) <= inputs(233);
    layer0_outputs(771) <= (inputs(199)) and not (inputs(116));
    layer0_outputs(772) <= not(inputs(72));
    layer0_outputs(773) <= not((inputs(237)) or (inputs(22)));
    layer0_outputs(774) <= not(inputs(92));
    layer0_outputs(775) <= inputs(241);
    layer0_outputs(776) <= not(inputs(29));
    layer0_outputs(777) <= not((inputs(99)) xor (inputs(133)));
    layer0_outputs(778) <= inputs(230);
    layer0_outputs(779) <= (inputs(26)) xor (inputs(19));
    layer0_outputs(780) <= inputs(73);
    layer0_outputs(781) <= not(inputs(247)) or (inputs(223));
    layer0_outputs(782) <= not((inputs(176)) or (inputs(191)));
    layer0_outputs(783) <= (inputs(243)) or (inputs(251));
    layer0_outputs(784) <= not((inputs(6)) xor (inputs(5)));
    layer0_outputs(785) <= inputs(99);
    layer0_outputs(786) <= inputs(168);
    layer0_outputs(787) <= inputs(115);
    layer0_outputs(788) <= not((inputs(167)) or (inputs(222)));
    layer0_outputs(789) <= '1';
    layer0_outputs(790) <= inputs(251);
    layer0_outputs(791) <= (inputs(177)) or (inputs(232));
    layer0_outputs(792) <= (inputs(233)) or (inputs(180));
    layer0_outputs(793) <= inputs(255);
    layer0_outputs(794) <= not(inputs(216));
    layer0_outputs(795) <= not((inputs(217)) and (inputs(225)));
    layer0_outputs(796) <= (inputs(99)) or (inputs(53));
    layer0_outputs(797) <= inputs(83);
    layer0_outputs(798) <= (inputs(158)) xor (inputs(114));
    layer0_outputs(799) <= inputs(215);
    layer0_outputs(800) <= not((inputs(182)) or (inputs(175)));
    layer0_outputs(801) <= (inputs(37)) and (inputs(42));
    layer0_outputs(802) <= inputs(169);
    layer0_outputs(803) <= '1';
    layer0_outputs(804) <= not((inputs(15)) or (inputs(29)));
    layer0_outputs(805) <= not(inputs(214)) or (inputs(238));
    layer0_outputs(806) <= not(inputs(67)) or (inputs(169));
    layer0_outputs(807) <= not(inputs(213));
    layer0_outputs(808) <= not(inputs(148));
    layer0_outputs(809) <= not(inputs(133));
    layer0_outputs(810) <= not(inputs(26));
    layer0_outputs(811) <= (inputs(24)) and not (inputs(144));
    layer0_outputs(812) <= not(inputs(106));
    layer0_outputs(813) <= (inputs(170)) or (inputs(84));
    layer0_outputs(814) <= (inputs(197)) and not (inputs(79));
    layer0_outputs(815) <= (inputs(102)) and not (inputs(159));
    layer0_outputs(816) <= not((inputs(252)) or (inputs(228)));
    layer0_outputs(817) <= not(inputs(68)) or (inputs(141));
    layer0_outputs(818) <= (inputs(119)) and not (inputs(240));
    layer0_outputs(819) <= (inputs(205)) and (inputs(250));
    layer0_outputs(820) <= not(inputs(38)) or (inputs(239));
    layer0_outputs(821) <= not((inputs(252)) or (inputs(198)));
    layer0_outputs(822) <= (inputs(104)) and not (inputs(70));
    layer0_outputs(823) <= inputs(19);
    layer0_outputs(824) <= inputs(60);
    layer0_outputs(825) <= not((inputs(142)) or (inputs(141)));
    layer0_outputs(826) <= '1';
    layer0_outputs(827) <= not(inputs(10));
    layer0_outputs(828) <= (inputs(34)) and not (inputs(202));
    layer0_outputs(829) <= (inputs(103)) and not (inputs(98));
    layer0_outputs(830) <= not(inputs(184)) or (inputs(78));
    layer0_outputs(831) <= not(inputs(224));
    layer0_outputs(832) <= not(inputs(189));
    layer0_outputs(833) <= inputs(101);
    layer0_outputs(834) <= inputs(10);
    layer0_outputs(835) <= not(inputs(42));
    layer0_outputs(836) <= not(inputs(237)) or (inputs(66));
    layer0_outputs(837) <= not((inputs(41)) and (inputs(230)));
    layer0_outputs(838) <= (inputs(190)) or (inputs(140));
    layer0_outputs(839) <= inputs(65);
    layer0_outputs(840) <= not(inputs(74)) or (inputs(74));
    layer0_outputs(841) <= not(inputs(134)) or (inputs(172));
    layer0_outputs(842) <= (inputs(229)) or (inputs(144));
    layer0_outputs(843) <= not(inputs(134));
    layer0_outputs(844) <= inputs(163);
    layer0_outputs(845) <= not(inputs(167)) or (inputs(180));
    layer0_outputs(846) <= not((inputs(159)) or (inputs(85)));
    layer0_outputs(847) <= inputs(24);
    layer0_outputs(848) <= (inputs(197)) or (inputs(157));
    layer0_outputs(849) <= not((inputs(75)) or (inputs(207)));
    layer0_outputs(850) <= (inputs(137)) or (inputs(243));
    layer0_outputs(851) <= (inputs(130)) and (inputs(162));
    layer0_outputs(852) <= not((inputs(111)) xor (inputs(160)));
    layer0_outputs(853) <= (inputs(42)) and (inputs(115));
    layer0_outputs(854) <= not(inputs(212)) or (inputs(253));
    layer0_outputs(855) <= inputs(114);
    layer0_outputs(856) <= inputs(9);
    layer0_outputs(857) <= not(inputs(139)) or (inputs(247));
    layer0_outputs(858) <= not(inputs(122));
    layer0_outputs(859) <= not(inputs(60));
    layer0_outputs(860) <= not(inputs(20)) or (inputs(131));
    layer0_outputs(861) <= inputs(109);
    layer0_outputs(862) <= not(inputs(42));
    layer0_outputs(863) <= not((inputs(212)) or (inputs(230)));
    layer0_outputs(864) <= (inputs(75)) or (inputs(92));
    layer0_outputs(865) <= not(inputs(70));
    layer0_outputs(866) <= (inputs(192)) or (inputs(46));
    layer0_outputs(867) <= inputs(148);
    layer0_outputs(868) <= not((inputs(95)) xor (inputs(173)));
    layer0_outputs(869) <= inputs(145);
    layer0_outputs(870) <= inputs(57);
    layer0_outputs(871) <= not(inputs(82));
    layer0_outputs(872) <= not(inputs(158)) or (inputs(223));
    layer0_outputs(873) <= inputs(254);
    layer0_outputs(874) <= not(inputs(135));
    layer0_outputs(875) <= (inputs(199)) and not (inputs(202));
    layer0_outputs(876) <= not(inputs(75));
    layer0_outputs(877) <= not(inputs(101));
    layer0_outputs(878) <= not(inputs(211)) or (inputs(182));
    layer0_outputs(879) <= not(inputs(133)) or (inputs(153));
    layer0_outputs(880) <= inputs(72);
    layer0_outputs(881) <= (inputs(22)) and not (inputs(221));
    layer0_outputs(882) <= not((inputs(106)) or (inputs(112)));
    layer0_outputs(883) <= not(inputs(90)) or (inputs(3));
    layer0_outputs(884) <= (inputs(171)) or (inputs(95));
    layer0_outputs(885) <= inputs(109);
    layer0_outputs(886) <= not(inputs(197));
    layer0_outputs(887) <= inputs(45);
    layer0_outputs(888) <= not(inputs(230)) or (inputs(72));
    layer0_outputs(889) <= (inputs(113)) and not (inputs(94));
    layer0_outputs(890) <= not(inputs(58)) or (inputs(192));
    layer0_outputs(891) <= not(inputs(139)) or (inputs(75));
    layer0_outputs(892) <= not((inputs(42)) xor (inputs(45)));
    layer0_outputs(893) <= inputs(155);
    layer0_outputs(894) <= not(inputs(163)) or (inputs(48));
    layer0_outputs(895) <= (inputs(3)) or (inputs(47));
    layer0_outputs(896) <= not(inputs(165));
    layer0_outputs(897) <= (inputs(54)) and not (inputs(235));
    layer0_outputs(898) <= not((inputs(146)) or (inputs(133)));
    layer0_outputs(899) <= not(inputs(28));
    layer0_outputs(900) <= inputs(131);
    layer0_outputs(901) <= inputs(88);
    layer0_outputs(902) <= not(inputs(87)) or (inputs(204));
    layer0_outputs(903) <= inputs(133);
    layer0_outputs(904) <= not((inputs(209)) xor (inputs(177)));
    layer0_outputs(905) <= not((inputs(37)) or (inputs(116)));
    layer0_outputs(906) <= inputs(77);
    layer0_outputs(907) <= not(inputs(38)) or (inputs(63));
    layer0_outputs(908) <= (inputs(217)) and not (inputs(222));
    layer0_outputs(909) <= (inputs(102)) and not (inputs(160));
    layer0_outputs(910) <= (inputs(87)) and not (inputs(206));
    layer0_outputs(911) <= (inputs(6)) or (inputs(21));
    layer0_outputs(912) <= not((inputs(147)) or (inputs(149)));
    layer0_outputs(913) <= (inputs(66)) or (inputs(58));
    layer0_outputs(914) <= (inputs(137)) and not (inputs(2));
    layer0_outputs(915) <= (inputs(228)) and not (inputs(0));
    layer0_outputs(916) <= (inputs(220)) xor (inputs(126));
    layer0_outputs(917) <= not(inputs(150));
    layer0_outputs(918) <= not(inputs(91)) or (inputs(41));
    layer0_outputs(919) <= (inputs(147)) or (inputs(245));
    layer0_outputs(920) <= not((inputs(208)) or (inputs(32)));
    layer0_outputs(921) <= inputs(201);
    layer0_outputs(922) <= not((inputs(116)) or (inputs(86)));
    layer0_outputs(923) <= not(inputs(192)) or (inputs(47));
    layer0_outputs(924) <= not(inputs(253)) or (inputs(17));
    layer0_outputs(925) <= inputs(165);
    layer0_outputs(926) <= not(inputs(27));
    layer0_outputs(927) <= not(inputs(246));
    layer0_outputs(928) <= (inputs(121)) and not (inputs(226));
    layer0_outputs(929) <= (inputs(146)) or (inputs(246));
    layer0_outputs(930) <= (inputs(121)) xor (inputs(78));
    layer0_outputs(931) <= (inputs(1)) or (inputs(48));
    layer0_outputs(932) <= '1';
    layer0_outputs(933) <= not(inputs(42));
    layer0_outputs(934) <= (inputs(202)) and not (inputs(95));
    layer0_outputs(935) <= '1';
    layer0_outputs(936) <= not((inputs(255)) or (inputs(75)));
    layer0_outputs(937) <= not(inputs(84));
    layer0_outputs(938) <= inputs(117);
    layer0_outputs(939) <= (inputs(49)) or (inputs(42));
    layer0_outputs(940) <= not((inputs(231)) xor (inputs(147)));
    layer0_outputs(941) <= not(inputs(140)) or (inputs(111));
    layer0_outputs(942) <= not(inputs(104));
    layer0_outputs(943) <= not((inputs(4)) and (inputs(17)));
    layer0_outputs(944) <= inputs(100);
    layer0_outputs(945) <= not(inputs(195));
    layer0_outputs(946) <= not((inputs(83)) and (inputs(137)));
    layer0_outputs(947) <= not(inputs(58)) or (inputs(196));
    layer0_outputs(948) <= not(inputs(37)) or (inputs(126));
    layer0_outputs(949) <= not(inputs(0));
    layer0_outputs(950) <= not((inputs(134)) xor (inputs(119)));
    layer0_outputs(951) <= not(inputs(230)) or (inputs(208));
    layer0_outputs(952) <= not(inputs(179));
    layer0_outputs(953) <= inputs(226);
    layer0_outputs(954) <= inputs(40);
    layer0_outputs(955) <= not(inputs(150));
    layer0_outputs(956) <= inputs(215);
    layer0_outputs(957) <= not(inputs(159));
    layer0_outputs(958) <= not(inputs(169)) or (inputs(121));
    layer0_outputs(959) <= not(inputs(235)) or (inputs(112));
    layer0_outputs(960) <= inputs(193);
    layer0_outputs(961) <= (inputs(20)) and not (inputs(143));
    layer0_outputs(962) <= inputs(196);
    layer0_outputs(963) <= not(inputs(189));
    layer0_outputs(964) <= (inputs(124)) or (inputs(126));
    layer0_outputs(965) <= (inputs(202)) and not (inputs(74));
    layer0_outputs(966) <= (inputs(247)) or (inputs(247));
    layer0_outputs(967) <= (inputs(168)) and not (inputs(43));
    layer0_outputs(968) <= not((inputs(164)) or (inputs(221)));
    layer0_outputs(969) <= not((inputs(100)) xor (inputs(178)));
    layer0_outputs(970) <= not((inputs(66)) xor (inputs(68)));
    layer0_outputs(971) <= inputs(12);
    layer0_outputs(972) <= not(inputs(90));
    layer0_outputs(973) <= (inputs(157)) or (inputs(194));
    layer0_outputs(974) <= not((inputs(97)) or (inputs(239)));
    layer0_outputs(975) <= not(inputs(21)) or (inputs(184));
    layer0_outputs(976) <= (inputs(196)) and not (inputs(65));
    layer0_outputs(977) <= not(inputs(196));
    layer0_outputs(978) <= not(inputs(218)) or (inputs(243));
    layer0_outputs(979) <= not(inputs(107)) or (inputs(0));
    layer0_outputs(980) <= (inputs(238)) and not (inputs(157));
    layer0_outputs(981) <= (inputs(155)) and not (inputs(28));
    layer0_outputs(982) <= not(inputs(61));
    layer0_outputs(983) <= not(inputs(169));
    layer0_outputs(984) <= inputs(123);
    layer0_outputs(985) <= (inputs(142)) and (inputs(62));
    layer0_outputs(986) <= '1';
    layer0_outputs(987) <= not(inputs(165));
    layer0_outputs(988) <= not(inputs(180));
    layer0_outputs(989) <= not(inputs(166));
    layer0_outputs(990) <= inputs(15);
    layer0_outputs(991) <= not(inputs(177));
    layer0_outputs(992) <= inputs(131);
    layer0_outputs(993) <= not((inputs(171)) or (inputs(234)));
    layer0_outputs(994) <= not(inputs(101));
    layer0_outputs(995) <= (inputs(158)) or (inputs(162));
    layer0_outputs(996) <= not(inputs(178)) or (inputs(170));
    layer0_outputs(997) <= inputs(130);
    layer0_outputs(998) <= (inputs(67)) or (inputs(52));
    layer0_outputs(999) <= (inputs(176)) or (inputs(162));
    layer0_outputs(1000) <= (inputs(9)) and not (inputs(227));
    layer0_outputs(1001) <= not(inputs(169));
    layer0_outputs(1002) <= (inputs(165)) xor (inputs(134));
    layer0_outputs(1003) <= not((inputs(36)) or (inputs(66)));
    layer0_outputs(1004) <= (inputs(200)) or (inputs(234));
    layer0_outputs(1005) <= not(inputs(183)) or (inputs(93));
    layer0_outputs(1006) <= inputs(213);
    layer0_outputs(1007) <= inputs(198);
    layer0_outputs(1008) <= (inputs(205)) and not (inputs(146));
    layer0_outputs(1009) <= inputs(150);
    layer0_outputs(1010) <= not((inputs(213)) or (inputs(125)));
    layer0_outputs(1011) <= not(inputs(74)) or (inputs(178));
    layer0_outputs(1012) <= inputs(162);
    layer0_outputs(1013) <= (inputs(53)) or (inputs(164));
    layer0_outputs(1014) <= (inputs(11)) and not (inputs(143));
    layer0_outputs(1015) <= not(inputs(111));
    layer0_outputs(1016) <= not(inputs(92));
    layer0_outputs(1017) <= not((inputs(45)) and (inputs(39)));
    layer0_outputs(1018) <= not((inputs(133)) xor (inputs(206)));
    layer0_outputs(1019) <= (inputs(197)) or (inputs(189));
    layer0_outputs(1020) <= (inputs(175)) or (inputs(68));
    layer0_outputs(1021) <= (inputs(249)) and not (inputs(101));
    layer0_outputs(1022) <= (inputs(123)) xor (inputs(141));
    layer0_outputs(1023) <= not(inputs(121));
    layer0_outputs(1024) <= not((inputs(182)) or (inputs(153)));
    layer0_outputs(1025) <= not(inputs(39)) or (inputs(165));
    layer0_outputs(1026) <= not(inputs(41));
    layer0_outputs(1027) <= not(inputs(149));
    layer0_outputs(1028) <= not(inputs(92)) or (inputs(252));
    layer0_outputs(1029) <= not(inputs(101));
    layer0_outputs(1030) <= not(inputs(102));
    layer0_outputs(1031) <= not(inputs(24)) or (inputs(183));
    layer0_outputs(1032) <= not(inputs(103));
    layer0_outputs(1033) <= not(inputs(131));
    layer0_outputs(1034) <= (inputs(38)) or (inputs(16));
    layer0_outputs(1035) <= not(inputs(19));
    layer0_outputs(1036) <= (inputs(242)) or (inputs(253));
    layer0_outputs(1037) <= inputs(106);
    layer0_outputs(1038) <= not(inputs(222));
    layer0_outputs(1039) <= inputs(117);
    layer0_outputs(1040) <= (inputs(91)) or (inputs(185));
    layer0_outputs(1041) <= not(inputs(152)) or (inputs(4));
    layer0_outputs(1042) <= (inputs(204)) and not (inputs(137));
    layer0_outputs(1043) <= (inputs(79)) and not (inputs(158));
    layer0_outputs(1044) <= (inputs(166)) and (inputs(198));
    layer0_outputs(1045) <= (inputs(179)) and not (inputs(129));
    layer0_outputs(1046) <= (inputs(254)) or (inputs(146));
    layer0_outputs(1047) <= not(inputs(14));
    layer0_outputs(1048) <= (inputs(33)) or (inputs(94));
    layer0_outputs(1049) <= not((inputs(207)) or (inputs(243)));
    layer0_outputs(1050) <= not(inputs(195)) or (inputs(93));
    layer0_outputs(1051) <= not((inputs(144)) xor (inputs(237)));
    layer0_outputs(1052) <= inputs(74);
    layer0_outputs(1053) <= not((inputs(168)) or (inputs(128)));
    layer0_outputs(1054) <= inputs(172);
    layer0_outputs(1055) <= not((inputs(238)) and (inputs(239)));
    layer0_outputs(1056) <= not(inputs(183)) or (inputs(31));
    layer0_outputs(1057) <= (inputs(27)) xor (inputs(126));
    layer0_outputs(1058) <= not((inputs(206)) or (inputs(41)));
    layer0_outputs(1059) <= (inputs(79)) and not (inputs(254));
    layer0_outputs(1060) <= inputs(164);
    layer0_outputs(1061) <= inputs(20);
    layer0_outputs(1062) <= (inputs(244)) xor (inputs(173));
    layer0_outputs(1063) <= not(inputs(154)) or (inputs(79));
    layer0_outputs(1064) <= (inputs(183)) and not (inputs(228));
    layer0_outputs(1065) <= inputs(12);
    layer0_outputs(1066) <= not((inputs(220)) or (inputs(239)));
    layer0_outputs(1067) <= (inputs(119)) and not (inputs(1));
    layer0_outputs(1068) <= not(inputs(132));
    layer0_outputs(1069) <= inputs(174);
    layer0_outputs(1070) <= (inputs(19)) and not (inputs(160));
    layer0_outputs(1071) <= inputs(246);
    layer0_outputs(1072) <= (inputs(52)) and not (inputs(161));
    layer0_outputs(1073) <= not(inputs(110)) or (inputs(48));
    layer0_outputs(1074) <= not(inputs(213));
    layer0_outputs(1075) <= (inputs(247)) or (inputs(44));
    layer0_outputs(1076) <= not((inputs(110)) or (inputs(11)));
    layer0_outputs(1077) <= not((inputs(32)) or (inputs(75)));
    layer0_outputs(1078) <= not(inputs(226));
    layer0_outputs(1079) <= inputs(231);
    layer0_outputs(1080) <= not(inputs(48));
    layer0_outputs(1081) <= not(inputs(97));
    layer0_outputs(1082) <= not(inputs(88));
    layer0_outputs(1083) <= not(inputs(180));
    layer0_outputs(1084) <= (inputs(1)) or (inputs(187));
    layer0_outputs(1085) <= not((inputs(124)) or (inputs(100)));
    layer0_outputs(1086) <= (inputs(20)) or (inputs(27));
    layer0_outputs(1087) <= (inputs(37)) and (inputs(247));
    layer0_outputs(1088) <= inputs(211);
    layer0_outputs(1089) <= inputs(105);
    layer0_outputs(1090) <= not(inputs(116));
    layer0_outputs(1091) <= not(inputs(100)) or (inputs(178));
    layer0_outputs(1092) <= inputs(149);
    layer0_outputs(1093) <= not(inputs(142));
    layer0_outputs(1094) <= not((inputs(94)) or (inputs(53)));
    layer0_outputs(1095) <= inputs(142);
    layer0_outputs(1096) <= not(inputs(61));
    layer0_outputs(1097) <= not(inputs(146));
    layer0_outputs(1098) <= not(inputs(39)) or (inputs(214));
    layer0_outputs(1099) <= (inputs(164)) and not (inputs(96));
    layer0_outputs(1100) <= not((inputs(161)) xor (inputs(5)));
    layer0_outputs(1101) <= not(inputs(214));
    layer0_outputs(1102) <= not(inputs(6)) or (inputs(255));
    layer0_outputs(1103) <= not(inputs(232)) or (inputs(47));
    layer0_outputs(1104) <= inputs(170);
    layer0_outputs(1105) <= (inputs(203)) or (inputs(194));
    layer0_outputs(1106) <= not(inputs(59)) or (inputs(112));
    layer0_outputs(1107) <= inputs(67);
    layer0_outputs(1108) <= inputs(183);
    layer0_outputs(1109) <= not(inputs(97)) or (inputs(215));
    layer0_outputs(1110) <= inputs(137);
    layer0_outputs(1111) <= not(inputs(234));
    layer0_outputs(1112) <= (inputs(59)) and not (inputs(255));
    layer0_outputs(1113) <= (inputs(192)) xor (inputs(79));
    layer0_outputs(1114) <= (inputs(24)) and not (inputs(255));
    layer0_outputs(1115) <= inputs(163);
    layer0_outputs(1116) <= inputs(130);
    layer0_outputs(1117) <= (inputs(34)) and not (inputs(9));
    layer0_outputs(1118) <= (inputs(108)) and not (inputs(98));
    layer0_outputs(1119) <= not((inputs(170)) and (inputs(55)));
    layer0_outputs(1120) <= inputs(20);
    layer0_outputs(1121) <= not((inputs(106)) and (inputs(76)));
    layer0_outputs(1122) <= (inputs(115)) xor (inputs(161));
    layer0_outputs(1123) <= not(inputs(60)) or (inputs(49));
    layer0_outputs(1124) <= inputs(149);
    layer0_outputs(1125) <= (inputs(132)) and not (inputs(73));
    layer0_outputs(1126) <= not((inputs(107)) xor (inputs(4)));
    layer0_outputs(1127) <= inputs(242);
    layer0_outputs(1128) <= not(inputs(235)) or (inputs(94));
    layer0_outputs(1129) <= not(inputs(61)) or (inputs(162));
    layer0_outputs(1130) <= (inputs(1)) and (inputs(240));
    layer0_outputs(1131) <= (inputs(45)) and not (inputs(255));
    layer0_outputs(1132) <= not(inputs(216)) or (inputs(3));
    layer0_outputs(1133) <= not(inputs(186));
    layer0_outputs(1134) <= (inputs(214)) and not (inputs(238));
    layer0_outputs(1135) <= not(inputs(61));
    layer0_outputs(1136) <= not((inputs(40)) xor (inputs(25)));
    layer0_outputs(1137) <= (inputs(17)) xor (inputs(108));
    layer0_outputs(1138) <= inputs(141);
    layer0_outputs(1139) <= inputs(8);
    layer0_outputs(1140) <= not(inputs(104)) or (inputs(17));
    layer0_outputs(1141) <= (inputs(105)) and not (inputs(3));
    layer0_outputs(1142) <= (inputs(32)) and not (inputs(108));
    layer0_outputs(1143) <= (inputs(126)) xor (inputs(157));
    layer0_outputs(1144) <= not(inputs(11)) or (inputs(160));
    layer0_outputs(1145) <= (inputs(86)) or (inputs(112));
    layer0_outputs(1146) <= not(inputs(57));
    layer0_outputs(1147) <= (inputs(160)) or (inputs(80));
    layer0_outputs(1148) <= (inputs(82)) xor (inputs(193));
    layer0_outputs(1149) <= not(inputs(59));
    layer0_outputs(1150) <= not(inputs(93));
    layer0_outputs(1151) <= not(inputs(200)) or (inputs(55));
    layer0_outputs(1152) <= not((inputs(211)) or (inputs(218)));
    layer0_outputs(1153) <= not(inputs(200)) or (inputs(106));
    layer0_outputs(1154) <= (inputs(220)) and not (inputs(36));
    layer0_outputs(1155) <= (inputs(207)) and (inputs(53));
    layer0_outputs(1156) <= inputs(220);
    layer0_outputs(1157) <= (inputs(226)) and not (inputs(147));
    layer0_outputs(1158) <= not((inputs(1)) xor (inputs(107)));
    layer0_outputs(1159) <= (inputs(183)) and not (inputs(124));
    layer0_outputs(1160) <= '0';
    layer0_outputs(1161) <= inputs(23);
    layer0_outputs(1162) <= not(inputs(200));
    layer0_outputs(1163) <= not(inputs(13));
    layer0_outputs(1164) <= inputs(222);
    layer0_outputs(1165) <= (inputs(107)) or (inputs(208));
    layer0_outputs(1166) <= not((inputs(170)) xor (inputs(169)));
    layer0_outputs(1167) <= (inputs(150)) and not (inputs(108));
    layer0_outputs(1168) <= inputs(116);
    layer0_outputs(1169) <= not(inputs(54));
    layer0_outputs(1170) <= not(inputs(217));
    layer0_outputs(1171) <= not(inputs(164));
    layer0_outputs(1172) <= (inputs(187)) or (inputs(97));
    layer0_outputs(1173) <= not(inputs(231));
    layer0_outputs(1174) <= not(inputs(58)) or (inputs(249));
    layer0_outputs(1175) <= inputs(190);
    layer0_outputs(1176) <= not(inputs(55));
    layer0_outputs(1177) <= inputs(56);
    layer0_outputs(1178) <= not(inputs(121));
    layer0_outputs(1179) <= inputs(120);
    layer0_outputs(1180) <= not((inputs(22)) or (inputs(36)));
    layer0_outputs(1181) <= inputs(190);
    layer0_outputs(1182) <= inputs(38);
    layer0_outputs(1183) <= not((inputs(135)) and (inputs(166)));
    layer0_outputs(1184) <= '1';
    layer0_outputs(1185) <= (inputs(186)) and not (inputs(17));
    layer0_outputs(1186) <= inputs(92);
    layer0_outputs(1187) <= not(inputs(65));
    layer0_outputs(1188) <= not(inputs(250));
    layer0_outputs(1189) <= not(inputs(208));
    layer0_outputs(1190) <= not((inputs(189)) or (inputs(206)));
    layer0_outputs(1191) <= not(inputs(215));
    layer0_outputs(1192) <= inputs(78);
    layer0_outputs(1193) <= not(inputs(33));
    layer0_outputs(1194) <= (inputs(124)) and not (inputs(132));
    layer0_outputs(1195) <= (inputs(24)) and (inputs(246));
    layer0_outputs(1196) <= not(inputs(33));
    layer0_outputs(1197) <= not((inputs(160)) or (inputs(84)));
    layer0_outputs(1198) <= not(inputs(156));
    layer0_outputs(1199) <= inputs(47);
    layer0_outputs(1200) <= not(inputs(198));
    layer0_outputs(1201) <= (inputs(119)) and not (inputs(80));
    layer0_outputs(1202) <= inputs(160);
    layer0_outputs(1203) <= inputs(66);
    layer0_outputs(1204) <= not((inputs(175)) or (inputs(22)));
    layer0_outputs(1205) <= not(inputs(28)) or (inputs(91));
    layer0_outputs(1206) <= inputs(197);
    layer0_outputs(1207) <= (inputs(148)) or (inputs(95));
    layer0_outputs(1208) <= not(inputs(213)) or (inputs(32));
    layer0_outputs(1209) <= not(inputs(45));
    layer0_outputs(1210) <= not(inputs(166));
    layer0_outputs(1211) <= not((inputs(164)) or (inputs(18)));
    layer0_outputs(1212) <= (inputs(58)) and not (inputs(216));
    layer0_outputs(1213) <= inputs(205);
    layer0_outputs(1214) <= (inputs(107)) and not (inputs(175));
    layer0_outputs(1215) <= not(inputs(181));
    layer0_outputs(1216) <= inputs(73);
    layer0_outputs(1217) <= not(inputs(130)) or (inputs(106));
    layer0_outputs(1218) <= (inputs(176)) or (inputs(85));
    layer0_outputs(1219) <= (inputs(145)) xor (inputs(211));
    layer0_outputs(1220) <= (inputs(98)) or (inputs(47));
    layer0_outputs(1221) <= not((inputs(201)) or (inputs(232)));
    layer0_outputs(1222) <= not(inputs(39));
    layer0_outputs(1223) <= not(inputs(106));
    layer0_outputs(1224) <= inputs(24);
    layer0_outputs(1225) <= not(inputs(22));
    layer0_outputs(1226) <= inputs(162);
    layer0_outputs(1227) <= (inputs(227)) or (inputs(226));
    layer0_outputs(1228) <= not((inputs(16)) or (inputs(48)));
    layer0_outputs(1229) <= not((inputs(121)) and (inputs(115)));
    layer0_outputs(1230) <= not(inputs(138)) or (inputs(207));
    layer0_outputs(1231) <= '0';
    layer0_outputs(1232) <= inputs(67);
    layer0_outputs(1233) <= (inputs(15)) or (inputs(2));
    layer0_outputs(1234) <= not((inputs(7)) xor (inputs(110)));
    layer0_outputs(1235) <= (inputs(153)) and (inputs(96));
    layer0_outputs(1236) <= not((inputs(184)) or (inputs(147)));
    layer0_outputs(1237) <= not(inputs(69)) or (inputs(157));
    layer0_outputs(1238) <= (inputs(120)) and not (inputs(191));
    layer0_outputs(1239) <= not(inputs(133));
    layer0_outputs(1240) <= not(inputs(214));
    layer0_outputs(1241) <= not((inputs(92)) or (inputs(36)));
    layer0_outputs(1242) <= not((inputs(78)) or (inputs(93)));
    layer0_outputs(1243) <= not((inputs(32)) or (inputs(104)));
    layer0_outputs(1244) <= not(inputs(125));
    layer0_outputs(1245) <= inputs(99);
    layer0_outputs(1246) <= not((inputs(117)) or (inputs(222)));
    layer0_outputs(1247) <= not(inputs(26));
    layer0_outputs(1248) <= '1';
    layer0_outputs(1249) <= not(inputs(165));
    layer0_outputs(1250) <= (inputs(136)) or (inputs(38));
    layer0_outputs(1251) <= not(inputs(31));
    layer0_outputs(1252) <= not(inputs(83)) or (inputs(203));
    layer0_outputs(1253) <= (inputs(245)) and not (inputs(244));
    layer0_outputs(1254) <= inputs(252);
    layer0_outputs(1255) <= inputs(236);
    layer0_outputs(1256) <= not((inputs(248)) or (inputs(70)));
    layer0_outputs(1257) <= not((inputs(71)) xor (inputs(66)));
    layer0_outputs(1258) <= '1';
    layer0_outputs(1259) <= (inputs(1)) or (inputs(83));
    layer0_outputs(1260) <= (inputs(108)) or (inputs(90));
    layer0_outputs(1261) <= (inputs(140)) and not (inputs(211));
    layer0_outputs(1262) <= not(inputs(92)) or (inputs(181));
    layer0_outputs(1263) <= not((inputs(72)) xor (inputs(155)));
    layer0_outputs(1264) <= inputs(248);
    layer0_outputs(1265) <= inputs(149);
    layer0_outputs(1266) <= not((inputs(193)) or (inputs(166)));
    layer0_outputs(1267) <= not(inputs(134)) or (inputs(18));
    layer0_outputs(1268) <= '1';
    layer0_outputs(1269) <= not((inputs(234)) or (inputs(191)));
    layer0_outputs(1270) <= inputs(47);
    layer0_outputs(1271) <= (inputs(95)) or (inputs(213));
    layer0_outputs(1272) <= (inputs(26)) or (inputs(191));
    layer0_outputs(1273) <= '0';
    layer0_outputs(1274) <= (inputs(60)) xor (inputs(73));
    layer0_outputs(1275) <= not((inputs(106)) or (inputs(142)));
    layer0_outputs(1276) <= (inputs(130)) or (inputs(155));
    layer0_outputs(1277) <= not(inputs(35));
    layer0_outputs(1278) <= not(inputs(170));
    layer0_outputs(1279) <= (inputs(23)) or (inputs(17));
    layer0_outputs(1280) <= (inputs(4)) or (inputs(23));
    layer0_outputs(1281) <= not((inputs(140)) or (inputs(108)));
    layer0_outputs(1282) <= not((inputs(233)) or (inputs(163)));
    layer0_outputs(1283) <= not(inputs(122)) or (inputs(255));
    layer0_outputs(1284) <= not((inputs(245)) or (inputs(72)));
    layer0_outputs(1285) <= not(inputs(47));
    layer0_outputs(1286) <= not((inputs(81)) or (inputs(70)));
    layer0_outputs(1287) <= not((inputs(125)) xor (inputs(191)));
    layer0_outputs(1288) <= not(inputs(130));
    layer0_outputs(1289) <= inputs(235);
    layer0_outputs(1290) <= '1';
    layer0_outputs(1291) <= inputs(73);
    layer0_outputs(1292) <= not(inputs(15));
    layer0_outputs(1293) <= not((inputs(220)) or (inputs(1)));
    layer0_outputs(1294) <= not(inputs(136)) or (inputs(178));
    layer0_outputs(1295) <= (inputs(173)) and not (inputs(239));
    layer0_outputs(1296) <= (inputs(141)) xor (inputs(110));
    layer0_outputs(1297) <= not((inputs(174)) or (inputs(115)));
    layer0_outputs(1298) <= not((inputs(123)) or (inputs(127)));
    layer0_outputs(1299) <= not(inputs(89));
    layer0_outputs(1300) <= (inputs(79)) or (inputs(195));
    layer0_outputs(1301) <= not((inputs(156)) or (inputs(145)));
    layer0_outputs(1302) <= not(inputs(43));
    layer0_outputs(1303) <= not((inputs(91)) and (inputs(213)));
    layer0_outputs(1304) <= (inputs(76)) or (inputs(127));
    layer0_outputs(1305) <= inputs(167);
    layer0_outputs(1306) <= not((inputs(183)) or (inputs(164)));
    layer0_outputs(1307) <= not(inputs(83)) or (inputs(131));
    layer0_outputs(1308) <= inputs(204);
    layer0_outputs(1309) <= not((inputs(32)) or (inputs(13)));
    layer0_outputs(1310) <= (inputs(159)) and (inputs(238));
    layer0_outputs(1311) <= not(inputs(83));
    layer0_outputs(1312) <= not((inputs(229)) or (inputs(198)));
    layer0_outputs(1313) <= inputs(146);
    layer0_outputs(1314) <= not(inputs(149)) or (inputs(208));
    layer0_outputs(1315) <= inputs(107);
    layer0_outputs(1316) <= not(inputs(59)) or (inputs(146));
    layer0_outputs(1317) <= not((inputs(30)) or (inputs(62)));
    layer0_outputs(1318) <= not(inputs(205));
    layer0_outputs(1319) <= not(inputs(83));
    layer0_outputs(1320) <= not(inputs(117));
    layer0_outputs(1321) <= (inputs(128)) or (inputs(43));
    layer0_outputs(1322) <= not((inputs(173)) xor (inputs(123)));
    layer0_outputs(1323) <= not(inputs(220));
    layer0_outputs(1324) <= not(inputs(46)) or (inputs(77));
    layer0_outputs(1325) <= (inputs(251)) xor (inputs(50));
    layer0_outputs(1326) <= not(inputs(36)) or (inputs(190));
    layer0_outputs(1327) <= inputs(198);
    layer0_outputs(1328) <= (inputs(120)) and not (inputs(114));
    layer0_outputs(1329) <= not(inputs(46));
    layer0_outputs(1330) <= (inputs(63)) or (inputs(85));
    layer0_outputs(1331) <= not((inputs(157)) or (inputs(3)));
    layer0_outputs(1332) <= (inputs(17)) or (inputs(45));
    layer0_outputs(1333) <= inputs(45);
    layer0_outputs(1334) <= inputs(125);
    layer0_outputs(1335) <= inputs(151);
    layer0_outputs(1336) <= not(inputs(122));
    layer0_outputs(1337) <= inputs(38);
    layer0_outputs(1338) <= not(inputs(217));
    layer0_outputs(1339) <= not(inputs(36));
    layer0_outputs(1340) <= not((inputs(152)) or (inputs(34)));
    layer0_outputs(1341) <= inputs(169);
    layer0_outputs(1342) <= inputs(47);
    layer0_outputs(1343) <= not((inputs(116)) xor (inputs(64)));
    layer0_outputs(1344) <= inputs(136);
    layer0_outputs(1345) <= (inputs(254)) xor (inputs(53));
    layer0_outputs(1346) <= not(inputs(157)) or (inputs(142));
    layer0_outputs(1347) <= (inputs(126)) or (inputs(225));
    layer0_outputs(1348) <= (inputs(143)) and not (inputs(213));
    layer0_outputs(1349) <= inputs(144);
    layer0_outputs(1350) <= not(inputs(198));
    layer0_outputs(1351) <= not(inputs(117));
    layer0_outputs(1352) <= inputs(239);
    layer0_outputs(1353) <= not((inputs(239)) xor (inputs(190)));
    layer0_outputs(1354) <= inputs(8);
    layer0_outputs(1355) <= not((inputs(153)) or (inputs(162)));
    layer0_outputs(1356) <= inputs(106);
    layer0_outputs(1357) <= not(inputs(9)) or (inputs(67));
    layer0_outputs(1358) <= not(inputs(149));
    layer0_outputs(1359) <= not(inputs(167)) or (inputs(27));
    layer0_outputs(1360) <= not(inputs(157)) or (inputs(17));
    layer0_outputs(1361) <= (inputs(177)) and not (inputs(28));
    layer0_outputs(1362) <= (inputs(38)) and not (inputs(97));
    layer0_outputs(1363) <= not(inputs(164));
    layer0_outputs(1364) <= (inputs(186)) or (inputs(172));
    layer0_outputs(1365) <= not((inputs(3)) or (inputs(130)));
    layer0_outputs(1366) <= not(inputs(87));
    layer0_outputs(1367) <= not((inputs(252)) or (inputs(193)));
    layer0_outputs(1368) <= (inputs(155)) and (inputs(215));
    layer0_outputs(1369) <= not(inputs(39));
    layer0_outputs(1370) <= not(inputs(230)) or (inputs(98));
    layer0_outputs(1371) <= '0';
    layer0_outputs(1372) <= inputs(79);
    layer0_outputs(1373) <= inputs(114);
    layer0_outputs(1374) <= (inputs(230)) or (inputs(127));
    layer0_outputs(1375) <= (inputs(176)) xor (inputs(166));
    layer0_outputs(1376) <= (inputs(22)) xor (inputs(88));
    layer0_outputs(1377) <= (inputs(233)) and (inputs(195));
    layer0_outputs(1378) <= inputs(78);
    layer0_outputs(1379) <= (inputs(20)) and not (inputs(112));
    layer0_outputs(1380) <= inputs(166);
    layer0_outputs(1381) <= not(inputs(63)) or (inputs(5));
    layer0_outputs(1382) <= not(inputs(83)) or (inputs(173));
    layer0_outputs(1383) <= (inputs(4)) or (inputs(216));
    layer0_outputs(1384) <= inputs(246);
    layer0_outputs(1385) <= not((inputs(220)) xor (inputs(127)));
    layer0_outputs(1386) <= (inputs(15)) or (inputs(192));
    layer0_outputs(1387) <= not(inputs(237)) or (inputs(32));
    layer0_outputs(1388) <= (inputs(242)) or (inputs(61));
    layer0_outputs(1389) <= inputs(100);
    layer0_outputs(1390) <= not(inputs(230));
    layer0_outputs(1391) <= inputs(90);
    layer0_outputs(1392) <= not((inputs(240)) xor (inputs(160)));
    layer0_outputs(1393) <= not(inputs(229));
    layer0_outputs(1394) <= inputs(107);
    layer0_outputs(1395) <= not((inputs(23)) xor (inputs(217)));
    layer0_outputs(1396) <= (inputs(211)) and not (inputs(166));
    layer0_outputs(1397) <= (inputs(206)) xor (inputs(194));
    layer0_outputs(1398) <= not(inputs(145));
    layer0_outputs(1399) <= not(inputs(64));
    layer0_outputs(1400) <= (inputs(51)) xor (inputs(39));
    layer0_outputs(1401) <= inputs(186);
    layer0_outputs(1402) <= not(inputs(91));
    layer0_outputs(1403) <= (inputs(28)) or (inputs(175));
    layer0_outputs(1404) <= not((inputs(82)) or (inputs(247)));
    layer0_outputs(1405) <= not((inputs(252)) or (inputs(97)));
    layer0_outputs(1406) <= (inputs(85)) and not (inputs(117));
    layer0_outputs(1407) <= not((inputs(63)) or (inputs(86)));
    layer0_outputs(1408) <= not(inputs(39));
    layer0_outputs(1409) <= not((inputs(80)) and (inputs(166)));
    layer0_outputs(1410) <= not((inputs(85)) or (inputs(192)));
    layer0_outputs(1411) <= not(inputs(185)) or (inputs(91));
    layer0_outputs(1412) <= inputs(101);
    layer0_outputs(1413) <= (inputs(55)) and not (inputs(17));
    layer0_outputs(1414) <= not(inputs(139)) or (inputs(191));
    layer0_outputs(1415) <= (inputs(206)) or (inputs(179));
    layer0_outputs(1416) <= not((inputs(55)) or (inputs(56)));
    layer0_outputs(1417) <= not(inputs(181)) or (inputs(64));
    layer0_outputs(1418) <= not(inputs(222));
    layer0_outputs(1419) <= inputs(243);
    layer0_outputs(1420) <= not(inputs(242)) or (inputs(141));
    layer0_outputs(1421) <= (inputs(237)) xor (inputs(137));
    layer0_outputs(1422) <= not(inputs(204));
    layer0_outputs(1423) <= (inputs(177)) xor (inputs(182));
    layer0_outputs(1424) <= not(inputs(212)) or (inputs(239));
    layer0_outputs(1425) <= not((inputs(183)) or (inputs(125)));
    layer0_outputs(1426) <= (inputs(89)) and not (inputs(176));
    layer0_outputs(1427) <= not((inputs(157)) xor (inputs(111)));
    layer0_outputs(1428) <= (inputs(145)) and not (inputs(254));
    layer0_outputs(1429) <= inputs(187);
    layer0_outputs(1430) <= inputs(233);
    layer0_outputs(1431) <= not(inputs(41)) or (inputs(173));
    layer0_outputs(1432) <= not(inputs(24));
    layer0_outputs(1433) <= inputs(231);
    layer0_outputs(1434) <= (inputs(221)) xor (inputs(32));
    layer0_outputs(1435) <= (inputs(133)) and not (inputs(171));
    layer0_outputs(1436) <= not((inputs(171)) or (inputs(235)));
    layer0_outputs(1437) <= inputs(245);
    layer0_outputs(1438) <= (inputs(211)) or (inputs(235));
    layer0_outputs(1439) <= (inputs(177)) and not (inputs(112));
    layer0_outputs(1440) <= (inputs(105)) and not (inputs(70));
    layer0_outputs(1441) <= not(inputs(179));
    layer0_outputs(1442) <= not(inputs(73)) or (inputs(166));
    layer0_outputs(1443) <= not(inputs(56)) or (inputs(253));
    layer0_outputs(1444) <= inputs(93);
    layer0_outputs(1445) <= not(inputs(203)) or (inputs(192));
    layer0_outputs(1446) <= (inputs(40)) or (inputs(234));
    layer0_outputs(1447) <= '0';
    layer0_outputs(1448) <= inputs(107);
    layer0_outputs(1449) <= not(inputs(92));
    layer0_outputs(1450) <= (inputs(114)) or (inputs(83));
    layer0_outputs(1451) <= (inputs(230)) or (inputs(175));
    layer0_outputs(1452) <= (inputs(106)) or (inputs(32));
    layer0_outputs(1453) <= (inputs(52)) and not (inputs(118));
    layer0_outputs(1454) <= (inputs(232)) or (inputs(230));
    layer0_outputs(1455) <= not((inputs(117)) or (inputs(111)));
    layer0_outputs(1456) <= not((inputs(171)) or (inputs(239)));
    layer0_outputs(1457) <= inputs(189);
    layer0_outputs(1458) <= not(inputs(32)) or (inputs(255));
    layer0_outputs(1459) <= inputs(26);
    layer0_outputs(1460) <= inputs(55);
    layer0_outputs(1461) <= inputs(236);
    layer0_outputs(1462) <= inputs(250);
    layer0_outputs(1463) <= not((inputs(123)) xor (inputs(75)));
    layer0_outputs(1464) <= (inputs(161)) or (inputs(127));
    layer0_outputs(1465) <= not(inputs(178));
    layer0_outputs(1466) <= not((inputs(62)) or (inputs(49)));
    layer0_outputs(1467) <= not(inputs(136)) or (inputs(10));
    layer0_outputs(1468) <= not((inputs(36)) xor (inputs(187)));
    layer0_outputs(1469) <= inputs(249);
    layer0_outputs(1470) <= not((inputs(137)) or (inputs(245)));
    layer0_outputs(1471) <= not(inputs(163));
    layer0_outputs(1472) <= (inputs(162)) or (inputs(56));
    layer0_outputs(1473) <= (inputs(251)) and (inputs(123));
    layer0_outputs(1474) <= (inputs(90)) and not (inputs(184));
    layer0_outputs(1475) <= '1';
    layer0_outputs(1476) <= inputs(81);
    layer0_outputs(1477) <= (inputs(216)) and not (inputs(9));
    layer0_outputs(1478) <= not(inputs(174));
    layer0_outputs(1479) <= (inputs(160)) xor (inputs(226));
    layer0_outputs(1480) <= (inputs(219)) or (inputs(188));
    layer0_outputs(1481) <= (inputs(163)) and not (inputs(238));
    layer0_outputs(1482) <= inputs(40);
    layer0_outputs(1483) <= not(inputs(25));
    layer0_outputs(1484) <= not(inputs(105)) or (inputs(53));
    layer0_outputs(1485) <= (inputs(7)) xor (inputs(29));
    layer0_outputs(1486) <= inputs(76);
    layer0_outputs(1487) <= '1';
    layer0_outputs(1488) <= not((inputs(210)) or (inputs(173)));
    layer0_outputs(1489) <= (inputs(150)) and not (inputs(159));
    layer0_outputs(1490) <= not(inputs(254)) or (inputs(236));
    layer0_outputs(1491) <= not(inputs(147));
    layer0_outputs(1492) <= not((inputs(9)) or (inputs(177)));
    layer0_outputs(1493) <= (inputs(214)) or (inputs(222));
    layer0_outputs(1494) <= (inputs(87)) and (inputs(50));
    layer0_outputs(1495) <= (inputs(232)) and not (inputs(102));
    layer0_outputs(1496) <= (inputs(45)) or (inputs(16));
    layer0_outputs(1497) <= not((inputs(208)) or (inputs(20)));
    layer0_outputs(1498) <= inputs(172);
    layer0_outputs(1499) <= not((inputs(240)) or (inputs(71)));
    layer0_outputs(1500) <= not((inputs(65)) or (inputs(56)));
    layer0_outputs(1501) <= (inputs(223)) xor (inputs(98));
    layer0_outputs(1502) <= inputs(232);
    layer0_outputs(1503) <= not(inputs(162));
    layer0_outputs(1504) <= not(inputs(85));
    layer0_outputs(1505) <= (inputs(66)) or (inputs(67));
    layer0_outputs(1506) <= not(inputs(141));
    layer0_outputs(1507) <= not((inputs(226)) xor (inputs(244)));
    layer0_outputs(1508) <= inputs(35);
    layer0_outputs(1509) <= inputs(152);
    layer0_outputs(1510) <= (inputs(163)) or (inputs(211));
    layer0_outputs(1511) <= not((inputs(63)) or (inputs(126)));
    layer0_outputs(1512) <= not((inputs(55)) xor (inputs(23)));
    layer0_outputs(1513) <= not(inputs(118));
    layer0_outputs(1514) <= inputs(137);
    layer0_outputs(1515) <= not(inputs(20)) or (inputs(146));
    layer0_outputs(1516) <= not(inputs(0)) or (inputs(224));
    layer0_outputs(1517) <= '1';
    layer0_outputs(1518) <= not(inputs(166));
    layer0_outputs(1519) <= (inputs(114)) or (inputs(84));
    layer0_outputs(1520) <= (inputs(11)) or (inputs(160));
    layer0_outputs(1521) <= not(inputs(98)) or (inputs(65));
    layer0_outputs(1522) <= inputs(100);
    layer0_outputs(1523) <= not((inputs(246)) xor (inputs(23)));
    layer0_outputs(1524) <= not(inputs(233));
    layer0_outputs(1525) <= (inputs(117)) and not (inputs(219));
    layer0_outputs(1526) <= (inputs(140)) and not (inputs(159));
    layer0_outputs(1527) <= (inputs(160)) xor (inputs(113));
    layer0_outputs(1528) <= (inputs(5)) and not (inputs(191));
    layer0_outputs(1529) <= not((inputs(176)) and (inputs(87)));
    layer0_outputs(1530) <= (inputs(251)) xor (inputs(174));
    layer0_outputs(1531) <= inputs(179);
    layer0_outputs(1532) <= (inputs(150)) or (inputs(196));
    layer0_outputs(1533) <= not(inputs(88)) or (inputs(48));
    layer0_outputs(1534) <= (inputs(189)) xor (inputs(236));
    layer0_outputs(1535) <= (inputs(171)) and not (inputs(253));
    layer0_outputs(1536) <= not((inputs(113)) or (inputs(227)));
    layer0_outputs(1537) <= not(inputs(12)) or (inputs(54));
    layer0_outputs(1538) <= not((inputs(81)) xor (inputs(124)));
    layer0_outputs(1539) <= inputs(71);
    layer0_outputs(1540) <= inputs(131);
    layer0_outputs(1541) <= (inputs(34)) or (inputs(4));
    layer0_outputs(1542) <= (inputs(35)) and not (inputs(28));
    layer0_outputs(1543) <= not((inputs(0)) or (inputs(149)));
    layer0_outputs(1544) <= inputs(24);
    layer0_outputs(1545) <= not((inputs(36)) and (inputs(42)));
    layer0_outputs(1546) <= not(inputs(128));
    layer0_outputs(1547) <= (inputs(56)) and not (inputs(64));
    layer0_outputs(1548) <= not((inputs(244)) or (inputs(86)));
    layer0_outputs(1549) <= (inputs(225)) or (inputs(235));
    layer0_outputs(1550) <= not(inputs(117)) or (inputs(50));
    layer0_outputs(1551) <= not((inputs(57)) and (inputs(91)));
    layer0_outputs(1552) <= not(inputs(58)) or (inputs(206));
    layer0_outputs(1553) <= '0';
    layer0_outputs(1554) <= not(inputs(87)) or (inputs(157));
    layer0_outputs(1555) <= inputs(183);
    layer0_outputs(1556) <= (inputs(250)) and not (inputs(47));
    layer0_outputs(1557) <= not(inputs(229)) or (inputs(181));
    layer0_outputs(1558) <= inputs(31);
    layer0_outputs(1559) <= not(inputs(44));
    layer0_outputs(1560) <= not(inputs(41));
    layer0_outputs(1561) <= (inputs(142)) and (inputs(128));
    layer0_outputs(1562) <= not(inputs(114));
    layer0_outputs(1563) <= inputs(195);
    layer0_outputs(1564) <= (inputs(187)) or (inputs(151));
    layer0_outputs(1565) <= not(inputs(118));
    layer0_outputs(1566) <= (inputs(133)) or (inputs(245));
    layer0_outputs(1567) <= not(inputs(138)) or (inputs(207));
    layer0_outputs(1568) <= not(inputs(59)) or (inputs(136));
    layer0_outputs(1569) <= not((inputs(194)) or (inputs(41)));
    layer0_outputs(1570) <= (inputs(38)) and not (inputs(207));
    layer0_outputs(1571) <= (inputs(140)) or (inputs(27));
    layer0_outputs(1572) <= not((inputs(119)) and (inputs(201)));
    layer0_outputs(1573) <= not(inputs(200)) or (inputs(111));
    layer0_outputs(1574) <= inputs(34);
    layer0_outputs(1575) <= not(inputs(166));
    layer0_outputs(1576) <= inputs(166);
    layer0_outputs(1577) <= inputs(166);
    layer0_outputs(1578) <= not(inputs(118));
    layer0_outputs(1579) <= not(inputs(79));
    layer0_outputs(1580) <= not(inputs(251)) or (inputs(206));
    layer0_outputs(1581) <= not(inputs(87));
    layer0_outputs(1582) <= not((inputs(146)) xor (inputs(151)));
    layer0_outputs(1583) <= inputs(128);
    layer0_outputs(1584) <= not((inputs(196)) or (inputs(213)));
    layer0_outputs(1585) <= (inputs(172)) or (inputs(253));
    layer0_outputs(1586) <= not((inputs(105)) or (inputs(189)));
    layer0_outputs(1587) <= not(inputs(106)) or (inputs(113));
    layer0_outputs(1588) <= '0';
    layer0_outputs(1589) <= inputs(230);
    layer0_outputs(1590) <= not((inputs(206)) or (inputs(19)));
    layer0_outputs(1591) <= (inputs(203)) xor (inputs(222));
    layer0_outputs(1592) <= not((inputs(129)) xor (inputs(117)));
    layer0_outputs(1593) <= not(inputs(16));
    layer0_outputs(1594) <= not(inputs(170)) or (inputs(87));
    layer0_outputs(1595) <= (inputs(36)) or (inputs(9));
    layer0_outputs(1596) <= (inputs(56)) or (inputs(77));
    layer0_outputs(1597) <= (inputs(34)) xor (inputs(76));
    layer0_outputs(1598) <= inputs(177);
    layer0_outputs(1599) <= (inputs(93)) or (inputs(110));
    layer0_outputs(1600) <= (inputs(215)) or (inputs(150));
    layer0_outputs(1601) <= not((inputs(253)) or (inputs(98)));
    layer0_outputs(1602) <= (inputs(225)) and not (inputs(60));
    layer0_outputs(1603) <= (inputs(169)) and not (inputs(132));
    layer0_outputs(1604) <= (inputs(207)) and not (inputs(129));
    layer0_outputs(1605) <= (inputs(174)) xor (inputs(194));
    layer0_outputs(1606) <= inputs(24);
    layer0_outputs(1607) <= (inputs(142)) or (inputs(164));
    layer0_outputs(1608) <= not((inputs(73)) or (inputs(42)));
    layer0_outputs(1609) <= not((inputs(199)) or (inputs(128)));
    layer0_outputs(1610) <= (inputs(209)) and (inputs(95));
    layer0_outputs(1611) <= not((inputs(140)) xor (inputs(97)));
    layer0_outputs(1612) <= inputs(27);
    layer0_outputs(1613) <= not((inputs(129)) or (inputs(179)));
    layer0_outputs(1614) <= (inputs(10)) or (inputs(126));
    layer0_outputs(1615) <= not((inputs(181)) or (inputs(205)));
    layer0_outputs(1616) <= not(inputs(160)) or (inputs(250));
    layer0_outputs(1617) <= (inputs(20)) or (inputs(29));
    layer0_outputs(1618) <= inputs(164);
    layer0_outputs(1619) <= inputs(100);
    layer0_outputs(1620) <= not(inputs(2));
    layer0_outputs(1621) <= (inputs(81)) and (inputs(194));
    layer0_outputs(1622) <= not(inputs(25));
    layer0_outputs(1623) <= (inputs(18)) and not (inputs(112));
    layer0_outputs(1624) <= not((inputs(171)) or (inputs(3)));
    layer0_outputs(1625) <= (inputs(99)) and not (inputs(206));
    layer0_outputs(1626) <= inputs(76);
    layer0_outputs(1627) <= '0';
    layer0_outputs(1628) <= not(inputs(98));
    layer0_outputs(1629) <= '0';
    layer0_outputs(1630) <= not(inputs(203));
    layer0_outputs(1631) <= (inputs(131)) or (inputs(179));
    layer0_outputs(1632) <= (inputs(57)) or (inputs(175));
    layer0_outputs(1633) <= not(inputs(21));
    layer0_outputs(1634) <= not(inputs(68));
    layer0_outputs(1635) <= not((inputs(45)) and (inputs(223)));
    layer0_outputs(1636) <= (inputs(157)) or (inputs(132));
    layer0_outputs(1637) <= inputs(233);
    layer0_outputs(1638) <= not((inputs(152)) or (inputs(221)));
    layer0_outputs(1639) <= (inputs(10)) and not (inputs(18));
    layer0_outputs(1640) <= not((inputs(110)) and (inputs(50)));
    layer0_outputs(1641) <= inputs(126);
    layer0_outputs(1642) <= (inputs(13)) or (inputs(181));
    layer0_outputs(1643) <= not(inputs(145));
    layer0_outputs(1644) <= not(inputs(25));
    layer0_outputs(1645) <= not(inputs(182));
    layer0_outputs(1646) <= (inputs(175)) or (inputs(181));
    layer0_outputs(1647) <= not(inputs(217));
    layer0_outputs(1648) <= not((inputs(206)) xor (inputs(211)));
    layer0_outputs(1649) <= (inputs(95)) xor (inputs(0));
    layer0_outputs(1650) <= not(inputs(56));
    layer0_outputs(1651) <= not(inputs(156)) or (inputs(169));
    layer0_outputs(1652) <= (inputs(204)) xor (inputs(20));
    layer0_outputs(1653) <= inputs(212);
    layer0_outputs(1654) <= not((inputs(69)) and (inputs(91)));
    layer0_outputs(1655) <= not(inputs(9));
    layer0_outputs(1656) <= not((inputs(245)) or (inputs(209)));
    layer0_outputs(1657) <= not(inputs(136));
    layer0_outputs(1658) <= not(inputs(120));
    layer0_outputs(1659) <= (inputs(130)) or (inputs(237));
    layer0_outputs(1660) <= not(inputs(117));
    layer0_outputs(1661) <= inputs(21);
    layer0_outputs(1662) <= inputs(229);
    layer0_outputs(1663) <= not(inputs(72)) or (inputs(184));
    layer0_outputs(1664) <= (inputs(116)) and not (inputs(188));
    layer0_outputs(1665) <= (inputs(156)) and not (inputs(255));
    layer0_outputs(1666) <= inputs(135);
    layer0_outputs(1667) <= not(inputs(21));
    layer0_outputs(1668) <= (inputs(251)) or (inputs(67));
    layer0_outputs(1669) <= inputs(71);
    layer0_outputs(1670) <= not(inputs(15)) or (inputs(236));
    layer0_outputs(1671) <= (inputs(94)) or (inputs(231));
    layer0_outputs(1672) <= inputs(99);
    layer0_outputs(1673) <= not(inputs(127));
    layer0_outputs(1674) <= '1';
    layer0_outputs(1675) <= not((inputs(108)) or (inputs(164)));
    layer0_outputs(1676) <= inputs(27);
    layer0_outputs(1677) <= not((inputs(8)) or (inputs(132)));
    layer0_outputs(1678) <= not((inputs(58)) or (inputs(253)));
    layer0_outputs(1679) <= inputs(185);
    layer0_outputs(1680) <= not(inputs(105));
    layer0_outputs(1681) <= (inputs(138)) and (inputs(69));
    layer0_outputs(1682) <= inputs(148);
    layer0_outputs(1683) <= not(inputs(194));
    layer0_outputs(1684) <= (inputs(211)) and not (inputs(81));
    layer0_outputs(1685) <= not(inputs(250));
    layer0_outputs(1686) <= (inputs(237)) xor (inputs(40));
    layer0_outputs(1687) <= not((inputs(45)) xor (inputs(49)));
    layer0_outputs(1688) <= '0';
    layer0_outputs(1689) <= not((inputs(143)) xor (inputs(31)));
    layer0_outputs(1690) <= inputs(163);
    layer0_outputs(1691) <= not((inputs(154)) or (inputs(175)));
    layer0_outputs(1692) <= not(inputs(88));
    layer0_outputs(1693) <= inputs(238);
    layer0_outputs(1694) <= (inputs(212)) xor (inputs(6));
    layer0_outputs(1695) <= inputs(106);
    layer0_outputs(1696) <= (inputs(4)) or (inputs(221));
    layer0_outputs(1697) <= (inputs(247)) or (inputs(30));
    layer0_outputs(1698) <= (inputs(118)) and (inputs(45));
    layer0_outputs(1699) <= not((inputs(231)) or (inputs(230)));
    layer0_outputs(1700) <= not(inputs(154)) or (inputs(70));
    layer0_outputs(1701) <= not((inputs(37)) xor (inputs(12)));
    layer0_outputs(1702) <= (inputs(105)) xor (inputs(183));
    layer0_outputs(1703) <= not(inputs(90)) or (inputs(47));
    layer0_outputs(1704) <= not(inputs(227)) or (inputs(149));
    layer0_outputs(1705) <= not((inputs(48)) or (inputs(229)));
    layer0_outputs(1706) <= not(inputs(144));
    layer0_outputs(1707) <= not((inputs(98)) or (inputs(23)));
    layer0_outputs(1708) <= not(inputs(192));
    layer0_outputs(1709) <= not((inputs(14)) or (inputs(91)));
    layer0_outputs(1710) <= not((inputs(38)) or (inputs(125)));
    layer0_outputs(1711) <= (inputs(202)) and not (inputs(59));
    layer0_outputs(1712) <= (inputs(78)) xor (inputs(7));
    layer0_outputs(1713) <= not((inputs(103)) xor (inputs(14)));
    layer0_outputs(1714) <= (inputs(252)) or (inputs(209));
    layer0_outputs(1715) <= not(inputs(135));
    layer0_outputs(1716) <= (inputs(79)) or (inputs(224));
    layer0_outputs(1717) <= inputs(74);
    layer0_outputs(1718) <= inputs(177);
    layer0_outputs(1719) <= not(inputs(60));
    layer0_outputs(1720) <= inputs(175);
    layer0_outputs(1721) <= not(inputs(223));
    layer0_outputs(1722) <= not(inputs(48)) or (inputs(218));
    layer0_outputs(1723) <= not(inputs(129)) or (inputs(20));
    layer0_outputs(1724) <= not((inputs(203)) xor (inputs(16)));
    layer0_outputs(1725) <= (inputs(5)) or (inputs(196));
    layer0_outputs(1726) <= inputs(193);
    layer0_outputs(1727) <= (inputs(105)) and not (inputs(10));
    layer0_outputs(1728) <= (inputs(133)) or (inputs(170));
    layer0_outputs(1729) <= not(inputs(20));
    layer0_outputs(1730) <= not((inputs(107)) or (inputs(223)));
    layer0_outputs(1731) <= inputs(124);
    layer0_outputs(1732) <= inputs(226);
    layer0_outputs(1733) <= not((inputs(144)) or (inputs(133)));
    layer0_outputs(1734) <= (inputs(238)) or (inputs(117));
    layer0_outputs(1735) <= (inputs(162)) or (inputs(81));
    layer0_outputs(1736) <= not(inputs(53)) or (inputs(92));
    layer0_outputs(1737) <= not((inputs(151)) and (inputs(35)));
    layer0_outputs(1738) <= (inputs(209)) or (inputs(227));
    layer0_outputs(1739) <= not(inputs(52));
    layer0_outputs(1740) <= not((inputs(50)) or (inputs(129)));
    layer0_outputs(1741) <= (inputs(202)) or (inputs(190));
    layer0_outputs(1742) <= not((inputs(80)) or (inputs(144)));
    layer0_outputs(1743) <= not((inputs(188)) and (inputs(132)));
    layer0_outputs(1744) <= inputs(118);
    layer0_outputs(1745) <= inputs(97);
    layer0_outputs(1746) <= not((inputs(55)) xor (inputs(1)));
    layer0_outputs(1747) <= not(inputs(147));
    layer0_outputs(1748) <= inputs(53);
    layer0_outputs(1749) <= (inputs(54)) or (inputs(209));
    layer0_outputs(1750) <= not(inputs(214)) or (inputs(66));
    layer0_outputs(1751) <= (inputs(63)) or (inputs(230));
    layer0_outputs(1752) <= not(inputs(107)) or (inputs(210));
    layer0_outputs(1753) <= (inputs(69)) and not (inputs(207));
    layer0_outputs(1754) <= inputs(100);
    layer0_outputs(1755) <= (inputs(104)) and not (inputs(2));
    layer0_outputs(1756) <= not((inputs(89)) or (inputs(61)));
    layer0_outputs(1757) <= inputs(123);
    layer0_outputs(1758) <= not(inputs(24));
    layer0_outputs(1759) <= (inputs(235)) or (inputs(69));
    layer0_outputs(1760) <= inputs(24);
    layer0_outputs(1761) <= (inputs(16)) xor (inputs(31));
    layer0_outputs(1762) <= not((inputs(190)) or (inputs(171)));
    layer0_outputs(1763) <= not((inputs(194)) xor (inputs(249)));
    layer0_outputs(1764) <= not(inputs(9));
    layer0_outputs(1765) <= not((inputs(147)) xor (inputs(180)));
    layer0_outputs(1766) <= not(inputs(179)) or (inputs(128));
    layer0_outputs(1767) <= inputs(229);
    layer0_outputs(1768) <= not((inputs(162)) or (inputs(146)));
    layer0_outputs(1769) <= not(inputs(82)) or (inputs(38));
    layer0_outputs(1770) <= inputs(229);
    layer0_outputs(1771) <= '0';
    layer0_outputs(1772) <= not((inputs(124)) or (inputs(251)));
    layer0_outputs(1773) <= not(inputs(178));
    layer0_outputs(1774) <= (inputs(158)) or (inputs(65));
    layer0_outputs(1775) <= inputs(248);
    layer0_outputs(1776) <= not(inputs(234));
    layer0_outputs(1777) <= not(inputs(167)) or (inputs(134));
    layer0_outputs(1778) <= not(inputs(128)) or (inputs(252));
    layer0_outputs(1779) <= '1';
    layer0_outputs(1780) <= inputs(69);
    layer0_outputs(1781) <= (inputs(92)) and not (inputs(2));
    layer0_outputs(1782) <= not(inputs(23));
    layer0_outputs(1783) <= not((inputs(237)) xor (inputs(223)));
    layer0_outputs(1784) <= inputs(29);
    layer0_outputs(1785) <= not((inputs(0)) or (inputs(48)));
    layer0_outputs(1786) <= not((inputs(157)) or (inputs(62)));
    layer0_outputs(1787) <= not(inputs(118));
    layer0_outputs(1788) <= inputs(241);
    layer0_outputs(1789) <= (inputs(1)) xor (inputs(31));
    layer0_outputs(1790) <= not((inputs(229)) or (inputs(178)));
    layer0_outputs(1791) <= not((inputs(178)) or (inputs(219)));
    layer0_outputs(1792) <= (inputs(60)) xor (inputs(49));
    layer0_outputs(1793) <= not((inputs(214)) or (inputs(200)));
    layer0_outputs(1794) <= not(inputs(50));
    layer0_outputs(1795) <= (inputs(246)) and not (inputs(31));
    layer0_outputs(1796) <= inputs(91);
    layer0_outputs(1797) <= inputs(24);
    layer0_outputs(1798) <= (inputs(84)) or (inputs(194));
    layer0_outputs(1799) <= not(inputs(88)) or (inputs(140));
    layer0_outputs(1800) <= inputs(165);
    layer0_outputs(1801) <= not(inputs(142)) or (inputs(175));
    layer0_outputs(1802) <= not((inputs(56)) xor (inputs(102)));
    layer0_outputs(1803) <= not((inputs(129)) or (inputs(244)));
    layer0_outputs(1804) <= inputs(100);
    layer0_outputs(1805) <= inputs(174);
    layer0_outputs(1806) <= not((inputs(182)) xor (inputs(222)));
    layer0_outputs(1807) <= (inputs(206)) and not (inputs(65));
    layer0_outputs(1808) <= not(inputs(164));
    layer0_outputs(1809) <= not(inputs(179));
    layer0_outputs(1810) <= not((inputs(147)) or (inputs(108)));
    layer0_outputs(1811) <= (inputs(169)) or (inputs(177));
    layer0_outputs(1812) <= not(inputs(102));
    layer0_outputs(1813) <= not((inputs(212)) or (inputs(173)));
    layer0_outputs(1814) <= not(inputs(30)) or (inputs(170));
    layer0_outputs(1815) <= not((inputs(161)) or (inputs(20)));
    layer0_outputs(1816) <= inputs(68);
    layer0_outputs(1817) <= not((inputs(21)) and (inputs(75)));
    layer0_outputs(1818) <= inputs(25);
    layer0_outputs(1819) <= not((inputs(218)) or (inputs(203)));
    layer0_outputs(1820) <= (inputs(137)) or (inputs(3));
    layer0_outputs(1821) <= not(inputs(204));
    layer0_outputs(1822) <= not(inputs(5)) or (inputs(130));
    layer0_outputs(1823) <= not(inputs(52));
    layer0_outputs(1824) <= inputs(73);
    layer0_outputs(1825) <= not(inputs(106));
    layer0_outputs(1826) <= (inputs(212)) and not (inputs(79));
    layer0_outputs(1827) <= not(inputs(226));
    layer0_outputs(1828) <= (inputs(93)) and not (inputs(99));
    layer0_outputs(1829) <= not((inputs(23)) xor (inputs(81)));
    layer0_outputs(1830) <= (inputs(142)) or (inputs(13));
    layer0_outputs(1831) <= (inputs(123)) or (inputs(31));
    layer0_outputs(1832) <= not((inputs(122)) xor (inputs(204)));
    layer0_outputs(1833) <= (inputs(46)) or (inputs(231));
    layer0_outputs(1834) <= not((inputs(46)) xor (inputs(176)));
    layer0_outputs(1835) <= (inputs(179)) or (inputs(210));
    layer0_outputs(1836) <= not(inputs(184)) or (inputs(104));
    layer0_outputs(1837) <= not(inputs(21));
    layer0_outputs(1838) <= '0';
    layer0_outputs(1839) <= inputs(40);
    layer0_outputs(1840) <= inputs(94);
    layer0_outputs(1841) <= (inputs(100)) or (inputs(92));
    layer0_outputs(1842) <= (inputs(8)) or (inputs(223));
    layer0_outputs(1843) <= (inputs(161)) or (inputs(150));
    layer0_outputs(1844) <= (inputs(233)) xor (inputs(228));
    layer0_outputs(1845) <= not(inputs(220)) or (inputs(80));
    layer0_outputs(1846) <= not((inputs(224)) or (inputs(190)));
    layer0_outputs(1847) <= not(inputs(152));
    layer0_outputs(1848) <= not((inputs(227)) or (inputs(239)));
    layer0_outputs(1849) <= not(inputs(50));
    layer0_outputs(1850) <= (inputs(76)) or (inputs(22));
    layer0_outputs(1851) <= inputs(130);
    layer0_outputs(1852) <= (inputs(139)) xor (inputs(149));
    layer0_outputs(1853) <= inputs(196);
    layer0_outputs(1854) <= not((inputs(62)) xor (inputs(181)));
    layer0_outputs(1855) <= (inputs(238)) or (inputs(203));
    layer0_outputs(1856) <= (inputs(161)) or (inputs(109));
    layer0_outputs(1857) <= (inputs(243)) xor (inputs(199));
    layer0_outputs(1858) <= not(inputs(183)) or (inputs(83));
    layer0_outputs(1859) <= (inputs(86)) and not (inputs(248));
    layer0_outputs(1860) <= not(inputs(166));
    layer0_outputs(1861) <= inputs(166);
    layer0_outputs(1862) <= (inputs(52)) or (inputs(209));
    layer0_outputs(1863) <= not((inputs(122)) or (inputs(2)));
    layer0_outputs(1864) <= inputs(120);
    layer0_outputs(1865) <= inputs(238);
    layer0_outputs(1866) <= (inputs(2)) or (inputs(139));
    layer0_outputs(1867) <= not(inputs(167));
    layer0_outputs(1868) <= not((inputs(46)) or (inputs(61)));
    layer0_outputs(1869) <= not(inputs(156));
    layer0_outputs(1870) <= (inputs(146)) or (inputs(176));
    layer0_outputs(1871) <= inputs(67);
    layer0_outputs(1872) <= not(inputs(151)) or (inputs(125));
    layer0_outputs(1873) <= not(inputs(205)) or (inputs(204));
    layer0_outputs(1874) <= inputs(44);
    layer0_outputs(1875) <= not((inputs(34)) xor (inputs(53)));
    layer0_outputs(1876) <= inputs(76);
    layer0_outputs(1877) <= not(inputs(213));
    layer0_outputs(1878) <= (inputs(183)) and not (inputs(222));
    layer0_outputs(1879) <= not(inputs(176)) or (inputs(251));
    layer0_outputs(1880) <= not(inputs(105));
    layer0_outputs(1881) <= (inputs(28)) and (inputs(217));
    layer0_outputs(1882) <= (inputs(196)) and not (inputs(76));
    layer0_outputs(1883) <= inputs(91);
    layer0_outputs(1884) <= (inputs(71)) xor (inputs(116));
    layer0_outputs(1885) <= not((inputs(143)) xor (inputs(25)));
    layer0_outputs(1886) <= (inputs(64)) and (inputs(73));
    layer0_outputs(1887) <= not((inputs(71)) or (inputs(165)));
    layer0_outputs(1888) <= (inputs(119)) and not (inputs(220));
    layer0_outputs(1889) <= not(inputs(37));
    layer0_outputs(1890) <= not(inputs(112));
    layer0_outputs(1891) <= (inputs(212)) and not (inputs(41));
    layer0_outputs(1892) <= inputs(131);
    layer0_outputs(1893) <= not(inputs(192));
    layer0_outputs(1894) <= not((inputs(104)) or (inputs(132)));
    layer0_outputs(1895) <= not(inputs(170));
    layer0_outputs(1896) <= not(inputs(131));
    layer0_outputs(1897) <= inputs(59);
    layer0_outputs(1898) <= not(inputs(44));
    layer0_outputs(1899) <= (inputs(231)) and not (inputs(223));
    layer0_outputs(1900) <= inputs(249);
    layer0_outputs(1901) <= inputs(210);
    layer0_outputs(1902) <= not(inputs(181));
    layer0_outputs(1903) <= not((inputs(152)) or (inputs(234)));
    layer0_outputs(1904) <= inputs(50);
    layer0_outputs(1905) <= inputs(135);
    layer0_outputs(1906) <= not(inputs(114));
    layer0_outputs(1907) <= inputs(59);
    layer0_outputs(1908) <= not(inputs(213)) or (inputs(128));
    layer0_outputs(1909) <= (inputs(199)) xor (inputs(49));
    layer0_outputs(1910) <= (inputs(121)) xor (inputs(165));
    layer0_outputs(1911) <= (inputs(152)) and not (inputs(249));
    layer0_outputs(1912) <= not((inputs(107)) or (inputs(88)));
    layer0_outputs(1913) <= not((inputs(244)) or (inputs(157)));
    layer0_outputs(1914) <= inputs(228);
    layer0_outputs(1915) <= (inputs(215)) xor (inputs(173));
    layer0_outputs(1916) <= not(inputs(73)) or (inputs(4));
    layer0_outputs(1917) <= not(inputs(189));
    layer0_outputs(1918) <= inputs(129);
    layer0_outputs(1919) <= not(inputs(231)) or (inputs(143));
    layer0_outputs(1920) <= not(inputs(112)) or (inputs(177));
    layer0_outputs(1921) <= inputs(228);
    layer0_outputs(1922) <= (inputs(1)) and not (inputs(248));
    layer0_outputs(1923) <= not((inputs(197)) or (inputs(131)));
    layer0_outputs(1924) <= not((inputs(233)) and (inputs(168)));
    layer0_outputs(1925) <= not(inputs(202));
    layer0_outputs(1926) <= (inputs(18)) and not (inputs(223));
    layer0_outputs(1927) <= (inputs(254)) or (inputs(1));
    layer0_outputs(1928) <= not(inputs(228));
    layer0_outputs(1929) <= inputs(194);
    layer0_outputs(1930) <= inputs(25);
    layer0_outputs(1931) <= '0';
    layer0_outputs(1932) <= not((inputs(33)) or (inputs(19)));
    layer0_outputs(1933) <= (inputs(163)) and not (inputs(62));
    layer0_outputs(1934) <= (inputs(158)) or (inputs(159));
    layer0_outputs(1935) <= inputs(139);
    layer0_outputs(1936) <= inputs(45);
    layer0_outputs(1937) <= not(inputs(165));
    layer0_outputs(1938) <= not(inputs(92));
    layer0_outputs(1939) <= (inputs(209)) and not (inputs(112));
    layer0_outputs(1940) <= (inputs(118)) or (inputs(202));
    layer0_outputs(1941) <= (inputs(8)) and not (inputs(110));
    layer0_outputs(1942) <= not(inputs(67));
    layer0_outputs(1943) <= not(inputs(147));
    layer0_outputs(1944) <= not((inputs(68)) xor (inputs(149)));
    layer0_outputs(1945) <= (inputs(52)) xor (inputs(132));
    layer0_outputs(1946) <= not(inputs(75));
    layer0_outputs(1947) <= not(inputs(212));
    layer0_outputs(1948) <= not((inputs(171)) or (inputs(168)));
    layer0_outputs(1949) <= not((inputs(237)) or (inputs(139)));
    layer0_outputs(1950) <= not((inputs(11)) xor (inputs(91)));
    layer0_outputs(1951) <= (inputs(196)) or (inputs(53));
    layer0_outputs(1952) <= not((inputs(240)) or (inputs(7)));
    layer0_outputs(1953) <= not(inputs(20));
    layer0_outputs(1954) <= not(inputs(233));
    layer0_outputs(1955) <= not((inputs(247)) or (inputs(249)));
    layer0_outputs(1956) <= not((inputs(194)) xor (inputs(201)));
    layer0_outputs(1957) <= not(inputs(85)) or (inputs(240));
    layer0_outputs(1958) <= (inputs(52)) and not (inputs(130));
    layer0_outputs(1959) <= not((inputs(115)) or (inputs(131)));
    layer0_outputs(1960) <= not(inputs(110));
    layer0_outputs(1961) <= not(inputs(168)) or (inputs(1));
    layer0_outputs(1962) <= inputs(83);
    layer0_outputs(1963) <= inputs(235);
    layer0_outputs(1964) <= (inputs(195)) or (inputs(115));
    layer0_outputs(1965) <= not(inputs(29));
    layer0_outputs(1966) <= '0';
    layer0_outputs(1967) <= inputs(53);
    layer0_outputs(1968) <= (inputs(84)) and not (inputs(30));
    layer0_outputs(1969) <= (inputs(93)) and not (inputs(207));
    layer0_outputs(1970) <= not((inputs(225)) or (inputs(68)));
    layer0_outputs(1971) <= not(inputs(151));
    layer0_outputs(1972) <= not(inputs(188)) or (inputs(67));
    layer0_outputs(1973) <= inputs(104);
    layer0_outputs(1974) <= inputs(146);
    layer0_outputs(1975) <= not((inputs(155)) or (inputs(35)));
    layer0_outputs(1976) <= inputs(9);
    layer0_outputs(1977) <= (inputs(189)) or (inputs(96));
    layer0_outputs(1978) <= not(inputs(89));
    layer0_outputs(1979) <= not(inputs(3));
    layer0_outputs(1980) <= (inputs(0)) or (inputs(94));
    layer0_outputs(1981) <= '1';
    layer0_outputs(1982) <= (inputs(33)) or (inputs(162));
    layer0_outputs(1983) <= (inputs(189)) xor (inputs(67));
    layer0_outputs(1984) <= not((inputs(70)) xor (inputs(89)));
    layer0_outputs(1985) <= not(inputs(99));
    layer0_outputs(1986) <= (inputs(190)) or (inputs(212));
    layer0_outputs(1987) <= inputs(247);
    layer0_outputs(1988) <= (inputs(204)) or (inputs(162));
    layer0_outputs(1989) <= not(inputs(64));
    layer0_outputs(1990) <= inputs(215);
    layer0_outputs(1991) <= not(inputs(180));
    layer0_outputs(1992) <= not(inputs(146));
    layer0_outputs(1993) <= inputs(179);
    layer0_outputs(1994) <= not(inputs(123)) or (inputs(193));
    layer0_outputs(1995) <= inputs(229);
    layer0_outputs(1996) <= inputs(169);
    layer0_outputs(1997) <= (inputs(130)) xor (inputs(86));
    layer0_outputs(1998) <= (inputs(10)) and not (inputs(15));
    layer0_outputs(1999) <= (inputs(5)) or (inputs(208));
    layer0_outputs(2000) <= not((inputs(206)) or (inputs(236)));
    layer0_outputs(2001) <= inputs(157);
    layer0_outputs(2002) <= inputs(155);
    layer0_outputs(2003) <= not(inputs(9)) or (inputs(51));
    layer0_outputs(2004) <= not((inputs(193)) and (inputs(133)));
    layer0_outputs(2005) <= (inputs(194)) and not (inputs(155));
    layer0_outputs(2006) <= not(inputs(86));
    layer0_outputs(2007) <= (inputs(166)) xor (inputs(136));
    layer0_outputs(2008) <= not(inputs(166));
    layer0_outputs(2009) <= not((inputs(32)) or (inputs(31)));
    layer0_outputs(2010) <= not(inputs(57));
    layer0_outputs(2011) <= not(inputs(68)) or (inputs(242));
    layer0_outputs(2012) <= not(inputs(121));
    layer0_outputs(2013) <= (inputs(190)) and not (inputs(223));
    layer0_outputs(2014) <= (inputs(225)) and not (inputs(234));
    layer0_outputs(2015) <= not((inputs(238)) or (inputs(199)));
    layer0_outputs(2016) <= not(inputs(166));
    layer0_outputs(2017) <= inputs(152);
    layer0_outputs(2018) <= (inputs(128)) or (inputs(165));
    layer0_outputs(2019) <= (inputs(199)) and not (inputs(161));
    layer0_outputs(2020) <= not(inputs(28)) or (inputs(87));
    layer0_outputs(2021) <= (inputs(223)) and (inputs(94));
    layer0_outputs(2022) <= not(inputs(131));
    layer0_outputs(2023) <= (inputs(105)) or (inputs(106));
    layer0_outputs(2024) <= (inputs(105)) xor (inputs(137));
    layer0_outputs(2025) <= not((inputs(113)) or (inputs(233)));
    layer0_outputs(2026) <= inputs(36);
    layer0_outputs(2027) <= (inputs(18)) xor (inputs(246));
    layer0_outputs(2028) <= inputs(245);
    layer0_outputs(2029) <= not((inputs(72)) or (inputs(171)));
    layer0_outputs(2030) <= not(inputs(136)) or (inputs(159));
    layer0_outputs(2031) <= not((inputs(221)) xor (inputs(54)));
    layer0_outputs(2032) <= not((inputs(47)) or (inputs(136)));
    layer0_outputs(2033) <= (inputs(135)) or (inputs(176));
    layer0_outputs(2034) <= not(inputs(230));
    layer0_outputs(2035) <= (inputs(74)) and not (inputs(233));
    layer0_outputs(2036) <= not(inputs(247));
    layer0_outputs(2037) <= (inputs(19)) and not (inputs(110));
    layer0_outputs(2038) <= (inputs(123)) and not (inputs(132));
    layer0_outputs(2039) <= (inputs(56)) or (inputs(113));
    layer0_outputs(2040) <= not(inputs(230));
    layer0_outputs(2041) <= not(inputs(25));
    layer0_outputs(2042) <= not(inputs(167)) or (inputs(1));
    layer0_outputs(2043) <= (inputs(129)) or (inputs(147));
    layer0_outputs(2044) <= not((inputs(159)) or (inputs(17)));
    layer0_outputs(2045) <= (inputs(140)) or (inputs(96));
    layer0_outputs(2046) <= (inputs(9)) and not (inputs(14));
    layer0_outputs(2047) <= not(inputs(176));
    layer0_outputs(2048) <= inputs(135);
    layer0_outputs(2049) <= (inputs(233)) and not (inputs(15));
    layer0_outputs(2050) <= inputs(123);
    layer0_outputs(2051) <= not(inputs(214)) or (inputs(190));
    layer0_outputs(2052) <= not(inputs(231));
    layer0_outputs(2053) <= inputs(161);
    layer0_outputs(2054) <= '0';
    layer0_outputs(2055) <= inputs(113);
    layer0_outputs(2056) <= not((inputs(73)) xor (inputs(119)));
    layer0_outputs(2057) <= (inputs(227)) xor (inputs(16));
    layer0_outputs(2058) <= not(inputs(179));
    layer0_outputs(2059) <= (inputs(23)) and not (inputs(112));
    layer0_outputs(2060) <= not(inputs(194)) or (inputs(49));
    layer0_outputs(2061) <= (inputs(162)) or (inputs(200));
    layer0_outputs(2062) <= not((inputs(142)) or (inputs(4)));
    layer0_outputs(2063) <= inputs(84);
    layer0_outputs(2064) <= not(inputs(215)) or (inputs(30));
    layer0_outputs(2065) <= not((inputs(178)) xor (inputs(82)));
    layer0_outputs(2066) <= not((inputs(179)) or (inputs(84)));
    layer0_outputs(2067) <= (inputs(125)) or (inputs(36));
    layer0_outputs(2068) <= (inputs(64)) or (inputs(63));
    layer0_outputs(2069) <= (inputs(54)) and not (inputs(234));
    layer0_outputs(2070) <= inputs(178);
    layer0_outputs(2071) <= not(inputs(187)) or (inputs(86));
    layer0_outputs(2072) <= inputs(152);
    layer0_outputs(2073) <= not(inputs(218));
    layer0_outputs(2074) <= (inputs(245)) xor (inputs(191));
    layer0_outputs(2075) <= (inputs(18)) and not (inputs(131));
    layer0_outputs(2076) <= (inputs(218)) or (inputs(172));
    layer0_outputs(2077) <= (inputs(247)) and not (inputs(95));
    layer0_outputs(2078) <= not(inputs(98));
    layer0_outputs(2079) <= not(inputs(173));
    layer0_outputs(2080) <= not(inputs(138)) or (inputs(230));
    layer0_outputs(2081) <= (inputs(178)) or (inputs(191));
    layer0_outputs(2082) <= (inputs(11)) and not (inputs(224));
    layer0_outputs(2083) <= (inputs(26)) and not (inputs(218));
    layer0_outputs(2084) <= inputs(103);
    layer0_outputs(2085) <= (inputs(152)) xor (inputs(145));
    layer0_outputs(2086) <= (inputs(173)) or (inputs(209));
    layer0_outputs(2087) <= not((inputs(114)) or (inputs(249)));
    layer0_outputs(2088) <= not(inputs(85));
    layer0_outputs(2089) <= not(inputs(202)) or (inputs(110));
    layer0_outputs(2090) <= (inputs(131)) and not (inputs(34));
    layer0_outputs(2091) <= not(inputs(25));
    layer0_outputs(2092) <= (inputs(51)) or (inputs(188));
    layer0_outputs(2093) <= not(inputs(197)) or (inputs(144));
    layer0_outputs(2094) <= not((inputs(64)) or (inputs(206)));
    layer0_outputs(2095) <= inputs(21);
    layer0_outputs(2096) <= inputs(85);
    layer0_outputs(2097) <= not((inputs(194)) or (inputs(75)));
    layer0_outputs(2098) <= not(inputs(253));
    layer0_outputs(2099) <= inputs(56);
    layer0_outputs(2100) <= (inputs(124)) or (inputs(160));
    layer0_outputs(2101) <= not(inputs(185)) or (inputs(25));
    layer0_outputs(2102) <= (inputs(14)) xor (inputs(243));
    layer0_outputs(2103) <= not((inputs(204)) xor (inputs(147)));
    layer0_outputs(2104) <= (inputs(54)) or (inputs(255));
    layer0_outputs(2105) <= inputs(194);
    layer0_outputs(2106) <= not(inputs(18));
    layer0_outputs(2107) <= not(inputs(100));
    layer0_outputs(2108) <= inputs(75);
    layer0_outputs(2109) <= not(inputs(99));
    layer0_outputs(2110) <= inputs(201);
    layer0_outputs(2111) <= (inputs(130)) or (inputs(152));
    layer0_outputs(2112) <= (inputs(41)) or (inputs(210));
    layer0_outputs(2113) <= not((inputs(53)) xor (inputs(115)));
    layer0_outputs(2114) <= (inputs(246)) or (inputs(187));
    layer0_outputs(2115) <= not(inputs(57));
    layer0_outputs(2116) <= (inputs(171)) or (inputs(6));
    layer0_outputs(2117) <= not(inputs(58));
    layer0_outputs(2118) <= inputs(205);
    layer0_outputs(2119) <= not(inputs(209));
    layer0_outputs(2120) <= not((inputs(210)) or (inputs(181)));
    layer0_outputs(2121) <= not((inputs(78)) or (inputs(38)));
    layer0_outputs(2122) <= not(inputs(231));
    layer0_outputs(2123) <= (inputs(6)) or (inputs(239));
    layer0_outputs(2124) <= (inputs(161)) or (inputs(33));
    layer0_outputs(2125) <= not((inputs(244)) or (inputs(129)));
    layer0_outputs(2126) <= (inputs(234)) or (inputs(130));
    layer0_outputs(2127) <= (inputs(227)) or (inputs(173));
    layer0_outputs(2128) <= (inputs(217)) or (inputs(159));
    layer0_outputs(2129) <= not((inputs(49)) or (inputs(173)));
    layer0_outputs(2130) <= inputs(60);
    layer0_outputs(2131) <= (inputs(69)) and not (inputs(205));
    layer0_outputs(2132) <= not((inputs(146)) or (inputs(225)));
    layer0_outputs(2133) <= not(inputs(19));
    layer0_outputs(2134) <= inputs(79);
    layer0_outputs(2135) <= (inputs(244)) and not (inputs(254));
    layer0_outputs(2136) <= not((inputs(62)) xor (inputs(227)));
    layer0_outputs(2137) <= (inputs(67)) or (inputs(101));
    layer0_outputs(2138) <= not((inputs(127)) or (inputs(155)));
    layer0_outputs(2139) <= not(inputs(218));
    layer0_outputs(2140) <= (inputs(40)) and not (inputs(129));
    layer0_outputs(2141) <= (inputs(227)) xor (inputs(14));
    layer0_outputs(2142) <= inputs(75);
    layer0_outputs(2143) <= not(inputs(26)) or (inputs(250));
    layer0_outputs(2144) <= not((inputs(43)) or (inputs(138)));
    layer0_outputs(2145) <= (inputs(85)) and not (inputs(223));
    layer0_outputs(2146) <= (inputs(227)) and not (inputs(137));
    layer0_outputs(2147) <= not(inputs(90));
    layer0_outputs(2148) <= not(inputs(4));
    layer0_outputs(2149) <= not(inputs(22));
    layer0_outputs(2150) <= (inputs(15)) and not (inputs(76));
    layer0_outputs(2151) <= not((inputs(16)) or (inputs(124)));
    layer0_outputs(2152) <= (inputs(79)) or (inputs(189));
    layer0_outputs(2153) <= (inputs(254)) or (inputs(68));
    layer0_outputs(2154) <= not(inputs(195));
    layer0_outputs(2155) <= '1';
    layer0_outputs(2156) <= (inputs(193)) or (inputs(205));
    layer0_outputs(2157) <= inputs(227);
    layer0_outputs(2158) <= (inputs(25)) and not (inputs(226));
    layer0_outputs(2159) <= (inputs(106)) and not (inputs(20));
    layer0_outputs(2160) <= inputs(51);
    layer0_outputs(2161) <= inputs(76);
    layer0_outputs(2162) <= not(inputs(168));
    layer0_outputs(2163) <= not(inputs(38));
    layer0_outputs(2164) <= (inputs(154)) or (inputs(57));
    layer0_outputs(2165) <= inputs(229);
    layer0_outputs(2166) <= inputs(137);
    layer0_outputs(2167) <= not(inputs(41)) or (inputs(117));
    layer0_outputs(2168) <= (inputs(94)) and not (inputs(158));
    layer0_outputs(2169) <= not(inputs(118)) or (inputs(18));
    layer0_outputs(2170) <= (inputs(137)) xor (inputs(29));
    layer0_outputs(2171) <= '1';
    layer0_outputs(2172) <= (inputs(60)) or (inputs(46));
    layer0_outputs(2173) <= not(inputs(208)) or (inputs(32));
    layer0_outputs(2174) <= (inputs(103)) and (inputs(167));
    layer0_outputs(2175) <= (inputs(59)) or (inputs(60));
    layer0_outputs(2176) <= (inputs(48)) or (inputs(179));
    layer0_outputs(2177) <= (inputs(87)) or (inputs(100));
    layer0_outputs(2178) <= (inputs(53)) and (inputs(78));
    layer0_outputs(2179) <= not((inputs(2)) or (inputs(121)));
    layer0_outputs(2180) <= (inputs(102)) xor (inputs(217));
    layer0_outputs(2181) <= not(inputs(111));
    layer0_outputs(2182) <= not((inputs(253)) or (inputs(187)));
    layer0_outputs(2183) <= not(inputs(123)) or (inputs(227));
    layer0_outputs(2184) <= not(inputs(116));
    layer0_outputs(2185) <= inputs(165);
    layer0_outputs(2186) <= not(inputs(74));
    layer0_outputs(2187) <= not((inputs(183)) or (inputs(252)));
    layer0_outputs(2188) <= inputs(138);
    layer0_outputs(2189) <= not(inputs(197)) or (inputs(29));
    layer0_outputs(2190) <= not(inputs(221)) or (inputs(177));
    layer0_outputs(2191) <= (inputs(64)) xor (inputs(88));
    layer0_outputs(2192) <= inputs(233);
    layer0_outputs(2193) <= not(inputs(27)) or (inputs(130));
    layer0_outputs(2194) <= not(inputs(21));
    layer0_outputs(2195) <= not(inputs(148));
    layer0_outputs(2196) <= not((inputs(114)) or (inputs(119)));
    layer0_outputs(2197) <= not((inputs(174)) or (inputs(243)));
    layer0_outputs(2198) <= not((inputs(137)) or (inputs(34)));
    layer0_outputs(2199) <= not((inputs(221)) xor (inputs(83)));
    layer0_outputs(2200) <= inputs(103);
    layer0_outputs(2201) <= inputs(93);
    layer0_outputs(2202) <= not((inputs(50)) or (inputs(214)));
    layer0_outputs(2203) <= (inputs(75)) and not (inputs(3));
    layer0_outputs(2204) <= (inputs(210)) or (inputs(156));
    layer0_outputs(2205) <= not(inputs(6)) or (inputs(83));
    layer0_outputs(2206) <= (inputs(219)) and not (inputs(22));
    layer0_outputs(2207) <= not(inputs(228));
    layer0_outputs(2208) <= (inputs(240)) xor (inputs(13));
    layer0_outputs(2209) <= not(inputs(224)) or (inputs(82));
    layer0_outputs(2210) <= not(inputs(105));
    layer0_outputs(2211) <= not(inputs(119));
    layer0_outputs(2212) <= inputs(35);
    layer0_outputs(2213) <= inputs(38);
    layer0_outputs(2214) <= not((inputs(124)) and (inputs(252)));
    layer0_outputs(2215) <= not(inputs(151)) or (inputs(224));
    layer0_outputs(2216) <= not(inputs(69));
    layer0_outputs(2217) <= not(inputs(252));
    layer0_outputs(2218) <= not(inputs(22));
    layer0_outputs(2219) <= (inputs(185)) and not (inputs(118));
    layer0_outputs(2220) <= (inputs(247)) and (inputs(234));
    layer0_outputs(2221) <= not((inputs(68)) xor (inputs(112)));
    layer0_outputs(2222) <= not(inputs(56)) or (inputs(224));
    layer0_outputs(2223) <= not((inputs(6)) and (inputs(23)));
    layer0_outputs(2224) <= (inputs(12)) xor (inputs(160));
    layer0_outputs(2225) <= inputs(7);
    layer0_outputs(2226) <= not((inputs(213)) and (inputs(41)));
    layer0_outputs(2227) <= (inputs(82)) xor (inputs(26));
    layer0_outputs(2228) <= (inputs(231)) and not (inputs(78));
    layer0_outputs(2229) <= not(inputs(103)) or (inputs(2));
    layer0_outputs(2230) <= not((inputs(133)) or (inputs(54)));
    layer0_outputs(2231) <= not((inputs(44)) or (inputs(112)));
    layer0_outputs(2232) <= not(inputs(176)) or (inputs(48));
    layer0_outputs(2233) <= not((inputs(182)) xor (inputs(161)));
    layer0_outputs(2234) <= (inputs(2)) or (inputs(148));
    layer0_outputs(2235) <= not(inputs(121)) or (inputs(253));
    layer0_outputs(2236) <= (inputs(245)) and not (inputs(52));
    layer0_outputs(2237) <= (inputs(194)) or (inputs(53));
    layer0_outputs(2238) <= (inputs(53)) and not (inputs(172));
    layer0_outputs(2239) <= not((inputs(38)) or (inputs(193)));
    layer0_outputs(2240) <= (inputs(152)) or (inputs(152));
    layer0_outputs(2241) <= not(inputs(38));
    layer0_outputs(2242) <= (inputs(0)) xor (inputs(195));
    layer0_outputs(2243) <= not(inputs(252));
    layer0_outputs(2244) <= (inputs(254)) or (inputs(44));
    layer0_outputs(2245) <= not((inputs(161)) or (inputs(132)));
    layer0_outputs(2246) <= inputs(162);
    layer0_outputs(2247) <= not(inputs(188));
    layer0_outputs(2248) <= not(inputs(235));
    layer0_outputs(2249) <= not((inputs(253)) xor (inputs(90)));
    layer0_outputs(2250) <= (inputs(50)) or (inputs(103));
    layer0_outputs(2251) <= not(inputs(77));
    layer0_outputs(2252) <= not((inputs(22)) xor (inputs(40)));
    layer0_outputs(2253) <= (inputs(198)) and not (inputs(45));
    layer0_outputs(2254) <= inputs(158);
    layer0_outputs(2255) <= inputs(150);
    layer0_outputs(2256) <= '0';
    layer0_outputs(2257) <= inputs(237);
    layer0_outputs(2258) <= (inputs(247)) and not (inputs(246));
    layer0_outputs(2259) <= inputs(179);
    layer0_outputs(2260) <= inputs(188);
    layer0_outputs(2261) <= (inputs(79)) or (inputs(122));
    layer0_outputs(2262) <= (inputs(80)) or (inputs(208));
    layer0_outputs(2263) <= not(inputs(225));
    layer0_outputs(2264) <= not((inputs(134)) and (inputs(226)));
    layer0_outputs(2265) <= not(inputs(147));
    layer0_outputs(2266) <= '0';
    layer0_outputs(2267) <= (inputs(222)) xor (inputs(55));
    layer0_outputs(2268) <= (inputs(63)) xor (inputs(39));
    layer0_outputs(2269) <= inputs(110);
    layer0_outputs(2270) <= (inputs(82)) and not (inputs(126));
    layer0_outputs(2271) <= inputs(115);
    layer0_outputs(2272) <= not((inputs(23)) or (inputs(75)));
    layer0_outputs(2273) <= not(inputs(184)) or (inputs(237));
    layer0_outputs(2274) <= not(inputs(107)) or (inputs(50));
    layer0_outputs(2275) <= not(inputs(106)) or (inputs(196));
    layer0_outputs(2276) <= not((inputs(97)) xor (inputs(85)));
    layer0_outputs(2277) <= (inputs(18)) or (inputs(139));
    layer0_outputs(2278) <= not(inputs(104)) or (inputs(35));
    layer0_outputs(2279) <= not(inputs(88)) or (inputs(15));
    layer0_outputs(2280) <= inputs(211);
    layer0_outputs(2281) <= not((inputs(208)) or (inputs(73)));
    layer0_outputs(2282) <= not(inputs(102));
    layer0_outputs(2283) <= inputs(8);
    layer0_outputs(2284) <= (inputs(120)) and not (inputs(5));
    layer0_outputs(2285) <= (inputs(4)) or (inputs(215));
    layer0_outputs(2286) <= not(inputs(193));
    layer0_outputs(2287) <= not(inputs(38)) or (inputs(215));
    layer0_outputs(2288) <= inputs(148);
    layer0_outputs(2289) <= not((inputs(201)) or (inputs(236)));
    layer0_outputs(2290) <= not(inputs(99)) or (inputs(226));
    layer0_outputs(2291) <= not(inputs(149)) or (inputs(221));
    layer0_outputs(2292) <= not((inputs(62)) or (inputs(61)));
    layer0_outputs(2293) <= inputs(207);
    layer0_outputs(2294) <= not(inputs(115));
    layer0_outputs(2295) <= not((inputs(166)) or (inputs(12)));
    layer0_outputs(2296) <= inputs(147);
    layer0_outputs(2297) <= (inputs(133)) and not (inputs(20));
    layer0_outputs(2298) <= not((inputs(136)) xor (inputs(246)));
    layer0_outputs(2299) <= not(inputs(197)) or (inputs(216));
    layer0_outputs(2300) <= (inputs(98)) and not (inputs(15));
    layer0_outputs(2301) <= (inputs(221)) or (inputs(177));
    layer0_outputs(2302) <= (inputs(95)) or (inputs(163));
    layer0_outputs(2303) <= inputs(154);
    layer0_outputs(2304) <= (inputs(141)) or (inputs(193));
    layer0_outputs(2305) <= not(inputs(36));
    layer0_outputs(2306) <= not(inputs(250));
    layer0_outputs(2307) <= not(inputs(120));
    layer0_outputs(2308) <= (inputs(146)) and not (inputs(0));
    layer0_outputs(2309) <= (inputs(134)) xor (inputs(120));
    layer0_outputs(2310) <= not(inputs(110));
    layer0_outputs(2311) <= (inputs(138)) or (inputs(184));
    layer0_outputs(2312) <= not(inputs(167)) or (inputs(253));
    layer0_outputs(2313) <= not((inputs(46)) xor (inputs(222)));
    layer0_outputs(2314) <= not(inputs(245));
    layer0_outputs(2315) <= not((inputs(40)) or (inputs(49)));
    layer0_outputs(2316) <= not(inputs(29));
    layer0_outputs(2317) <= not((inputs(71)) or (inputs(102)));
    layer0_outputs(2318) <= not((inputs(56)) or (inputs(162)));
    layer0_outputs(2319) <= not(inputs(181)) or (inputs(58));
    layer0_outputs(2320) <= (inputs(21)) and not (inputs(224));
    layer0_outputs(2321) <= (inputs(112)) or (inputs(154));
    layer0_outputs(2322) <= not((inputs(70)) or (inputs(14)));
    layer0_outputs(2323) <= inputs(13);
    layer0_outputs(2324) <= (inputs(155)) or (inputs(116));
    layer0_outputs(2325) <= (inputs(100)) and not (inputs(120));
    layer0_outputs(2326) <= not((inputs(195)) xor (inputs(212)));
    layer0_outputs(2327) <= not((inputs(117)) or (inputs(243)));
    layer0_outputs(2328) <= not(inputs(142));
    layer0_outputs(2329) <= (inputs(143)) and not (inputs(253));
    layer0_outputs(2330) <= (inputs(79)) xor (inputs(173));
    layer0_outputs(2331) <= (inputs(129)) or (inputs(132));
    layer0_outputs(2332) <= (inputs(157)) or (inputs(191));
    layer0_outputs(2333) <= not(inputs(57)) or (inputs(15));
    layer0_outputs(2334) <= not(inputs(38));
    layer0_outputs(2335) <= (inputs(66)) or (inputs(123));
    layer0_outputs(2336) <= not(inputs(32));
    layer0_outputs(2337) <= not((inputs(193)) or (inputs(180)));
    layer0_outputs(2338) <= inputs(210);
    layer0_outputs(2339) <= inputs(73);
    layer0_outputs(2340) <= not(inputs(51));
    layer0_outputs(2341) <= (inputs(164)) or (inputs(74));
    layer0_outputs(2342) <= inputs(190);
    layer0_outputs(2343) <= not((inputs(64)) xor (inputs(74)));
    layer0_outputs(2344) <= not(inputs(49)) or (inputs(154));
    layer0_outputs(2345) <= not((inputs(206)) xor (inputs(112)));
    layer0_outputs(2346) <= inputs(223);
    layer0_outputs(2347) <= inputs(91);
    layer0_outputs(2348) <= (inputs(53)) or (inputs(66));
    layer0_outputs(2349) <= not(inputs(91));
    layer0_outputs(2350) <= not(inputs(60));
    layer0_outputs(2351) <= not(inputs(169));
    layer0_outputs(2352) <= not(inputs(26)) or (inputs(177));
    layer0_outputs(2353) <= not(inputs(124)) or (inputs(78));
    layer0_outputs(2354) <= (inputs(91)) and not (inputs(50));
    layer0_outputs(2355) <= inputs(247);
    layer0_outputs(2356) <= not((inputs(54)) or (inputs(14)));
    layer0_outputs(2357) <= not((inputs(141)) or (inputs(249)));
    layer0_outputs(2358) <= (inputs(250)) xor (inputs(244));
    layer0_outputs(2359) <= (inputs(237)) and (inputs(112));
    layer0_outputs(2360) <= (inputs(58)) and not (inputs(239));
    layer0_outputs(2361) <= not((inputs(52)) or (inputs(97)));
    layer0_outputs(2362) <= not(inputs(211));
    layer0_outputs(2363) <= inputs(180);
    layer0_outputs(2364) <= (inputs(247)) or (inputs(145));
    layer0_outputs(2365) <= (inputs(168)) xor (inputs(61));
    layer0_outputs(2366) <= not((inputs(220)) or (inputs(186)));
    layer0_outputs(2367) <= not(inputs(213));
    layer0_outputs(2368) <= (inputs(199)) and (inputs(39));
    layer0_outputs(2369) <= not((inputs(234)) or (inputs(163)));
    layer0_outputs(2370) <= not((inputs(199)) or (inputs(74)));
    layer0_outputs(2371) <= (inputs(224)) or (inputs(192));
    layer0_outputs(2372) <= not((inputs(206)) xor (inputs(255)));
    layer0_outputs(2373) <= not(inputs(157));
    layer0_outputs(2374) <= (inputs(29)) and not (inputs(15));
    layer0_outputs(2375) <= not(inputs(25));
    layer0_outputs(2376) <= (inputs(45)) or (inputs(179));
    layer0_outputs(2377) <= inputs(238);
    layer0_outputs(2378) <= (inputs(249)) or (inputs(128));
    layer0_outputs(2379) <= inputs(84);
    layer0_outputs(2380) <= not(inputs(187));
    layer0_outputs(2381) <= inputs(147);
    layer0_outputs(2382) <= (inputs(65)) or (inputs(226));
    layer0_outputs(2383) <= not(inputs(73)) or (inputs(151));
    layer0_outputs(2384) <= not(inputs(202)) or (inputs(141));
    layer0_outputs(2385) <= not((inputs(22)) or (inputs(17)));
    layer0_outputs(2386) <= inputs(153);
    layer0_outputs(2387) <= not(inputs(150)) or (inputs(67));
    layer0_outputs(2388) <= not(inputs(229));
    layer0_outputs(2389) <= not(inputs(77));
    layer0_outputs(2390) <= (inputs(171)) xor (inputs(220));
    layer0_outputs(2391) <= (inputs(24)) and not (inputs(253));
    layer0_outputs(2392) <= inputs(235);
    layer0_outputs(2393) <= not(inputs(194));
    layer0_outputs(2394) <= inputs(163);
    layer0_outputs(2395) <= '0';
    layer0_outputs(2396) <= not((inputs(202)) or (inputs(227)));
    layer0_outputs(2397) <= not(inputs(178));
    layer0_outputs(2398) <= not(inputs(122)) or (inputs(19));
    layer0_outputs(2399) <= (inputs(243)) xor (inputs(62));
    layer0_outputs(2400) <= (inputs(67)) or (inputs(14));
    layer0_outputs(2401) <= not((inputs(192)) or (inputs(101)));
    layer0_outputs(2402) <= (inputs(129)) or (inputs(222));
    layer0_outputs(2403) <= '1';
    layer0_outputs(2404) <= not(inputs(153));
    layer0_outputs(2405) <= not((inputs(93)) xor (inputs(60)));
    layer0_outputs(2406) <= inputs(5);
    layer0_outputs(2407) <= not((inputs(55)) xor (inputs(253)));
    layer0_outputs(2408) <= '0';
    layer0_outputs(2409) <= '1';
    layer0_outputs(2410) <= inputs(229);
    layer0_outputs(2411) <= (inputs(116)) xor (inputs(175));
    layer0_outputs(2412) <= inputs(140);
    layer0_outputs(2413) <= (inputs(5)) or (inputs(60));
    layer0_outputs(2414) <= (inputs(241)) or (inputs(198));
    layer0_outputs(2415) <= not((inputs(80)) or (inputs(98)));
    layer0_outputs(2416) <= (inputs(89)) and (inputs(40));
    layer0_outputs(2417) <= inputs(202);
    layer0_outputs(2418) <= (inputs(126)) or (inputs(31));
    layer0_outputs(2419) <= inputs(33);
    layer0_outputs(2420) <= not(inputs(10)) or (inputs(253));
    layer0_outputs(2421) <= inputs(132);
    layer0_outputs(2422) <= (inputs(179)) or (inputs(147));
    layer0_outputs(2423) <= not(inputs(202)) or (inputs(103));
    layer0_outputs(2424) <= not((inputs(141)) or (inputs(188)));
    layer0_outputs(2425) <= not(inputs(106)) or (inputs(246));
    layer0_outputs(2426) <= (inputs(217)) or (inputs(201));
    layer0_outputs(2427) <= inputs(197);
    layer0_outputs(2428) <= not(inputs(213));
    layer0_outputs(2429) <= inputs(205);
    layer0_outputs(2430) <= (inputs(154)) or (inputs(0));
    layer0_outputs(2431) <= not(inputs(231));
    layer0_outputs(2432) <= not(inputs(101));
    layer0_outputs(2433) <= inputs(127);
    layer0_outputs(2434) <= inputs(104);
    layer0_outputs(2435) <= not(inputs(57)) or (inputs(146));
    layer0_outputs(2436) <= not(inputs(84)) or (inputs(55));
    layer0_outputs(2437) <= (inputs(199)) and not (inputs(117));
    layer0_outputs(2438) <= inputs(168);
    layer0_outputs(2439) <= (inputs(3)) or (inputs(43));
    layer0_outputs(2440) <= inputs(104);
    layer0_outputs(2441) <= (inputs(244)) or (inputs(229));
    layer0_outputs(2442) <= not(inputs(102));
    layer0_outputs(2443) <= not(inputs(161));
    layer0_outputs(2444) <= not(inputs(133));
    layer0_outputs(2445) <= not((inputs(9)) or (inputs(25)));
    layer0_outputs(2446) <= (inputs(146)) or (inputs(63));
    layer0_outputs(2447) <= not((inputs(3)) or (inputs(169)));
    layer0_outputs(2448) <= (inputs(206)) and not (inputs(109));
    layer0_outputs(2449) <= not(inputs(16)) or (inputs(255));
    layer0_outputs(2450) <= inputs(29);
    layer0_outputs(2451) <= (inputs(215)) or (inputs(200));
    layer0_outputs(2452) <= not(inputs(191)) or (inputs(162));
    layer0_outputs(2453) <= (inputs(87)) and not (inputs(98));
    layer0_outputs(2454) <= (inputs(2)) and not (inputs(15));
    layer0_outputs(2455) <= (inputs(125)) and not (inputs(21));
    layer0_outputs(2456) <= not((inputs(45)) and (inputs(95)));
    layer0_outputs(2457) <= (inputs(164)) or (inputs(101));
    layer0_outputs(2458) <= (inputs(105)) xor (inputs(173));
    layer0_outputs(2459) <= not((inputs(62)) or (inputs(92)));
    layer0_outputs(2460) <= (inputs(124)) and not (inputs(255));
    layer0_outputs(2461) <= not(inputs(197));
    layer0_outputs(2462) <= not((inputs(5)) xor (inputs(127)));
    layer0_outputs(2463) <= not((inputs(32)) xor (inputs(86)));
    layer0_outputs(2464) <= (inputs(77)) xor (inputs(151));
    layer0_outputs(2465) <= not((inputs(66)) or (inputs(184)));
    layer0_outputs(2466) <= inputs(215);
    layer0_outputs(2467) <= (inputs(247)) or (inputs(213));
    layer0_outputs(2468) <= not(inputs(148));
    layer0_outputs(2469) <= not(inputs(8));
    layer0_outputs(2470) <= (inputs(233)) or (inputs(0));
    layer0_outputs(2471) <= (inputs(221)) and not (inputs(59));
    layer0_outputs(2472) <= not((inputs(244)) or (inputs(206)));
    layer0_outputs(2473) <= '1';
    layer0_outputs(2474) <= '0';
    layer0_outputs(2475) <= not((inputs(76)) or (inputs(20)));
    layer0_outputs(2476) <= (inputs(153)) or (inputs(163));
    layer0_outputs(2477) <= (inputs(167)) and not (inputs(37));
    layer0_outputs(2478) <= not(inputs(195));
    layer0_outputs(2479) <= (inputs(81)) or (inputs(94));
    layer0_outputs(2480) <= '1';
    layer0_outputs(2481) <= not((inputs(70)) or (inputs(144)));
    layer0_outputs(2482) <= (inputs(88)) and (inputs(125));
    layer0_outputs(2483) <= inputs(239);
    layer0_outputs(2484) <= (inputs(140)) xor (inputs(107));
    layer0_outputs(2485) <= not((inputs(198)) or (inputs(70)));
    layer0_outputs(2486) <= (inputs(29)) xor (inputs(124));
    layer0_outputs(2487) <= inputs(37);
    layer0_outputs(2488) <= inputs(160);
    layer0_outputs(2489) <= not(inputs(55));
    layer0_outputs(2490) <= not((inputs(126)) or (inputs(250)));
    layer0_outputs(2491) <= inputs(188);
    layer0_outputs(2492) <= inputs(181);
    layer0_outputs(2493) <= (inputs(164)) or (inputs(181));
    layer0_outputs(2494) <= (inputs(136)) and not (inputs(57));
    layer0_outputs(2495) <= (inputs(72)) and not (inputs(211));
    layer0_outputs(2496) <= '0';
    layer0_outputs(2497) <= inputs(125);
    layer0_outputs(2498) <= not(inputs(33)) or (inputs(94));
    layer0_outputs(2499) <= not(inputs(96));
    layer0_outputs(2500) <= not(inputs(224));
    layer0_outputs(2501) <= inputs(147);
    layer0_outputs(2502) <= (inputs(76)) and not (inputs(239));
    layer0_outputs(2503) <= (inputs(146)) or (inputs(231));
    layer0_outputs(2504) <= (inputs(102)) or (inputs(95));
    layer0_outputs(2505) <= (inputs(187)) and not (inputs(61));
    layer0_outputs(2506) <= (inputs(188)) and not (inputs(94));
    layer0_outputs(2507) <= not(inputs(59)) or (inputs(89));
    layer0_outputs(2508) <= not((inputs(35)) xor (inputs(7)));
    layer0_outputs(2509) <= (inputs(165)) or (inputs(135));
    layer0_outputs(2510) <= inputs(81);
    layer0_outputs(2511) <= inputs(5);
    layer0_outputs(2512) <= not(inputs(184));
    layer0_outputs(2513) <= not(inputs(172));
    layer0_outputs(2514) <= inputs(148);
    layer0_outputs(2515) <= not((inputs(213)) or (inputs(151)));
    layer0_outputs(2516) <= (inputs(231)) or (inputs(178));
    layer0_outputs(2517) <= not(inputs(31)) or (inputs(234));
    layer0_outputs(2518) <= not((inputs(1)) xor (inputs(11)));
    layer0_outputs(2519) <= not(inputs(46)) or (inputs(193));
    layer0_outputs(2520) <= (inputs(30)) or (inputs(64));
    layer0_outputs(2521) <= inputs(116);
    layer0_outputs(2522) <= inputs(245);
    layer0_outputs(2523) <= not(inputs(199)) or (inputs(35));
    layer0_outputs(2524) <= not((inputs(74)) or (inputs(91)));
    layer0_outputs(2525) <= not(inputs(48)) or (inputs(131));
    layer0_outputs(2526) <= not(inputs(213));
    layer0_outputs(2527) <= inputs(103);
    layer0_outputs(2528) <= not(inputs(98));
    layer0_outputs(2529) <= inputs(151);
    layer0_outputs(2530) <= (inputs(217)) and not (inputs(18));
    layer0_outputs(2531) <= not((inputs(111)) xor (inputs(63)));
    layer0_outputs(2532) <= not(inputs(248)) or (inputs(59));
    layer0_outputs(2533) <= inputs(5);
    layer0_outputs(2534) <= inputs(103);
    layer0_outputs(2535) <= (inputs(148)) and not (inputs(17));
    layer0_outputs(2536) <= not(inputs(182));
    layer0_outputs(2537) <= (inputs(31)) or (inputs(173));
    layer0_outputs(2538) <= (inputs(170)) or (inputs(21));
    layer0_outputs(2539) <= not(inputs(214));
    layer0_outputs(2540) <= not(inputs(13)) or (inputs(42));
    layer0_outputs(2541) <= not((inputs(62)) or (inputs(159)));
    layer0_outputs(2542) <= inputs(99);
    layer0_outputs(2543) <= not(inputs(156));
    layer0_outputs(2544) <= not((inputs(229)) and (inputs(125)));
    layer0_outputs(2545) <= not(inputs(183)) or (inputs(88));
    layer0_outputs(2546) <= (inputs(104)) and not (inputs(36));
    layer0_outputs(2547) <= not(inputs(165));
    layer0_outputs(2548) <= (inputs(220)) and not (inputs(109));
    layer0_outputs(2549) <= not((inputs(225)) or (inputs(174)));
    layer0_outputs(2550) <= (inputs(209)) and not (inputs(9));
    layer0_outputs(2551) <= not(inputs(135)) or (inputs(178));
    layer0_outputs(2552) <= inputs(204);
    layer0_outputs(2553) <= (inputs(23)) or (inputs(128));
    layer0_outputs(2554) <= not((inputs(198)) and (inputs(137)));
    layer0_outputs(2555) <= inputs(230);
    layer0_outputs(2556) <= not((inputs(221)) or (inputs(219)));
    layer0_outputs(2557) <= not(inputs(22));
    layer0_outputs(2558) <= (inputs(111)) or (inputs(161));
    layer0_outputs(2559) <= (inputs(167)) and (inputs(105));
    layer0_outputs(2560) <= not(inputs(90));
    layer0_outputs(2561) <= (inputs(221)) or (inputs(145));
    layer0_outputs(2562) <= (inputs(105)) and not (inputs(130));
    layer0_outputs(2563) <= inputs(27);
    layer0_outputs(2564) <= '0';
    layer0_outputs(2565) <= not(inputs(100));
    layer0_outputs(2566) <= not(inputs(231));
    layer0_outputs(2567) <= not((inputs(76)) or (inputs(34)));
    layer0_outputs(2568) <= not(inputs(85));
    layer0_outputs(2569) <= (inputs(194)) or (inputs(198));
    layer0_outputs(2570) <= (inputs(161)) or (inputs(48));
    layer0_outputs(2571) <= not(inputs(101)) or (inputs(88));
    layer0_outputs(2572) <= (inputs(180)) or (inputs(70));
    layer0_outputs(2573) <= (inputs(230)) or (inputs(96));
    layer0_outputs(2574) <= (inputs(59)) xor (inputs(9));
    layer0_outputs(2575) <= not((inputs(45)) or (inputs(12)));
    layer0_outputs(2576) <= not((inputs(202)) or (inputs(79)));
    layer0_outputs(2577) <= inputs(21);
    layer0_outputs(2578) <= (inputs(19)) or (inputs(207));
    layer0_outputs(2579) <= (inputs(219)) and (inputs(244));
    layer0_outputs(2580) <= not(inputs(39)) or (inputs(143));
    layer0_outputs(2581) <= (inputs(56)) xor (inputs(29));
    layer0_outputs(2582) <= not(inputs(234));
    layer0_outputs(2583) <= inputs(208);
    layer0_outputs(2584) <= not(inputs(66));
    layer0_outputs(2585) <= (inputs(39)) and not (inputs(208));
    layer0_outputs(2586) <= (inputs(214)) and not (inputs(33));
    layer0_outputs(2587) <= not(inputs(232)) or (inputs(73));
    layer0_outputs(2588) <= not(inputs(72));
    layer0_outputs(2589) <= (inputs(89)) and not (inputs(64));
    layer0_outputs(2590) <= not(inputs(26));
    layer0_outputs(2591) <= not((inputs(77)) xor (inputs(86)));
    layer0_outputs(2592) <= not(inputs(31)) or (inputs(12));
    layer0_outputs(2593) <= not(inputs(0)) or (inputs(171));
    layer0_outputs(2594) <= inputs(101);
    layer0_outputs(2595) <= inputs(23);
    layer0_outputs(2596) <= not((inputs(126)) or (inputs(239)));
    layer0_outputs(2597) <= '1';
    layer0_outputs(2598) <= (inputs(88)) and (inputs(136));
    layer0_outputs(2599) <= (inputs(59)) xor (inputs(121));
    layer0_outputs(2600) <= not(inputs(34));
    layer0_outputs(2601) <= not(inputs(32));
    layer0_outputs(2602) <= (inputs(118)) and not (inputs(242));
    layer0_outputs(2603) <= inputs(196);
    layer0_outputs(2604) <= (inputs(182)) and not (inputs(132));
    layer0_outputs(2605) <= inputs(0);
    layer0_outputs(2606) <= (inputs(56)) and (inputs(184));
    layer0_outputs(2607) <= not(inputs(197));
    layer0_outputs(2608) <= (inputs(251)) and not (inputs(200));
    layer0_outputs(2609) <= (inputs(23)) and not (inputs(14));
    layer0_outputs(2610) <= not(inputs(14));
    layer0_outputs(2611) <= inputs(46);
    layer0_outputs(2612) <= (inputs(94)) or (inputs(54));
    layer0_outputs(2613) <= not((inputs(73)) xor (inputs(251)));
    layer0_outputs(2614) <= (inputs(219)) and not (inputs(45));
    layer0_outputs(2615) <= not((inputs(198)) and (inputs(54)));
    layer0_outputs(2616) <= not(inputs(229));
    layer0_outputs(2617) <= not((inputs(215)) or (inputs(8)));
    layer0_outputs(2618) <= (inputs(51)) and not (inputs(127));
    layer0_outputs(2619) <= not((inputs(246)) or (inputs(205)));
    layer0_outputs(2620) <= (inputs(141)) xor (inputs(207));
    layer0_outputs(2621) <= not((inputs(189)) xor (inputs(220)));
    layer0_outputs(2622) <= (inputs(137)) xor (inputs(221));
    layer0_outputs(2623) <= (inputs(41)) and not (inputs(217));
    layer0_outputs(2624) <= inputs(68);
    layer0_outputs(2625) <= not(inputs(151));
    layer0_outputs(2626) <= inputs(85);
    layer0_outputs(2627) <= not(inputs(75)) or (inputs(243));
    layer0_outputs(2628) <= (inputs(129)) xor (inputs(116));
    layer0_outputs(2629) <= not(inputs(46)) or (inputs(255));
    layer0_outputs(2630) <= not(inputs(213));
    layer0_outputs(2631) <= not(inputs(80));
    layer0_outputs(2632) <= not((inputs(194)) or (inputs(133)));
    layer0_outputs(2633) <= '1';
    layer0_outputs(2634) <= (inputs(159)) and not (inputs(98));
    layer0_outputs(2635) <= (inputs(127)) or (inputs(100));
    layer0_outputs(2636) <= not(inputs(97)) or (inputs(133));
    layer0_outputs(2637) <= not(inputs(146));
    layer0_outputs(2638) <= not(inputs(68)) or (inputs(20));
    layer0_outputs(2639) <= inputs(18);
    layer0_outputs(2640) <= not((inputs(25)) or (inputs(126)));
    layer0_outputs(2641) <= (inputs(115)) or (inputs(246));
    layer0_outputs(2642) <= inputs(19);
    layer0_outputs(2643) <= not((inputs(0)) or (inputs(145)));
    layer0_outputs(2644) <= not((inputs(127)) or (inputs(227)));
    layer0_outputs(2645) <= not(inputs(227));
    layer0_outputs(2646) <= inputs(162);
    layer0_outputs(2647) <= (inputs(91)) xor (inputs(174));
    layer0_outputs(2648) <= (inputs(108)) or (inputs(82));
    layer0_outputs(2649) <= not(inputs(103));
    layer0_outputs(2650) <= not(inputs(55));
    layer0_outputs(2651) <= inputs(99);
    layer0_outputs(2652) <= (inputs(72)) or (inputs(218));
    layer0_outputs(2653) <= not((inputs(131)) or (inputs(116)));
    layer0_outputs(2654) <= inputs(99);
    layer0_outputs(2655) <= (inputs(7)) and not (inputs(114));
    layer0_outputs(2656) <= not(inputs(225)) or (inputs(159));
    layer0_outputs(2657) <= not((inputs(203)) or (inputs(190)));
    layer0_outputs(2658) <= (inputs(26)) and not (inputs(198));
    layer0_outputs(2659) <= inputs(90);
    layer0_outputs(2660) <= not(inputs(165));
    layer0_outputs(2661) <= not((inputs(192)) or (inputs(165)));
    layer0_outputs(2662) <= (inputs(75)) xor (inputs(199));
    layer0_outputs(2663) <= inputs(246);
    layer0_outputs(2664) <= (inputs(80)) or (inputs(227));
    layer0_outputs(2665) <= inputs(9);
    layer0_outputs(2666) <= not(inputs(39));
    layer0_outputs(2667) <= not((inputs(93)) or (inputs(219)));
    layer0_outputs(2668) <= not((inputs(111)) or (inputs(78)));
    layer0_outputs(2669) <= not(inputs(230));
    layer0_outputs(2670) <= not(inputs(119));
    layer0_outputs(2671) <= not((inputs(158)) or (inputs(130)));
    layer0_outputs(2672) <= not((inputs(248)) or (inputs(217)));
    layer0_outputs(2673) <= inputs(156);
    layer0_outputs(2674) <= inputs(120);
    layer0_outputs(2675) <= (inputs(27)) and not (inputs(150));
    layer0_outputs(2676) <= not(inputs(199)) or (inputs(56));
    layer0_outputs(2677) <= not((inputs(50)) or (inputs(168)));
    layer0_outputs(2678) <= not(inputs(42));
    layer0_outputs(2679) <= not((inputs(191)) and (inputs(147)));
    layer0_outputs(2680) <= (inputs(97)) or (inputs(161));
    layer0_outputs(2681) <= (inputs(123)) and not (inputs(36));
    layer0_outputs(2682) <= inputs(122);
    layer0_outputs(2683) <= inputs(26);
    layer0_outputs(2684) <= not((inputs(221)) xor (inputs(32)));
    layer0_outputs(2685) <= (inputs(100)) or (inputs(167));
    layer0_outputs(2686) <= not(inputs(233)) or (inputs(145));
    layer0_outputs(2687) <= inputs(209);
    layer0_outputs(2688) <= not(inputs(231));
    layer0_outputs(2689) <= (inputs(206)) and not (inputs(62));
    layer0_outputs(2690) <= not(inputs(102));
    layer0_outputs(2691) <= not(inputs(246)) or (inputs(77));
    layer0_outputs(2692) <= not(inputs(73));
    layer0_outputs(2693) <= inputs(20);
    layer0_outputs(2694) <= '0';
    layer0_outputs(2695) <= not((inputs(125)) xor (inputs(64)));
    layer0_outputs(2696) <= not((inputs(200)) or (inputs(203)));
    layer0_outputs(2697) <= inputs(248);
    layer0_outputs(2698) <= not(inputs(19)) or (inputs(113));
    layer0_outputs(2699) <= inputs(174);
    layer0_outputs(2700) <= (inputs(51)) or (inputs(244));
    layer0_outputs(2701) <= '0';
    layer0_outputs(2702) <= not(inputs(158)) or (inputs(253));
    layer0_outputs(2703) <= not(inputs(134));
    layer0_outputs(2704) <= (inputs(122)) and not (inputs(128));
    layer0_outputs(2705) <= not(inputs(129));
    layer0_outputs(2706) <= (inputs(86)) or (inputs(111));
    layer0_outputs(2707) <= inputs(143);
    layer0_outputs(2708) <= not(inputs(99));
    layer0_outputs(2709) <= (inputs(36)) xor (inputs(136));
    layer0_outputs(2710) <= (inputs(176)) or (inputs(187));
    layer0_outputs(2711) <= not(inputs(236)) or (inputs(2));
    layer0_outputs(2712) <= inputs(138);
    layer0_outputs(2713) <= inputs(82);
    layer0_outputs(2714) <= (inputs(42)) or (inputs(107));
    layer0_outputs(2715) <= not((inputs(34)) xor (inputs(61)));
    layer0_outputs(2716) <= not(inputs(151));
    layer0_outputs(2717) <= not(inputs(160));
    layer0_outputs(2718) <= (inputs(252)) and not (inputs(244));
    layer0_outputs(2719) <= not((inputs(224)) or (inputs(234)));
    layer0_outputs(2720) <= not((inputs(135)) or (inputs(18)));
    layer0_outputs(2721) <= (inputs(123)) or (inputs(66));
    layer0_outputs(2722) <= not(inputs(166));
    layer0_outputs(2723) <= not(inputs(68)) or (inputs(131));
    layer0_outputs(2724) <= (inputs(27)) and not (inputs(150));
    layer0_outputs(2725) <= (inputs(239)) or (inputs(52));
    layer0_outputs(2726) <= (inputs(81)) or (inputs(8));
    layer0_outputs(2727) <= not((inputs(236)) or (inputs(163)));
    layer0_outputs(2728) <= (inputs(233)) or (inputs(144));
    layer0_outputs(2729) <= not(inputs(85));
    layer0_outputs(2730) <= (inputs(51)) and not (inputs(234));
    layer0_outputs(2731) <= not(inputs(186)) or (inputs(66));
    layer0_outputs(2732) <= (inputs(7)) or (inputs(85));
    layer0_outputs(2733) <= not((inputs(199)) and (inputs(127)));
    layer0_outputs(2734) <= (inputs(174)) xor (inputs(27));
    layer0_outputs(2735) <= (inputs(16)) or (inputs(185));
    layer0_outputs(2736) <= not(inputs(136));
    layer0_outputs(2737) <= not(inputs(106));
    layer0_outputs(2738) <= (inputs(163)) or (inputs(94));
    layer0_outputs(2739) <= (inputs(96)) xor (inputs(86));
    layer0_outputs(2740) <= (inputs(139)) xor (inputs(170));
    layer0_outputs(2741) <= (inputs(95)) or (inputs(152));
    layer0_outputs(2742) <= (inputs(101)) or (inputs(12));
    layer0_outputs(2743) <= (inputs(78)) or (inputs(46));
    layer0_outputs(2744) <= not(inputs(138));
    layer0_outputs(2745) <= (inputs(11)) xor (inputs(35));
    layer0_outputs(2746) <= not((inputs(7)) or (inputs(156)));
    layer0_outputs(2747) <= not(inputs(204)) or (inputs(109));
    layer0_outputs(2748) <= not(inputs(199)) or (inputs(213));
    layer0_outputs(2749) <= inputs(63);
    layer0_outputs(2750) <= not((inputs(111)) or (inputs(252)));
    layer0_outputs(2751) <= not((inputs(116)) or (inputs(190)));
    layer0_outputs(2752) <= not(inputs(59));
    layer0_outputs(2753) <= not(inputs(215)) or (inputs(132));
    layer0_outputs(2754) <= not(inputs(29));
    layer0_outputs(2755) <= not(inputs(26));
    layer0_outputs(2756) <= not(inputs(211));
    layer0_outputs(2757) <= inputs(137);
    layer0_outputs(2758) <= (inputs(100)) or (inputs(116));
    layer0_outputs(2759) <= inputs(213);
    layer0_outputs(2760) <= not(inputs(26));
    layer0_outputs(2761) <= not(inputs(101));
    layer0_outputs(2762) <= inputs(150);
    layer0_outputs(2763) <= not((inputs(163)) or (inputs(176)));
    layer0_outputs(2764) <= not((inputs(127)) or (inputs(6)));
    layer0_outputs(2765) <= (inputs(170)) and not (inputs(115));
    layer0_outputs(2766) <= not(inputs(220));
    layer0_outputs(2767) <= inputs(27);
    layer0_outputs(2768) <= (inputs(37)) and not (inputs(88));
    layer0_outputs(2769) <= (inputs(17)) xor (inputs(204));
    layer0_outputs(2770) <= '0';
    layer0_outputs(2771) <= inputs(129);
    layer0_outputs(2772) <= not((inputs(16)) or (inputs(234)));
    layer0_outputs(2773) <= inputs(147);
    layer0_outputs(2774) <= not((inputs(148)) or (inputs(232)));
    layer0_outputs(2775) <= not((inputs(32)) or (inputs(218)));
    layer0_outputs(2776) <= (inputs(162)) and not (inputs(47));
    layer0_outputs(2777) <= not(inputs(108)) or (inputs(1));
    layer0_outputs(2778) <= not((inputs(33)) and (inputs(19)));
    layer0_outputs(2779) <= not(inputs(109)) or (inputs(109));
    layer0_outputs(2780) <= (inputs(199)) and not (inputs(17));
    layer0_outputs(2781) <= inputs(131);
    layer0_outputs(2782) <= inputs(48);
    layer0_outputs(2783) <= not(inputs(164));
    layer0_outputs(2784) <= (inputs(185)) xor (inputs(172));
    layer0_outputs(2785) <= inputs(133);
    layer0_outputs(2786) <= (inputs(235)) and not (inputs(254));
    layer0_outputs(2787) <= not(inputs(198)) or (inputs(66));
    layer0_outputs(2788) <= not(inputs(134)) or (inputs(140));
    layer0_outputs(2789) <= (inputs(213)) and not (inputs(119));
    layer0_outputs(2790) <= not(inputs(107));
    layer0_outputs(2791) <= inputs(5);
    layer0_outputs(2792) <= not(inputs(104)) or (inputs(16));
    layer0_outputs(2793) <= not(inputs(161));
    layer0_outputs(2794) <= not(inputs(167)) or (inputs(31));
    layer0_outputs(2795) <= (inputs(184)) or (inputs(76));
    layer0_outputs(2796) <= not(inputs(7)) or (inputs(233));
    layer0_outputs(2797) <= (inputs(108)) or (inputs(78));
    layer0_outputs(2798) <= inputs(237);
    layer0_outputs(2799) <= inputs(227);
    layer0_outputs(2800) <= (inputs(58)) and not (inputs(215));
    layer0_outputs(2801) <= not((inputs(52)) or (inputs(252)));
    layer0_outputs(2802) <= (inputs(4)) or (inputs(239));
    layer0_outputs(2803) <= inputs(115);
    layer0_outputs(2804) <= not((inputs(61)) xor (inputs(250)));
    layer0_outputs(2805) <= (inputs(34)) or (inputs(149));
    layer0_outputs(2806) <= not((inputs(152)) xor (inputs(213)));
    layer0_outputs(2807) <= (inputs(105)) and not (inputs(229));
    layer0_outputs(2808) <= (inputs(105)) and not (inputs(119));
    layer0_outputs(2809) <= (inputs(20)) or (inputs(34));
    layer0_outputs(2810) <= not(inputs(122));
    layer0_outputs(2811) <= inputs(110);
    layer0_outputs(2812) <= (inputs(42)) or (inputs(95));
    layer0_outputs(2813) <= not(inputs(35));
    layer0_outputs(2814) <= inputs(146);
    layer0_outputs(2815) <= (inputs(22)) and not (inputs(29));
    layer0_outputs(2816) <= not((inputs(142)) and (inputs(47)));
    layer0_outputs(2817) <= not((inputs(164)) xor (inputs(155)));
    layer0_outputs(2818) <= not((inputs(93)) or (inputs(69)));
    layer0_outputs(2819) <= (inputs(246)) xor (inputs(4));
    layer0_outputs(2820) <= not(inputs(39)) or (inputs(175));
    layer0_outputs(2821) <= inputs(164);
    layer0_outputs(2822) <= not((inputs(48)) xor (inputs(189)));
    layer0_outputs(2823) <= inputs(93);
    layer0_outputs(2824) <= not(inputs(206));
    layer0_outputs(2825) <= inputs(181);
    layer0_outputs(2826) <= (inputs(76)) xor (inputs(105));
    layer0_outputs(2827) <= not(inputs(49));
    layer0_outputs(2828) <= not(inputs(23));
    layer0_outputs(2829) <= not((inputs(99)) or (inputs(113)));
    layer0_outputs(2830) <= inputs(44);
    layer0_outputs(2831) <= not(inputs(102));
    layer0_outputs(2832) <= inputs(105);
    layer0_outputs(2833) <= (inputs(113)) or (inputs(144));
    layer0_outputs(2834) <= not((inputs(3)) and (inputs(134)));
    layer0_outputs(2835) <= inputs(102);
    layer0_outputs(2836) <= inputs(121);
    layer0_outputs(2837) <= inputs(77);
    layer0_outputs(2838) <= not(inputs(146));
    layer0_outputs(2839) <= inputs(5);
    layer0_outputs(2840) <= not(inputs(183)) or (inputs(77));
    layer0_outputs(2841) <= not((inputs(64)) or (inputs(169)));
    layer0_outputs(2842) <= '0';
    layer0_outputs(2843) <= not((inputs(73)) and (inputs(105)));
    layer0_outputs(2844) <= not(inputs(19)) or (inputs(140));
    layer0_outputs(2845) <= (inputs(210)) or (inputs(102));
    layer0_outputs(2846) <= (inputs(36)) and (inputs(117));
    layer0_outputs(2847) <= not((inputs(225)) or (inputs(197)));
    layer0_outputs(2848) <= not(inputs(90)) or (inputs(159));
    layer0_outputs(2849) <= not((inputs(106)) or (inputs(185)));
    layer0_outputs(2850) <= '1';
    layer0_outputs(2851) <= (inputs(214)) or (inputs(2));
    layer0_outputs(2852) <= not((inputs(122)) or (inputs(163)));
    layer0_outputs(2853) <= not((inputs(204)) xor (inputs(121)));
    layer0_outputs(2854) <= not(inputs(222)) or (inputs(71));
    layer0_outputs(2855) <= inputs(242);
    layer0_outputs(2856) <= inputs(240);
    layer0_outputs(2857) <= not((inputs(176)) xor (inputs(0)));
    layer0_outputs(2858) <= (inputs(149)) and not (inputs(36));
    layer0_outputs(2859) <= not(inputs(105)) or (inputs(207));
    layer0_outputs(2860) <= '1';
    layer0_outputs(2861) <= not(inputs(69));
    layer0_outputs(2862) <= inputs(52);
    layer0_outputs(2863) <= not((inputs(156)) and (inputs(156)));
    layer0_outputs(2864) <= (inputs(144)) xor (inputs(165));
    layer0_outputs(2865) <= not(inputs(89));
    layer0_outputs(2866) <= (inputs(150)) and not (inputs(157));
    layer0_outputs(2867) <= (inputs(108)) or (inputs(175));
    layer0_outputs(2868) <= (inputs(218)) and not (inputs(75));
    layer0_outputs(2869) <= not((inputs(148)) or (inputs(189)));
    layer0_outputs(2870) <= not(inputs(186)) or (inputs(36));
    layer0_outputs(2871) <= not(inputs(241)) or (inputs(75));
    layer0_outputs(2872) <= not(inputs(75));
    layer0_outputs(2873) <= '0';
    layer0_outputs(2874) <= (inputs(68)) or (inputs(145));
    layer0_outputs(2875) <= (inputs(157)) or (inputs(150));
    layer0_outputs(2876) <= not(inputs(173)) or (inputs(27));
    layer0_outputs(2877) <= inputs(105);
    layer0_outputs(2878) <= not(inputs(166));
    layer0_outputs(2879) <= not(inputs(135));
    layer0_outputs(2880) <= not(inputs(157)) or (inputs(170));
    layer0_outputs(2881) <= not((inputs(157)) or (inputs(23)));
    layer0_outputs(2882) <= not((inputs(64)) or (inputs(163)));
    layer0_outputs(2883) <= (inputs(85)) and not (inputs(251));
    layer0_outputs(2884) <= inputs(182);
    layer0_outputs(2885) <= inputs(26);
    layer0_outputs(2886) <= inputs(82);
    layer0_outputs(2887) <= '1';
    layer0_outputs(2888) <= not(inputs(214));
    layer0_outputs(2889) <= (inputs(210)) and not (inputs(156));
    layer0_outputs(2890) <= (inputs(78)) or (inputs(49));
    layer0_outputs(2891) <= inputs(110);
    layer0_outputs(2892) <= (inputs(158)) or (inputs(247));
    layer0_outputs(2893) <= inputs(34);
    layer0_outputs(2894) <= inputs(18);
    layer0_outputs(2895) <= inputs(104);
    layer0_outputs(2896) <= not(inputs(196));
    layer0_outputs(2897) <= not(inputs(100));
    layer0_outputs(2898) <= (inputs(250)) and not (inputs(137));
    layer0_outputs(2899) <= not((inputs(96)) xor (inputs(7)));
    layer0_outputs(2900) <= not(inputs(83)) or (inputs(157));
    layer0_outputs(2901) <= (inputs(187)) or (inputs(39));
    layer0_outputs(2902) <= not(inputs(103)) or (inputs(200));
    layer0_outputs(2903) <= not(inputs(210));
    layer0_outputs(2904) <= (inputs(248)) or (inputs(45));
    layer0_outputs(2905) <= not(inputs(11)) or (inputs(80));
    layer0_outputs(2906) <= not(inputs(150)) or (inputs(228));
    layer0_outputs(2907) <= not((inputs(240)) xor (inputs(66)));
    layer0_outputs(2908) <= (inputs(75)) or (inputs(155));
    layer0_outputs(2909) <= not(inputs(205));
    layer0_outputs(2910) <= (inputs(249)) or (inputs(102));
    layer0_outputs(2911) <= (inputs(228)) or (inputs(137));
    layer0_outputs(2912) <= '0';
    layer0_outputs(2913) <= not((inputs(55)) xor (inputs(12)));
    layer0_outputs(2914) <= not(inputs(150));
    layer0_outputs(2915) <= (inputs(54)) xor (inputs(189));
    layer0_outputs(2916) <= inputs(167);
    layer0_outputs(2917) <= inputs(25);
    layer0_outputs(2918) <= (inputs(231)) and not (inputs(254));
    layer0_outputs(2919) <= (inputs(196)) or (inputs(18));
    layer0_outputs(2920) <= (inputs(51)) xor (inputs(5));
    layer0_outputs(2921) <= not((inputs(58)) or (inputs(121)));
    layer0_outputs(2922) <= not(inputs(141)) or (inputs(233));
    layer0_outputs(2923) <= not(inputs(201)) or (inputs(39));
    layer0_outputs(2924) <= inputs(136);
    layer0_outputs(2925) <= not((inputs(14)) or (inputs(142)));
    layer0_outputs(2926) <= not(inputs(25));
    layer0_outputs(2927) <= inputs(229);
    layer0_outputs(2928) <= inputs(110);
    layer0_outputs(2929) <= (inputs(181)) and not (inputs(241));
    layer0_outputs(2930) <= (inputs(183)) and not (inputs(142));
    layer0_outputs(2931) <= not(inputs(73));
    layer0_outputs(2932) <= not(inputs(106));
    layer0_outputs(2933) <= inputs(33);
    layer0_outputs(2934) <= inputs(147);
    layer0_outputs(2935) <= not(inputs(151));
    layer0_outputs(2936) <= not(inputs(6)) or (inputs(145));
    layer0_outputs(2937) <= (inputs(47)) and (inputs(201));
    layer0_outputs(2938) <= not(inputs(228));
    layer0_outputs(2939) <= not(inputs(159));
    layer0_outputs(2940) <= not(inputs(116));
    layer0_outputs(2941) <= not(inputs(116));
    layer0_outputs(2942) <= not((inputs(168)) or (inputs(121)));
    layer0_outputs(2943) <= (inputs(9)) and not (inputs(196));
    layer0_outputs(2944) <= (inputs(243)) or (inputs(137));
    layer0_outputs(2945) <= (inputs(71)) and not (inputs(44));
    layer0_outputs(2946) <= (inputs(238)) or (inputs(67));
    layer0_outputs(2947) <= inputs(253);
    layer0_outputs(2948) <= not(inputs(125)) or (inputs(225));
    layer0_outputs(2949) <= '1';
    layer0_outputs(2950) <= inputs(248);
    layer0_outputs(2951) <= not(inputs(32));
    layer0_outputs(2952) <= inputs(94);
    layer0_outputs(2953) <= inputs(248);
    layer0_outputs(2954) <= (inputs(132)) or (inputs(207));
    layer0_outputs(2955) <= inputs(119);
    layer0_outputs(2956) <= inputs(72);
    layer0_outputs(2957) <= (inputs(48)) or (inputs(24));
    layer0_outputs(2958) <= (inputs(54)) or (inputs(247));
    layer0_outputs(2959) <= inputs(111);
    layer0_outputs(2960) <= not(inputs(61));
    layer0_outputs(2961) <= (inputs(26)) and not (inputs(237));
    layer0_outputs(2962) <= inputs(60);
    layer0_outputs(2963) <= inputs(87);
    layer0_outputs(2964) <= not((inputs(245)) or (inputs(193)));
    layer0_outputs(2965) <= (inputs(233)) xor (inputs(241));
    layer0_outputs(2966) <= not(inputs(108)) or (inputs(208));
    layer0_outputs(2967) <= (inputs(72)) or (inputs(224));
    layer0_outputs(2968) <= (inputs(67)) and not (inputs(3));
    layer0_outputs(2969) <= inputs(219);
    layer0_outputs(2970) <= inputs(180);
    layer0_outputs(2971) <= (inputs(255)) or (inputs(4));
    layer0_outputs(2972) <= (inputs(125)) or (inputs(90));
    layer0_outputs(2973) <= not(inputs(93));
    layer0_outputs(2974) <= not(inputs(40));
    layer0_outputs(2975) <= inputs(155);
    layer0_outputs(2976) <= inputs(45);
    layer0_outputs(2977) <= '0';
    layer0_outputs(2978) <= (inputs(4)) and not (inputs(41));
    layer0_outputs(2979) <= inputs(67);
    layer0_outputs(2980) <= (inputs(231)) and not (inputs(207));
    layer0_outputs(2981) <= not((inputs(214)) xor (inputs(225)));
    layer0_outputs(2982) <= not((inputs(205)) or (inputs(149)));
    layer0_outputs(2983) <= not((inputs(158)) or (inputs(9)));
    layer0_outputs(2984) <= not(inputs(248));
    layer0_outputs(2985) <= inputs(158);
    layer0_outputs(2986) <= not(inputs(217));
    layer0_outputs(2987) <= '0';
    layer0_outputs(2988) <= inputs(217);
    layer0_outputs(2989) <= (inputs(73)) and not (inputs(111));
    layer0_outputs(2990) <= (inputs(226)) or (inputs(234));
    layer0_outputs(2991) <= (inputs(227)) and not (inputs(255));
    layer0_outputs(2992) <= not((inputs(153)) xor (inputs(184)));
    layer0_outputs(2993) <= not(inputs(26)) or (inputs(208));
    layer0_outputs(2994) <= (inputs(89)) or (inputs(153));
    layer0_outputs(2995) <= (inputs(238)) and not (inputs(54));
    layer0_outputs(2996) <= inputs(23);
    layer0_outputs(2997) <= not(inputs(122));
    layer0_outputs(2998) <= (inputs(39)) and not (inputs(148));
    layer0_outputs(2999) <= '1';
    layer0_outputs(3000) <= (inputs(26)) or (inputs(41));
    layer0_outputs(3001) <= inputs(152);
    layer0_outputs(3002) <= inputs(82);
    layer0_outputs(3003) <= (inputs(224)) or (inputs(86));
    layer0_outputs(3004) <= not(inputs(13));
    layer0_outputs(3005) <= (inputs(8)) and not (inputs(147));
    layer0_outputs(3006) <= not(inputs(189)) or (inputs(252));
    layer0_outputs(3007) <= (inputs(136)) and not (inputs(30));
    layer0_outputs(3008) <= not(inputs(42));
    layer0_outputs(3009) <= (inputs(123)) and not (inputs(47));
    layer0_outputs(3010) <= not(inputs(167)) or (inputs(142));
    layer0_outputs(3011) <= not(inputs(178));
    layer0_outputs(3012) <= not(inputs(246));
    layer0_outputs(3013) <= (inputs(193)) and not (inputs(223));
    layer0_outputs(3014) <= inputs(195);
    layer0_outputs(3015) <= inputs(168);
    layer0_outputs(3016) <= (inputs(4)) or (inputs(144));
    layer0_outputs(3017) <= not(inputs(245));
    layer0_outputs(3018) <= inputs(122);
    layer0_outputs(3019) <= (inputs(212)) or (inputs(82));
    layer0_outputs(3020) <= not(inputs(88)) or (inputs(160));
    layer0_outputs(3021) <= (inputs(57)) and (inputs(42));
    layer0_outputs(3022) <= '0';
    layer0_outputs(3023) <= not(inputs(149));
    layer0_outputs(3024) <= inputs(130);
    layer0_outputs(3025) <= not((inputs(202)) or (inputs(178)));
    layer0_outputs(3026) <= not((inputs(170)) or (inputs(130)));
    layer0_outputs(3027) <= inputs(84);
    layer0_outputs(3028) <= inputs(101);
    layer0_outputs(3029) <= not((inputs(22)) or (inputs(239)));
    layer0_outputs(3030) <= not((inputs(243)) xor (inputs(238)));
    layer0_outputs(3031) <= not((inputs(55)) xor (inputs(165)));
    layer0_outputs(3032) <= inputs(92);
    layer0_outputs(3033) <= inputs(29);
    layer0_outputs(3034) <= not((inputs(161)) or (inputs(41)));
    layer0_outputs(3035) <= inputs(124);
    layer0_outputs(3036) <= inputs(9);
    layer0_outputs(3037) <= inputs(196);
    layer0_outputs(3038) <= (inputs(153)) xor (inputs(28));
    layer0_outputs(3039) <= (inputs(62)) and (inputs(42));
    layer0_outputs(3040) <= inputs(211);
    layer0_outputs(3041) <= inputs(18);
    layer0_outputs(3042) <= inputs(177);
    layer0_outputs(3043) <= (inputs(19)) and not (inputs(14));
    layer0_outputs(3044) <= (inputs(15)) or (inputs(120));
    layer0_outputs(3045) <= not(inputs(115));
    layer0_outputs(3046) <= not(inputs(230));
    layer0_outputs(3047) <= (inputs(179)) and not (inputs(42));
    layer0_outputs(3048) <= not((inputs(10)) or (inputs(197)));
    layer0_outputs(3049) <= (inputs(24)) or (inputs(160));
    layer0_outputs(3050) <= (inputs(37)) or (inputs(175));
    layer0_outputs(3051) <= not((inputs(252)) or (inputs(151)));
    layer0_outputs(3052) <= (inputs(197)) xor (inputs(231));
    layer0_outputs(3053) <= inputs(127);
    layer0_outputs(3054) <= inputs(142);
    layer0_outputs(3055) <= not(inputs(93));
    layer0_outputs(3056) <= (inputs(65)) xor (inputs(25));
    layer0_outputs(3057) <= not((inputs(254)) or (inputs(126)));
    layer0_outputs(3058) <= not(inputs(76));
    layer0_outputs(3059) <= (inputs(235)) xor (inputs(95));
    layer0_outputs(3060) <= inputs(121);
    layer0_outputs(3061) <= (inputs(122)) and not (inputs(223));
    layer0_outputs(3062) <= not((inputs(33)) or (inputs(204)));
    layer0_outputs(3063) <= (inputs(140)) or (inputs(156));
    layer0_outputs(3064) <= (inputs(161)) and (inputs(186));
    layer0_outputs(3065) <= (inputs(23)) and not (inputs(222));
    layer0_outputs(3066) <= inputs(79);
    layer0_outputs(3067) <= inputs(138);
    layer0_outputs(3068) <= not(inputs(7));
    layer0_outputs(3069) <= not(inputs(23));
    layer0_outputs(3070) <= (inputs(141)) or (inputs(132));
    layer0_outputs(3071) <= not((inputs(181)) xor (inputs(77)));
    layer0_outputs(3072) <= not((inputs(49)) xor (inputs(71)));
    layer0_outputs(3073) <= (inputs(141)) and not (inputs(245));
    layer0_outputs(3074) <= not((inputs(103)) and (inputs(140)));
    layer0_outputs(3075) <= not((inputs(45)) xor (inputs(187)));
    layer0_outputs(3076) <= not(inputs(72));
    layer0_outputs(3077) <= not((inputs(215)) or (inputs(166)));
    layer0_outputs(3078) <= (inputs(83)) or (inputs(156));
    layer0_outputs(3079) <= (inputs(114)) or (inputs(113));
    layer0_outputs(3080) <= not((inputs(106)) or (inputs(131)));
    layer0_outputs(3081) <= not(inputs(45));
    layer0_outputs(3082) <= not(inputs(204));
    layer0_outputs(3083) <= inputs(105);
    layer0_outputs(3084) <= (inputs(13)) or (inputs(103));
    layer0_outputs(3085) <= not((inputs(225)) or (inputs(0)));
    layer0_outputs(3086) <= not((inputs(102)) or (inputs(118)));
    layer0_outputs(3087) <= not(inputs(180));
    layer0_outputs(3088) <= not((inputs(197)) or (inputs(159)));
    layer0_outputs(3089) <= inputs(8);
    layer0_outputs(3090) <= inputs(19);
    layer0_outputs(3091) <= inputs(73);
    layer0_outputs(3092) <= not((inputs(198)) and (inputs(5)));
    layer0_outputs(3093) <= (inputs(169)) or (inputs(221));
    layer0_outputs(3094) <= not((inputs(144)) or (inputs(178)));
    layer0_outputs(3095) <= (inputs(100)) or (inputs(246));
    layer0_outputs(3096) <= (inputs(241)) or (inputs(161));
    layer0_outputs(3097) <= inputs(129);
    layer0_outputs(3098) <= not(inputs(28)) or (inputs(223));
    layer0_outputs(3099) <= inputs(182);
    layer0_outputs(3100) <= (inputs(96)) and not (inputs(254));
    layer0_outputs(3101) <= (inputs(154)) xor (inputs(187));
    layer0_outputs(3102) <= '1';
    layer0_outputs(3103) <= inputs(46);
    layer0_outputs(3104) <= inputs(124);
    layer0_outputs(3105) <= not(inputs(206));
    layer0_outputs(3106) <= (inputs(144)) or (inputs(109));
    layer0_outputs(3107) <= inputs(68);
    layer0_outputs(3108) <= inputs(10);
    layer0_outputs(3109) <= not((inputs(55)) or (inputs(142)));
    layer0_outputs(3110) <= not((inputs(87)) or (inputs(226)));
    layer0_outputs(3111) <= not((inputs(181)) and (inputs(181)));
    layer0_outputs(3112) <= not(inputs(218));
    layer0_outputs(3113) <= (inputs(241)) and not (inputs(223));
    layer0_outputs(3114) <= (inputs(171)) and not (inputs(37));
    layer0_outputs(3115) <= (inputs(3)) or (inputs(35));
    layer0_outputs(3116) <= not(inputs(163)) or (inputs(32));
    layer0_outputs(3117) <= (inputs(117)) and not (inputs(79));
    layer0_outputs(3118) <= not(inputs(3));
    layer0_outputs(3119) <= (inputs(50)) xor (inputs(18));
    layer0_outputs(3120) <= inputs(14);
    layer0_outputs(3121) <= not(inputs(135)) or (inputs(110));
    layer0_outputs(3122) <= not((inputs(104)) or (inputs(81)));
    layer0_outputs(3123) <= not(inputs(164));
    layer0_outputs(3124) <= not(inputs(88));
    layer0_outputs(3125) <= (inputs(86)) and not (inputs(157));
    layer0_outputs(3126) <= (inputs(117)) or (inputs(208));
    layer0_outputs(3127) <= not(inputs(38));
    layer0_outputs(3128) <= (inputs(10)) and not (inputs(19));
    layer0_outputs(3129) <= not(inputs(167));
    layer0_outputs(3130) <= not(inputs(148));
    layer0_outputs(3131) <= inputs(137);
    layer0_outputs(3132) <= not(inputs(61));
    layer0_outputs(3133) <= not((inputs(246)) or (inputs(126)));
    layer0_outputs(3134) <= not((inputs(154)) or (inputs(7)));
    layer0_outputs(3135) <= inputs(34);
    layer0_outputs(3136) <= (inputs(57)) xor (inputs(36));
    layer0_outputs(3137) <= inputs(101);
    layer0_outputs(3138) <= (inputs(96)) and (inputs(71));
    layer0_outputs(3139) <= (inputs(67)) and not (inputs(143));
    layer0_outputs(3140) <= not(inputs(74));
    layer0_outputs(3141) <= not(inputs(150)) or (inputs(98));
    layer0_outputs(3142) <= not(inputs(226)) or (inputs(101));
    layer0_outputs(3143) <= not((inputs(64)) xor (inputs(16)));
    layer0_outputs(3144) <= not(inputs(120));
    layer0_outputs(3145) <= not((inputs(193)) or (inputs(178)));
    layer0_outputs(3146) <= not((inputs(135)) and (inputs(185)));
    layer0_outputs(3147) <= inputs(27);
    layer0_outputs(3148) <= inputs(115);
    layer0_outputs(3149) <= not(inputs(203));
    layer0_outputs(3150) <= (inputs(76)) or (inputs(143));
    layer0_outputs(3151) <= not(inputs(150)) or (inputs(172));
    layer0_outputs(3152) <= inputs(38);
    layer0_outputs(3153) <= (inputs(241)) or (inputs(239));
    layer0_outputs(3154) <= (inputs(239)) xor (inputs(234));
    layer0_outputs(3155) <= not(inputs(132));
    layer0_outputs(3156) <= not(inputs(89)) or (inputs(63));
    layer0_outputs(3157) <= not((inputs(7)) or (inputs(71)));
    layer0_outputs(3158) <= (inputs(163)) xor (inputs(179));
    layer0_outputs(3159) <= (inputs(114)) or (inputs(160));
    layer0_outputs(3160) <= (inputs(184)) or (inputs(200));
    layer0_outputs(3161) <= (inputs(39)) or (inputs(253));
    layer0_outputs(3162) <= not(inputs(19));
    layer0_outputs(3163) <= not(inputs(89));
    layer0_outputs(3164) <= inputs(110);
    layer0_outputs(3165) <= not(inputs(205));
    layer0_outputs(3166) <= not((inputs(126)) or (inputs(187)));
    layer0_outputs(3167) <= (inputs(208)) xor (inputs(241));
    layer0_outputs(3168) <= not(inputs(254)) or (inputs(160));
    layer0_outputs(3169) <= not(inputs(59));
    layer0_outputs(3170) <= (inputs(118)) and not (inputs(186));
    layer0_outputs(3171) <= (inputs(195)) or (inputs(204));
    layer0_outputs(3172) <= not((inputs(23)) or (inputs(95)));
    layer0_outputs(3173) <= not(inputs(55));
    layer0_outputs(3174) <= (inputs(201)) xor (inputs(74));
    layer0_outputs(3175) <= not(inputs(247));
    layer0_outputs(3176) <= (inputs(104)) xor (inputs(27));
    layer0_outputs(3177) <= not((inputs(166)) xor (inputs(233)));
    layer0_outputs(3178) <= (inputs(9)) and not (inputs(247));
    layer0_outputs(3179) <= (inputs(101)) and not (inputs(108));
    layer0_outputs(3180) <= not(inputs(92)) or (inputs(224));
    layer0_outputs(3181) <= not((inputs(245)) or (inputs(32)));
    layer0_outputs(3182) <= (inputs(65)) and (inputs(159));
    layer0_outputs(3183) <= (inputs(231)) and not (inputs(238));
    layer0_outputs(3184) <= inputs(245);
    layer0_outputs(3185) <= not((inputs(242)) or (inputs(26)));
    layer0_outputs(3186) <= inputs(85);
    layer0_outputs(3187) <= not(inputs(75));
    layer0_outputs(3188) <= not((inputs(43)) xor (inputs(201)));
    layer0_outputs(3189) <= (inputs(29)) xor (inputs(62));
    layer0_outputs(3190) <= not((inputs(126)) or (inputs(162)));
    layer0_outputs(3191) <= inputs(24);
    layer0_outputs(3192) <= not(inputs(71)) or (inputs(223));
    layer0_outputs(3193) <= not(inputs(240));
    layer0_outputs(3194) <= not((inputs(239)) or (inputs(51)));
    layer0_outputs(3195) <= inputs(230);
    layer0_outputs(3196) <= (inputs(153)) or (inputs(180));
    layer0_outputs(3197) <= not(inputs(121));
    layer0_outputs(3198) <= (inputs(77)) and not (inputs(184));
    layer0_outputs(3199) <= not(inputs(189));
    layer0_outputs(3200) <= inputs(139);
    layer0_outputs(3201) <= inputs(59);
    layer0_outputs(3202) <= not((inputs(167)) xor (inputs(37)));
    layer0_outputs(3203) <= (inputs(242)) or (inputs(122));
    layer0_outputs(3204) <= (inputs(159)) xor (inputs(71));
    layer0_outputs(3205) <= not(inputs(150));
    layer0_outputs(3206) <= not(inputs(22));
    layer0_outputs(3207) <= not((inputs(254)) or (inputs(49)));
    layer0_outputs(3208) <= not(inputs(151)) or (inputs(208));
    layer0_outputs(3209) <= (inputs(21)) and not (inputs(203));
    layer0_outputs(3210) <= (inputs(138)) and (inputs(153));
    layer0_outputs(3211) <= not((inputs(215)) and (inputs(3)));
    layer0_outputs(3212) <= not(inputs(46));
    layer0_outputs(3213) <= (inputs(217)) xor (inputs(201));
    layer0_outputs(3214) <= inputs(177);
    layer0_outputs(3215) <= (inputs(168)) or (inputs(136));
    layer0_outputs(3216) <= not(inputs(232));
    layer0_outputs(3217) <= inputs(63);
    layer0_outputs(3218) <= not((inputs(14)) or (inputs(70)));
    layer0_outputs(3219) <= (inputs(182)) and not (inputs(140));
    layer0_outputs(3220) <= inputs(163);
    layer0_outputs(3221) <= (inputs(167)) and not (inputs(239));
    layer0_outputs(3222) <= (inputs(121)) and not (inputs(159));
    layer0_outputs(3223) <= not((inputs(129)) or (inputs(114)));
    layer0_outputs(3224) <= '0';
    layer0_outputs(3225) <= not((inputs(255)) or (inputs(252)));
    layer0_outputs(3226) <= not(inputs(182));
    layer0_outputs(3227) <= not((inputs(47)) or (inputs(156)));
    layer0_outputs(3228) <= inputs(93);
    layer0_outputs(3229) <= not((inputs(116)) or (inputs(18)));
    layer0_outputs(3230) <= not(inputs(115));
    layer0_outputs(3231) <= not(inputs(122));
    layer0_outputs(3232) <= not((inputs(80)) or (inputs(227)));
    layer0_outputs(3233) <= inputs(76);
    layer0_outputs(3234) <= not(inputs(54));
    layer0_outputs(3235) <= not(inputs(96));
    layer0_outputs(3236) <= inputs(130);
    layer0_outputs(3237) <= not(inputs(32));
    layer0_outputs(3238) <= (inputs(234)) xor (inputs(53));
    layer0_outputs(3239) <= not((inputs(84)) or (inputs(131)));
    layer0_outputs(3240) <= not((inputs(12)) xor (inputs(76)));
    layer0_outputs(3241) <= (inputs(69)) and not (inputs(166));
    layer0_outputs(3242) <= inputs(203);
    layer0_outputs(3243) <= (inputs(144)) or (inputs(217));
    layer0_outputs(3244) <= not((inputs(176)) xor (inputs(22)));
    layer0_outputs(3245) <= not((inputs(86)) or (inputs(69)));
    layer0_outputs(3246) <= (inputs(86)) or (inputs(214));
    layer0_outputs(3247) <= (inputs(36)) or (inputs(176));
    layer0_outputs(3248) <= inputs(246);
    layer0_outputs(3249) <= not(inputs(84));
    layer0_outputs(3250) <= not(inputs(155));
    layer0_outputs(3251) <= (inputs(154)) xor (inputs(169));
    layer0_outputs(3252) <= not(inputs(106));
    layer0_outputs(3253) <= not((inputs(80)) xor (inputs(68)));
    layer0_outputs(3254) <= inputs(69);
    layer0_outputs(3255) <= not((inputs(96)) or (inputs(249)));
    layer0_outputs(3256) <= '0';
    layer0_outputs(3257) <= not(inputs(135)) or (inputs(65));
    layer0_outputs(3258) <= not(inputs(133));
    layer0_outputs(3259) <= not(inputs(199)) or (inputs(47));
    layer0_outputs(3260) <= not(inputs(117)) or (inputs(93));
    layer0_outputs(3261) <= not((inputs(76)) or (inputs(90)));
    layer0_outputs(3262) <= not(inputs(51));
    layer0_outputs(3263) <= not(inputs(206)) or (inputs(132));
    layer0_outputs(3264) <= '0';
    layer0_outputs(3265) <= not(inputs(82)) or (inputs(129));
    layer0_outputs(3266) <= not((inputs(179)) xor (inputs(254)));
    layer0_outputs(3267) <= (inputs(171)) and not (inputs(247));
    layer0_outputs(3268) <= not(inputs(201)) or (inputs(55));
    layer0_outputs(3269) <= not((inputs(61)) or (inputs(2)));
    layer0_outputs(3270) <= not(inputs(183)) or (inputs(198));
    layer0_outputs(3271) <= (inputs(66)) or (inputs(207));
    layer0_outputs(3272) <= (inputs(68)) and not (inputs(145));
    layer0_outputs(3273) <= not(inputs(165));
    layer0_outputs(3274) <= inputs(132);
    layer0_outputs(3275) <= inputs(44);
    layer0_outputs(3276) <= not(inputs(219)) or (inputs(35));
    layer0_outputs(3277) <= not((inputs(207)) xor (inputs(172)));
    layer0_outputs(3278) <= not(inputs(22));
    layer0_outputs(3279) <= inputs(109);
    layer0_outputs(3280) <= not((inputs(187)) or (inputs(222)));
    layer0_outputs(3281) <= not((inputs(55)) or (inputs(67)));
    layer0_outputs(3282) <= inputs(6);
    layer0_outputs(3283) <= (inputs(201)) and not (inputs(192));
    layer0_outputs(3284) <= (inputs(72)) and not (inputs(75));
    layer0_outputs(3285) <= inputs(232);
    layer0_outputs(3286) <= (inputs(150)) and (inputs(243));
    layer0_outputs(3287) <= not((inputs(16)) or (inputs(135)));
    layer0_outputs(3288) <= (inputs(56)) or (inputs(3));
    layer0_outputs(3289) <= inputs(21);
    layer0_outputs(3290) <= not(inputs(229)) or (inputs(62));
    layer0_outputs(3291) <= inputs(41);
    layer0_outputs(3292) <= (inputs(105)) and not (inputs(125));
    layer0_outputs(3293) <= (inputs(213)) and not (inputs(79));
    layer0_outputs(3294) <= inputs(181);
    layer0_outputs(3295) <= inputs(109);
    layer0_outputs(3296) <= not((inputs(224)) or (inputs(151)));
    layer0_outputs(3297) <= not(inputs(74)) or (inputs(210));
    layer0_outputs(3298) <= (inputs(105)) and not (inputs(19));
    layer0_outputs(3299) <= (inputs(132)) or (inputs(143));
    layer0_outputs(3300) <= (inputs(5)) xor (inputs(191));
    layer0_outputs(3301) <= (inputs(103)) or (inputs(110));
    layer0_outputs(3302) <= inputs(180);
    layer0_outputs(3303) <= not((inputs(77)) xor (inputs(45)));
    layer0_outputs(3304) <= not(inputs(203));
    layer0_outputs(3305) <= not(inputs(106)) or (inputs(141));
    layer0_outputs(3306) <= not((inputs(182)) or (inputs(131)));
    layer0_outputs(3307) <= not(inputs(88));
    layer0_outputs(3308) <= inputs(194);
    layer0_outputs(3309) <= inputs(249);
    layer0_outputs(3310) <= (inputs(145)) or (inputs(239));
    layer0_outputs(3311) <= inputs(246);
    layer0_outputs(3312) <= (inputs(13)) and not (inputs(161));
    layer0_outputs(3313) <= (inputs(243)) and (inputs(106));
    layer0_outputs(3314) <= inputs(70);
    layer0_outputs(3315) <= (inputs(86)) xor (inputs(70));
    layer0_outputs(3316) <= not((inputs(192)) or (inputs(122)));
    layer0_outputs(3317) <= not((inputs(223)) xor (inputs(150)));
    layer0_outputs(3318) <= not(inputs(103)) or (inputs(59));
    layer0_outputs(3319) <= '1';
    layer0_outputs(3320) <= not(inputs(187)) or (inputs(72));
    layer0_outputs(3321) <= not(inputs(193));
    layer0_outputs(3322) <= not(inputs(119));
    layer0_outputs(3323) <= (inputs(103)) and not (inputs(83));
    layer0_outputs(3324) <= (inputs(41)) and not (inputs(28));
    layer0_outputs(3325) <= inputs(233);
    layer0_outputs(3326) <= (inputs(171)) or (inputs(179));
    layer0_outputs(3327) <= not((inputs(190)) or (inputs(199)));
    layer0_outputs(3328) <= inputs(189);
    layer0_outputs(3329) <= (inputs(90)) or (inputs(165));
    layer0_outputs(3330) <= inputs(170);
    layer0_outputs(3331) <= not(inputs(139));
    layer0_outputs(3332) <= (inputs(120)) or (inputs(212));
    layer0_outputs(3333) <= inputs(89);
    layer0_outputs(3334) <= (inputs(87)) and not (inputs(49));
    layer0_outputs(3335) <= (inputs(168)) and (inputs(152));
    layer0_outputs(3336) <= inputs(210);
    layer0_outputs(3337) <= not(inputs(120));
    layer0_outputs(3338) <= not((inputs(174)) or (inputs(180)));
    layer0_outputs(3339) <= (inputs(205)) and not (inputs(98));
    layer0_outputs(3340) <= not(inputs(166));
    layer0_outputs(3341) <= inputs(40);
    layer0_outputs(3342) <= (inputs(4)) or (inputs(33));
    layer0_outputs(3343) <= not(inputs(150));
    layer0_outputs(3344) <= inputs(240);
    layer0_outputs(3345) <= not(inputs(40)) or (inputs(13));
    layer0_outputs(3346) <= not(inputs(129));
    layer0_outputs(3347) <= not(inputs(216));
    layer0_outputs(3348) <= inputs(135);
    layer0_outputs(3349) <= inputs(51);
    layer0_outputs(3350) <= inputs(52);
    layer0_outputs(3351) <= (inputs(114)) xor (inputs(89));
    layer0_outputs(3352) <= inputs(104);
    layer0_outputs(3353) <= not(inputs(138));
    layer0_outputs(3354) <= (inputs(117)) and (inputs(246));
    layer0_outputs(3355) <= (inputs(148)) and (inputs(132));
    layer0_outputs(3356) <= '0';
    layer0_outputs(3357) <= inputs(138);
    layer0_outputs(3358) <= (inputs(229)) or (inputs(55));
    layer0_outputs(3359) <= (inputs(58)) or (inputs(18));
    layer0_outputs(3360) <= not(inputs(130));
    layer0_outputs(3361) <= '1';
    layer0_outputs(3362) <= inputs(101);
    layer0_outputs(3363) <= not((inputs(102)) or (inputs(11)));
    layer0_outputs(3364) <= (inputs(58)) or (inputs(158));
    layer0_outputs(3365) <= inputs(203);
    layer0_outputs(3366) <= not((inputs(54)) or (inputs(53)));
    layer0_outputs(3367) <= inputs(183);
    layer0_outputs(3368) <= (inputs(124)) and not (inputs(194));
    layer0_outputs(3369) <= inputs(93);
    layer0_outputs(3370) <= not(inputs(24)) or (inputs(32));
    layer0_outputs(3371) <= inputs(226);
    layer0_outputs(3372) <= inputs(198);
    layer0_outputs(3373) <= not(inputs(247)) or (inputs(192));
    layer0_outputs(3374) <= not(inputs(29));
    layer0_outputs(3375) <= inputs(35);
    layer0_outputs(3376) <= (inputs(0)) and (inputs(164));
    layer0_outputs(3377) <= (inputs(195)) or (inputs(57));
    layer0_outputs(3378) <= inputs(217);
    layer0_outputs(3379) <= not(inputs(106)) or (inputs(100));
    layer0_outputs(3380) <= inputs(220);
    layer0_outputs(3381) <= inputs(249);
    layer0_outputs(3382) <= (inputs(220)) or (inputs(217));
    layer0_outputs(3383) <= not(inputs(192)) or (inputs(143));
    layer0_outputs(3384) <= (inputs(204)) and not (inputs(234));
    layer0_outputs(3385) <= inputs(157);
    layer0_outputs(3386) <= not(inputs(217)) or (inputs(136));
    layer0_outputs(3387) <= (inputs(210)) xor (inputs(112));
    layer0_outputs(3388) <= not((inputs(223)) xor (inputs(140)));
    layer0_outputs(3389) <= inputs(43);
    layer0_outputs(3390) <= (inputs(155)) or (inputs(107));
    layer0_outputs(3391) <= (inputs(206)) and (inputs(35));
    layer0_outputs(3392) <= not((inputs(224)) xor (inputs(201)));
    layer0_outputs(3393) <= '0';
    layer0_outputs(3394) <= not((inputs(232)) or (inputs(31)));
    layer0_outputs(3395) <= inputs(86);
    layer0_outputs(3396) <= not((inputs(242)) xor (inputs(227)));
    layer0_outputs(3397) <= (inputs(189)) or (inputs(65));
    layer0_outputs(3398) <= not((inputs(173)) or (inputs(197)));
    layer0_outputs(3399) <= not((inputs(252)) or (inputs(254)));
    layer0_outputs(3400) <= inputs(159);
    layer0_outputs(3401) <= not((inputs(252)) xor (inputs(37)));
    layer0_outputs(3402) <= not((inputs(168)) xor (inputs(168)));
    layer0_outputs(3403) <= inputs(123);
    layer0_outputs(3404) <= (inputs(251)) xor (inputs(171));
    layer0_outputs(3405) <= not(inputs(213)) or (inputs(11));
    layer0_outputs(3406) <= (inputs(151)) and not (inputs(242));
    layer0_outputs(3407) <= not(inputs(250));
    layer0_outputs(3408) <= not(inputs(21));
    layer0_outputs(3409) <= not((inputs(170)) or (inputs(142)));
    layer0_outputs(3410) <= inputs(187);
    layer0_outputs(3411) <= inputs(164);
    layer0_outputs(3412) <= '1';
    layer0_outputs(3413) <= not((inputs(71)) xor (inputs(25)));
    layer0_outputs(3414) <= not(inputs(178));
    layer0_outputs(3415) <= (inputs(218)) or (inputs(157));
    layer0_outputs(3416) <= not(inputs(205)) or (inputs(108));
    layer0_outputs(3417) <= (inputs(106)) and not (inputs(173));
    layer0_outputs(3418) <= (inputs(183)) or (inputs(82));
    layer0_outputs(3419) <= not((inputs(99)) or (inputs(88)));
    layer0_outputs(3420) <= inputs(90);
    layer0_outputs(3421) <= not((inputs(7)) or (inputs(95)));
    layer0_outputs(3422) <= inputs(114);
    layer0_outputs(3423) <= not(inputs(121));
    layer0_outputs(3424) <= not(inputs(37)) or (inputs(45));
    layer0_outputs(3425) <= not(inputs(159)) or (inputs(240));
    layer0_outputs(3426) <= not(inputs(105)) or (inputs(40));
    layer0_outputs(3427) <= (inputs(118)) or (inputs(211));
    layer0_outputs(3428) <= (inputs(212)) and not (inputs(53));
    layer0_outputs(3429) <= (inputs(169)) or (inputs(189));
    layer0_outputs(3430) <= (inputs(246)) or (inputs(220));
    layer0_outputs(3431) <= inputs(156);
    layer0_outputs(3432) <= inputs(165);
    layer0_outputs(3433) <= not((inputs(5)) xor (inputs(69)));
    layer0_outputs(3434) <= not((inputs(223)) or (inputs(148)));
    layer0_outputs(3435) <= not((inputs(172)) or (inputs(171)));
    layer0_outputs(3436) <= (inputs(179)) or (inputs(108));
    layer0_outputs(3437) <= not(inputs(237));
    layer0_outputs(3438) <= not(inputs(168));
    layer0_outputs(3439) <= (inputs(106)) xor (inputs(129));
    layer0_outputs(3440) <= not((inputs(160)) or (inputs(245)));
    layer0_outputs(3441) <= not(inputs(224)) or (inputs(157));
    layer0_outputs(3442) <= not(inputs(110));
    layer0_outputs(3443) <= inputs(26);
    layer0_outputs(3444) <= not((inputs(66)) or (inputs(9)));
    layer0_outputs(3445) <= not((inputs(190)) or (inputs(32)));
    layer0_outputs(3446) <= not((inputs(110)) xor (inputs(33)));
    layer0_outputs(3447) <= not((inputs(248)) or (inputs(190)));
    layer0_outputs(3448) <= not((inputs(190)) or (inputs(194)));
    layer0_outputs(3449) <= not((inputs(157)) and (inputs(173)));
    layer0_outputs(3450) <= not((inputs(126)) or (inputs(211)));
    layer0_outputs(3451) <= (inputs(103)) or (inputs(207));
    layer0_outputs(3452) <= not((inputs(69)) and (inputs(26)));
    layer0_outputs(3453) <= not(inputs(26));
    layer0_outputs(3454) <= not(inputs(180)) or (inputs(59));
    layer0_outputs(3455) <= not(inputs(98));
    layer0_outputs(3456) <= not((inputs(38)) xor (inputs(143)));
    layer0_outputs(3457) <= not(inputs(114)) or (inputs(5));
    layer0_outputs(3458) <= not(inputs(24));
    layer0_outputs(3459) <= (inputs(6)) and not (inputs(158));
    layer0_outputs(3460) <= (inputs(80)) xor (inputs(251));
    layer0_outputs(3461) <= (inputs(228)) and (inputs(231));
    layer0_outputs(3462) <= not(inputs(217));
    layer0_outputs(3463) <= not(inputs(216)) or (inputs(255));
    layer0_outputs(3464) <= not(inputs(231)) or (inputs(33));
    layer0_outputs(3465) <= not(inputs(109));
    layer0_outputs(3466) <= not(inputs(243));
    layer0_outputs(3467) <= not(inputs(193)) or (inputs(109));
    layer0_outputs(3468) <= not((inputs(167)) xor (inputs(95)));
    layer0_outputs(3469) <= (inputs(46)) or (inputs(204));
    layer0_outputs(3470) <= inputs(166);
    layer0_outputs(3471) <= (inputs(138)) or (inputs(9));
    layer0_outputs(3472) <= not((inputs(179)) xor (inputs(192)));
    layer0_outputs(3473) <= (inputs(149)) and not (inputs(53));
    layer0_outputs(3474) <= (inputs(153)) or (inputs(65));
    layer0_outputs(3475) <= (inputs(59)) or (inputs(114));
    layer0_outputs(3476) <= inputs(100);
    layer0_outputs(3477) <= '1';
    layer0_outputs(3478) <= not(inputs(9));
    layer0_outputs(3479) <= (inputs(239)) and not (inputs(15));
    layer0_outputs(3480) <= not(inputs(218)) or (inputs(108));
    layer0_outputs(3481) <= (inputs(200)) or (inputs(216));
    layer0_outputs(3482) <= not(inputs(137)) or (inputs(49));
    layer0_outputs(3483) <= inputs(16);
    layer0_outputs(3484) <= not((inputs(70)) or (inputs(221)));
    layer0_outputs(3485) <= (inputs(204)) or (inputs(150));
    layer0_outputs(3486) <= not((inputs(116)) or (inputs(100)));
    layer0_outputs(3487) <= inputs(143);
    layer0_outputs(3488) <= (inputs(128)) or (inputs(113));
    layer0_outputs(3489) <= (inputs(149)) and not (inputs(79));
    layer0_outputs(3490) <= not((inputs(58)) or (inputs(211)));
    layer0_outputs(3491) <= (inputs(148)) and not (inputs(20));
    layer0_outputs(3492) <= (inputs(164)) and not (inputs(240));
    layer0_outputs(3493) <= not((inputs(223)) or (inputs(54)));
    layer0_outputs(3494) <= (inputs(127)) or (inputs(3));
    layer0_outputs(3495) <= (inputs(84)) and not (inputs(194));
    layer0_outputs(3496) <= not(inputs(233)) or (inputs(45));
    layer0_outputs(3497) <= (inputs(54)) or (inputs(175));
    layer0_outputs(3498) <= not(inputs(198)) or (inputs(209));
    layer0_outputs(3499) <= (inputs(74)) or (inputs(254));
    layer0_outputs(3500) <= not(inputs(196)) or (inputs(175));
    layer0_outputs(3501) <= not(inputs(208)) or (inputs(5));
    layer0_outputs(3502) <= (inputs(50)) or (inputs(118));
    layer0_outputs(3503) <= (inputs(168)) or (inputs(69));
    layer0_outputs(3504) <= not(inputs(40));
    layer0_outputs(3505) <= not(inputs(212));
    layer0_outputs(3506) <= (inputs(138)) and not (inputs(114));
    layer0_outputs(3507) <= not((inputs(112)) or (inputs(44)));
    layer0_outputs(3508) <= not(inputs(44)) or (inputs(208));
    layer0_outputs(3509) <= not((inputs(75)) xor (inputs(149)));
    layer0_outputs(3510) <= not(inputs(210)) or (inputs(2));
    layer0_outputs(3511) <= not(inputs(167)) or (inputs(21));
    layer0_outputs(3512) <= (inputs(178)) and not (inputs(48));
    layer0_outputs(3513) <= not(inputs(79));
    layer0_outputs(3514) <= inputs(9);
    layer0_outputs(3515) <= (inputs(108)) or (inputs(126));
    layer0_outputs(3516) <= (inputs(246)) or (inputs(194));
    layer0_outputs(3517) <= (inputs(220)) or (inputs(238));
    layer0_outputs(3518) <= '0';
    layer0_outputs(3519) <= not(inputs(163));
    layer0_outputs(3520) <= inputs(77);
    layer0_outputs(3521) <= not((inputs(191)) or (inputs(156)));
    layer0_outputs(3522) <= inputs(129);
    layer0_outputs(3523) <= not(inputs(13)) or (inputs(252));
    layer0_outputs(3524) <= not(inputs(90)) or (inputs(40));
    layer0_outputs(3525) <= not((inputs(98)) or (inputs(93)));
    layer0_outputs(3526) <= inputs(148);
    layer0_outputs(3527) <= not(inputs(217)) or (inputs(120));
    layer0_outputs(3528) <= not((inputs(218)) and (inputs(165)));
    layer0_outputs(3529) <= (inputs(166)) and not (inputs(83));
    layer0_outputs(3530) <= (inputs(16)) or (inputs(183));
    layer0_outputs(3531) <= (inputs(170)) or (inputs(37));
    layer0_outputs(3532) <= not((inputs(109)) or (inputs(122)));
    layer0_outputs(3533) <= (inputs(139)) and not (inputs(162));
    layer0_outputs(3534) <= (inputs(43)) or (inputs(96));
    layer0_outputs(3535) <= '1';
    layer0_outputs(3536) <= not(inputs(224)) or (inputs(0));
    layer0_outputs(3537) <= not(inputs(30));
    layer0_outputs(3538) <= not(inputs(21));
    layer0_outputs(3539) <= not((inputs(75)) or (inputs(80)));
    layer0_outputs(3540) <= not(inputs(233));
    layer0_outputs(3541) <= inputs(116);
    layer0_outputs(3542) <= (inputs(74)) or (inputs(3));
    layer0_outputs(3543) <= (inputs(188)) and not (inputs(15));
    layer0_outputs(3544) <= (inputs(136)) or (inputs(242));
    layer0_outputs(3545) <= (inputs(6)) xor (inputs(219));
    layer0_outputs(3546) <= (inputs(245)) or (inputs(183));
    layer0_outputs(3547) <= not(inputs(206));
    layer0_outputs(3548) <= '0';
    layer0_outputs(3549) <= not(inputs(177)) or (inputs(203));
    layer0_outputs(3550) <= (inputs(116)) or (inputs(86));
    layer0_outputs(3551) <= inputs(140);
    layer0_outputs(3552) <= inputs(216);
    layer0_outputs(3553) <= inputs(20);
    layer0_outputs(3554) <= not((inputs(209)) or (inputs(25)));
    layer0_outputs(3555) <= not((inputs(121)) xor (inputs(154)));
    layer0_outputs(3556) <= not(inputs(47)) or (inputs(188));
    layer0_outputs(3557) <= (inputs(129)) or (inputs(198));
    layer0_outputs(3558) <= (inputs(182)) and not (inputs(112));
    layer0_outputs(3559) <= not((inputs(196)) and (inputs(193)));
    layer0_outputs(3560) <= inputs(35);
    layer0_outputs(3561) <= not((inputs(186)) xor (inputs(189)));
    layer0_outputs(3562) <= inputs(156);
    layer0_outputs(3563) <= (inputs(8)) and not (inputs(129));
    layer0_outputs(3564) <= not(inputs(214)) or (inputs(47));
    layer0_outputs(3565) <= inputs(115);
    layer0_outputs(3566) <= (inputs(104)) and not (inputs(160));
    layer0_outputs(3567) <= not((inputs(185)) xor (inputs(220)));
    layer0_outputs(3568) <= not(inputs(22));
    layer0_outputs(3569) <= not((inputs(33)) or (inputs(1)));
    layer0_outputs(3570) <= (inputs(213)) and not (inputs(3));
    layer0_outputs(3571) <= not(inputs(67));
    layer0_outputs(3572) <= inputs(162);
    layer0_outputs(3573) <= not(inputs(56)) or (inputs(9));
    layer0_outputs(3574) <= not(inputs(212));
    layer0_outputs(3575) <= (inputs(113)) or (inputs(210));
    layer0_outputs(3576) <= (inputs(35)) or (inputs(84));
    layer0_outputs(3577) <= (inputs(172)) and not (inputs(237));
    layer0_outputs(3578) <= inputs(234);
    layer0_outputs(3579) <= not(inputs(167)) or (inputs(17));
    layer0_outputs(3580) <= '0';
    layer0_outputs(3581) <= not(inputs(206));
    layer0_outputs(3582) <= not(inputs(196)) or (inputs(97));
    layer0_outputs(3583) <= (inputs(52)) or (inputs(91));
    layer0_outputs(3584) <= (inputs(110)) and not (inputs(63));
    layer0_outputs(3585) <= not((inputs(47)) or (inputs(100)));
    layer0_outputs(3586) <= inputs(139);
    layer0_outputs(3587) <= (inputs(249)) or (inputs(24));
    layer0_outputs(3588) <= inputs(146);
    layer0_outputs(3589) <= inputs(173);
    layer0_outputs(3590) <= not(inputs(103)) or (inputs(112));
    layer0_outputs(3591) <= (inputs(190)) xor (inputs(157));
    layer0_outputs(3592) <= not(inputs(219));
    layer0_outputs(3593) <= not(inputs(133));
    layer0_outputs(3594) <= not((inputs(177)) xor (inputs(233)));
    layer0_outputs(3595) <= inputs(194);
    layer0_outputs(3596) <= (inputs(38)) and not (inputs(16));
    layer0_outputs(3597) <= inputs(3);
    layer0_outputs(3598) <= (inputs(243)) or (inputs(175));
    layer0_outputs(3599) <= inputs(209);
    layer0_outputs(3600) <= inputs(83);
    layer0_outputs(3601) <= not(inputs(113));
    layer0_outputs(3602) <= not(inputs(183));
    layer0_outputs(3603) <= inputs(212);
    layer0_outputs(3604) <= inputs(182);
    layer0_outputs(3605) <= not(inputs(145));
    layer0_outputs(3606) <= (inputs(117)) or (inputs(31));
    layer0_outputs(3607) <= (inputs(8)) or (inputs(77));
    layer0_outputs(3608) <= not(inputs(3));
    layer0_outputs(3609) <= (inputs(8)) or (inputs(61));
    layer0_outputs(3610) <= (inputs(10)) and not (inputs(248));
    layer0_outputs(3611) <= not(inputs(42));
    layer0_outputs(3612) <= not(inputs(152));
    layer0_outputs(3613) <= not(inputs(68)) or (inputs(108));
    layer0_outputs(3614) <= not((inputs(200)) xor (inputs(180)));
    layer0_outputs(3615) <= inputs(207);
    layer0_outputs(3616) <= not((inputs(113)) or (inputs(107)));
    layer0_outputs(3617) <= inputs(196);
    layer0_outputs(3618) <= (inputs(235)) or (inputs(208));
    layer0_outputs(3619) <= (inputs(5)) xor (inputs(9));
    layer0_outputs(3620) <= inputs(180);
    layer0_outputs(3621) <= inputs(173);
    layer0_outputs(3622) <= not((inputs(7)) or (inputs(46)));
    layer0_outputs(3623) <= (inputs(178)) and not (inputs(130));
    layer0_outputs(3624) <= not((inputs(0)) and (inputs(94)));
    layer0_outputs(3625) <= not((inputs(205)) and (inputs(186)));
    layer0_outputs(3626) <= (inputs(17)) or (inputs(237));
    layer0_outputs(3627) <= (inputs(128)) or (inputs(125));
    layer0_outputs(3628) <= not(inputs(188)) or (inputs(49));
    layer0_outputs(3629) <= inputs(136);
    layer0_outputs(3630) <= inputs(217);
    layer0_outputs(3631) <= not((inputs(53)) or (inputs(57)));
    layer0_outputs(3632) <= (inputs(123)) and not (inputs(13));
    layer0_outputs(3633) <= '0';
    layer0_outputs(3634) <= inputs(91);
    layer0_outputs(3635) <= not(inputs(195)) or (inputs(166));
    layer0_outputs(3636) <= not((inputs(15)) or (inputs(136)));
    layer0_outputs(3637) <= inputs(92);
    layer0_outputs(3638) <= not(inputs(89)) or (inputs(30));
    layer0_outputs(3639) <= inputs(18);
    layer0_outputs(3640) <= (inputs(61)) and not (inputs(141));
    layer0_outputs(3641) <= not(inputs(22)) or (inputs(179));
    layer0_outputs(3642) <= (inputs(161)) or (inputs(46));
    layer0_outputs(3643) <= (inputs(110)) or (inputs(227));
    layer0_outputs(3644) <= not(inputs(200));
    layer0_outputs(3645) <= not(inputs(105));
    layer0_outputs(3646) <= (inputs(199)) or (inputs(239));
    layer0_outputs(3647) <= inputs(225);
    layer0_outputs(3648) <= '0';
    layer0_outputs(3649) <= (inputs(184)) and not (inputs(243));
    layer0_outputs(3650) <= not((inputs(52)) or (inputs(46)));
    layer0_outputs(3651) <= inputs(201);
    layer0_outputs(3652) <= not((inputs(238)) or (inputs(25)));
    layer0_outputs(3653) <= (inputs(247)) and not (inputs(199));
    layer0_outputs(3654) <= not(inputs(143));
    layer0_outputs(3655) <= inputs(182);
    layer0_outputs(3656) <= inputs(185);
    layer0_outputs(3657) <= inputs(103);
    layer0_outputs(3658) <= not(inputs(111)) or (inputs(214));
    layer0_outputs(3659) <= not((inputs(148)) xor (inputs(51)));
    layer0_outputs(3660) <= not((inputs(132)) or (inputs(86)));
    layer0_outputs(3661) <= not(inputs(198));
    layer0_outputs(3662) <= inputs(90);
    layer0_outputs(3663) <= not((inputs(43)) or (inputs(249)));
    layer0_outputs(3664) <= not(inputs(217)) or (inputs(77));
    layer0_outputs(3665) <= not(inputs(28)) or (inputs(209));
    layer0_outputs(3666) <= not(inputs(164));
    layer0_outputs(3667) <= '1';
    layer0_outputs(3668) <= (inputs(80)) or (inputs(243));
    layer0_outputs(3669) <= (inputs(129)) xor (inputs(118));
    layer0_outputs(3670) <= (inputs(104)) and not (inputs(224));
    layer0_outputs(3671) <= not((inputs(29)) or (inputs(79)));
    layer0_outputs(3672) <= (inputs(175)) or (inputs(176));
    layer0_outputs(3673) <= not((inputs(202)) or (inputs(96)));
    layer0_outputs(3674) <= not(inputs(130)) or (inputs(35));
    layer0_outputs(3675) <= (inputs(143)) or (inputs(234));
    layer0_outputs(3676) <= inputs(237);
    layer0_outputs(3677) <= inputs(77);
    layer0_outputs(3678) <= (inputs(205)) or (inputs(161));
    layer0_outputs(3679) <= not((inputs(240)) or (inputs(56)));
    layer0_outputs(3680) <= '1';
    layer0_outputs(3681) <= (inputs(19)) and not (inputs(236));
    layer0_outputs(3682) <= not(inputs(212));
    layer0_outputs(3683) <= (inputs(189)) or (inputs(186));
    layer0_outputs(3684) <= not((inputs(49)) and (inputs(195)));
    layer0_outputs(3685) <= (inputs(26)) and not (inputs(142));
    layer0_outputs(3686) <= not(inputs(235)) or (inputs(254));
    layer0_outputs(3687) <= (inputs(174)) or (inputs(216));
    layer0_outputs(3688) <= not((inputs(30)) or (inputs(190)));
    layer0_outputs(3689) <= not(inputs(130));
    layer0_outputs(3690) <= inputs(189);
    layer0_outputs(3691) <= (inputs(19)) and not (inputs(44));
    layer0_outputs(3692) <= not((inputs(177)) or (inputs(67)));
    layer0_outputs(3693) <= not(inputs(35));
    layer0_outputs(3694) <= (inputs(10)) and not (inputs(86));
    layer0_outputs(3695) <= not(inputs(181));
    layer0_outputs(3696) <= not(inputs(67));
    layer0_outputs(3697) <= (inputs(122)) or (inputs(145));
    layer0_outputs(3698) <= not(inputs(198)) or (inputs(82));
    layer0_outputs(3699) <= (inputs(247)) or (inputs(225));
    layer0_outputs(3700) <= (inputs(92)) or (inputs(188));
    layer0_outputs(3701) <= not((inputs(108)) or (inputs(199)));
    layer0_outputs(3702) <= not((inputs(95)) and (inputs(123)));
    layer0_outputs(3703) <= not(inputs(239)) or (inputs(13));
    layer0_outputs(3704) <= not((inputs(11)) xor (inputs(176)));
    layer0_outputs(3705) <= inputs(166);
    layer0_outputs(3706) <= not(inputs(93));
    layer0_outputs(3707) <= not(inputs(17));
    layer0_outputs(3708) <= '1';
    layer0_outputs(3709) <= not((inputs(237)) and (inputs(225)));
    layer0_outputs(3710) <= not((inputs(67)) or (inputs(59)));
    layer0_outputs(3711) <= inputs(110);
    layer0_outputs(3712) <= not(inputs(182));
    layer0_outputs(3713) <= not((inputs(158)) or (inputs(16)));
    layer0_outputs(3714) <= not((inputs(171)) and (inputs(50)));
    layer0_outputs(3715) <= inputs(218);
    layer0_outputs(3716) <= (inputs(246)) xor (inputs(63));
    layer0_outputs(3717) <= not((inputs(143)) or (inputs(254)));
    layer0_outputs(3718) <= not(inputs(227));
    layer0_outputs(3719) <= inputs(8);
    layer0_outputs(3720) <= not(inputs(21));
    layer0_outputs(3721) <= (inputs(245)) and not (inputs(19));
    layer0_outputs(3722) <= '1';
    layer0_outputs(3723) <= inputs(165);
    layer0_outputs(3724) <= not((inputs(247)) or (inputs(27)));
    layer0_outputs(3725) <= '0';
    layer0_outputs(3726) <= (inputs(244)) or (inputs(103));
    layer0_outputs(3727) <= not((inputs(9)) or (inputs(232)));
    layer0_outputs(3728) <= (inputs(209)) or (inputs(120));
    layer0_outputs(3729) <= not((inputs(162)) or (inputs(104)));
    layer0_outputs(3730) <= not(inputs(97));
    layer0_outputs(3731) <= not((inputs(117)) or (inputs(214)));
    layer0_outputs(3732) <= not((inputs(243)) or (inputs(78)));
    layer0_outputs(3733) <= not((inputs(13)) or (inputs(153)));
    layer0_outputs(3734) <= not((inputs(202)) xor (inputs(33)));
    layer0_outputs(3735) <= not(inputs(23)) or (inputs(14));
    layer0_outputs(3736) <= (inputs(41)) or (inputs(143));
    layer0_outputs(3737) <= not((inputs(238)) or (inputs(122)));
    layer0_outputs(3738) <= inputs(204);
    layer0_outputs(3739) <= not(inputs(85)) or (inputs(1));
    layer0_outputs(3740) <= not(inputs(87)) or (inputs(33));
    layer0_outputs(3741) <= not(inputs(57)) or (inputs(188));
    layer0_outputs(3742) <= not(inputs(153));
    layer0_outputs(3743) <= inputs(69);
    layer0_outputs(3744) <= not(inputs(228)) or (inputs(107));
    layer0_outputs(3745) <= not(inputs(148));
    layer0_outputs(3746) <= not(inputs(120)) or (inputs(115));
    layer0_outputs(3747) <= not((inputs(166)) or (inputs(30)));
    layer0_outputs(3748) <= inputs(214);
    layer0_outputs(3749) <= not((inputs(233)) xor (inputs(186)));
    layer0_outputs(3750) <= inputs(149);
    layer0_outputs(3751) <= inputs(61);
    layer0_outputs(3752) <= not((inputs(50)) or (inputs(145)));
    layer0_outputs(3753) <= not((inputs(30)) xor (inputs(145)));
    layer0_outputs(3754) <= (inputs(27)) and not (inputs(219));
    layer0_outputs(3755) <= (inputs(68)) or (inputs(54));
    layer0_outputs(3756) <= inputs(188);
    layer0_outputs(3757) <= inputs(219);
    layer0_outputs(3758) <= not(inputs(26));
    layer0_outputs(3759) <= (inputs(89)) and not (inputs(81));
    layer0_outputs(3760) <= not(inputs(240));
    layer0_outputs(3761) <= not((inputs(178)) xor (inputs(8)));
    layer0_outputs(3762) <= (inputs(108)) and not (inputs(209));
    layer0_outputs(3763) <= inputs(232);
    layer0_outputs(3764) <= (inputs(80)) and (inputs(52));
    layer0_outputs(3765) <= not(inputs(204)) or (inputs(129));
    layer0_outputs(3766) <= not(inputs(209)) or (inputs(20));
    layer0_outputs(3767) <= not(inputs(73));
    layer0_outputs(3768) <= (inputs(177)) or (inputs(145));
    layer0_outputs(3769) <= (inputs(43)) xor (inputs(74));
    layer0_outputs(3770) <= not((inputs(150)) and (inputs(197)));
    layer0_outputs(3771) <= (inputs(218)) or (inputs(151));
    layer0_outputs(3772) <= not(inputs(73));
    layer0_outputs(3773) <= not(inputs(24)) or (inputs(82));
    layer0_outputs(3774) <= inputs(112);
    layer0_outputs(3775) <= not((inputs(58)) or (inputs(205)));
    layer0_outputs(3776) <= not(inputs(162));
    layer0_outputs(3777) <= not((inputs(98)) xor (inputs(70)));
    layer0_outputs(3778) <= inputs(149);
    layer0_outputs(3779) <= not(inputs(238));
    layer0_outputs(3780) <= inputs(231);
    layer0_outputs(3781) <= not((inputs(52)) xor (inputs(231)));
    layer0_outputs(3782) <= inputs(183);
    layer0_outputs(3783) <= inputs(122);
    layer0_outputs(3784) <= inputs(95);
    layer0_outputs(3785) <= (inputs(114)) and not (inputs(253));
    layer0_outputs(3786) <= not((inputs(139)) xor (inputs(235)));
    layer0_outputs(3787) <= not(inputs(92));
    layer0_outputs(3788) <= (inputs(212)) or (inputs(190));
    layer0_outputs(3789) <= not(inputs(235));
    layer0_outputs(3790) <= not(inputs(126));
    layer0_outputs(3791) <= not((inputs(21)) or (inputs(14)));
    layer0_outputs(3792) <= not(inputs(155));
    layer0_outputs(3793) <= (inputs(212)) or (inputs(7));
    layer0_outputs(3794) <= not(inputs(152));
    layer0_outputs(3795) <= not((inputs(17)) or (inputs(104)));
    layer0_outputs(3796) <= not(inputs(109)) or (inputs(191));
    layer0_outputs(3797) <= inputs(84);
    layer0_outputs(3798) <= inputs(25);
    layer0_outputs(3799) <= not((inputs(207)) or (inputs(70)));
    layer0_outputs(3800) <= not((inputs(90)) or (inputs(3)));
    layer0_outputs(3801) <= not(inputs(68));
    layer0_outputs(3802) <= (inputs(29)) xor (inputs(2));
    layer0_outputs(3803) <= not(inputs(199)) or (inputs(135));
    layer0_outputs(3804) <= not((inputs(41)) or (inputs(172)));
    layer0_outputs(3805) <= inputs(82);
    layer0_outputs(3806) <= not((inputs(203)) and (inputs(152)));
    layer0_outputs(3807) <= not(inputs(119));
    layer0_outputs(3808) <= '0';
    layer0_outputs(3809) <= not(inputs(120)) or (inputs(248));
    layer0_outputs(3810) <= inputs(169);
    layer0_outputs(3811) <= not((inputs(192)) or (inputs(211)));
    layer0_outputs(3812) <= not(inputs(234)) or (inputs(74));
    layer0_outputs(3813) <= (inputs(37)) and not (inputs(161));
    layer0_outputs(3814) <= not((inputs(110)) or (inputs(114)));
    layer0_outputs(3815) <= not(inputs(115));
    layer0_outputs(3816) <= (inputs(80)) or (inputs(185));
    layer0_outputs(3817) <= inputs(68);
    layer0_outputs(3818) <= not(inputs(104));
    layer0_outputs(3819) <= (inputs(62)) xor (inputs(119));
    layer0_outputs(3820) <= not(inputs(112));
    layer0_outputs(3821) <= not(inputs(22));
    layer0_outputs(3822) <= not(inputs(143));
    layer0_outputs(3823) <= not(inputs(198));
    layer0_outputs(3824) <= (inputs(38)) xor (inputs(247));
    layer0_outputs(3825) <= inputs(242);
    layer0_outputs(3826) <= (inputs(12)) and not (inputs(111));
    layer0_outputs(3827) <= inputs(178);
    layer0_outputs(3828) <= (inputs(207)) xor (inputs(162));
    layer0_outputs(3829) <= (inputs(185)) or (inputs(76));
    layer0_outputs(3830) <= inputs(221);
    layer0_outputs(3831) <= not(inputs(93));
    layer0_outputs(3832) <= (inputs(255)) or (inputs(189));
    layer0_outputs(3833) <= inputs(27);
    layer0_outputs(3834) <= not(inputs(74));
    layer0_outputs(3835) <= inputs(91);
    layer0_outputs(3836) <= not(inputs(130));
    layer0_outputs(3837) <= (inputs(103)) and (inputs(135));
    layer0_outputs(3838) <= not(inputs(155)) or (inputs(18));
    layer0_outputs(3839) <= inputs(228);
    layer0_outputs(3840) <= (inputs(70)) xor (inputs(172));
    layer0_outputs(3841) <= not(inputs(115));
    layer0_outputs(3842) <= not((inputs(134)) or (inputs(87)));
    layer0_outputs(3843) <= not(inputs(197));
    layer0_outputs(3844) <= not(inputs(209));
    layer0_outputs(3845) <= inputs(77);
    layer0_outputs(3846) <= (inputs(246)) or (inputs(174));
    layer0_outputs(3847) <= not(inputs(29));
    layer0_outputs(3848) <= not((inputs(234)) or (inputs(236)));
    layer0_outputs(3849) <= not(inputs(135)) or (inputs(2));
    layer0_outputs(3850) <= not((inputs(212)) or (inputs(177)));
    layer0_outputs(3851) <= (inputs(228)) and not (inputs(0));
    layer0_outputs(3852) <= (inputs(111)) or (inputs(40));
    layer0_outputs(3853) <= inputs(147);
    layer0_outputs(3854) <= (inputs(61)) and not (inputs(155));
    layer0_outputs(3855) <= inputs(225);
    layer0_outputs(3856) <= inputs(232);
    layer0_outputs(3857) <= not((inputs(156)) xor (inputs(137)));
    layer0_outputs(3858) <= (inputs(6)) and not (inputs(109));
    layer0_outputs(3859) <= (inputs(87)) and not (inputs(206));
    layer0_outputs(3860) <= (inputs(188)) xor (inputs(168));
    layer0_outputs(3861) <= not(inputs(102)) or (inputs(110));
    layer0_outputs(3862) <= (inputs(123)) or (inputs(59));
    layer0_outputs(3863) <= inputs(37);
    layer0_outputs(3864) <= not(inputs(178));
    layer0_outputs(3865) <= not(inputs(7));
    layer0_outputs(3866) <= (inputs(253)) and not (inputs(158));
    layer0_outputs(3867) <= not(inputs(34)) or (inputs(97));
    layer0_outputs(3868) <= not(inputs(59));
    layer0_outputs(3869) <= (inputs(124)) or (inputs(116));
    layer0_outputs(3870) <= inputs(90);
    layer0_outputs(3871) <= (inputs(226)) or (inputs(208));
    layer0_outputs(3872) <= not((inputs(139)) or (inputs(63)));
    layer0_outputs(3873) <= (inputs(119)) and not (inputs(177));
    layer0_outputs(3874) <= (inputs(48)) xor (inputs(19));
    layer0_outputs(3875) <= not(inputs(197));
    layer0_outputs(3876) <= (inputs(170)) xor (inputs(153));
    layer0_outputs(3877) <= not(inputs(84));
    layer0_outputs(3878) <= not((inputs(52)) or (inputs(126)));
    layer0_outputs(3879) <= inputs(99);
    layer0_outputs(3880) <= not((inputs(105)) xor (inputs(254)));
    layer0_outputs(3881) <= (inputs(240)) xor (inputs(107));
    layer0_outputs(3882) <= (inputs(8)) and not (inputs(230));
    layer0_outputs(3883) <= (inputs(158)) or (inputs(249));
    layer0_outputs(3884) <= not(inputs(75));
    layer0_outputs(3885) <= not((inputs(254)) and (inputs(50)));
    layer0_outputs(3886) <= not((inputs(222)) or (inputs(186)));
    layer0_outputs(3887) <= inputs(67);
    layer0_outputs(3888) <= (inputs(7)) and not (inputs(81));
    layer0_outputs(3889) <= not(inputs(228)) or (inputs(131));
    layer0_outputs(3890) <= not(inputs(8));
    layer0_outputs(3891) <= not(inputs(184)) or (inputs(97));
    layer0_outputs(3892) <= not(inputs(109));
    layer0_outputs(3893) <= inputs(151);
    layer0_outputs(3894) <= not((inputs(232)) xor (inputs(242)));
    layer0_outputs(3895) <= inputs(151);
    layer0_outputs(3896) <= (inputs(219)) xor (inputs(158));
    layer0_outputs(3897) <= (inputs(236)) or (inputs(131));
    layer0_outputs(3898) <= (inputs(41)) or (inputs(206));
    layer0_outputs(3899) <= (inputs(112)) and not (inputs(64));
    layer0_outputs(3900) <= (inputs(26)) or (inputs(99));
    layer0_outputs(3901) <= (inputs(174)) or (inputs(197));
    layer0_outputs(3902) <= not((inputs(94)) or (inputs(228)));
    layer0_outputs(3903) <= '0';
    layer0_outputs(3904) <= not(inputs(228));
    layer0_outputs(3905) <= not(inputs(95));
    layer0_outputs(3906) <= not(inputs(254));
    layer0_outputs(3907) <= not((inputs(33)) or (inputs(73)));
    layer0_outputs(3908) <= not(inputs(57));
    layer0_outputs(3909) <= (inputs(39)) xor (inputs(24));
    layer0_outputs(3910) <= (inputs(253)) or (inputs(94));
    layer0_outputs(3911) <= (inputs(119)) and not (inputs(241));
    layer0_outputs(3912) <= (inputs(25)) or (inputs(0));
    layer0_outputs(3913) <= inputs(226);
    layer0_outputs(3914) <= not((inputs(204)) or (inputs(194)));
    layer0_outputs(3915) <= (inputs(40)) or (inputs(1));
    layer0_outputs(3916) <= inputs(235);
    layer0_outputs(3917) <= not((inputs(51)) and (inputs(87)));
    layer0_outputs(3918) <= not((inputs(244)) xor (inputs(42)));
    layer0_outputs(3919) <= (inputs(65)) and (inputs(6));
    layer0_outputs(3920) <= inputs(102);
    layer0_outputs(3921) <= not(inputs(136)) or (inputs(30));
    layer0_outputs(3922) <= (inputs(5)) xor (inputs(79));
    layer0_outputs(3923) <= not(inputs(123)) or (inputs(184));
    layer0_outputs(3924) <= not((inputs(205)) or (inputs(92)));
    layer0_outputs(3925) <= (inputs(141)) or (inputs(145));
    layer0_outputs(3926) <= (inputs(127)) or (inputs(157));
    layer0_outputs(3927) <= not(inputs(119));
    layer0_outputs(3928) <= not(inputs(91)) or (inputs(32));
    layer0_outputs(3929) <= not(inputs(207)) or (inputs(142));
    layer0_outputs(3930) <= (inputs(224)) or (inputs(26));
    layer0_outputs(3931) <= not((inputs(214)) or (inputs(192)));
    layer0_outputs(3932) <= not((inputs(96)) xor (inputs(147)));
    layer0_outputs(3933) <= not(inputs(200)) or (inputs(63));
    layer0_outputs(3934) <= (inputs(177)) xor (inputs(248));
    layer0_outputs(3935) <= not((inputs(122)) or (inputs(155)));
    layer0_outputs(3936) <= not((inputs(196)) or (inputs(37)));
    layer0_outputs(3937) <= (inputs(111)) or (inputs(62));
    layer0_outputs(3938) <= inputs(147);
    layer0_outputs(3939) <= inputs(52);
    layer0_outputs(3940) <= (inputs(166)) and (inputs(141));
    layer0_outputs(3941) <= '0';
    layer0_outputs(3942) <= not((inputs(135)) and (inputs(233)));
    layer0_outputs(3943) <= not(inputs(115));
    layer0_outputs(3944) <= not(inputs(36));
    layer0_outputs(3945) <= (inputs(146)) or (inputs(219));
    layer0_outputs(3946) <= not(inputs(111)) or (inputs(1));
    layer0_outputs(3947) <= (inputs(195)) or (inputs(38));
    layer0_outputs(3948) <= not(inputs(114));
    layer0_outputs(3949) <= (inputs(25)) and not (inputs(225));
    layer0_outputs(3950) <= not((inputs(112)) and (inputs(158)));
    layer0_outputs(3951) <= not(inputs(108)) or (inputs(222));
    layer0_outputs(3952) <= not(inputs(238));
    layer0_outputs(3953) <= (inputs(25)) or (inputs(16));
    layer0_outputs(3954) <= not(inputs(49));
    layer0_outputs(3955) <= (inputs(226)) or (inputs(80));
    layer0_outputs(3956) <= not(inputs(238));
    layer0_outputs(3957) <= not((inputs(224)) xor (inputs(160)));
    layer0_outputs(3958) <= not(inputs(79));
    layer0_outputs(3959) <= (inputs(131)) or (inputs(55));
    layer0_outputs(3960) <= not(inputs(29)) or (inputs(138));
    layer0_outputs(3961) <= (inputs(200)) xor (inputs(44));
    layer0_outputs(3962) <= (inputs(125)) or (inputs(92));
    layer0_outputs(3963) <= not((inputs(54)) and (inputs(171)));
    layer0_outputs(3964) <= (inputs(83)) or (inputs(170));
    layer0_outputs(3965) <= not(inputs(190));
    layer0_outputs(3966) <= (inputs(195)) and (inputs(168));
    layer0_outputs(3967) <= not(inputs(124)) or (inputs(30));
    layer0_outputs(3968) <= (inputs(117)) and not (inputs(39));
    layer0_outputs(3969) <= (inputs(231)) and not (inputs(145));
    layer0_outputs(3970) <= not(inputs(52));
    layer0_outputs(3971) <= inputs(190);
    layer0_outputs(3972) <= not((inputs(47)) or (inputs(223)));
    layer0_outputs(3973) <= (inputs(174)) and not (inputs(243));
    layer0_outputs(3974) <= not(inputs(133));
    layer0_outputs(3975) <= (inputs(41)) or (inputs(189));
    layer0_outputs(3976) <= not((inputs(32)) or (inputs(213)));
    layer0_outputs(3977) <= not((inputs(21)) or (inputs(95)));
    layer0_outputs(3978) <= not((inputs(205)) or (inputs(159)));
    layer0_outputs(3979) <= not(inputs(86));
    layer0_outputs(3980) <= (inputs(210)) or (inputs(87));
    layer0_outputs(3981) <= (inputs(63)) or (inputs(0));
    layer0_outputs(3982) <= not(inputs(75)) or (inputs(251));
    layer0_outputs(3983) <= not((inputs(120)) xor (inputs(89)));
    layer0_outputs(3984) <= not(inputs(148));
    layer0_outputs(3985) <= (inputs(5)) or (inputs(47));
    layer0_outputs(3986) <= (inputs(115)) or (inputs(113));
    layer0_outputs(3987) <= not(inputs(122));
    layer0_outputs(3988) <= not(inputs(230)) or (inputs(156));
    layer0_outputs(3989) <= (inputs(152)) or (inputs(81));
    layer0_outputs(3990) <= '0';
    layer0_outputs(3991) <= (inputs(203)) xor (inputs(188));
    layer0_outputs(3992) <= not(inputs(25));
    layer0_outputs(3993) <= not((inputs(62)) xor (inputs(126)));
    layer0_outputs(3994) <= not((inputs(81)) or (inputs(10)));
    layer0_outputs(3995) <= not(inputs(132)) or (inputs(142));
    layer0_outputs(3996) <= not((inputs(193)) or (inputs(178)));
    layer0_outputs(3997) <= inputs(65);
    layer0_outputs(3998) <= not((inputs(116)) xor (inputs(152)));
    layer0_outputs(3999) <= not(inputs(91));
    layer0_outputs(4000) <= not(inputs(177));
    layer0_outputs(4001) <= inputs(96);
    layer0_outputs(4002) <= not((inputs(250)) and (inputs(51)));
    layer0_outputs(4003) <= (inputs(33)) or (inputs(37));
    layer0_outputs(4004) <= (inputs(65)) or (inputs(195));
    layer0_outputs(4005) <= inputs(50);
    layer0_outputs(4006) <= (inputs(80)) xor (inputs(90));
    layer0_outputs(4007) <= inputs(235);
    layer0_outputs(4008) <= not((inputs(176)) xor (inputs(225)));
    layer0_outputs(4009) <= (inputs(130)) and (inputs(125));
    layer0_outputs(4010) <= not((inputs(186)) or (inputs(217)));
    layer0_outputs(4011) <= not(inputs(132)) or (inputs(1));
    layer0_outputs(4012) <= '0';
    layer0_outputs(4013) <= (inputs(249)) xor (inputs(178));
    layer0_outputs(4014) <= not(inputs(85));
    layer0_outputs(4015) <= inputs(181);
    layer0_outputs(4016) <= inputs(76);
    layer0_outputs(4017) <= not((inputs(186)) or (inputs(201)));
    layer0_outputs(4018) <= '0';
    layer0_outputs(4019) <= inputs(47);
    layer0_outputs(4020) <= not((inputs(10)) or (inputs(223)));
    layer0_outputs(4021) <= (inputs(43)) or (inputs(125));
    layer0_outputs(4022) <= not((inputs(107)) or (inputs(176)));
    layer0_outputs(4023) <= not(inputs(58)) or (inputs(15));
    layer0_outputs(4024) <= inputs(195);
    layer0_outputs(4025) <= not(inputs(118));
    layer0_outputs(4026) <= (inputs(83)) and not (inputs(78));
    layer0_outputs(4027) <= (inputs(132)) or (inputs(193));
    layer0_outputs(4028) <= inputs(146);
    layer0_outputs(4029) <= (inputs(149)) and (inputs(167));
    layer0_outputs(4030) <= (inputs(39)) and not (inputs(155));
    layer0_outputs(4031) <= not(inputs(52));
    layer0_outputs(4032) <= not(inputs(220)) or (inputs(109));
    layer0_outputs(4033) <= inputs(218);
    layer0_outputs(4034) <= inputs(89);
    layer0_outputs(4035) <= not(inputs(230)) or (inputs(50));
    layer0_outputs(4036) <= (inputs(98)) and not (inputs(65));
    layer0_outputs(4037) <= not(inputs(91));
    layer0_outputs(4038) <= not((inputs(170)) and (inputs(135)));
    layer0_outputs(4039) <= (inputs(118)) and not (inputs(201));
    layer0_outputs(4040) <= inputs(238);
    layer0_outputs(4041) <= not((inputs(203)) and (inputs(148)));
    layer0_outputs(4042) <= not((inputs(235)) or (inputs(156)));
    layer0_outputs(4043) <= (inputs(249)) or (inputs(189));
    layer0_outputs(4044) <= (inputs(182)) and not (inputs(208));
    layer0_outputs(4045) <= (inputs(144)) or (inputs(1));
    layer0_outputs(4046) <= not(inputs(187));
    layer0_outputs(4047) <= not((inputs(255)) or (inputs(79)));
    layer0_outputs(4048) <= inputs(98);
    layer0_outputs(4049) <= not(inputs(172));
    layer0_outputs(4050) <= inputs(195);
    layer0_outputs(4051) <= (inputs(232)) or (inputs(71));
    layer0_outputs(4052) <= (inputs(222)) or (inputs(136));
    layer0_outputs(4053) <= (inputs(221)) or (inputs(251));
    layer0_outputs(4054) <= not(inputs(101)) or (inputs(62));
    layer0_outputs(4055) <= not(inputs(210));
    layer0_outputs(4056) <= not(inputs(230));
    layer0_outputs(4057) <= not(inputs(151));
    layer0_outputs(4058) <= not((inputs(27)) or (inputs(122)));
    layer0_outputs(4059) <= not(inputs(60)) or (inputs(178));
    layer0_outputs(4060) <= not(inputs(84));
    layer0_outputs(4061) <= not(inputs(113));
    layer0_outputs(4062) <= (inputs(225)) or (inputs(109));
    layer0_outputs(4063) <= not(inputs(183)) or (inputs(96));
    layer0_outputs(4064) <= not((inputs(245)) xor (inputs(244)));
    layer0_outputs(4065) <= not(inputs(10));
    layer0_outputs(4066) <= (inputs(99)) and not (inputs(45));
    layer0_outputs(4067) <= not((inputs(33)) or (inputs(236)));
    layer0_outputs(4068) <= (inputs(116)) and (inputs(1));
    layer0_outputs(4069) <= not((inputs(234)) xor (inputs(50)));
    layer0_outputs(4070) <= (inputs(64)) or (inputs(144));
    layer0_outputs(4071) <= inputs(180);
    layer0_outputs(4072) <= not(inputs(39));
    layer0_outputs(4073) <= not((inputs(191)) or (inputs(103)));
    layer0_outputs(4074) <= inputs(175);
    layer0_outputs(4075) <= inputs(116);
    layer0_outputs(4076) <= not(inputs(94)) or (inputs(175));
    layer0_outputs(4077) <= not(inputs(84));
    layer0_outputs(4078) <= inputs(214);
    layer0_outputs(4079) <= (inputs(160)) or (inputs(247));
    layer0_outputs(4080) <= inputs(66);
    layer0_outputs(4081) <= inputs(245);
    layer0_outputs(4082) <= (inputs(165)) xor (inputs(103));
    layer0_outputs(4083) <= not(inputs(149));
    layer0_outputs(4084) <= not(inputs(193));
    layer0_outputs(4085) <= not(inputs(165));
    layer0_outputs(4086) <= not((inputs(14)) or (inputs(78)));
    layer0_outputs(4087) <= not((inputs(124)) or (inputs(255)));
    layer0_outputs(4088) <= not(inputs(43)) or (inputs(228));
    layer0_outputs(4089) <= not((inputs(110)) or (inputs(182)));
    layer0_outputs(4090) <= (inputs(129)) and (inputs(129));
    layer0_outputs(4091) <= (inputs(81)) or (inputs(4));
    layer0_outputs(4092) <= (inputs(218)) or (inputs(193));
    layer0_outputs(4093) <= (inputs(98)) or (inputs(179));
    layer0_outputs(4094) <= (inputs(90)) and not (inputs(216));
    layer0_outputs(4095) <= (inputs(239)) xor (inputs(135));
    layer0_outputs(4096) <= not(inputs(134));
    layer0_outputs(4097) <= not(inputs(176));
    layer0_outputs(4098) <= inputs(78);
    layer0_outputs(4099) <= (inputs(120)) and not (inputs(252));
    layer0_outputs(4100) <= not(inputs(52)) or (inputs(213));
    layer0_outputs(4101) <= not(inputs(208));
    layer0_outputs(4102) <= inputs(200);
    layer0_outputs(4103) <= (inputs(51)) or (inputs(48));
    layer0_outputs(4104) <= not(inputs(23));
    layer0_outputs(4105) <= (inputs(93)) or (inputs(42));
    layer0_outputs(4106) <= not(inputs(23)) or (inputs(147));
    layer0_outputs(4107) <= not(inputs(58));
    layer0_outputs(4108) <= inputs(21);
    layer0_outputs(4109) <= not((inputs(48)) or (inputs(4)));
    layer0_outputs(4110) <= not((inputs(178)) xor (inputs(229)));
    layer0_outputs(4111) <= '1';
    layer0_outputs(4112) <= not(inputs(176)) or (inputs(111));
    layer0_outputs(4113) <= not((inputs(103)) or (inputs(77)));
    layer0_outputs(4114) <= (inputs(122)) or (inputs(221));
    layer0_outputs(4115) <= (inputs(17)) xor (inputs(84));
    layer0_outputs(4116) <= (inputs(220)) and not (inputs(72));
    layer0_outputs(4117) <= not((inputs(148)) and (inputs(23)));
    layer0_outputs(4118) <= (inputs(13)) and not (inputs(162));
    layer0_outputs(4119) <= not(inputs(213)) or (inputs(51));
    layer0_outputs(4120) <= (inputs(102)) and not (inputs(219));
    layer0_outputs(4121) <= not(inputs(31));
    layer0_outputs(4122) <= not((inputs(53)) xor (inputs(250)));
    layer0_outputs(4123) <= (inputs(149)) or (inputs(41));
    layer0_outputs(4124) <= (inputs(180)) and not (inputs(47));
    layer0_outputs(4125) <= (inputs(193)) or (inputs(151));
    layer0_outputs(4126) <= inputs(226);
    layer0_outputs(4127) <= not(inputs(70));
    layer0_outputs(4128) <= not((inputs(138)) or (inputs(194)));
    layer0_outputs(4129) <= not((inputs(131)) xor (inputs(100)));
    layer0_outputs(4130) <= inputs(89);
    layer0_outputs(4131) <= not(inputs(85));
    layer0_outputs(4132) <= not(inputs(248)) or (inputs(237));
    layer0_outputs(4133) <= not(inputs(200)) or (inputs(73));
    layer0_outputs(4134) <= inputs(94);
    layer0_outputs(4135) <= (inputs(249)) or (inputs(208));
    layer0_outputs(4136) <= (inputs(83)) and not (inputs(64));
    layer0_outputs(4137) <= inputs(217);
    layer0_outputs(4138) <= not(inputs(84)) or (inputs(111));
    layer0_outputs(4139) <= (inputs(68)) xor (inputs(143));
    layer0_outputs(4140) <= (inputs(74)) and not (inputs(204));
    layer0_outputs(4141) <= not((inputs(228)) or (inputs(207)));
    layer0_outputs(4142) <= not(inputs(74)) or (inputs(203));
    layer0_outputs(4143) <= inputs(133);
    layer0_outputs(4144) <= not(inputs(68)) or (inputs(147));
    layer0_outputs(4145) <= not((inputs(80)) or (inputs(193)));
    layer0_outputs(4146) <= not((inputs(150)) or (inputs(251)));
    layer0_outputs(4147) <= (inputs(69)) or (inputs(50));
    layer0_outputs(4148) <= not((inputs(224)) xor (inputs(135)));
    layer0_outputs(4149) <= not((inputs(186)) or (inputs(4)));
    layer0_outputs(4150) <= '1';
    layer0_outputs(4151) <= (inputs(169)) xor (inputs(185));
    layer0_outputs(4152) <= not(inputs(89));
    layer0_outputs(4153) <= not((inputs(227)) or (inputs(165)));
    layer0_outputs(4154) <= not(inputs(183));
    layer0_outputs(4155) <= not(inputs(6)) or (inputs(156));
    layer0_outputs(4156) <= not((inputs(4)) or (inputs(240)));
    layer0_outputs(4157) <= not(inputs(132)) or (inputs(206));
    layer0_outputs(4158) <= not((inputs(188)) xor (inputs(122)));
    layer0_outputs(4159) <= not((inputs(188)) and (inputs(228)));
    layer0_outputs(4160) <= not(inputs(58));
    layer0_outputs(4161) <= (inputs(77)) or (inputs(244));
    layer0_outputs(4162) <= (inputs(189)) or (inputs(214));
    layer0_outputs(4163) <= not(inputs(219)) or (inputs(37));
    layer0_outputs(4164) <= not(inputs(218)) or (inputs(49));
    layer0_outputs(4165) <= (inputs(226)) and not (inputs(131));
    layer0_outputs(4166) <= inputs(154);
    layer0_outputs(4167) <= not(inputs(97));
    layer0_outputs(4168) <= inputs(24);
    layer0_outputs(4169) <= inputs(204);
    layer0_outputs(4170) <= (inputs(182)) or (inputs(19));
    layer0_outputs(4171) <= (inputs(218)) xor (inputs(124));
    layer0_outputs(4172) <= (inputs(144)) or (inputs(247));
    layer0_outputs(4173) <= inputs(63);
    layer0_outputs(4174) <= not(inputs(242)) or (inputs(16));
    layer0_outputs(4175) <= not(inputs(28)) or (inputs(103));
    layer0_outputs(4176) <= (inputs(86)) xor (inputs(22));
    layer0_outputs(4177) <= not(inputs(62));
    layer0_outputs(4178) <= (inputs(39)) xor (inputs(2));
    layer0_outputs(4179) <= (inputs(2)) xor (inputs(216));
    layer0_outputs(4180) <= not(inputs(166));
    layer0_outputs(4181) <= not(inputs(252)) or (inputs(123));
    layer0_outputs(4182) <= not(inputs(197));
    layer0_outputs(4183) <= (inputs(169)) and (inputs(183));
    layer0_outputs(4184) <= '0';
    layer0_outputs(4185) <= inputs(90);
    layer0_outputs(4186) <= '0';
    layer0_outputs(4187) <= not(inputs(108)) or (inputs(45));
    layer0_outputs(4188) <= inputs(180);
    layer0_outputs(4189) <= not((inputs(16)) or (inputs(90)));
    layer0_outputs(4190) <= (inputs(12)) xor (inputs(94));
    layer0_outputs(4191) <= (inputs(165)) and not (inputs(81));
    layer0_outputs(4192) <= not((inputs(221)) and (inputs(253)));
    layer0_outputs(4193) <= not((inputs(65)) or (inputs(203)));
    layer0_outputs(4194) <= not(inputs(82));
    layer0_outputs(4195) <= not((inputs(117)) or (inputs(156)));
    layer0_outputs(4196) <= (inputs(125)) or (inputs(7));
    layer0_outputs(4197) <= not(inputs(144));
    layer0_outputs(4198) <= not(inputs(120)) or (inputs(255));
    layer0_outputs(4199) <= not((inputs(221)) or (inputs(135)));
    layer0_outputs(4200) <= not((inputs(172)) or (inputs(209)));
    layer0_outputs(4201) <= inputs(103);
    layer0_outputs(4202) <= not((inputs(109)) xor (inputs(176)));
    layer0_outputs(4203) <= not(inputs(5));
    layer0_outputs(4204) <= not(inputs(153)) or (inputs(28));
    layer0_outputs(4205) <= not((inputs(32)) or (inputs(20)));
    layer0_outputs(4206) <= inputs(154);
    layer0_outputs(4207) <= inputs(72);
    layer0_outputs(4208) <= inputs(70);
    layer0_outputs(4209) <= not(inputs(227)) or (inputs(121));
    layer0_outputs(4210) <= inputs(70);
    layer0_outputs(4211) <= '1';
    layer0_outputs(4212) <= not(inputs(130));
    layer0_outputs(4213) <= (inputs(46)) and not (inputs(91));
    layer0_outputs(4214) <= not(inputs(115)) or (inputs(43));
    layer0_outputs(4215) <= inputs(151);
    layer0_outputs(4216) <= inputs(23);
    layer0_outputs(4217) <= (inputs(48)) or (inputs(7));
    layer0_outputs(4218) <= (inputs(143)) or (inputs(34));
    layer0_outputs(4219) <= (inputs(129)) or (inputs(178));
    layer0_outputs(4220) <= (inputs(204)) and not (inputs(125));
    layer0_outputs(4221) <= not(inputs(167)) or (inputs(177));
    layer0_outputs(4222) <= (inputs(179)) and not (inputs(90));
    layer0_outputs(4223) <= not((inputs(6)) or (inputs(155)));
    layer0_outputs(4224) <= inputs(20);
    layer0_outputs(4225) <= (inputs(28)) and not (inputs(182));
    layer0_outputs(4226) <= not(inputs(212)) or (inputs(159));
    layer0_outputs(4227) <= not((inputs(103)) xor (inputs(196)));
    layer0_outputs(4228) <= not(inputs(144)) or (inputs(242));
    layer0_outputs(4229) <= inputs(228);
    layer0_outputs(4230) <= inputs(124);
    layer0_outputs(4231) <= (inputs(177)) and not (inputs(91));
    layer0_outputs(4232) <= (inputs(202)) xor (inputs(205));
    layer0_outputs(4233) <= not(inputs(177)) or (inputs(251));
    layer0_outputs(4234) <= not((inputs(169)) xor (inputs(166)));
    layer0_outputs(4235) <= inputs(30);
    layer0_outputs(4236) <= not(inputs(104));
    layer0_outputs(4237) <= (inputs(131)) xor (inputs(134));
    layer0_outputs(4238) <= not(inputs(69));
    layer0_outputs(4239) <= (inputs(95)) and not (inputs(48));
    layer0_outputs(4240) <= not((inputs(48)) or (inputs(9)));
    layer0_outputs(4241) <= not(inputs(51)) or (inputs(108));
    layer0_outputs(4242) <= not(inputs(21));
    layer0_outputs(4243) <= not(inputs(58));
    layer0_outputs(4244) <= inputs(95);
    layer0_outputs(4245) <= '1';
    layer0_outputs(4246) <= (inputs(101)) and (inputs(27));
    layer0_outputs(4247) <= not(inputs(22)) or (inputs(113));
    layer0_outputs(4248) <= not((inputs(191)) xor (inputs(198)));
    layer0_outputs(4249) <= not(inputs(233));
    layer0_outputs(4250) <= '0';
    layer0_outputs(4251) <= not(inputs(42));
    layer0_outputs(4252) <= not((inputs(64)) or (inputs(203)));
    layer0_outputs(4253) <= not(inputs(228));
    layer0_outputs(4254) <= not(inputs(21)) or (inputs(176));
    layer0_outputs(4255) <= not(inputs(143));
    layer0_outputs(4256) <= not(inputs(2));
    layer0_outputs(4257) <= '0';
    layer0_outputs(4258) <= '0';
    layer0_outputs(4259) <= inputs(144);
    layer0_outputs(4260) <= (inputs(40)) and (inputs(89));
    layer0_outputs(4261) <= (inputs(16)) xor (inputs(154));
    layer0_outputs(4262) <= (inputs(146)) xor (inputs(212));
    layer0_outputs(4263) <= not(inputs(29)) or (inputs(34));
    layer0_outputs(4264) <= not(inputs(182));
    layer0_outputs(4265) <= (inputs(205)) and not (inputs(109));
    layer0_outputs(4266) <= inputs(165);
    layer0_outputs(4267) <= (inputs(208)) and not (inputs(111));
    layer0_outputs(4268) <= inputs(125);
    layer0_outputs(4269) <= inputs(85);
    layer0_outputs(4270) <= not(inputs(85));
    layer0_outputs(4271) <= not(inputs(139)) or (inputs(224));
    layer0_outputs(4272) <= inputs(131);
    layer0_outputs(4273) <= not(inputs(173)) or (inputs(79));
    layer0_outputs(4274) <= (inputs(192)) or (inputs(236));
    layer0_outputs(4275) <= not(inputs(177));
    layer0_outputs(4276) <= not((inputs(200)) or (inputs(184)));
    layer0_outputs(4277) <= (inputs(67)) and not (inputs(0));
    layer0_outputs(4278) <= (inputs(118)) and not (inputs(221));
    layer0_outputs(4279) <= not(inputs(199)) or (inputs(216));
    layer0_outputs(4280) <= (inputs(28)) or (inputs(218));
    layer0_outputs(4281) <= (inputs(145)) or (inputs(44));
    layer0_outputs(4282) <= not((inputs(14)) or (inputs(80)));
    layer0_outputs(4283) <= not(inputs(24));
    layer0_outputs(4284) <= not(inputs(65));
    layer0_outputs(4285) <= inputs(181);
    layer0_outputs(4286) <= inputs(232);
    layer0_outputs(4287) <= (inputs(25)) and not (inputs(4));
    layer0_outputs(4288) <= inputs(232);
    layer0_outputs(4289) <= not(inputs(152)) or (inputs(170));
    layer0_outputs(4290) <= not(inputs(66));
    layer0_outputs(4291) <= inputs(247);
    layer0_outputs(4292) <= '1';
    layer0_outputs(4293) <= inputs(219);
    layer0_outputs(4294) <= inputs(231);
    layer0_outputs(4295) <= not((inputs(208)) and (inputs(251)));
    layer0_outputs(4296) <= (inputs(181)) or (inputs(32));
    layer0_outputs(4297) <= not(inputs(92)) or (inputs(248));
    layer0_outputs(4298) <= inputs(231);
    layer0_outputs(4299) <= '1';
    layer0_outputs(4300) <= (inputs(108)) and not (inputs(160));
    layer0_outputs(4301) <= not((inputs(142)) or (inputs(131)));
    layer0_outputs(4302) <= not(inputs(69));
    layer0_outputs(4303) <= not(inputs(133));
    layer0_outputs(4304) <= (inputs(215)) and not (inputs(43));
    layer0_outputs(4305) <= (inputs(242)) and not (inputs(128));
    layer0_outputs(4306) <= not(inputs(238));
    layer0_outputs(4307) <= not(inputs(2)) or (inputs(238));
    layer0_outputs(4308) <= (inputs(156)) and not (inputs(19));
    layer0_outputs(4309) <= (inputs(64)) or (inputs(204));
    layer0_outputs(4310) <= not(inputs(77));
    layer0_outputs(4311) <= not(inputs(8));
    layer0_outputs(4312) <= not((inputs(22)) xor (inputs(66)));
    layer0_outputs(4313) <= (inputs(66)) and not (inputs(158));
    layer0_outputs(4314) <= not((inputs(56)) xor (inputs(20)));
    layer0_outputs(4315) <= (inputs(31)) and (inputs(28));
    layer0_outputs(4316) <= not(inputs(254)) or (inputs(79));
    layer0_outputs(4317) <= not(inputs(123));
    layer0_outputs(4318) <= not(inputs(209));
    layer0_outputs(4319) <= not((inputs(37)) or (inputs(51)));
    layer0_outputs(4320) <= (inputs(85)) and not (inputs(127));
    layer0_outputs(4321) <= not((inputs(44)) or (inputs(42)));
    layer0_outputs(4322) <= (inputs(80)) or (inputs(232));
    layer0_outputs(4323) <= not(inputs(63)) or (inputs(13));
    layer0_outputs(4324) <= (inputs(52)) and not (inputs(207));
    layer0_outputs(4325) <= not((inputs(200)) or (inputs(224)));
    layer0_outputs(4326) <= not((inputs(16)) or (inputs(61)));
    layer0_outputs(4327) <= (inputs(136)) xor (inputs(239));
    layer0_outputs(4328) <= (inputs(71)) and (inputs(80));
    layer0_outputs(4329) <= not(inputs(184)) or (inputs(71));
    layer0_outputs(4330) <= inputs(90);
    layer0_outputs(4331) <= not(inputs(189));
    layer0_outputs(4332) <= inputs(57);
    layer0_outputs(4333) <= not(inputs(88)) or (inputs(96));
    layer0_outputs(4334) <= not(inputs(54)) or (inputs(1));
    layer0_outputs(4335) <= (inputs(154)) and not (inputs(5));
    layer0_outputs(4336) <= inputs(194);
    layer0_outputs(4337) <= not((inputs(191)) or (inputs(199)));
    layer0_outputs(4338) <= not((inputs(75)) or (inputs(175)));
    layer0_outputs(4339) <= not(inputs(29));
    layer0_outputs(4340) <= not((inputs(175)) or (inputs(227)));
    layer0_outputs(4341) <= not(inputs(116)) or (inputs(126));
    layer0_outputs(4342) <= not((inputs(61)) xor (inputs(141)));
    layer0_outputs(4343) <= (inputs(226)) or (inputs(241));
    layer0_outputs(4344) <= not((inputs(168)) and (inputs(22)));
    layer0_outputs(4345) <= not(inputs(69)) or (inputs(176));
    layer0_outputs(4346) <= not(inputs(120)) or (inputs(149));
    layer0_outputs(4347) <= (inputs(30)) or (inputs(11));
    layer0_outputs(4348) <= not(inputs(115)) or (inputs(48));
    layer0_outputs(4349) <= (inputs(210)) and not (inputs(35));
    layer0_outputs(4350) <= inputs(67);
    layer0_outputs(4351) <= inputs(228);
    layer0_outputs(4352) <= (inputs(164)) xor (inputs(114));
    layer0_outputs(4353) <= not(inputs(24));
    layer0_outputs(4354) <= (inputs(44)) and not (inputs(219));
    layer0_outputs(4355) <= (inputs(46)) and not (inputs(109));
    layer0_outputs(4356) <= (inputs(83)) or (inputs(47));
    layer0_outputs(4357) <= not(inputs(68)) or (inputs(1));
    layer0_outputs(4358) <= inputs(89);
    layer0_outputs(4359) <= not((inputs(185)) or (inputs(232)));
    layer0_outputs(4360) <= not((inputs(171)) xor (inputs(222)));
    layer0_outputs(4361) <= (inputs(123)) and (inputs(76));
    layer0_outputs(4362) <= not((inputs(6)) or (inputs(243)));
    layer0_outputs(4363) <= '0';
    layer0_outputs(4364) <= not((inputs(186)) or (inputs(2)));
    layer0_outputs(4365) <= (inputs(1)) or (inputs(254));
    layer0_outputs(4366) <= inputs(195);
    layer0_outputs(4367) <= (inputs(38)) and not (inputs(220));
    layer0_outputs(4368) <= (inputs(156)) xor (inputs(127));
    layer0_outputs(4369) <= not(inputs(131)) or (inputs(241));
    layer0_outputs(4370) <= inputs(91);
    layer0_outputs(4371) <= not(inputs(131));
    layer0_outputs(4372) <= not(inputs(151));
    layer0_outputs(4373) <= inputs(93);
    layer0_outputs(4374) <= not(inputs(181));
    layer0_outputs(4375) <= (inputs(48)) and (inputs(195));
    layer0_outputs(4376) <= (inputs(97)) and not (inputs(218));
    layer0_outputs(4377) <= not((inputs(228)) or (inputs(123)));
    layer0_outputs(4378) <= not(inputs(77));
    layer0_outputs(4379) <= '1';
    layer0_outputs(4380) <= not((inputs(218)) and (inputs(12)));
    layer0_outputs(4381) <= not((inputs(47)) xor (inputs(15)));
    layer0_outputs(4382) <= (inputs(160)) or (inputs(202));
    layer0_outputs(4383) <= not((inputs(179)) or (inputs(244)));
    layer0_outputs(4384) <= not(inputs(230));
    layer0_outputs(4385) <= not(inputs(32));
    layer0_outputs(4386) <= (inputs(97)) or (inputs(213));
    layer0_outputs(4387) <= inputs(90);
    layer0_outputs(4388) <= not(inputs(237));
    layer0_outputs(4389) <= not((inputs(161)) xor (inputs(111)));
    layer0_outputs(4390) <= not((inputs(4)) or (inputs(196)));
    layer0_outputs(4391) <= not(inputs(134)) or (inputs(155));
    layer0_outputs(4392) <= (inputs(246)) and not (inputs(114));
    layer0_outputs(4393) <= not((inputs(243)) or (inputs(209)));
    layer0_outputs(4394) <= not(inputs(212));
    layer0_outputs(4395) <= not((inputs(135)) xor (inputs(127)));
    layer0_outputs(4396) <= inputs(108);
    layer0_outputs(4397) <= inputs(118);
    layer0_outputs(4398) <= (inputs(154)) xor (inputs(199));
    layer0_outputs(4399) <= not((inputs(47)) xor (inputs(176)));
    layer0_outputs(4400) <= not((inputs(147)) or (inputs(150)));
    layer0_outputs(4401) <= inputs(229);
    layer0_outputs(4402) <= not((inputs(3)) xor (inputs(141)));
    layer0_outputs(4403) <= not(inputs(21)) or (inputs(42));
    layer0_outputs(4404) <= inputs(94);
    layer0_outputs(4405) <= (inputs(101)) or (inputs(133));
    layer0_outputs(4406) <= not(inputs(86));
    layer0_outputs(4407) <= '1';
    layer0_outputs(4408) <= inputs(36);
    layer0_outputs(4409) <= inputs(89);
    layer0_outputs(4410) <= not((inputs(131)) or (inputs(255)));
    layer0_outputs(4411) <= not((inputs(235)) xor (inputs(162)));
    layer0_outputs(4412) <= not(inputs(135));
    layer0_outputs(4413) <= (inputs(222)) xor (inputs(192));
    layer0_outputs(4414) <= not(inputs(190));
    layer0_outputs(4415) <= not(inputs(134)) or (inputs(188));
    layer0_outputs(4416) <= (inputs(77)) and not (inputs(96));
    layer0_outputs(4417) <= not(inputs(168));
    layer0_outputs(4418) <= not(inputs(164)) or (inputs(160));
    layer0_outputs(4419) <= (inputs(193)) and not (inputs(253));
    layer0_outputs(4420) <= (inputs(117)) xor (inputs(113));
    layer0_outputs(4421) <= (inputs(189)) and not (inputs(117));
    layer0_outputs(4422) <= not(inputs(119)) or (inputs(83));
    layer0_outputs(4423) <= not((inputs(4)) xor (inputs(125)));
    layer0_outputs(4424) <= not(inputs(230)) or (inputs(116));
    layer0_outputs(4425) <= not(inputs(48));
    layer0_outputs(4426) <= not(inputs(58)) or (inputs(173));
    layer0_outputs(4427) <= (inputs(243)) and not (inputs(150));
    layer0_outputs(4428) <= (inputs(83)) or (inputs(10));
    layer0_outputs(4429) <= (inputs(234)) xor (inputs(175));
    layer0_outputs(4430) <= (inputs(137)) and not (inputs(82));
    layer0_outputs(4431) <= (inputs(144)) or (inputs(202));
    layer0_outputs(4432) <= (inputs(226)) or (inputs(150));
    layer0_outputs(4433) <= not(inputs(44)) or (inputs(69));
    layer0_outputs(4434) <= (inputs(26)) and not (inputs(65));
    layer0_outputs(4435) <= not(inputs(35));
    layer0_outputs(4436) <= (inputs(76)) or (inputs(165));
    layer0_outputs(4437) <= (inputs(85)) and not (inputs(109));
    layer0_outputs(4438) <= not((inputs(134)) or (inputs(148)));
    layer0_outputs(4439) <= (inputs(167)) or (inputs(17));
    layer0_outputs(4440) <= inputs(126);
    layer0_outputs(4441) <= (inputs(24)) or (inputs(40));
    layer0_outputs(4442) <= not(inputs(205)) or (inputs(31));
    layer0_outputs(4443) <= not(inputs(153));
    layer0_outputs(4444) <= (inputs(116)) and not (inputs(14));
    layer0_outputs(4445) <= (inputs(128)) or (inputs(168));
    layer0_outputs(4446) <= (inputs(8)) or (inputs(194));
    layer0_outputs(4447) <= inputs(181);
    layer0_outputs(4448) <= inputs(193);
    layer0_outputs(4449) <= inputs(164);
    layer0_outputs(4450) <= not((inputs(211)) or (inputs(252)));
    layer0_outputs(4451) <= not((inputs(1)) or (inputs(160)));
    layer0_outputs(4452) <= (inputs(229)) and not (inputs(207));
    layer0_outputs(4453) <= (inputs(81)) and not (inputs(97));
    layer0_outputs(4454) <= inputs(129);
    layer0_outputs(4455) <= (inputs(134)) or (inputs(197));
    layer0_outputs(4456) <= not(inputs(196)) or (inputs(215));
    layer0_outputs(4457) <= not(inputs(92));
    layer0_outputs(4458) <= not(inputs(119)) or (inputs(63));
    layer0_outputs(4459) <= (inputs(52)) xor (inputs(99));
    layer0_outputs(4460) <= not(inputs(99)) or (inputs(46));
    layer0_outputs(4461) <= inputs(60);
    layer0_outputs(4462) <= (inputs(8)) and (inputs(8));
    layer0_outputs(4463) <= not(inputs(32));
    layer0_outputs(4464) <= (inputs(242)) or (inputs(20));
    layer0_outputs(4465) <= not(inputs(176)) or (inputs(108));
    layer0_outputs(4466) <= inputs(2);
    layer0_outputs(4467) <= not((inputs(11)) and (inputs(217)));
    layer0_outputs(4468) <= (inputs(154)) xor (inputs(34));
    layer0_outputs(4469) <= not(inputs(84)) or (inputs(142));
    layer0_outputs(4470) <= not(inputs(96));
    layer0_outputs(4471) <= inputs(214);
    layer0_outputs(4472) <= inputs(226);
    layer0_outputs(4473) <= not((inputs(212)) and (inputs(215)));
    layer0_outputs(4474) <= not(inputs(101));
    layer0_outputs(4475) <= not((inputs(81)) or (inputs(195)));
    layer0_outputs(4476) <= (inputs(47)) xor (inputs(7));
    layer0_outputs(4477) <= (inputs(170)) or (inputs(219));
    layer0_outputs(4478) <= not((inputs(154)) or (inputs(9)));
    layer0_outputs(4479) <= not(inputs(24));
    layer0_outputs(4480) <= inputs(83);
    layer0_outputs(4481) <= (inputs(88)) and not (inputs(223));
    layer0_outputs(4482) <= (inputs(59)) xor (inputs(177));
    layer0_outputs(4483) <= inputs(244);
    layer0_outputs(4484) <= not((inputs(172)) xor (inputs(32)));
    layer0_outputs(4485) <= not((inputs(172)) or (inputs(43)));
    layer0_outputs(4486) <= not(inputs(141)) or (inputs(255));
    layer0_outputs(4487) <= not((inputs(2)) or (inputs(61)));
    layer0_outputs(4488) <= not((inputs(220)) or (inputs(236)));
    layer0_outputs(4489) <= (inputs(83)) and not (inputs(191));
    layer0_outputs(4490) <= not(inputs(145));
    layer0_outputs(4491) <= not(inputs(152)) or (inputs(48));
    layer0_outputs(4492) <= '0';
    layer0_outputs(4493) <= (inputs(153)) xor (inputs(123));
    layer0_outputs(4494) <= inputs(123);
    layer0_outputs(4495) <= inputs(174);
    layer0_outputs(4496) <= not((inputs(187)) or (inputs(200)));
    layer0_outputs(4497) <= not(inputs(211)) or (inputs(182));
    layer0_outputs(4498) <= not((inputs(167)) or (inputs(150)));
    layer0_outputs(4499) <= (inputs(50)) and not (inputs(179));
    layer0_outputs(4500) <= not(inputs(196));
    layer0_outputs(4501) <= (inputs(18)) and not (inputs(113));
    layer0_outputs(4502) <= not(inputs(245));
    layer0_outputs(4503) <= '0';
    layer0_outputs(4504) <= not(inputs(121));
    layer0_outputs(4505) <= (inputs(132)) xor (inputs(128));
    layer0_outputs(4506) <= (inputs(125)) xor (inputs(158));
    layer0_outputs(4507) <= (inputs(111)) or (inputs(92));
    layer0_outputs(4508) <= not((inputs(157)) or (inputs(115)));
    layer0_outputs(4509) <= (inputs(229)) and not (inputs(156));
    layer0_outputs(4510) <= not(inputs(142)) or (inputs(18));
    layer0_outputs(4511) <= (inputs(212)) xor (inputs(209));
    layer0_outputs(4512) <= inputs(140);
    layer0_outputs(4513) <= not(inputs(21)) or (inputs(221));
    layer0_outputs(4514) <= (inputs(192)) or (inputs(141));
    layer0_outputs(4515) <= inputs(139);
    layer0_outputs(4516) <= (inputs(139)) or (inputs(77));
    layer0_outputs(4517) <= not((inputs(165)) or (inputs(85)));
    layer0_outputs(4518) <= not(inputs(108));
    layer0_outputs(4519) <= not((inputs(214)) or (inputs(114)));
    layer0_outputs(4520) <= not(inputs(248)) or (inputs(44));
    layer0_outputs(4521) <= (inputs(230)) and not (inputs(207));
    layer0_outputs(4522) <= not(inputs(146));
    layer0_outputs(4523) <= not(inputs(246));
    layer0_outputs(4524) <= inputs(216);
    layer0_outputs(4525) <= not((inputs(122)) or (inputs(94)));
    layer0_outputs(4526) <= inputs(14);
    layer0_outputs(4527) <= (inputs(37)) and not (inputs(54));
    layer0_outputs(4528) <= not(inputs(170)) or (inputs(240));
    layer0_outputs(4529) <= inputs(17);
    layer0_outputs(4530) <= (inputs(49)) or (inputs(185));
    layer0_outputs(4531) <= inputs(102);
    layer0_outputs(4532) <= not((inputs(47)) or (inputs(128)));
    layer0_outputs(4533) <= not((inputs(161)) xor (inputs(181)));
    layer0_outputs(4534) <= not(inputs(203)) or (inputs(160));
    layer0_outputs(4535) <= (inputs(60)) and not (inputs(255));
    layer0_outputs(4536) <= inputs(77);
    layer0_outputs(4537) <= not(inputs(231)) or (inputs(141));
    layer0_outputs(4538) <= not(inputs(125));
    layer0_outputs(4539) <= (inputs(136)) and not (inputs(238));
    layer0_outputs(4540) <= not(inputs(68));
    layer0_outputs(4541) <= not(inputs(8));
    layer0_outputs(4542) <= inputs(148);
    layer0_outputs(4543) <= not((inputs(232)) or (inputs(154)));
    layer0_outputs(4544) <= inputs(44);
    layer0_outputs(4545) <= not((inputs(47)) or (inputs(165)));
    layer0_outputs(4546) <= inputs(254);
    layer0_outputs(4547) <= (inputs(118)) and not (inputs(8));
    layer0_outputs(4548) <= not((inputs(15)) and (inputs(28)));
    layer0_outputs(4549) <= not(inputs(38)) or (inputs(226));
    layer0_outputs(4550) <= inputs(154);
    layer0_outputs(4551) <= (inputs(2)) and (inputs(21));
    layer0_outputs(4552) <= not((inputs(184)) xor (inputs(13)));
    layer0_outputs(4553) <= (inputs(84)) or (inputs(147));
    layer0_outputs(4554) <= not((inputs(214)) or (inputs(228)));
    layer0_outputs(4555) <= not(inputs(100)) or (inputs(10));
    layer0_outputs(4556) <= inputs(110);
    layer0_outputs(4557) <= not(inputs(146));
    layer0_outputs(4558) <= not(inputs(246));
    layer0_outputs(4559) <= not(inputs(82));
    layer0_outputs(4560) <= inputs(162);
    layer0_outputs(4561) <= not(inputs(78));
    layer0_outputs(4562) <= not(inputs(75));
    layer0_outputs(4563) <= not(inputs(102));
    layer0_outputs(4564) <= not(inputs(72)) or (inputs(44));
    layer0_outputs(4565) <= not((inputs(23)) xor (inputs(225)));
    layer0_outputs(4566) <= not(inputs(255)) or (inputs(14));
    layer0_outputs(4567) <= inputs(26);
    layer0_outputs(4568) <= not((inputs(210)) or (inputs(65)));
    layer0_outputs(4569) <= not(inputs(136)) or (inputs(249));
    layer0_outputs(4570) <= not((inputs(145)) or (inputs(230)));
    layer0_outputs(4571) <= inputs(59);
    layer0_outputs(4572) <= inputs(231);
    layer0_outputs(4573) <= not(inputs(28));
    layer0_outputs(4574) <= (inputs(42)) and not (inputs(191));
    layer0_outputs(4575) <= not(inputs(104));
    layer0_outputs(4576) <= not((inputs(101)) and (inputs(180)));
    layer0_outputs(4577) <= inputs(85);
    layer0_outputs(4578) <= (inputs(80)) or (inputs(192));
    layer0_outputs(4579) <= not(inputs(146)) or (inputs(1));
    layer0_outputs(4580) <= not(inputs(226));
    layer0_outputs(4581) <= (inputs(86)) xor (inputs(5));
    layer0_outputs(4582) <= inputs(120);
    layer0_outputs(4583) <= not((inputs(74)) or (inputs(74)));
    layer0_outputs(4584) <= (inputs(34)) and not (inputs(44));
    layer0_outputs(4585) <= inputs(164);
    layer0_outputs(4586) <= (inputs(25)) xor (inputs(245));
    layer0_outputs(4587) <= not(inputs(50));
    layer0_outputs(4588) <= not(inputs(81)) or (inputs(108));
    layer0_outputs(4589) <= inputs(199);
    layer0_outputs(4590) <= not((inputs(58)) or (inputs(175)));
    layer0_outputs(4591) <= not(inputs(128));
    layer0_outputs(4592) <= (inputs(85)) and not (inputs(220));
    layer0_outputs(4593) <= not(inputs(115));
    layer0_outputs(4594) <= (inputs(43)) and not (inputs(16));
    layer0_outputs(4595) <= not((inputs(133)) xor (inputs(158)));
    layer0_outputs(4596) <= (inputs(69)) and not (inputs(244));
    layer0_outputs(4597) <= not(inputs(138));
    layer0_outputs(4598) <= (inputs(76)) and not (inputs(14));
    layer0_outputs(4599) <= (inputs(41)) and (inputs(211));
    layer0_outputs(4600) <= not((inputs(36)) or (inputs(172)));
    layer0_outputs(4601) <= inputs(192);
    layer0_outputs(4602) <= not(inputs(135)) or (inputs(1));
    layer0_outputs(4603) <= inputs(146);
    layer0_outputs(4604) <= not((inputs(48)) or (inputs(172)));
    layer0_outputs(4605) <= (inputs(236)) and not (inputs(41));
    layer0_outputs(4606) <= not((inputs(53)) or (inputs(127)));
    layer0_outputs(4607) <= not((inputs(192)) xor (inputs(16)));
    layer0_outputs(4608) <= inputs(218);
    layer0_outputs(4609) <= inputs(131);
    layer0_outputs(4610) <= (inputs(133)) and (inputs(108));
    layer0_outputs(4611) <= (inputs(174)) and not (inputs(86));
    layer0_outputs(4612) <= not(inputs(82));
    layer0_outputs(4613) <= not(inputs(106));
    layer0_outputs(4614) <= inputs(181);
    layer0_outputs(4615) <= not(inputs(240));
    layer0_outputs(4616) <= (inputs(53)) or (inputs(54));
    layer0_outputs(4617) <= (inputs(77)) and (inputs(3));
    layer0_outputs(4618) <= inputs(101);
    layer0_outputs(4619) <= not(inputs(254));
    layer0_outputs(4620) <= inputs(80);
    layer0_outputs(4621) <= not(inputs(92)) or (inputs(255));
    layer0_outputs(4622) <= not((inputs(162)) or (inputs(179)));
    layer0_outputs(4623) <= not((inputs(206)) xor (inputs(226)));
    layer0_outputs(4624) <= '0';
    layer0_outputs(4625) <= inputs(215);
    layer0_outputs(4626) <= not(inputs(72));
    layer0_outputs(4627) <= not((inputs(8)) or (inputs(210)));
    layer0_outputs(4628) <= (inputs(203)) xor (inputs(237));
    layer0_outputs(4629) <= not((inputs(176)) xor (inputs(247)));
    layer0_outputs(4630) <= inputs(180);
    layer0_outputs(4631) <= inputs(146);
    layer0_outputs(4632) <= (inputs(245)) and not (inputs(255));
    layer0_outputs(4633) <= not((inputs(212)) xor (inputs(214)));
    layer0_outputs(4634) <= not(inputs(102));
    layer0_outputs(4635) <= not((inputs(2)) or (inputs(11)));
    layer0_outputs(4636) <= (inputs(13)) and not (inputs(77));
    layer0_outputs(4637) <= inputs(187);
    layer0_outputs(4638) <= not(inputs(176));
    layer0_outputs(4639) <= not((inputs(129)) xor (inputs(83)));
    layer0_outputs(4640) <= (inputs(192)) and not (inputs(17));
    layer0_outputs(4641) <= (inputs(7)) and not (inputs(12));
    layer0_outputs(4642) <= not(inputs(43));
    layer0_outputs(4643) <= inputs(124);
    layer0_outputs(4644) <= not((inputs(86)) or (inputs(174)));
    layer0_outputs(4645) <= not((inputs(127)) xor (inputs(71)));
    layer0_outputs(4646) <= (inputs(99)) and not (inputs(207));
    layer0_outputs(4647) <= not(inputs(228));
    layer0_outputs(4648) <= (inputs(52)) or (inputs(33));
    layer0_outputs(4649) <= (inputs(61)) or (inputs(65));
    layer0_outputs(4650) <= not((inputs(15)) or (inputs(0)));
    layer0_outputs(4651) <= (inputs(35)) and not (inputs(250));
    layer0_outputs(4652) <= (inputs(116)) xor (inputs(129));
    layer0_outputs(4653) <= (inputs(10)) xor (inputs(45));
    layer0_outputs(4654) <= inputs(28);
    layer0_outputs(4655) <= not((inputs(53)) and (inputs(55)));
    layer0_outputs(4656) <= not((inputs(21)) or (inputs(62)));
    layer0_outputs(4657) <= (inputs(70)) xor (inputs(18));
    layer0_outputs(4658) <= not((inputs(59)) and (inputs(23)));
    layer0_outputs(4659) <= not(inputs(84));
    layer0_outputs(4660) <= not(inputs(18));
    layer0_outputs(4661) <= not(inputs(221)) or (inputs(139));
    layer0_outputs(4662) <= not((inputs(209)) or (inputs(40)));
    layer0_outputs(4663) <= inputs(247);
    layer0_outputs(4664) <= inputs(128);
    layer0_outputs(4665) <= not(inputs(14));
    layer0_outputs(4666) <= (inputs(234)) and not (inputs(193));
    layer0_outputs(4667) <= inputs(186);
    layer0_outputs(4668) <= not((inputs(90)) xor (inputs(95)));
    layer0_outputs(4669) <= not(inputs(132)) or (inputs(78));
    layer0_outputs(4670) <= inputs(118);
    layer0_outputs(4671) <= (inputs(238)) or (inputs(108));
    layer0_outputs(4672) <= not(inputs(207));
    layer0_outputs(4673) <= (inputs(85)) and not (inputs(143));
    layer0_outputs(4674) <= not(inputs(250)) or (inputs(92));
    layer0_outputs(4675) <= not(inputs(186)) or (inputs(33));
    layer0_outputs(4676) <= (inputs(36)) or (inputs(236));
    layer0_outputs(4677) <= (inputs(194)) and not (inputs(55));
    layer0_outputs(4678) <= not((inputs(138)) or (inputs(102)));
    layer0_outputs(4679) <= not(inputs(135)) or (inputs(74));
    layer0_outputs(4680) <= inputs(171);
    layer0_outputs(4681) <= (inputs(237)) or (inputs(52));
    layer0_outputs(4682) <= inputs(119);
    layer0_outputs(4683) <= not(inputs(69)) or (inputs(63));
    layer0_outputs(4684) <= not((inputs(183)) xor (inputs(246)));
    layer0_outputs(4685) <= not((inputs(119)) or (inputs(27)));
    layer0_outputs(4686) <= not(inputs(230)) or (inputs(3));
    layer0_outputs(4687) <= not((inputs(151)) or (inputs(110)));
    layer0_outputs(4688) <= not((inputs(194)) or (inputs(174)));
    layer0_outputs(4689) <= not(inputs(98));
    layer0_outputs(4690) <= inputs(53);
    layer0_outputs(4691) <= not((inputs(75)) or (inputs(91)));
    layer0_outputs(4692) <= (inputs(145)) or (inputs(173));
    layer0_outputs(4693) <= not(inputs(2));
    layer0_outputs(4694) <= inputs(94);
    layer0_outputs(4695) <= not(inputs(105));
    layer0_outputs(4696) <= not(inputs(201)) or (inputs(98));
    layer0_outputs(4697) <= inputs(27);
    layer0_outputs(4698) <= (inputs(198)) or (inputs(149));
    layer0_outputs(4699) <= not((inputs(233)) xor (inputs(102)));
    layer0_outputs(4700) <= not(inputs(100)) or (inputs(35));
    layer0_outputs(4701) <= (inputs(97)) or (inputs(51));
    layer0_outputs(4702) <= not(inputs(39));
    layer0_outputs(4703) <= (inputs(122)) and not (inputs(207));
    layer0_outputs(4704) <= (inputs(245)) or (inputs(124));
    layer0_outputs(4705) <= (inputs(178)) xor (inputs(247));
    layer0_outputs(4706) <= inputs(174);
    layer0_outputs(4707) <= not(inputs(25));
    layer0_outputs(4708) <= not(inputs(67)) or (inputs(94));
    layer0_outputs(4709) <= inputs(156);
    layer0_outputs(4710) <= (inputs(208)) or (inputs(201));
    layer0_outputs(4711) <= not(inputs(81));
    layer0_outputs(4712) <= inputs(229);
    layer0_outputs(4713) <= (inputs(210)) or (inputs(216));
    layer0_outputs(4714) <= not(inputs(152));
    layer0_outputs(4715) <= not((inputs(130)) or (inputs(144)));
    layer0_outputs(4716) <= not(inputs(143)) or (inputs(111));
    layer0_outputs(4717) <= not(inputs(169)) or (inputs(49));
    layer0_outputs(4718) <= (inputs(162)) or (inputs(218));
    layer0_outputs(4719) <= inputs(99);
    layer0_outputs(4720) <= (inputs(11)) xor (inputs(250));
    layer0_outputs(4721) <= not((inputs(252)) or (inputs(128)));
    layer0_outputs(4722) <= inputs(123);
    layer0_outputs(4723) <= inputs(126);
    layer0_outputs(4724) <= (inputs(255)) or (inputs(68));
    layer0_outputs(4725) <= inputs(68);
    layer0_outputs(4726) <= not((inputs(93)) or (inputs(17)));
    layer0_outputs(4727) <= inputs(199);
    layer0_outputs(4728) <= (inputs(98)) and not (inputs(210));
    layer0_outputs(4729) <= (inputs(145)) and not (inputs(57));
    layer0_outputs(4730) <= (inputs(115)) or (inputs(96));
    layer0_outputs(4731) <= (inputs(163)) or (inputs(102));
    layer0_outputs(4732) <= (inputs(37)) or (inputs(62));
    layer0_outputs(4733) <= inputs(130);
    layer0_outputs(4734) <= not((inputs(17)) xor (inputs(92)));
    layer0_outputs(4735) <= not(inputs(218));
    layer0_outputs(4736) <= not(inputs(100));
    layer0_outputs(4737) <= not(inputs(232));
    layer0_outputs(4738) <= inputs(119);
    layer0_outputs(4739) <= inputs(85);
    layer0_outputs(4740) <= (inputs(147)) and not (inputs(2));
    layer0_outputs(4741) <= (inputs(211)) or (inputs(176));
    layer0_outputs(4742) <= (inputs(60)) or (inputs(2));
    layer0_outputs(4743) <= not(inputs(56));
    layer0_outputs(4744) <= inputs(2);
    layer0_outputs(4745) <= not(inputs(66));
    layer0_outputs(4746) <= (inputs(37)) and not (inputs(141));
    layer0_outputs(4747) <= not(inputs(248)) or (inputs(143));
    layer0_outputs(4748) <= inputs(97);
    layer0_outputs(4749) <= not(inputs(119));
    layer0_outputs(4750) <= (inputs(230)) and (inputs(231));
    layer0_outputs(4751) <= (inputs(117)) and not (inputs(8));
    layer0_outputs(4752) <= not((inputs(173)) xor (inputs(185)));
    layer0_outputs(4753) <= '1';
    layer0_outputs(4754) <= not(inputs(23));
    layer0_outputs(4755) <= not((inputs(69)) xor (inputs(87)));
    layer0_outputs(4756) <= not(inputs(129));
    layer0_outputs(4757) <= not((inputs(66)) and (inputs(254)));
    layer0_outputs(4758) <= not(inputs(168));
    layer0_outputs(4759) <= (inputs(55)) xor (inputs(30));
    layer0_outputs(4760) <= (inputs(99)) or (inputs(82));
    layer0_outputs(4761) <= inputs(25);
    layer0_outputs(4762) <= not((inputs(226)) xor (inputs(183)));
    layer0_outputs(4763) <= not(inputs(154)) or (inputs(240));
    layer0_outputs(4764) <= inputs(22);
    layer0_outputs(4765) <= (inputs(49)) and not (inputs(123));
    layer0_outputs(4766) <= not(inputs(91));
    layer0_outputs(4767) <= inputs(134);
    layer0_outputs(4768) <= inputs(93);
    layer0_outputs(4769) <= (inputs(197)) and not (inputs(42));
    layer0_outputs(4770) <= not(inputs(81)) or (inputs(56));
    layer0_outputs(4771) <= (inputs(252)) and not (inputs(31));
    layer0_outputs(4772) <= not(inputs(155));
    layer0_outputs(4773) <= inputs(227);
    layer0_outputs(4774) <= not(inputs(52));
    layer0_outputs(4775) <= (inputs(127)) or (inputs(199));
    layer0_outputs(4776) <= not(inputs(85));
    layer0_outputs(4777) <= not(inputs(50)) or (inputs(2));
    layer0_outputs(4778) <= (inputs(188)) and not (inputs(12));
    layer0_outputs(4779) <= not(inputs(141));
    layer0_outputs(4780) <= inputs(150);
    layer0_outputs(4781) <= (inputs(17)) or (inputs(230));
    layer0_outputs(4782) <= not(inputs(163));
    layer0_outputs(4783) <= not((inputs(125)) or (inputs(96)));
    layer0_outputs(4784) <= not((inputs(130)) or (inputs(172)));
    layer0_outputs(4785) <= (inputs(62)) and (inputs(30));
    layer0_outputs(4786) <= not(inputs(247)) or (inputs(239));
    layer0_outputs(4787) <= not(inputs(143));
    layer0_outputs(4788) <= not((inputs(198)) xor (inputs(195)));
    layer0_outputs(4789) <= not(inputs(109)) or (inputs(49));
    layer0_outputs(4790) <= not((inputs(80)) or (inputs(201)));
    layer0_outputs(4791) <= not((inputs(167)) or (inputs(109)));
    layer0_outputs(4792) <= (inputs(173)) and (inputs(58));
    layer0_outputs(4793) <= not(inputs(38));
    layer0_outputs(4794) <= (inputs(79)) or (inputs(141));
    layer0_outputs(4795) <= not(inputs(120)) or (inputs(14));
    layer0_outputs(4796) <= not(inputs(167));
    layer0_outputs(4797) <= not((inputs(62)) or (inputs(206)));
    layer0_outputs(4798) <= not(inputs(38)) or (inputs(191));
    layer0_outputs(4799) <= inputs(114);
    layer0_outputs(4800) <= not(inputs(170));
    layer0_outputs(4801) <= (inputs(21)) and not (inputs(232));
    layer0_outputs(4802) <= not(inputs(231));
    layer0_outputs(4803) <= not(inputs(219)) or (inputs(149));
    layer0_outputs(4804) <= (inputs(63)) and (inputs(48));
    layer0_outputs(4805) <= not((inputs(28)) or (inputs(130)));
    layer0_outputs(4806) <= not(inputs(56));
    layer0_outputs(4807) <= (inputs(237)) or (inputs(135));
    layer0_outputs(4808) <= not(inputs(229));
    layer0_outputs(4809) <= not((inputs(191)) xor (inputs(24)));
    layer0_outputs(4810) <= not(inputs(160));
    layer0_outputs(4811) <= (inputs(134)) and not (inputs(254));
    layer0_outputs(4812) <= not((inputs(252)) or (inputs(193)));
    layer0_outputs(4813) <= not(inputs(88));
    layer0_outputs(4814) <= (inputs(49)) or (inputs(90));
    layer0_outputs(4815) <= inputs(74);
    layer0_outputs(4816) <= not((inputs(160)) or (inputs(237)));
    layer0_outputs(4817) <= inputs(98);
    layer0_outputs(4818) <= not((inputs(194)) or (inputs(232)));
    layer0_outputs(4819) <= inputs(142);
    layer0_outputs(4820) <= (inputs(175)) or (inputs(216));
    layer0_outputs(4821) <= (inputs(46)) or (inputs(76));
    layer0_outputs(4822) <= not(inputs(88)) or (inputs(65));
    layer0_outputs(4823) <= not(inputs(179)) or (inputs(172));
    layer0_outputs(4824) <= not((inputs(105)) or (inputs(194)));
    layer0_outputs(4825) <= not(inputs(27)) or (inputs(110));
    layer0_outputs(4826) <= not(inputs(112)) or (inputs(95));
    layer0_outputs(4827) <= (inputs(92)) and not (inputs(225));
    layer0_outputs(4828) <= not(inputs(216));
    layer0_outputs(4829) <= not(inputs(202)) or (inputs(112));
    layer0_outputs(4830) <= inputs(214);
    layer0_outputs(4831) <= not(inputs(92));
    layer0_outputs(4832) <= not(inputs(107));
    layer0_outputs(4833) <= (inputs(195)) or (inputs(10));
    layer0_outputs(4834) <= (inputs(68)) xor (inputs(49));
    layer0_outputs(4835) <= not((inputs(41)) xor (inputs(37)));
    layer0_outputs(4836) <= inputs(97);
    layer0_outputs(4837) <= inputs(82);
    layer0_outputs(4838) <= not(inputs(104));
    layer0_outputs(4839) <= inputs(140);
    layer0_outputs(4840) <= (inputs(9)) or (inputs(219));
    layer0_outputs(4841) <= not(inputs(167)) or (inputs(110));
    layer0_outputs(4842) <= not(inputs(191));
    layer0_outputs(4843) <= inputs(144);
    layer0_outputs(4844) <= not(inputs(229));
    layer0_outputs(4845) <= (inputs(97)) xor (inputs(85));
    layer0_outputs(4846) <= (inputs(11)) and not (inputs(242));
    layer0_outputs(4847) <= (inputs(177)) or (inputs(81));
    layer0_outputs(4848) <= not(inputs(84));
    layer0_outputs(4849) <= not((inputs(220)) or (inputs(224)));
    layer0_outputs(4850) <= not((inputs(117)) or (inputs(98)));
    layer0_outputs(4851) <= not((inputs(55)) or (inputs(6)));
    layer0_outputs(4852) <= (inputs(238)) or (inputs(205));
    layer0_outputs(4853) <= inputs(211);
    layer0_outputs(4854) <= (inputs(104)) xor (inputs(1));
    layer0_outputs(4855) <= not(inputs(62)) or (inputs(240));
    layer0_outputs(4856) <= not(inputs(72));
    layer0_outputs(4857) <= (inputs(242)) xor (inputs(214));
    layer0_outputs(4858) <= not((inputs(169)) xor (inputs(154)));
    layer0_outputs(4859) <= (inputs(73)) or (inputs(16));
    layer0_outputs(4860) <= (inputs(121)) and not (inputs(140));
    layer0_outputs(4861) <= not((inputs(170)) xor (inputs(196)));
    layer0_outputs(4862) <= (inputs(192)) or (inputs(5));
    layer0_outputs(4863) <= not((inputs(68)) or (inputs(127)));
    layer0_outputs(4864) <= (inputs(120)) and not (inputs(229));
    layer0_outputs(4865) <= (inputs(218)) xor (inputs(122));
    layer0_outputs(4866) <= not((inputs(48)) or (inputs(231)));
    layer0_outputs(4867) <= (inputs(249)) or (inputs(67));
    layer0_outputs(4868) <= not(inputs(10)) or (inputs(129));
    layer0_outputs(4869) <= not(inputs(255));
    layer0_outputs(4870) <= not(inputs(170)) or (inputs(229));
    layer0_outputs(4871) <= not(inputs(168)) or (inputs(174));
    layer0_outputs(4872) <= not((inputs(250)) xor (inputs(196)));
    layer0_outputs(4873) <= (inputs(20)) xor (inputs(111));
    layer0_outputs(4874) <= inputs(82);
    layer0_outputs(4875) <= not((inputs(217)) or (inputs(123)));
    layer0_outputs(4876) <= inputs(179);
    layer0_outputs(4877) <= inputs(43);
    layer0_outputs(4878) <= (inputs(151)) and (inputs(135));
    layer0_outputs(4879) <= not(inputs(138)) or (inputs(232));
    layer0_outputs(4880) <= not((inputs(160)) or (inputs(85)));
    layer0_outputs(4881) <= not((inputs(162)) or (inputs(236)));
    layer0_outputs(4882) <= (inputs(183)) and not (inputs(140));
    layer0_outputs(4883) <= inputs(173);
    layer0_outputs(4884) <= not(inputs(76));
    layer0_outputs(4885) <= not((inputs(127)) xor (inputs(5)));
    layer0_outputs(4886) <= (inputs(124)) xor (inputs(110));
    layer0_outputs(4887) <= inputs(181);
    layer0_outputs(4888) <= not(inputs(153)) or (inputs(240));
    layer0_outputs(4889) <= (inputs(120)) and not (inputs(7));
    layer0_outputs(4890) <= not(inputs(153));
    layer0_outputs(4891) <= (inputs(98)) and not (inputs(78));
    layer0_outputs(4892) <= (inputs(5)) and not (inputs(159));
    layer0_outputs(4893) <= not(inputs(250)) or (inputs(58));
    layer0_outputs(4894) <= not((inputs(218)) or (inputs(56)));
    layer0_outputs(4895) <= not(inputs(213));
    layer0_outputs(4896) <= not((inputs(84)) or (inputs(99)));
    layer0_outputs(4897) <= (inputs(229)) and not (inputs(135));
    layer0_outputs(4898) <= not((inputs(210)) or (inputs(5)));
    layer0_outputs(4899) <= (inputs(134)) and not (inputs(95));
    layer0_outputs(4900) <= inputs(92);
    layer0_outputs(4901) <= (inputs(227)) or (inputs(176));
    layer0_outputs(4902) <= (inputs(180)) and not (inputs(159));
    layer0_outputs(4903) <= '1';
    layer0_outputs(4904) <= (inputs(244)) or (inputs(187));
    layer0_outputs(4905) <= not((inputs(34)) or (inputs(140)));
    layer0_outputs(4906) <= not(inputs(217));
    layer0_outputs(4907) <= not((inputs(242)) xor (inputs(31)));
    layer0_outputs(4908) <= (inputs(240)) xor (inputs(7));
    layer0_outputs(4909) <= not(inputs(41));
    layer0_outputs(4910) <= '1';
    layer0_outputs(4911) <= not((inputs(2)) or (inputs(89)));
    layer0_outputs(4912) <= not((inputs(236)) or (inputs(248)));
    layer0_outputs(4913) <= not((inputs(21)) or (inputs(84)));
    layer0_outputs(4914) <= not((inputs(186)) or (inputs(159)));
    layer0_outputs(4915) <= not((inputs(83)) xor (inputs(211)));
    layer0_outputs(4916) <= (inputs(101)) xor (inputs(49));
    layer0_outputs(4917) <= not((inputs(71)) and (inputs(199)));
    layer0_outputs(4918) <= (inputs(20)) and not (inputs(253));
    layer0_outputs(4919) <= not((inputs(115)) or (inputs(239)));
    layer0_outputs(4920) <= not(inputs(92));
    layer0_outputs(4921) <= not((inputs(248)) or (inputs(112)));
    layer0_outputs(4922) <= not(inputs(66)) or (inputs(17));
    layer0_outputs(4923) <= not(inputs(216)) or (inputs(110));
    layer0_outputs(4924) <= (inputs(184)) and not (inputs(171));
    layer0_outputs(4925) <= not(inputs(59)) or (inputs(236));
    layer0_outputs(4926) <= inputs(67);
    layer0_outputs(4927) <= inputs(32);
    layer0_outputs(4928) <= (inputs(214)) xor (inputs(160));
    layer0_outputs(4929) <= not((inputs(151)) or (inputs(150)));
    layer0_outputs(4930) <= (inputs(11)) or (inputs(245));
    layer0_outputs(4931) <= '1';
    layer0_outputs(4932) <= inputs(45);
    layer0_outputs(4933) <= not((inputs(129)) xor (inputs(87)));
    layer0_outputs(4934) <= (inputs(209)) xor (inputs(88));
    layer0_outputs(4935) <= not(inputs(206)) or (inputs(97));
    layer0_outputs(4936) <= not(inputs(214));
    layer0_outputs(4937) <= not((inputs(154)) xor (inputs(54)));
    layer0_outputs(4938) <= not((inputs(12)) or (inputs(70)));
    layer0_outputs(4939) <= inputs(121);
    layer0_outputs(4940) <= inputs(121);
    layer0_outputs(4941) <= inputs(97);
    layer0_outputs(4942) <= (inputs(69)) or (inputs(84));
    layer0_outputs(4943) <= not(inputs(70)) or (inputs(94));
    layer0_outputs(4944) <= not(inputs(243)) or (inputs(177));
    layer0_outputs(4945) <= (inputs(40)) and not (inputs(77));
    layer0_outputs(4946) <= (inputs(244)) and (inputs(155));
    layer0_outputs(4947) <= (inputs(240)) or (inputs(168));
    layer0_outputs(4948) <= not((inputs(193)) or (inputs(88)));
    layer0_outputs(4949) <= not((inputs(74)) xor (inputs(0)));
    layer0_outputs(4950) <= (inputs(173)) xor (inputs(231));
    layer0_outputs(4951) <= (inputs(109)) or (inputs(179));
    layer0_outputs(4952) <= (inputs(36)) or (inputs(208));
    layer0_outputs(4953) <= not((inputs(253)) or (inputs(44)));
    layer0_outputs(4954) <= inputs(105);
    layer0_outputs(4955) <= not(inputs(118));
    layer0_outputs(4956) <= not(inputs(192)) or (inputs(156));
    layer0_outputs(4957) <= not(inputs(124));
    layer0_outputs(4958) <= not((inputs(12)) or (inputs(233)));
    layer0_outputs(4959) <= (inputs(84)) and not (inputs(165));
    layer0_outputs(4960) <= (inputs(253)) or (inputs(9));
    layer0_outputs(4961) <= not(inputs(46)) or (inputs(241));
    layer0_outputs(4962) <= not(inputs(240)) or (inputs(238));
    layer0_outputs(4963) <= not(inputs(120)) or (inputs(113));
    layer0_outputs(4964) <= inputs(34);
    layer0_outputs(4965) <= (inputs(229)) and not (inputs(63));
    layer0_outputs(4966) <= inputs(115);
    layer0_outputs(4967) <= not(inputs(218));
    layer0_outputs(4968) <= not((inputs(158)) or (inputs(220)));
    layer0_outputs(4969) <= not(inputs(179)) or (inputs(238));
    layer0_outputs(4970) <= (inputs(148)) or (inputs(116));
    layer0_outputs(4971) <= (inputs(167)) and not (inputs(91));
    layer0_outputs(4972) <= not((inputs(127)) or (inputs(98)));
    layer0_outputs(4973) <= not(inputs(215)) or (inputs(15));
    layer0_outputs(4974) <= not((inputs(218)) or (inputs(93)));
    layer0_outputs(4975) <= (inputs(128)) or (inputs(32));
    layer0_outputs(4976) <= not(inputs(201));
    layer0_outputs(4977) <= inputs(229);
    layer0_outputs(4978) <= (inputs(216)) and not (inputs(123));
    layer0_outputs(4979) <= not((inputs(204)) xor (inputs(30)));
    layer0_outputs(4980) <= inputs(226);
    layer0_outputs(4981) <= (inputs(87)) and not (inputs(207));
    layer0_outputs(4982) <= (inputs(122)) and not (inputs(193));
    layer0_outputs(4983) <= (inputs(27)) and not (inputs(244));
    layer0_outputs(4984) <= not((inputs(186)) or (inputs(239)));
    layer0_outputs(4985) <= not((inputs(238)) or (inputs(40)));
    layer0_outputs(4986) <= (inputs(241)) xor (inputs(164));
    layer0_outputs(4987) <= (inputs(96)) or (inputs(81));
    layer0_outputs(4988) <= not((inputs(171)) or (inputs(162)));
    layer0_outputs(4989) <= (inputs(8)) or (inputs(221));
    layer0_outputs(4990) <= not(inputs(134));
    layer0_outputs(4991) <= not(inputs(134)) or (inputs(127));
    layer0_outputs(4992) <= not(inputs(220));
    layer0_outputs(4993) <= inputs(217);
    layer0_outputs(4994) <= inputs(119);
    layer0_outputs(4995) <= inputs(23);
    layer0_outputs(4996) <= not((inputs(99)) and (inputs(133)));
    layer0_outputs(4997) <= inputs(58);
    layer0_outputs(4998) <= not((inputs(54)) or (inputs(116)));
    layer0_outputs(4999) <= (inputs(180)) or (inputs(64));
    layer0_outputs(5000) <= (inputs(82)) xor (inputs(96));
    layer0_outputs(5001) <= (inputs(164)) or (inputs(158));
    layer0_outputs(5002) <= (inputs(158)) or (inputs(130));
    layer0_outputs(5003) <= not((inputs(29)) or (inputs(3)));
    layer0_outputs(5004) <= not(inputs(153)) or (inputs(47));
    layer0_outputs(5005) <= not((inputs(23)) xor (inputs(174)));
    layer0_outputs(5006) <= not(inputs(73)) or (inputs(64));
    layer0_outputs(5007) <= not((inputs(205)) or (inputs(15)));
    layer0_outputs(5008) <= (inputs(105)) and not (inputs(210));
    layer0_outputs(5009) <= inputs(178);
    layer0_outputs(5010) <= not((inputs(192)) or (inputs(227)));
    layer0_outputs(5011) <= inputs(83);
    layer0_outputs(5012) <= (inputs(174)) xor (inputs(191));
    layer0_outputs(5013) <= not(inputs(119));
    layer0_outputs(5014) <= inputs(118);
    layer0_outputs(5015) <= inputs(107);
    layer0_outputs(5016) <= not((inputs(49)) or (inputs(249)));
    layer0_outputs(5017) <= (inputs(197)) and not (inputs(146));
    layer0_outputs(5018) <= (inputs(105)) and not (inputs(53));
    layer0_outputs(5019) <= not(inputs(209));
    layer0_outputs(5020) <= not((inputs(68)) or (inputs(52)));
    layer0_outputs(5021) <= inputs(75);
    layer0_outputs(5022) <= not(inputs(238));
    layer0_outputs(5023) <= not(inputs(246));
    layer0_outputs(5024) <= (inputs(106)) and not (inputs(216));
    layer0_outputs(5025) <= inputs(86);
    layer0_outputs(5026) <= inputs(40);
    layer0_outputs(5027) <= not((inputs(82)) xor (inputs(3)));
    layer0_outputs(5028) <= not((inputs(246)) or (inputs(161)));
    layer0_outputs(5029) <= not(inputs(165));
    layer0_outputs(5030) <= inputs(209);
    layer0_outputs(5031) <= (inputs(182)) and not (inputs(31));
    layer0_outputs(5032) <= inputs(125);
    layer0_outputs(5033) <= (inputs(120)) and not (inputs(36));
    layer0_outputs(5034) <= not((inputs(16)) xor (inputs(77)));
    layer0_outputs(5035) <= (inputs(68)) or (inputs(1));
    layer0_outputs(5036) <= (inputs(149)) xor (inputs(130));
    layer0_outputs(5037) <= not((inputs(56)) xor (inputs(75)));
    layer0_outputs(5038) <= not((inputs(248)) or (inputs(230)));
    layer0_outputs(5039) <= (inputs(27)) or (inputs(19));
    layer0_outputs(5040) <= not((inputs(97)) or (inputs(119)));
    layer0_outputs(5041) <= inputs(25);
    layer0_outputs(5042) <= (inputs(20)) xor (inputs(12));
    layer0_outputs(5043) <= '1';
    layer0_outputs(5044) <= (inputs(61)) or (inputs(164));
    layer0_outputs(5045) <= (inputs(133)) and (inputs(64));
    layer0_outputs(5046) <= (inputs(223)) or (inputs(222));
    layer0_outputs(5047) <= not(inputs(50));
    layer0_outputs(5048) <= not(inputs(162)) or (inputs(68));
    layer0_outputs(5049) <= not(inputs(182));
    layer0_outputs(5050) <= (inputs(202)) or (inputs(208));
    layer0_outputs(5051) <= (inputs(145)) and not (inputs(192));
    layer0_outputs(5052) <= (inputs(115)) or (inputs(69));
    layer0_outputs(5053) <= not(inputs(95));
    layer0_outputs(5054) <= (inputs(102)) xor (inputs(71));
    layer0_outputs(5055) <= (inputs(231)) and not (inputs(110));
    layer0_outputs(5056) <= inputs(179);
    layer0_outputs(5057) <= not(inputs(58)) or (inputs(222));
    layer0_outputs(5058) <= (inputs(242)) and not (inputs(161));
    layer0_outputs(5059) <= not(inputs(228));
    layer0_outputs(5060) <= (inputs(215)) and not (inputs(159));
    layer0_outputs(5061) <= inputs(207);
    layer0_outputs(5062) <= not(inputs(14));
    layer0_outputs(5063) <= inputs(176);
    layer0_outputs(5064) <= not(inputs(60));
    layer0_outputs(5065) <= inputs(249);
    layer0_outputs(5066) <= not((inputs(100)) or (inputs(141)));
    layer0_outputs(5067) <= (inputs(241)) or (inputs(111));
    layer0_outputs(5068) <= not(inputs(21)) or (inputs(128));
    layer0_outputs(5069) <= not(inputs(115));
    layer0_outputs(5070) <= not((inputs(51)) or (inputs(60)));
    layer0_outputs(5071) <= (inputs(196)) and not (inputs(58));
    layer0_outputs(5072) <= not((inputs(2)) or (inputs(183)));
    layer0_outputs(5073) <= inputs(150);
    layer0_outputs(5074) <= not(inputs(98));
    layer0_outputs(5075) <= not(inputs(197)) or (inputs(192));
    layer0_outputs(5076) <= not(inputs(52));
    layer0_outputs(5077) <= (inputs(60)) and not (inputs(210));
    layer0_outputs(5078) <= (inputs(255)) or (inputs(225));
    layer0_outputs(5079) <= (inputs(5)) and not (inputs(66));
    layer0_outputs(5080) <= not((inputs(6)) xor (inputs(71)));
    layer0_outputs(5081) <= inputs(134);
    layer0_outputs(5082) <= (inputs(196)) xor (inputs(38));
    layer0_outputs(5083) <= not(inputs(42));
    layer0_outputs(5084) <= not(inputs(184));
    layer0_outputs(5085) <= (inputs(1)) xor (inputs(163));
    layer0_outputs(5086) <= not(inputs(100)) or (inputs(33));
    layer0_outputs(5087) <= (inputs(182)) and not (inputs(128));
    layer0_outputs(5088) <= not(inputs(245));
    layer0_outputs(5089) <= not(inputs(123));
    layer0_outputs(5090) <= inputs(227);
    layer0_outputs(5091) <= not(inputs(228)) or (inputs(2));
    layer0_outputs(5092) <= not((inputs(14)) or (inputs(185)));
    layer0_outputs(5093) <= '0';
    layer0_outputs(5094) <= (inputs(17)) or (inputs(118));
    layer0_outputs(5095) <= inputs(18);
    layer0_outputs(5096) <= not(inputs(162));
    layer0_outputs(5097) <= not(inputs(74));
    layer0_outputs(5098) <= (inputs(60)) and (inputs(64));
    layer0_outputs(5099) <= (inputs(167)) and not (inputs(252));
    layer0_outputs(5100) <= (inputs(250)) or (inputs(163));
    layer0_outputs(5101) <= not(inputs(43)) or (inputs(186));
    layer0_outputs(5102) <= not(inputs(119));
    layer0_outputs(5103) <= inputs(195);
    layer0_outputs(5104) <= inputs(137);
    layer0_outputs(5105) <= not(inputs(94)) or (inputs(33));
    layer0_outputs(5106) <= (inputs(42)) or (inputs(40));
    layer0_outputs(5107) <= not(inputs(185));
    layer0_outputs(5108) <= not(inputs(104)) or (inputs(208));
    layer0_outputs(5109) <= not(inputs(164));
    layer0_outputs(5110) <= not(inputs(80));
    layer0_outputs(5111) <= '0';
    layer0_outputs(5112) <= (inputs(175)) xor (inputs(109));
    layer0_outputs(5113) <= inputs(11);
    layer0_outputs(5114) <= not(inputs(195)) or (inputs(233));
    layer0_outputs(5115) <= not((inputs(106)) or (inputs(233)));
    layer0_outputs(5116) <= not((inputs(104)) or (inputs(223)));
    layer0_outputs(5117) <= not(inputs(51));
    layer0_outputs(5118) <= (inputs(225)) xor (inputs(187));
    layer0_outputs(5119) <= not(inputs(204)) or (inputs(139));
    outputs(0) <= layer0_outputs(2927);
    outputs(1) <= (layer0_outputs(3917)) and (layer0_outputs(4511));
    outputs(2) <= (layer0_outputs(1860)) and not (layer0_outputs(2765));
    outputs(3) <= not(layer0_outputs(2333));
    outputs(4) <= not(layer0_outputs(3517)) or (layer0_outputs(4079));
    outputs(5) <= (layer0_outputs(4264)) and not (layer0_outputs(1696));
    outputs(6) <= not(layer0_outputs(3465));
    outputs(7) <= (layer0_outputs(1407)) xor (layer0_outputs(2785));
    outputs(8) <= (layer0_outputs(4760)) and (layer0_outputs(2625));
    outputs(9) <= layer0_outputs(4312);
    outputs(10) <= layer0_outputs(2090);
    outputs(11) <= not(layer0_outputs(1551));
    outputs(12) <= (layer0_outputs(3291)) and (layer0_outputs(4154));
    outputs(13) <= (layer0_outputs(2513)) xor (layer0_outputs(3165));
    outputs(14) <= not((layer0_outputs(686)) and (layer0_outputs(636)));
    outputs(15) <= not(layer0_outputs(2181)) or (layer0_outputs(5044));
    outputs(16) <= layer0_outputs(234);
    outputs(17) <= not((layer0_outputs(2861)) and (layer0_outputs(3132)));
    outputs(18) <= (layer0_outputs(408)) and not (layer0_outputs(1488));
    outputs(19) <= (layer0_outputs(1063)) and not (layer0_outputs(2097));
    outputs(20) <= not((layer0_outputs(1462)) or (layer0_outputs(4546)));
    outputs(21) <= (layer0_outputs(586)) and (layer0_outputs(4306));
    outputs(22) <= (layer0_outputs(3794)) and not (layer0_outputs(153));
    outputs(23) <= not((layer0_outputs(3300)) or (layer0_outputs(3394)));
    outputs(24) <= (layer0_outputs(1920)) and not (layer0_outputs(5083));
    outputs(25) <= not(layer0_outputs(409)) or (layer0_outputs(2069));
    outputs(26) <= layer0_outputs(1138);
    outputs(27) <= not((layer0_outputs(1656)) or (layer0_outputs(2565)));
    outputs(28) <= not(layer0_outputs(2414)) or (layer0_outputs(2518));
    outputs(29) <= layer0_outputs(3880);
    outputs(30) <= layer0_outputs(861);
    outputs(31) <= (layer0_outputs(672)) or (layer0_outputs(3483));
    outputs(32) <= not((layer0_outputs(1916)) and (layer0_outputs(3158)));
    outputs(33) <= not((layer0_outputs(5006)) and (layer0_outputs(5053)));
    outputs(34) <= not(layer0_outputs(1093));
    outputs(35) <= not(layer0_outputs(3357));
    outputs(36) <= (layer0_outputs(3340)) and not (layer0_outputs(4029));
    outputs(37) <= layer0_outputs(2201);
    outputs(38) <= not((layer0_outputs(3452)) and (layer0_outputs(656)));
    outputs(39) <= layer0_outputs(2032);
    outputs(40) <= layer0_outputs(1313);
    outputs(41) <= layer0_outputs(6);
    outputs(42) <= (layer0_outputs(2677)) and not (layer0_outputs(4116));
    outputs(43) <= not((layer0_outputs(4895)) or (layer0_outputs(3460)));
    outputs(44) <= not(layer0_outputs(4082));
    outputs(45) <= (layer0_outputs(3794)) and not (layer0_outputs(4914));
    outputs(46) <= not(layer0_outputs(961));
    outputs(47) <= layer0_outputs(1276);
    outputs(48) <= layer0_outputs(611);
    outputs(49) <= (layer0_outputs(4552)) and not (layer0_outputs(2533));
    outputs(50) <= (layer0_outputs(5022)) and not (layer0_outputs(4881));
    outputs(51) <= not(layer0_outputs(2257));
    outputs(52) <= not(layer0_outputs(30));
    outputs(53) <= (layer0_outputs(791)) and not (layer0_outputs(4780));
    outputs(54) <= (layer0_outputs(1192)) or (layer0_outputs(4815));
    outputs(55) <= layer0_outputs(4180);
    outputs(56) <= not(layer0_outputs(4302));
    outputs(57) <= layer0_outputs(1518);
    outputs(58) <= layer0_outputs(4332);
    outputs(59) <= layer0_outputs(2573);
    outputs(60) <= (layer0_outputs(2883)) and (layer0_outputs(2592));
    outputs(61) <= layer0_outputs(4176);
    outputs(62) <= layer0_outputs(4613);
    outputs(63) <= (layer0_outputs(1540)) and not (layer0_outputs(3090));
    outputs(64) <= not(layer0_outputs(3442));
    outputs(65) <= (layer0_outputs(3078)) and not (layer0_outputs(4974));
    outputs(66) <= not(layer0_outputs(474));
    outputs(67) <= not((layer0_outputs(2697)) xor (layer0_outputs(621)));
    outputs(68) <= not(layer0_outputs(1905));
    outputs(69) <= (layer0_outputs(5062)) and (layer0_outputs(4236));
    outputs(70) <= (layer0_outputs(4720)) or (layer0_outputs(764));
    outputs(71) <= not(layer0_outputs(120));
    outputs(72) <= (layer0_outputs(1783)) and (layer0_outputs(4597));
    outputs(73) <= not(layer0_outputs(4215));
    outputs(74) <= (layer0_outputs(3212)) and (layer0_outputs(2841));
    outputs(75) <= not(layer0_outputs(1132)) or (layer0_outputs(1020));
    outputs(76) <= not(layer0_outputs(63));
    outputs(77) <= layer0_outputs(3901);
    outputs(78) <= (layer0_outputs(853)) or (layer0_outputs(2130));
    outputs(79) <= layer0_outputs(542);
    outputs(80) <= not((layer0_outputs(1809)) and (layer0_outputs(4787)));
    outputs(81) <= not(layer0_outputs(2653));
    outputs(82) <= (layer0_outputs(2723)) and not (layer0_outputs(1719));
    outputs(83) <= (layer0_outputs(2012)) and not (layer0_outputs(2293));
    outputs(84) <= (layer0_outputs(2517)) and (layer0_outputs(4838));
    outputs(85) <= (layer0_outputs(4191)) xor (layer0_outputs(4083));
    outputs(86) <= (layer0_outputs(4792)) or (layer0_outputs(1639));
    outputs(87) <= not(layer0_outputs(2829));
    outputs(88) <= not(layer0_outputs(190));
    outputs(89) <= not(layer0_outputs(1611)) or (layer0_outputs(1220));
    outputs(90) <= not(layer0_outputs(2122));
    outputs(91) <= (layer0_outputs(460)) and (layer0_outputs(2360));
    outputs(92) <= (layer0_outputs(272)) or (layer0_outputs(205));
    outputs(93) <= (layer0_outputs(586)) and (layer0_outputs(537));
    outputs(94) <= layer0_outputs(1134);
    outputs(95) <= not(layer0_outputs(1108));
    outputs(96) <= layer0_outputs(3024);
    outputs(97) <= layer0_outputs(4236);
    outputs(98) <= layer0_outputs(2162);
    outputs(99) <= not(layer0_outputs(1861));
    outputs(100) <= layer0_outputs(338);
    outputs(101) <= not((layer0_outputs(3371)) xor (layer0_outputs(1417)));
    outputs(102) <= (layer0_outputs(3487)) or (layer0_outputs(1497));
    outputs(103) <= (layer0_outputs(4672)) and not (layer0_outputs(3433));
    outputs(104) <= (layer0_outputs(3711)) or (layer0_outputs(2325));
    outputs(105) <= not(layer0_outputs(3734)) or (layer0_outputs(723));
    outputs(106) <= (layer0_outputs(95)) or (layer0_outputs(1444));
    outputs(107) <= not((layer0_outputs(3745)) and (layer0_outputs(996)));
    outputs(108) <= (layer0_outputs(2991)) or (layer0_outputs(1519));
    outputs(109) <= not((layer0_outputs(3001)) xor (layer0_outputs(1886)));
    outputs(110) <= not(layer0_outputs(1960));
    outputs(111) <= not((layer0_outputs(4523)) and (layer0_outputs(11)));
    outputs(112) <= not((layer0_outputs(394)) and (layer0_outputs(5105)));
    outputs(113) <= layer0_outputs(5116);
    outputs(114) <= not((layer0_outputs(1487)) and (layer0_outputs(3133)));
    outputs(115) <= layer0_outputs(2817);
    outputs(116) <= not(layer0_outputs(1031));
    outputs(117) <= not(layer0_outputs(5104));
    outputs(118) <= not(layer0_outputs(1608));
    outputs(119) <= layer0_outputs(4239);
    outputs(120) <= (layer0_outputs(1645)) and not (layer0_outputs(3472));
    outputs(121) <= not(layer0_outputs(3710));
    outputs(122) <= not((layer0_outputs(1756)) xor (layer0_outputs(4462)));
    outputs(123) <= (layer0_outputs(1291)) or (layer0_outputs(764));
    outputs(124) <= layer0_outputs(4146);
    outputs(125) <= not(layer0_outputs(3166));
    outputs(126) <= (layer0_outputs(670)) xor (layer0_outputs(1034));
    outputs(127) <= not(layer0_outputs(2310));
    outputs(128) <= (layer0_outputs(3929)) and not (layer0_outputs(165));
    outputs(129) <= layer0_outputs(2530);
    outputs(130) <= not(layer0_outputs(5075)) or (layer0_outputs(439));
    outputs(131) <= (layer0_outputs(1252)) and (layer0_outputs(2501));
    outputs(132) <= layer0_outputs(4391);
    outputs(133) <= not(layer0_outputs(4233));
    outputs(134) <= not((layer0_outputs(1581)) xor (layer0_outputs(3430)));
    outputs(135) <= not((layer0_outputs(3945)) xor (layer0_outputs(2244)));
    outputs(136) <= not((layer0_outputs(3126)) and (layer0_outputs(3375)));
    outputs(137) <= (layer0_outputs(1589)) and (layer0_outputs(1825));
    outputs(138) <= not(layer0_outputs(3946));
    outputs(139) <= layer0_outputs(2840);
    outputs(140) <= not(layer0_outputs(3822));
    outputs(141) <= not(layer0_outputs(3676));
    outputs(142) <= not(layer0_outputs(961));
    outputs(143) <= not(layer0_outputs(3530)) or (layer0_outputs(2014));
    outputs(144) <= not(layer0_outputs(4789));
    outputs(145) <= not(layer0_outputs(3951));
    outputs(146) <= layer0_outputs(3324);
    outputs(147) <= layer0_outputs(4877);
    outputs(148) <= (layer0_outputs(324)) and not (layer0_outputs(2315));
    outputs(149) <= layer0_outputs(4749);
    outputs(150) <= not((layer0_outputs(3913)) xor (layer0_outputs(4227)));
    outputs(151) <= (layer0_outputs(3260)) and (layer0_outputs(4929));
    outputs(152) <= (layer0_outputs(4136)) and not (layer0_outputs(2445));
    outputs(153) <= not(layer0_outputs(31));
    outputs(154) <= layer0_outputs(4507);
    outputs(155) <= layer0_outputs(4176);
    outputs(156) <= not(layer0_outputs(3489)) or (layer0_outputs(2876));
    outputs(157) <= not(layer0_outputs(876));
    outputs(158) <= (layer0_outputs(1196)) and (layer0_outputs(2249));
    outputs(159) <= (layer0_outputs(1721)) and (layer0_outputs(3581));
    outputs(160) <= not((layer0_outputs(2738)) xor (layer0_outputs(1635)));
    outputs(161) <= layer0_outputs(1321);
    outputs(162) <= layer0_outputs(1715);
    outputs(163) <= not((layer0_outputs(3621)) xor (layer0_outputs(4604)));
    outputs(164) <= not(layer0_outputs(1455));
    outputs(165) <= not(layer0_outputs(72));
    outputs(166) <= not(layer0_outputs(1651)) or (layer0_outputs(3053));
    outputs(167) <= not(layer0_outputs(4275)) or (layer0_outputs(1437));
    outputs(168) <= (layer0_outputs(2209)) and not (layer0_outputs(3782));
    outputs(169) <= not((layer0_outputs(2640)) and (layer0_outputs(4921)));
    outputs(170) <= layer0_outputs(4758);
    outputs(171) <= not(layer0_outputs(4565));
    outputs(172) <= layer0_outputs(2404);
    outputs(173) <= layer0_outputs(1300);
    outputs(174) <= not((layer0_outputs(4529)) or (layer0_outputs(1169)));
    outputs(175) <= not(layer0_outputs(1398)) or (layer0_outputs(1253));
    outputs(176) <= not(layer0_outputs(4780));
    outputs(177) <= layer0_outputs(3572);
    outputs(178) <= layer0_outputs(3037);
    outputs(179) <= (layer0_outputs(4928)) or (layer0_outputs(1428));
    outputs(180) <= not(layer0_outputs(2022)) or (layer0_outputs(238));
    outputs(181) <= not(layer0_outputs(4767));
    outputs(182) <= (layer0_outputs(2748)) and not (layer0_outputs(1492));
    outputs(183) <= layer0_outputs(1860);
    outputs(184) <= (layer0_outputs(1792)) and not (layer0_outputs(3991));
    outputs(185) <= layer0_outputs(3106);
    outputs(186) <= layer0_outputs(3925);
    outputs(187) <= layer0_outputs(1918);
    outputs(188) <= layer0_outputs(4051);
    outputs(189) <= layer0_outputs(4825);
    outputs(190) <= not(layer0_outputs(3928));
    outputs(191) <= not(layer0_outputs(1973));
    outputs(192) <= (layer0_outputs(4911)) and not (layer0_outputs(127));
    outputs(193) <= (layer0_outputs(707)) or (layer0_outputs(717));
    outputs(194) <= not(layer0_outputs(4615)) or (layer0_outputs(4062));
    outputs(195) <= layer0_outputs(1428);
    outputs(196) <= layer0_outputs(2628);
    outputs(197) <= not(layer0_outputs(3215));
    outputs(198) <= not(layer0_outputs(1562));
    outputs(199) <= layer0_outputs(434);
    outputs(200) <= (layer0_outputs(2009)) and (layer0_outputs(908));
    outputs(201) <= (layer0_outputs(3800)) xor (layer0_outputs(574));
    outputs(202) <= not((layer0_outputs(2947)) or (layer0_outputs(4423)));
    outputs(203) <= layer0_outputs(3742);
    outputs(204) <= not(layer0_outputs(2674));
    outputs(205) <= not(layer0_outputs(462));
    outputs(206) <= layer0_outputs(1547);
    outputs(207) <= not(layer0_outputs(9)) or (layer0_outputs(2510));
    outputs(208) <= layer0_outputs(2519);
    outputs(209) <= (layer0_outputs(3404)) and not (layer0_outputs(1090));
    outputs(210) <= not(layer0_outputs(136));
    outputs(211) <= (layer0_outputs(2413)) and not (layer0_outputs(3384));
    outputs(212) <= layer0_outputs(4063);
    outputs(213) <= not(layer0_outputs(1342)) or (layer0_outputs(3922));
    outputs(214) <= not((layer0_outputs(3069)) and (layer0_outputs(2232)));
    outputs(215) <= layer0_outputs(132);
    outputs(216) <= (layer0_outputs(4592)) and not (layer0_outputs(2730));
    outputs(217) <= layer0_outputs(2677);
    outputs(218) <= (layer0_outputs(2980)) and (layer0_outputs(572));
    outputs(219) <= not((layer0_outputs(3355)) xor (layer0_outputs(311)));
    outputs(220) <= not(layer0_outputs(1123));
    outputs(221) <= layer0_outputs(1012);
    outputs(222) <= not(layer0_outputs(3894));
    outputs(223) <= not(layer0_outputs(1244)) or (layer0_outputs(4950));
    outputs(224) <= not((layer0_outputs(303)) xor (layer0_outputs(4837)));
    outputs(225) <= not((layer0_outputs(4925)) and (layer0_outputs(4557)));
    outputs(226) <= (layer0_outputs(38)) and (layer0_outputs(4412));
    outputs(227) <= layer0_outputs(747);
    outputs(228) <= not(layer0_outputs(3281));
    outputs(229) <= layer0_outputs(119);
    outputs(230) <= not(layer0_outputs(957)) or (layer0_outputs(780));
    outputs(231) <= not(layer0_outputs(2529));
    outputs(232) <= (layer0_outputs(382)) and (layer0_outputs(2720));
    outputs(233) <= not(layer0_outputs(4510));
    outputs(234) <= (layer0_outputs(2405)) and not (layer0_outputs(4182));
    outputs(235) <= not((layer0_outputs(2764)) xor (layer0_outputs(161)));
    outputs(236) <= layer0_outputs(444);
    outputs(237) <= (layer0_outputs(4951)) and not (layer0_outputs(3635));
    outputs(238) <= not((layer0_outputs(1025)) xor (layer0_outputs(73)));
    outputs(239) <= (layer0_outputs(2203)) and not (layer0_outputs(5109));
    outputs(240) <= not(layer0_outputs(4158));
    outputs(241) <= not(layer0_outputs(364));
    outputs(242) <= (layer0_outputs(1024)) and not (layer0_outputs(771));
    outputs(243) <= (layer0_outputs(451)) and not (layer0_outputs(3659));
    outputs(244) <= (layer0_outputs(257)) xor (layer0_outputs(2636));
    outputs(245) <= layer0_outputs(3588);
    outputs(246) <= not((layer0_outputs(3814)) and (layer0_outputs(1808)));
    outputs(247) <= (layer0_outputs(2797)) and not (layer0_outputs(1194));
    outputs(248) <= not((layer0_outputs(651)) or (layer0_outputs(1002)));
    outputs(249) <= layer0_outputs(3231);
    outputs(250) <= layer0_outputs(1075);
    outputs(251) <= (layer0_outputs(1871)) and (layer0_outputs(1787));
    outputs(252) <= (layer0_outputs(3861)) and not (layer0_outputs(3682));
    outputs(253) <= not(layer0_outputs(1089));
    outputs(254) <= layer0_outputs(371);
    outputs(255) <= not(layer0_outputs(2870)) or (layer0_outputs(1042));
    outputs(256) <= (layer0_outputs(1107)) or (layer0_outputs(13));
    outputs(257) <= not(layer0_outputs(2023));
    outputs(258) <= layer0_outputs(2555);
    outputs(259) <= (layer0_outputs(2380)) xor (layer0_outputs(1278));
    outputs(260) <= layer0_outputs(4454);
    outputs(261) <= not(layer0_outputs(5014));
    outputs(262) <= not(layer0_outputs(1864));
    outputs(263) <= (layer0_outputs(695)) xor (layer0_outputs(2746));
    outputs(264) <= (layer0_outputs(2384)) and not (layer0_outputs(1356));
    outputs(265) <= layer0_outputs(2146);
    outputs(266) <= layer0_outputs(2179);
    outputs(267) <= layer0_outputs(2535);
    outputs(268) <= not((layer0_outputs(3750)) xor (layer0_outputs(473)));
    outputs(269) <= (layer0_outputs(4273)) xor (layer0_outputs(3501));
    outputs(270) <= not(layer0_outputs(1854));
    outputs(271) <= not((layer0_outputs(1552)) or (layer0_outputs(4108)));
    outputs(272) <= not(layer0_outputs(2226)) or (layer0_outputs(4036));
    outputs(273) <= (layer0_outputs(3184)) or (layer0_outputs(4966));
    outputs(274) <= not((layer0_outputs(3895)) or (layer0_outputs(894)));
    outputs(275) <= not(layer0_outputs(863));
    outputs(276) <= layer0_outputs(2932);
    outputs(277) <= layer0_outputs(3318);
    outputs(278) <= (layer0_outputs(4587)) and not (layer0_outputs(2423));
    outputs(279) <= layer0_outputs(842);
    outputs(280) <= (layer0_outputs(3983)) and (layer0_outputs(2810));
    outputs(281) <= layer0_outputs(282);
    outputs(282) <= (layer0_outputs(1088)) and not (layer0_outputs(4387));
    outputs(283) <= layer0_outputs(5032);
    outputs(284) <= (layer0_outputs(1700)) and not (layer0_outputs(2930));
    outputs(285) <= layer0_outputs(1575);
    outputs(286) <= (layer0_outputs(2182)) xor (layer0_outputs(3644));
    outputs(287) <= (layer0_outputs(212)) xor (layer0_outputs(1563));
    outputs(288) <= not(layer0_outputs(1360)) or (layer0_outputs(4950));
    outputs(289) <= (layer0_outputs(2736)) and not (layer0_outputs(1461));
    outputs(290) <= layer0_outputs(844);
    outputs(291) <= not(layer0_outputs(1773)) or (layer0_outputs(1349));
    outputs(292) <= not(layer0_outputs(3654));
    outputs(293) <= not(layer0_outputs(489)) or (layer0_outputs(4020));
    outputs(294) <= (layer0_outputs(848)) and (layer0_outputs(1309));
    outputs(295) <= not(layer0_outputs(1983)) or (layer0_outputs(1597));
    outputs(296) <= not(layer0_outputs(2389)) or (layer0_outputs(235));
    outputs(297) <= not(layer0_outputs(3190));
    outputs(298) <= (layer0_outputs(2271)) and (layer0_outputs(3930));
    outputs(299) <= not(layer0_outputs(3781)) or (layer0_outputs(2352));
    outputs(300) <= not(layer0_outputs(1073));
    outputs(301) <= not((layer0_outputs(4972)) xor (layer0_outputs(2354)));
    outputs(302) <= (layer0_outputs(840)) xor (layer0_outputs(2702));
    outputs(303) <= (layer0_outputs(2676)) and not (layer0_outputs(4807));
    outputs(304) <= layer0_outputs(1023);
    outputs(305) <= not(layer0_outputs(2870)) or (layer0_outputs(2460));
    outputs(306) <= not(layer0_outputs(455));
    outputs(307) <= not(layer0_outputs(927));
    outputs(308) <= (layer0_outputs(3514)) or (layer0_outputs(735));
    outputs(309) <= (layer0_outputs(1515)) and not (layer0_outputs(1473));
    outputs(310) <= not((layer0_outputs(4766)) and (layer0_outputs(4000)));
    outputs(311) <= not(layer0_outputs(3321));
    outputs(312) <= not((layer0_outputs(3601)) xor (layer0_outputs(3354)));
    outputs(313) <= layer0_outputs(657);
    outputs(314) <= not(layer0_outputs(449));
    outputs(315) <= layer0_outputs(4552);
    outputs(316) <= not(layer0_outputs(4160)) or (layer0_outputs(1373));
    outputs(317) <= not(layer0_outputs(1944));
    outputs(318) <= layer0_outputs(2172);
    outputs(319) <= not(layer0_outputs(1441));
    outputs(320) <= not(layer0_outputs(3245)) or (layer0_outputs(557));
    outputs(321) <= layer0_outputs(160);
    outputs(322) <= (layer0_outputs(2525)) and not (layer0_outputs(3790));
    outputs(323) <= (layer0_outputs(2001)) or (layer0_outputs(22));
    outputs(324) <= not((layer0_outputs(3834)) or (layer0_outputs(895)));
    outputs(325) <= layer0_outputs(700);
    outputs(326) <= not(layer0_outputs(5114)) or (layer0_outputs(1851));
    outputs(327) <= not((layer0_outputs(125)) xor (layer0_outputs(2274)));
    outputs(328) <= not(layer0_outputs(777));
    outputs(329) <= not(layer0_outputs(2588)) or (layer0_outputs(367));
    outputs(330) <= layer0_outputs(29);
    outputs(331) <= not((layer0_outputs(3345)) or (layer0_outputs(3694)));
    outputs(332) <= not((layer0_outputs(5105)) or (layer0_outputs(1154)));
    outputs(333) <= layer0_outputs(4443);
    outputs(334) <= layer0_outputs(3927);
    outputs(335) <= not((layer0_outputs(709)) and (layer0_outputs(4913)));
    outputs(336) <= not((layer0_outputs(3401)) xor (layer0_outputs(5005)));
    outputs(337) <= layer0_outputs(1271);
    outputs(338) <= not(layer0_outputs(1568)) or (layer0_outputs(441));
    outputs(339) <= (layer0_outputs(625)) or (layer0_outputs(3784));
    outputs(340) <= layer0_outputs(2020);
    outputs(341) <= (layer0_outputs(1340)) and (layer0_outputs(744));
    outputs(342) <= not(layer0_outputs(781));
    outputs(343) <= layer0_outputs(2194);
    outputs(344) <= not(layer0_outputs(1097));
    outputs(345) <= layer0_outputs(4051);
    outputs(346) <= not(layer0_outputs(4103)) or (layer0_outputs(1871));
    outputs(347) <= (layer0_outputs(1697)) and not (layer0_outputs(573));
    outputs(348) <= not(layer0_outputs(239)) or (layer0_outputs(2901));
    outputs(349) <= (layer0_outputs(1840)) or (layer0_outputs(870));
    outputs(350) <= layer0_outputs(521);
    outputs(351) <= not((layer0_outputs(4258)) or (layer0_outputs(1124)));
    outputs(352) <= layer0_outputs(3343);
    outputs(353) <= not(layer0_outputs(4779));
    outputs(354) <= not(layer0_outputs(1201));
    outputs(355) <= not(layer0_outputs(4327));
    outputs(356) <= not(layer0_outputs(4451));
    outputs(357) <= not(layer0_outputs(5088));
    outputs(358) <= not((layer0_outputs(218)) and (layer0_outputs(3366)));
    outputs(359) <= layer0_outputs(3423);
    outputs(360) <= not(layer0_outputs(3418));
    outputs(361) <= not(layer0_outputs(92));
    outputs(362) <= (layer0_outputs(3480)) and (layer0_outputs(4762));
    outputs(363) <= (layer0_outputs(2269)) and not (layer0_outputs(400));
    outputs(364) <= (layer0_outputs(1808)) xor (layer0_outputs(1935));
    outputs(365) <= not(layer0_outputs(267));
    outputs(366) <= layer0_outputs(725);
    outputs(367) <= not(layer0_outputs(2762));
    outputs(368) <= layer0_outputs(4598);
    outputs(369) <= (layer0_outputs(3644)) or (layer0_outputs(5007));
    outputs(370) <= layer0_outputs(4446);
    outputs(371) <= (layer0_outputs(4714)) and (layer0_outputs(2043));
    outputs(372) <= (layer0_outputs(2902)) and not (layer0_outputs(2188));
    outputs(373) <= (layer0_outputs(1084)) or (layer0_outputs(113));
    outputs(374) <= not(layer0_outputs(4691));
    outputs(375) <= (layer0_outputs(4050)) and not (layer0_outputs(1233));
    outputs(376) <= not(layer0_outputs(3811));
    outputs(377) <= layer0_outputs(575);
    outputs(378) <= not(layer0_outputs(587)) or (layer0_outputs(2784));
    outputs(379) <= (layer0_outputs(948)) and not (layer0_outputs(3655));
    outputs(380) <= not((layer0_outputs(2836)) or (layer0_outputs(2386)));
    outputs(381) <= (layer0_outputs(229)) or (layer0_outputs(4723));
    outputs(382) <= not((layer0_outputs(716)) or (layer0_outputs(584)));
    outputs(383) <= (layer0_outputs(4680)) and not (layer0_outputs(1950));
    outputs(384) <= not((layer0_outputs(3744)) and (layer0_outputs(14)));
    outputs(385) <= not((layer0_outputs(1093)) and (layer0_outputs(553)));
    outputs(386) <= not(layer0_outputs(1452));
    outputs(387) <= not(layer0_outputs(4700));
    outputs(388) <= layer0_outputs(5009);
    outputs(389) <= layer0_outputs(1293);
    outputs(390) <= not(layer0_outputs(951)) or (layer0_outputs(2959));
    outputs(391) <= layer0_outputs(5036);
    outputs(392) <= layer0_outputs(2737);
    outputs(393) <= not(layer0_outputs(1322));
    outputs(394) <= not(layer0_outputs(2539));
    outputs(395) <= (layer0_outputs(2918)) and not (layer0_outputs(295));
    outputs(396) <= not(layer0_outputs(346));
    outputs(397) <= (layer0_outputs(918)) and not (layer0_outputs(3490));
    outputs(398) <= (layer0_outputs(3703)) and not (layer0_outputs(1028));
    outputs(399) <= not(layer0_outputs(626));
    outputs(400) <= not(layer0_outputs(393)) or (layer0_outputs(1565));
    outputs(401) <= (layer0_outputs(1676)) and (layer0_outputs(5007));
    outputs(402) <= not(layer0_outputs(2793));
    outputs(403) <= layer0_outputs(4352);
    outputs(404) <= not(layer0_outputs(2884));
    outputs(405) <= not((layer0_outputs(1503)) and (layer0_outputs(4917)));
    outputs(406) <= layer0_outputs(1207);
    outputs(407) <= not((layer0_outputs(907)) xor (layer0_outputs(3137)));
    outputs(408) <= not(layer0_outputs(612)) or (layer0_outputs(3827));
    outputs(409) <= (layer0_outputs(2280)) or (layer0_outputs(2821));
    outputs(410) <= not(layer0_outputs(4233)) or (layer0_outputs(2714));
    outputs(411) <= (layer0_outputs(4640)) or (layer0_outputs(37));
    outputs(412) <= layer0_outputs(1899);
    outputs(413) <= (layer0_outputs(1083)) xor (layer0_outputs(3605));
    outputs(414) <= not((layer0_outputs(4466)) or (layer0_outputs(4752)));
    outputs(415) <= (layer0_outputs(4431)) and (layer0_outputs(2306));
    outputs(416) <= layer0_outputs(3231);
    outputs(417) <= (layer0_outputs(4886)) and (layer0_outputs(2722));
    outputs(418) <= layer0_outputs(2970);
    outputs(419) <= layer0_outputs(396);
    outputs(420) <= not(layer0_outputs(455));
    outputs(421) <= not((layer0_outputs(2604)) or (layer0_outputs(141)));
    outputs(422) <= not(layer0_outputs(3561)) or (layer0_outputs(99));
    outputs(423) <= not(layer0_outputs(837)) or (layer0_outputs(2781));
    outputs(424) <= not(layer0_outputs(2964));
    outputs(425) <= not(layer0_outputs(3558));
    outputs(426) <= (layer0_outputs(4714)) and not (layer0_outputs(4947));
    outputs(427) <= layer0_outputs(4067);
    outputs(428) <= not((layer0_outputs(5094)) or (layer0_outputs(646)));
    outputs(429) <= (layer0_outputs(152)) xor (layer0_outputs(655));
    outputs(430) <= (layer0_outputs(833)) or (layer0_outputs(4231));
    outputs(431) <= layer0_outputs(4009);
    outputs(432) <= not((layer0_outputs(2856)) or (layer0_outputs(4939)));
    outputs(433) <= (layer0_outputs(2479)) or (layer0_outputs(3355));
    outputs(434) <= layer0_outputs(2519);
    outputs(435) <= layer0_outputs(3475);
    outputs(436) <= not(layer0_outputs(4891)) or (layer0_outputs(3436));
    outputs(437) <= (layer0_outputs(1949)) and not (layer0_outputs(1108));
    outputs(438) <= (layer0_outputs(1974)) and not (layer0_outputs(493));
    outputs(439) <= (layer0_outputs(4063)) or (layer0_outputs(2035));
    outputs(440) <= (layer0_outputs(906)) and (layer0_outputs(2840));
    outputs(441) <= not((layer0_outputs(1928)) and (layer0_outputs(4347)));
    outputs(442) <= layer0_outputs(1657);
    outputs(443) <= not(layer0_outputs(2166));
    outputs(444) <= not(layer0_outputs(3251));
    outputs(445) <= not(layer0_outputs(2861));
    outputs(446) <= (layer0_outputs(3250)) xor (layer0_outputs(2451));
    outputs(447) <= not(layer0_outputs(4261));
    outputs(448) <= layer0_outputs(3340);
    outputs(449) <= (layer0_outputs(2631)) and not (layer0_outputs(193));
    outputs(450) <= not(layer0_outputs(1623));
    outputs(451) <= not(layer0_outputs(3631)) or (layer0_outputs(2713));
    outputs(452) <= not(layer0_outputs(1509));
    outputs(453) <= not(layer0_outputs(878));
    outputs(454) <= layer0_outputs(706);
    outputs(455) <= layer0_outputs(2812);
    outputs(456) <= not(layer0_outputs(4497)) or (layer0_outputs(256));
    outputs(457) <= layer0_outputs(5056);
    outputs(458) <= (layer0_outputs(3688)) and not (layer0_outputs(4989));
    outputs(459) <= not((layer0_outputs(4787)) and (layer0_outputs(1217)));
    outputs(460) <= (layer0_outputs(4286)) and (layer0_outputs(3949));
    outputs(461) <= not(layer0_outputs(507));
    outputs(462) <= not(layer0_outputs(931));
    outputs(463) <= (layer0_outputs(2229)) and not (layer0_outputs(2311));
    outputs(464) <= layer0_outputs(1892);
    outputs(465) <= (layer0_outputs(2101)) or (layer0_outputs(3066));
    outputs(466) <= not((layer0_outputs(1303)) and (layer0_outputs(3958)));
    outputs(467) <= not((layer0_outputs(751)) xor (layer0_outputs(4782)));
    outputs(468) <= not(layer0_outputs(2717)) or (layer0_outputs(2673));
    outputs(469) <= layer0_outputs(4246);
    outputs(470) <= not(layer0_outputs(878));
    outputs(471) <= layer0_outputs(4417);
    outputs(472) <= (layer0_outputs(4660)) and not (layer0_outputs(3446));
    outputs(473) <= (layer0_outputs(3602)) and (layer0_outputs(2210));
    outputs(474) <= not(layer0_outputs(194)) or (layer0_outputs(2086));
    outputs(475) <= (layer0_outputs(548)) and not (layer0_outputs(3094));
    outputs(476) <= layer0_outputs(3512);
    outputs(477) <= (layer0_outputs(2625)) and not (layer0_outputs(4497));
    outputs(478) <= not(layer0_outputs(4884));
    outputs(479) <= (layer0_outputs(3714)) and not (layer0_outputs(4698));
    outputs(480) <= layer0_outputs(929);
    outputs(481) <= not(layer0_outputs(1778)) or (layer0_outputs(2676));
    outputs(482) <= layer0_outputs(2307);
    outputs(483) <= layer0_outputs(4505);
    outputs(484) <= not(layer0_outputs(684));
    outputs(485) <= layer0_outputs(983);
    outputs(486) <= layer0_outputs(2410);
    outputs(487) <= (layer0_outputs(561)) and (layer0_outputs(3627));
    outputs(488) <= (layer0_outputs(4488)) and (layer0_outputs(2900));
    outputs(489) <= not((layer0_outputs(2752)) and (layer0_outputs(3771)));
    outputs(490) <= layer0_outputs(540);
    outputs(491) <= layer0_outputs(3645);
    outputs(492) <= (layer0_outputs(3236)) or (layer0_outputs(1206));
    outputs(493) <= layer0_outputs(2935);
    outputs(494) <= not((layer0_outputs(4143)) or (layer0_outputs(3776)));
    outputs(495) <= (layer0_outputs(1145)) xor (layer0_outputs(2220));
    outputs(496) <= not(layer0_outputs(4738));
    outputs(497) <= not((layer0_outputs(4783)) or (layer0_outputs(3940)));
    outputs(498) <= not(layer0_outputs(300)) or (layer0_outputs(2242));
    outputs(499) <= not(layer0_outputs(5034));
    outputs(500) <= (layer0_outputs(4959)) and not (layer0_outputs(2091));
    outputs(501) <= layer0_outputs(3736);
    outputs(502) <= not(layer0_outputs(432)) or (layer0_outputs(4618));
    outputs(503) <= (layer0_outputs(3684)) and not (layer0_outputs(4576));
    outputs(504) <= not(layer0_outputs(3018));
    outputs(505) <= not((layer0_outputs(275)) or (layer0_outputs(4854)));
    outputs(506) <= not(layer0_outputs(48));
    outputs(507) <= layer0_outputs(4897);
    outputs(508) <= not(layer0_outputs(3673));
    outputs(509) <= (layer0_outputs(3353)) and not (layer0_outputs(1508));
    outputs(510) <= (layer0_outputs(2329)) or (layer0_outputs(4106));
    outputs(511) <= (layer0_outputs(3653)) and (layer0_outputs(3363));
    outputs(512) <= not((layer0_outputs(1421)) xor (layer0_outputs(2450)));
    outputs(513) <= '0';
    outputs(514) <= (layer0_outputs(2790)) and not (layer0_outputs(2435));
    outputs(515) <= (layer0_outputs(4855)) and not (layer0_outputs(286));
    outputs(516) <= not((layer0_outputs(186)) xor (layer0_outputs(226)));
    outputs(517) <= not(layer0_outputs(4944));
    outputs(518) <= (layer0_outputs(3316)) and not (layer0_outputs(3829));
    outputs(519) <= (layer0_outputs(1817)) and (layer0_outputs(487));
    outputs(520) <= (layer0_outputs(5059)) and not (layer0_outputs(89));
    outputs(521) <= (layer0_outputs(4842)) xor (layer0_outputs(3498));
    outputs(522) <= (layer0_outputs(4338)) and (layer0_outputs(4994));
    outputs(523) <= not((layer0_outputs(3033)) or (layer0_outputs(4958)));
    outputs(524) <= not((layer0_outputs(4930)) or (layer0_outputs(1554)));
    outputs(525) <= not((layer0_outputs(3308)) or (layer0_outputs(1806)));
    outputs(526) <= (layer0_outputs(102)) xor (layer0_outputs(1077));
    outputs(527) <= (layer0_outputs(2909)) and (layer0_outputs(829));
    outputs(528) <= (layer0_outputs(846)) and not (layer0_outputs(1510));
    outputs(529) <= (layer0_outputs(1736)) and not (layer0_outputs(5039));
    outputs(530) <= not((layer0_outputs(2304)) or (layer0_outputs(1070)));
    outputs(531) <= (layer0_outputs(554)) and not (layer0_outputs(3562));
    outputs(532) <= (layer0_outputs(1250)) and not (layer0_outputs(2512));
    outputs(533) <= (layer0_outputs(3084)) and not (layer0_outputs(2726));
    outputs(534) <= (layer0_outputs(4566)) and (layer0_outputs(3245));
    outputs(535) <= (layer0_outputs(1839)) xor (layer0_outputs(1014));
    outputs(536) <= (layer0_outputs(2983)) and not (layer0_outputs(1071));
    outputs(537) <= not((layer0_outputs(2400)) or (layer0_outputs(1793)));
    outputs(538) <= not((layer0_outputs(2212)) or (layer0_outputs(4575)));
    outputs(539) <= not((layer0_outputs(3191)) or (layer0_outputs(3093)));
    outputs(540) <= layer0_outputs(2546);
    outputs(541) <= not((layer0_outputs(1857)) xor (layer0_outputs(312)));
    outputs(542) <= (layer0_outputs(1785)) and (layer0_outputs(2556));
    outputs(543) <= not((layer0_outputs(3126)) or (layer0_outputs(4333)));
    outputs(544) <= not((layer0_outputs(2246)) or (layer0_outputs(4213)));
    outputs(545) <= (layer0_outputs(36)) and not (layer0_outputs(4300));
    outputs(546) <= (layer0_outputs(3811)) and not (layer0_outputs(2711));
    outputs(547) <= (layer0_outputs(3706)) and not (layer0_outputs(3410));
    outputs(548) <= not((layer0_outputs(1330)) or (layer0_outputs(189)));
    outputs(549) <= (layer0_outputs(330)) and not (layer0_outputs(4856));
    outputs(550) <= layer0_outputs(3692);
    outputs(551) <= layer0_outputs(3206);
    outputs(552) <= (layer0_outputs(5117)) and not (layer0_outputs(2693));
    outputs(553) <= (layer0_outputs(754)) and not (layer0_outputs(4883));
    outputs(554) <= (layer0_outputs(1773)) and (layer0_outputs(2294));
    outputs(555) <= (layer0_outputs(3046)) and not (layer0_outputs(4847));
    outputs(556) <= layer0_outputs(4905);
    outputs(557) <= not((layer0_outputs(602)) or (layer0_outputs(1300)));
    outputs(558) <= not((layer0_outputs(3746)) or (layer0_outputs(1002)));
    outputs(559) <= not((layer0_outputs(3856)) xor (layer0_outputs(307)));
    outputs(560) <= (layer0_outputs(4653)) and not (layer0_outputs(4218));
    outputs(561) <= not((layer0_outputs(24)) or (layer0_outputs(1750)));
    outputs(562) <= not((layer0_outputs(2523)) or (layer0_outputs(2748)));
    outputs(563) <= layer0_outputs(5033);
    outputs(564) <= (layer0_outputs(3567)) and not (layer0_outputs(1034));
    outputs(565) <= (layer0_outputs(3689)) and not (layer0_outputs(2027));
    outputs(566) <= (layer0_outputs(3873)) and not (layer0_outputs(3653));
    outputs(567) <= (layer0_outputs(2292)) and not (layer0_outputs(1853));
    outputs(568) <= not((layer0_outputs(2613)) or (layer0_outputs(2680)));
    outputs(569) <= '0';
    outputs(570) <= not((layer0_outputs(3307)) or (layer0_outputs(761)));
    outputs(571) <= layer0_outputs(2751);
    outputs(572) <= (layer0_outputs(888)) and not (layer0_outputs(2042));
    outputs(573) <= (layer0_outputs(1890)) and not (layer0_outputs(3531));
    outputs(574) <= (layer0_outputs(4490)) and not (layer0_outputs(4239));
    outputs(575) <= (layer0_outputs(3162)) and not (layer0_outputs(1798));
    outputs(576) <= '0';
    outputs(577) <= not(layer0_outputs(5044));
    outputs(578) <= (layer0_outputs(1035)) and not (layer0_outputs(893));
    outputs(579) <= not((layer0_outputs(3534)) or (layer0_outputs(4218)));
    outputs(580) <= not((layer0_outputs(4883)) or (layer0_outputs(2540)));
    outputs(581) <= not(layer0_outputs(3614));
    outputs(582) <= (layer0_outputs(1246)) and not (layer0_outputs(3909));
    outputs(583) <= (layer0_outputs(2645)) xor (layer0_outputs(1951));
    outputs(584) <= layer0_outputs(4528);
    outputs(585) <= not((layer0_outputs(998)) or (layer0_outputs(179)));
    outputs(586) <= (layer0_outputs(59)) and not (layer0_outputs(1799));
    outputs(587) <= (layer0_outputs(2857)) and not (layer0_outputs(3177));
    outputs(588) <= not((layer0_outputs(669)) or (layer0_outputs(108)));
    outputs(589) <= (layer0_outputs(3456)) and not (layer0_outputs(372));
    outputs(590) <= not((layer0_outputs(1222)) xor (layer0_outputs(978)));
    outputs(591) <= not(layer0_outputs(4289));
    outputs(592) <= (layer0_outputs(5018)) and not (layer0_outputs(1668));
    outputs(593) <= not((layer0_outputs(4127)) xor (layer0_outputs(3417)));
    outputs(594) <= (layer0_outputs(3130)) and (layer0_outputs(2240));
    outputs(595) <= not((layer0_outputs(4748)) or (layer0_outputs(3683)));
    outputs(596) <= layer0_outputs(1932);
    outputs(597) <= not((layer0_outputs(2050)) or (layer0_outputs(2634)));
    outputs(598) <= (layer0_outputs(681)) and (layer0_outputs(4310));
    outputs(599) <= (layer0_outputs(4688)) and not (layer0_outputs(3579));
    outputs(600) <= (layer0_outputs(4563)) and not (layer0_outputs(2273));
    outputs(601) <= (layer0_outputs(2904)) and not (layer0_outputs(2500));
    outputs(602) <= not((layer0_outputs(4652)) or (layer0_outputs(1795)));
    outputs(603) <= layer0_outputs(1085);
    outputs(604) <= layer0_outputs(326);
    outputs(605) <= not((layer0_outputs(4671)) or (layer0_outputs(2491)));
    outputs(606) <= (layer0_outputs(4402)) and (layer0_outputs(628));
    outputs(607) <= not((layer0_outputs(615)) xor (layer0_outputs(734)));
    outputs(608) <= not(layer0_outputs(2883));
    outputs(609) <= not((layer0_outputs(3188)) or (layer0_outputs(6)));
    outputs(610) <= (layer0_outputs(2936)) and not (layer0_outputs(2787));
    outputs(611) <= not(layer0_outputs(1585));
    outputs(612) <= (layer0_outputs(1262)) and not (layer0_outputs(1798));
    outputs(613) <= (layer0_outputs(4042)) and not (layer0_outputs(4372));
    outputs(614) <= (layer0_outputs(3726)) and not (layer0_outputs(5012));
    outputs(615) <= (layer0_outputs(1234)) and not (layer0_outputs(3620));
    outputs(616) <= not((layer0_outputs(534)) or (layer0_outputs(2686)));
    outputs(617) <= layer0_outputs(3444);
    outputs(618) <= layer0_outputs(3284);
    outputs(619) <= (layer0_outputs(2094)) and (layer0_outputs(937));
    outputs(620) <= not(layer0_outputs(3152));
    outputs(621) <= not(layer0_outputs(2538));
    outputs(622) <= (layer0_outputs(2213)) xor (layer0_outputs(2306));
    outputs(623) <= (layer0_outputs(3965)) and (layer0_outputs(3401));
    outputs(624) <= (layer0_outputs(2280)) xor (layer0_outputs(4030));
    outputs(625) <= layer0_outputs(1085);
    outputs(626) <= (layer0_outputs(2751)) and not (layer0_outputs(4066));
    outputs(627) <= (layer0_outputs(508)) and not (layer0_outputs(2422));
    outputs(628) <= (layer0_outputs(2956)) and not (layer0_outputs(3177));
    outputs(629) <= (layer0_outputs(3758)) xor (layer0_outputs(3542));
    outputs(630) <= (layer0_outputs(4785)) and (layer0_outputs(4647));
    outputs(631) <= (layer0_outputs(2667)) and (layer0_outputs(1302));
    outputs(632) <= (layer0_outputs(1768)) and not (layer0_outputs(271));
    outputs(633) <= layer0_outputs(2495);
    outputs(634) <= (layer0_outputs(1064)) and not (layer0_outputs(4970));
    outputs(635) <= not((layer0_outputs(291)) or (layer0_outputs(3998)));
    outputs(636) <= layer0_outputs(2653);
    outputs(637) <= (layer0_outputs(1764)) and (layer0_outputs(4095));
    outputs(638) <= not(layer0_outputs(3436));
    outputs(639) <= (layer0_outputs(2531)) and (layer0_outputs(4809));
    outputs(640) <= not((layer0_outputs(2554)) or (layer0_outputs(84)));
    outputs(641) <= (layer0_outputs(1584)) and not (layer0_outputs(678));
    outputs(642) <= not(layer0_outputs(3430));
    outputs(643) <= not((layer0_outputs(446)) or (layer0_outputs(90)));
    outputs(644) <= not(layer0_outputs(986));
    outputs(645) <= not(layer0_outputs(641));
    outputs(646) <= not(layer0_outputs(2734)) or (layer0_outputs(3298));
    outputs(647) <= not((layer0_outputs(1750)) xor (layer0_outputs(364)));
    outputs(648) <= layer0_outputs(1815);
    outputs(649) <= (layer0_outputs(2909)) and not (layer0_outputs(4151));
    outputs(650) <= not(layer0_outputs(2227));
    outputs(651) <= not((layer0_outputs(4704)) or (layer0_outputs(2254)));
    outputs(652) <= (layer0_outputs(2415)) and not (layer0_outputs(532));
    outputs(653) <= (layer0_outputs(1627)) xor (layer0_outputs(2453));
    outputs(654) <= (layer0_outputs(3923)) and not (layer0_outputs(1728));
    outputs(655) <= (layer0_outputs(4112)) and not (layer0_outputs(254));
    outputs(656) <= (layer0_outputs(232)) and (layer0_outputs(3928));
    outputs(657) <= (layer0_outputs(812)) and (layer0_outputs(1588));
    outputs(658) <= (layer0_outputs(3174)) and (layer0_outputs(2169));
    outputs(659) <= (layer0_outputs(739)) and not (layer0_outputs(1887));
    outputs(660) <= not((layer0_outputs(2419)) or (layer0_outputs(3817)));
    outputs(661) <= layer0_outputs(1611);
    outputs(662) <= (layer0_outputs(2507)) and not (layer0_outputs(2063));
    outputs(663) <= not((layer0_outputs(2919)) or (layer0_outputs(81)));
    outputs(664) <= (layer0_outputs(1707)) and (layer0_outputs(782));
    outputs(665) <= (layer0_outputs(2632)) and (layer0_outputs(3450));
    outputs(666) <= layer0_outputs(967);
    outputs(667) <= (layer0_outputs(3821)) and (layer0_outputs(1205));
    outputs(668) <= not(layer0_outputs(4092));
    outputs(669) <= (layer0_outputs(3111)) and not (layer0_outputs(1276));
    outputs(670) <= (layer0_outputs(3538)) and (layer0_outputs(3143));
    outputs(671) <= (layer0_outputs(1660)) and (layer0_outputs(565));
    outputs(672) <= (layer0_outputs(675)) and not (layer0_outputs(1606));
    outputs(673) <= (layer0_outputs(2041)) and not (layer0_outputs(1473));
    outputs(674) <= not((layer0_outputs(2551)) or (layer0_outputs(1261)));
    outputs(675) <= not(layer0_outputs(4382));
    outputs(676) <= not((layer0_outputs(3299)) or (layer0_outputs(2533)));
    outputs(677) <= (layer0_outputs(2369)) and not (layer0_outputs(3574));
    outputs(678) <= (layer0_outputs(2671)) and (layer0_outputs(4238));
    outputs(679) <= not(layer0_outputs(3953));
    outputs(680) <= (layer0_outputs(2499)) and not (layer0_outputs(3515));
    outputs(681) <= (layer0_outputs(1003)) and not (layer0_outputs(5041));
    outputs(682) <= (layer0_outputs(2715)) and (layer0_outputs(329));
    outputs(683) <= (layer0_outputs(2199)) and not (layer0_outputs(5037));
    outputs(684) <= (layer0_outputs(580)) and not (layer0_outputs(1048));
    outputs(685) <= (layer0_outputs(497)) xor (layer0_outputs(4367));
    outputs(686) <= not((layer0_outputs(4229)) or (layer0_outputs(2446)));
    outputs(687) <= '0';
    outputs(688) <= not((layer0_outputs(2406)) or (layer0_outputs(3032)));
    outputs(689) <= (layer0_outputs(807)) xor (layer0_outputs(1416));
    outputs(690) <= (layer0_outputs(1051)) and not (layer0_outputs(4781));
    outputs(691) <= (layer0_outputs(1298)) and (layer0_outputs(1829));
    outputs(692) <= (layer0_outputs(2388)) and not (layer0_outputs(787));
    outputs(693) <= (layer0_outputs(3819)) and not (layer0_outputs(3117));
    outputs(694) <= not(layer0_outputs(4762));
    outputs(695) <= (layer0_outputs(2385)) and not (layer0_outputs(4822));
    outputs(696) <= (layer0_outputs(1286)) and not (layer0_outputs(4865));
    outputs(697) <= not((layer0_outputs(3315)) or (layer0_outputs(3785)));
    outputs(698) <= (layer0_outputs(4519)) and (layer0_outputs(4797));
    outputs(699) <= (layer0_outputs(4699)) and (layer0_outputs(3207));
    outputs(700) <= layer0_outputs(4629);
    outputs(701) <= not((layer0_outputs(2885)) or (layer0_outputs(2045)));
    outputs(702) <= (layer0_outputs(213)) and (layer0_outputs(4774));
    outputs(703) <= (layer0_outputs(3844)) and not (layer0_outputs(2024));
    outputs(704) <= not((layer0_outputs(4006)) xor (layer0_outputs(2502)));
    outputs(705) <= layer0_outputs(3413);
    outputs(706) <= (layer0_outputs(1275)) and not (layer0_outputs(4527));
    outputs(707) <= (layer0_outputs(2849)) and not (layer0_outputs(2321));
    outputs(708) <= not(layer0_outputs(1818));
    outputs(709) <= (layer0_outputs(4661)) and not (layer0_outputs(4234));
    outputs(710) <= (layer0_outputs(4707)) and (layer0_outputs(4532));
    outputs(711) <= not((layer0_outputs(2126)) or (layer0_outputs(4213)));
    outputs(712) <= (layer0_outputs(4882)) and not (layer0_outputs(1715));
    outputs(713) <= (layer0_outputs(4020)) and not (layer0_outputs(2635));
    outputs(714) <= (layer0_outputs(4824)) and (layer0_outputs(3601));
    outputs(715) <= not(layer0_outputs(2067));
    outputs(716) <= layer0_outputs(1044);
    outputs(717) <= (layer0_outputs(1677)) and (layer0_outputs(3074));
    outputs(718) <= (layer0_outputs(2443)) and not (layer0_outputs(4746));
    outputs(719) <= (layer0_outputs(5027)) and not (layer0_outputs(4514));
    outputs(720) <= (layer0_outputs(515)) and not (layer0_outputs(3881));
    outputs(721) <= (layer0_outputs(2361)) and not (layer0_outputs(4458));
    outputs(722) <= not((layer0_outputs(1059)) or (layer0_outputs(4428)));
    outputs(723) <= (layer0_outputs(2600)) and (layer0_outputs(3229));
    outputs(724) <= (layer0_outputs(360)) and (layer0_outputs(4000));
    outputs(725) <= not((layer0_outputs(3378)) xor (layer0_outputs(142)));
    outputs(726) <= (layer0_outputs(4860)) and not (layer0_outputs(4091));
    outputs(727) <= (layer0_outputs(1358)) and (layer0_outputs(1159));
    outputs(728) <= not(layer0_outputs(2137));
    outputs(729) <= (layer0_outputs(2922)) and not (layer0_outputs(3664));
    outputs(730) <= layer0_outputs(3538);
    outputs(731) <= (layer0_outputs(2623)) and not (layer0_outputs(2703));
    outputs(732) <= not((layer0_outputs(2170)) or (layer0_outputs(2136)));
    outputs(733) <= (layer0_outputs(1064)) and not (layer0_outputs(2222));
    outputs(734) <= not((layer0_outputs(4732)) or (layer0_outputs(4091)));
    outputs(735) <= (layer0_outputs(5028)) and not (layer0_outputs(65));
    outputs(736) <= layer0_outputs(1351);
    outputs(737) <= (layer0_outputs(4364)) and not (layer0_outputs(2371));
    outputs(738) <= (layer0_outputs(1709)) and not (layer0_outputs(1092));
    outputs(739) <= (layer0_outputs(728)) and not (layer0_outputs(1369));
    outputs(740) <= (layer0_outputs(300)) and not (layer0_outputs(4657));
    outputs(741) <= not((layer0_outputs(4535)) or (layer0_outputs(3257)));
    outputs(742) <= (layer0_outputs(182)) and (layer0_outputs(4988));
    outputs(743) <= (layer0_outputs(3229)) and not (layer0_outputs(3511));
    outputs(744) <= (layer0_outputs(2226)) and not (layer0_outputs(486));
    outputs(745) <= (layer0_outputs(2287)) and (layer0_outputs(2014));
    outputs(746) <= not((layer0_outputs(715)) or (layer0_outputs(2641)));
    outputs(747) <= not(layer0_outputs(336));
    outputs(748) <= (layer0_outputs(3693)) and not (layer0_outputs(2124));
    outputs(749) <= (layer0_outputs(4863)) and not (layer0_outputs(2655));
    outputs(750) <= (layer0_outputs(4545)) and not (layer0_outputs(4674));
    outputs(751) <= (layer0_outputs(2436)) and (layer0_outputs(4467));
    outputs(752) <= (layer0_outputs(4321)) and not (layer0_outputs(1876));
    outputs(753) <= not(layer0_outputs(1040));
    outputs(754) <= (layer0_outputs(2276)) and not (layer0_outputs(4705));
    outputs(755) <= not((layer0_outputs(2470)) or (layer0_outputs(405)));
    outputs(756) <= (layer0_outputs(225)) and not (layer0_outputs(2140));
    outputs(757) <= (layer0_outputs(5020)) and not (layer0_outputs(2234));
    outputs(758) <= not((layer0_outputs(518)) or (layer0_outputs(4529)));
    outputs(759) <= not(layer0_outputs(3703));
    outputs(760) <= (layer0_outputs(978)) and (layer0_outputs(2643));
    outputs(761) <= not(layer0_outputs(4276));
    outputs(762) <= not(layer0_outputs(3772));
    outputs(763) <= not(layer0_outputs(5108));
    outputs(764) <= not((layer0_outputs(2413)) or (layer0_outputs(3076)));
    outputs(765) <= not((layer0_outputs(2324)) or (layer0_outputs(4989)));
    outputs(766) <= not(layer0_outputs(2299)) or (layer0_outputs(2174));
    outputs(767) <= (layer0_outputs(2219)) xor (layer0_outputs(3219));
    outputs(768) <= (layer0_outputs(4879)) and not (layer0_outputs(192));
    outputs(769) <= not((layer0_outputs(2635)) or (layer0_outputs(1272)));
    outputs(770) <= (layer0_outputs(4128)) and not (layer0_outputs(4679));
    outputs(771) <= not(layer0_outputs(1086));
    outputs(772) <= (layer0_outputs(467)) and (layer0_outputs(1844));
    outputs(773) <= not(layer0_outputs(3797));
    outputs(774) <= (layer0_outputs(609)) or (layer0_outputs(5058));
    outputs(775) <= not((layer0_outputs(3214)) or (layer0_outputs(4681)));
    outputs(776) <= (layer0_outputs(1274)) xor (layer0_outputs(1383));
    outputs(777) <= not(layer0_outputs(4687)) or (layer0_outputs(376));
    outputs(778) <= (layer0_outputs(1747)) and not (layer0_outputs(245));
    outputs(779) <= not((layer0_outputs(4230)) or (layer0_outputs(779)));
    outputs(780) <= (layer0_outputs(27)) and not (layer0_outputs(3047));
    outputs(781) <= not((layer0_outputs(1958)) or (layer0_outputs(3553)));
    outputs(782) <= (layer0_outputs(1217)) and not (layer0_outputs(390));
    outputs(783) <= not((layer0_outputs(2211)) or (layer0_outputs(3104)));
    outputs(784) <= (layer0_outputs(1328)) and not (layer0_outputs(3712));
    outputs(785) <= (layer0_outputs(922)) and not (layer0_outputs(4274));
    outputs(786) <= (layer0_outputs(475)) and (layer0_outputs(1190));
    outputs(787) <= (layer0_outputs(904)) and (layer0_outputs(4863));
    outputs(788) <= (layer0_outputs(1743)) and not (layer0_outputs(3809));
    outputs(789) <= not(layer0_outputs(219));
    outputs(790) <= not((layer0_outputs(2794)) or (layer0_outputs(3415)));
    outputs(791) <= not((layer0_outputs(2268)) or (layer0_outputs(2624)));
    outputs(792) <= not((layer0_outputs(3304)) xor (layer0_outputs(1516)));
    outputs(793) <= (layer0_outputs(4440)) and (layer0_outputs(262));
    outputs(794) <= not((layer0_outputs(4021)) or (layer0_outputs(2376)));
    outputs(795) <= (layer0_outputs(1331)) and not (layer0_outputs(1597));
    outputs(796) <= not(layer0_outputs(1685));
    outputs(797) <= not((layer0_outputs(3500)) xor (layer0_outputs(4340)));
    outputs(798) <= (layer0_outputs(2437)) and (layer0_outputs(2827));
    outputs(799) <= (layer0_outputs(613)) and not (layer0_outputs(1098));
    outputs(800) <= not((layer0_outputs(2828)) xor (layer0_outputs(69)));
    outputs(801) <= layer0_outputs(1440);
    outputs(802) <= (layer0_outputs(2326)) and not (layer0_outputs(2261));
    outputs(803) <= '0';
    outputs(804) <= (layer0_outputs(1539)) and (layer0_outputs(2202));
    outputs(805) <= (layer0_outputs(1567)) and not (layer0_outputs(2862));
    outputs(806) <= (layer0_outputs(974)) and not (layer0_outputs(2843));
    outputs(807) <= (layer0_outputs(1238)) and (layer0_outputs(2727));
    outputs(808) <= (layer0_outputs(1644)) and not (layer0_outputs(884));
    outputs(809) <= not((layer0_outputs(4608)) or (layer0_outputs(3397)));
    outputs(810) <= (layer0_outputs(3942)) xor (layer0_outputs(605));
    outputs(811) <= (layer0_outputs(733)) and not (layer0_outputs(1042));
    outputs(812) <= (layer0_outputs(4145)) and not (layer0_outputs(2728));
    outputs(813) <= (layer0_outputs(696)) and not (layer0_outputs(4923));
    outputs(814) <= (layer0_outputs(3269)) and not (layer0_outputs(3049));
    outputs(815) <= (layer0_outputs(4508)) and not (layer0_outputs(3135));
    outputs(816) <= not((layer0_outputs(4680)) or (layer0_outputs(1842)));
    outputs(817) <= (layer0_outputs(3657)) and (layer0_outputs(4800));
    outputs(818) <= (layer0_outputs(4726)) and not (layer0_outputs(3512));
    outputs(819) <= (layer0_outputs(1180)) and not (layer0_outputs(283));
    outputs(820) <= not((layer0_outputs(804)) or (layer0_outputs(4504)));
    outputs(821) <= (layer0_outputs(1663)) and (layer0_outputs(3652));
    outputs(822) <= (layer0_outputs(4427)) xor (layer0_outputs(3918));
    outputs(823) <= not((layer0_outputs(1345)) or (layer0_outputs(1859)));
    outputs(824) <= (layer0_outputs(3775)) xor (layer0_outputs(2589));
    outputs(825) <= (layer0_outputs(3166)) and not (layer0_outputs(2260));
    outputs(826) <= (layer0_outputs(1504)) and (layer0_outputs(1076));
    outputs(827) <= (layer0_outputs(2019)) xor (layer0_outputs(4999));
    outputs(828) <= not((layer0_outputs(2599)) or (layer0_outputs(2180)));
    outputs(829) <= not(layer0_outputs(2303));
    outputs(830) <= '0';
    outputs(831) <= (layer0_outputs(3868)) and not (layer0_outputs(170));
    outputs(832) <= (layer0_outputs(4179)) and not (layer0_outputs(1294));
    outputs(833) <= not(layer0_outputs(772)) or (layer0_outputs(2445));
    outputs(834) <= not(layer0_outputs(2648));
    outputs(835) <= not((layer0_outputs(1286)) or (layer0_outputs(1956)));
    outputs(836) <= (layer0_outputs(2586)) and (layer0_outputs(33));
    outputs(837) <= (layer0_outputs(4998)) and not (layer0_outputs(3587));
    outputs(838) <= not((layer0_outputs(669)) or (layer0_outputs(2142)));
    outputs(839) <= (layer0_outputs(746)) and not (layer0_outputs(599));
    outputs(840) <= (layer0_outputs(2397)) and not (layer0_outputs(3898));
    outputs(841) <= (layer0_outputs(2900)) and not (layer0_outputs(4703));
    outputs(842) <= not((layer0_outputs(562)) xor (layer0_outputs(1112)));
    outputs(843) <= (layer0_outputs(44)) and not (layer0_outputs(2736));
    outputs(844) <= (layer0_outputs(439)) and (layer0_outputs(3635));
    outputs(845) <= not((layer0_outputs(4999)) or (layer0_outputs(2347)));
    outputs(846) <= (layer0_outputs(1463)) and (layer0_outputs(459));
    outputs(847) <= not(layer0_outputs(502));
    outputs(848) <= not(layer0_outputs(2043));
    outputs(849) <= (layer0_outputs(4777)) and not (layer0_outputs(2237));
    outputs(850) <= (layer0_outputs(1466)) and (layer0_outputs(4790));
    outputs(851) <= (layer0_outputs(3804)) and (layer0_outputs(4672));
    outputs(852) <= not((layer0_outputs(3359)) or (layer0_outputs(145)));
    outputs(853) <= (layer0_outputs(728)) and not (layer0_outputs(915));
    outputs(854) <= not((layer0_outputs(3139)) or (layer0_outputs(4781)));
    outputs(855) <= (layer0_outputs(3509)) and (layer0_outputs(3873));
    outputs(856) <= layer0_outputs(1211);
    outputs(857) <= (layer0_outputs(4190)) and not (layer0_outputs(5043));
    outputs(858) <= (layer0_outputs(4559)) and not (layer0_outputs(1636));
    outputs(859) <= not((layer0_outputs(3184)) or (layer0_outputs(2170)));
    outputs(860) <= (layer0_outputs(3034)) and (layer0_outputs(50));
    outputs(861) <= (layer0_outputs(4076)) and not (layer0_outputs(4609));
    outputs(862) <= (layer0_outputs(2899)) and not (layer0_outputs(2100));
    outputs(863) <= (layer0_outputs(2992)) and not (layer0_outputs(3908));
    outputs(864) <= not((layer0_outputs(1945)) or (layer0_outputs(197)));
    outputs(865) <= (layer0_outputs(4915)) and not (layer0_outputs(4946));
    outputs(866) <= layer0_outputs(2432);
    outputs(867) <= layer0_outputs(3837);
    outputs(868) <= (layer0_outputs(5003)) and not (layer0_outputs(1294));
    outputs(869) <= (layer0_outputs(2746)) and not (layer0_outputs(1748));
    outputs(870) <= not((layer0_outputs(2976)) or (layer0_outputs(4578)));
    outputs(871) <= (layer0_outputs(1385)) and not (layer0_outputs(2204));
    outputs(872) <= not(layer0_outputs(4027));
    outputs(873) <= '0';
    outputs(874) <= not((layer0_outputs(2595)) or (layer0_outputs(1968)));
    outputs(875) <= not((layer0_outputs(3213)) or (layer0_outputs(1855)));
    outputs(876) <= not((layer0_outputs(0)) or (layer0_outputs(1671)));
    outputs(877) <= (layer0_outputs(3316)) and not (layer0_outputs(1267));
    outputs(878) <= layer0_outputs(1975);
    outputs(879) <= (layer0_outputs(3850)) and not (layer0_outputs(3882));
    outputs(880) <= (layer0_outputs(381)) and (layer0_outputs(2173));
    outputs(881) <= (layer0_outputs(3878)) and not (layer0_outputs(3238));
    outputs(882) <= (layer0_outputs(3455)) and (layer0_outputs(2924));
    outputs(883) <= not((layer0_outputs(1013)) or (layer0_outputs(2782)));
    outputs(884) <= layer0_outputs(993);
    outputs(885) <= (layer0_outputs(3693)) and (layer0_outputs(1179));
    outputs(886) <= (layer0_outputs(494)) and (layer0_outputs(4485));
    outputs(887) <= (layer0_outputs(1869)) and not (layer0_outputs(711));
    outputs(888) <= not((layer0_outputs(1280)) or (layer0_outputs(2212)));
    outputs(889) <= (layer0_outputs(1600)) and not (layer0_outputs(4760));
    outputs(890) <= (layer0_outputs(4947)) and (layer0_outputs(1497));
    outputs(891) <= layer0_outputs(4889);
    outputs(892) <= (layer0_outputs(4155)) and (layer0_outputs(3529));
    outputs(893) <= (layer0_outputs(2669)) and (layer0_outputs(4980));
    outputs(894) <= not(layer0_outputs(2726));
    outputs(895) <= (layer0_outputs(1436)) and not (layer0_outputs(842));
    outputs(896) <= layer0_outputs(466);
    outputs(897) <= (layer0_outputs(5028)) and not (layer0_outputs(4970));
    outputs(898) <= (layer0_outputs(249)) and (layer0_outputs(683));
    outputs(899) <= (layer0_outputs(703)) and not (layer0_outputs(769));
    outputs(900) <= (layer0_outputs(3739)) and not (layer0_outputs(1882));
    outputs(901) <= not((layer0_outputs(3050)) or (layer0_outputs(541)));
    outputs(902) <= (layer0_outputs(2780)) and (layer0_outputs(3118));
    outputs(903) <= layer0_outputs(4627);
    outputs(904) <= (layer0_outputs(2637)) and not (layer0_outputs(4901));
    outputs(905) <= not((layer0_outputs(4834)) or (layer0_outputs(3031)));
    outputs(906) <= (layer0_outputs(4857)) and not (layer0_outputs(2759));
    outputs(907) <= (layer0_outputs(4913)) and not (layer0_outputs(3636));
    outputs(908) <= not((layer0_outputs(2935)) or (layer0_outputs(3518)));
    outputs(909) <= (layer0_outputs(5033)) and not (layer0_outputs(542));
    outputs(910) <= not((layer0_outputs(773)) xor (layer0_outputs(517)));
    outputs(911) <= (layer0_outputs(4606)) and not (layer0_outputs(4750));
    outputs(912) <= (layer0_outputs(2102)) and (layer0_outputs(1471));
    outputs(913) <= (layer0_outputs(4875)) and (layer0_outputs(1634));
    outputs(914) <= (layer0_outputs(3752)) and not (layer0_outputs(3642));
    outputs(915) <= (layer0_outputs(5076)) and not (layer0_outputs(1359));
    outputs(916) <= (layer0_outputs(1197)) and (layer0_outputs(458));
    outputs(917) <= not((layer0_outputs(2502)) or (layer0_outputs(3818)));
    outputs(918) <= (layer0_outputs(4104)) and not (layer0_outputs(2612));
    outputs(919) <= not(layer0_outputs(2180));
    outputs(920) <= (layer0_outputs(3180)) and (layer0_outputs(816));
    outputs(921) <= (layer0_outputs(2964)) and (layer0_outputs(2459));
    outputs(922) <= not((layer0_outputs(3927)) or (layer0_outputs(813)));
    outputs(923) <= (layer0_outputs(3707)) and not (layer0_outputs(1984));
    outputs(924) <= not((layer0_outputs(3191)) or (layer0_outputs(3488)));
    outputs(925) <= not((layer0_outputs(5103)) or (layer0_outputs(576)));
    outputs(926) <= (layer0_outputs(4484)) and not (layer0_outputs(3247));
    outputs(927) <= (layer0_outputs(4406)) and (layer0_outputs(2477));
    outputs(928) <= '0';
    outputs(929) <= not((layer0_outputs(3845)) or (layer0_outputs(90)));
    outputs(930) <= not((layer0_outputs(2411)) or (layer0_outputs(4277)));
    outputs(931) <= layer0_outputs(4726);
    outputs(932) <= (layer0_outputs(3525)) and (layer0_outputs(894));
    outputs(933) <= (layer0_outputs(3957)) and (layer0_outputs(1076));
    outputs(934) <= layer0_outputs(1512);
    outputs(935) <= layer0_outputs(3652);
    outputs(936) <= (layer0_outputs(5023)) and not (layer0_outputs(2092));
    outputs(937) <= (layer0_outputs(3872)) and (layer0_outputs(3433));
    outputs(938) <= not((layer0_outputs(3326)) or (layer0_outputs(1519)));
    outputs(939) <= (layer0_outputs(2775)) and not (layer0_outputs(4413));
    outputs(940) <= not((layer0_outputs(362)) or (layer0_outputs(1420)));
    outputs(941) <= (layer0_outputs(5099)) and (layer0_outputs(381));
    outputs(942) <= (layer0_outputs(2924)) and (layer0_outputs(452));
    outputs(943) <= (layer0_outputs(4223)) and (layer0_outputs(1411));
    outputs(944) <= not(layer0_outputs(1218));
    outputs(945) <= layer0_outputs(1395);
    outputs(946) <= not((layer0_outputs(2558)) or (layer0_outputs(966)));
    outputs(947) <= (layer0_outputs(3974)) and not (layer0_outputs(3835));
    outputs(948) <= layer0_outputs(155);
    outputs(949) <= (layer0_outputs(963)) and not (layer0_outputs(549));
    outputs(950) <= (layer0_outputs(1879)) and not (layer0_outputs(1670));
    outputs(951) <= (layer0_outputs(3048)) and (layer0_outputs(4570));
    outputs(952) <= (layer0_outputs(1001)) and (layer0_outputs(4600));
    outputs(953) <= not((layer0_outputs(3597)) or (layer0_outputs(2700)));
    outputs(954) <= (layer0_outputs(1925)) and (layer0_outputs(374));
    outputs(955) <= (layer0_outputs(4013)) and (layer0_outputs(4969));
    outputs(956) <= not((layer0_outputs(4225)) or (layer0_outputs(2721)));
    outputs(957) <= not(layer0_outputs(3755));
    outputs(958) <= (layer0_outputs(4729)) and not (layer0_outputs(2834));
    outputs(959) <= not((layer0_outputs(2281)) or (layer0_outputs(796)));
    outputs(960) <= (layer0_outputs(4849)) and (layer0_outputs(3670));
    outputs(961) <= (layer0_outputs(3658)) and not (layer0_outputs(212));
    outputs(962) <= layer0_outputs(2103);
    outputs(963) <= (layer0_outputs(4549)) and not (layer0_outputs(1219));
    outputs(964) <= (layer0_outputs(1297)) and not (layer0_outputs(3678));
    outputs(965) <= layer0_outputs(4848);
    outputs(966) <= (layer0_outputs(2337)) and not (layer0_outputs(4045));
    outputs(967) <= (layer0_outputs(342)) and not (layer0_outputs(3981));
    outputs(968) <= (layer0_outputs(348)) and not (layer0_outputs(3285));
    outputs(969) <= (layer0_outputs(1616)) and not (layer0_outputs(4649));
    outputs(970) <= (layer0_outputs(3924)) and (layer0_outputs(4195));
    outputs(971) <= (layer0_outputs(590)) and not (layer0_outputs(1652));
    outputs(972) <= layer0_outputs(2576);
    outputs(973) <= (layer0_outputs(1849)) and not (layer0_outputs(4892));
    outputs(974) <= not((layer0_outputs(1796)) or (layer0_outputs(4709)));
    outputs(975) <= (layer0_outputs(2684)) and (layer0_outputs(4961));
    outputs(976) <= (layer0_outputs(406)) and (layer0_outputs(685));
    outputs(977) <= (layer0_outputs(1846)) and not (layer0_outputs(4347));
    outputs(978) <= (layer0_outputs(172)) and not (layer0_outputs(3964));
    outputs(979) <= not((layer0_outputs(2453)) xor (layer0_outputs(2553)));
    outputs(980) <= (layer0_outputs(3735)) and (layer0_outputs(127));
    outputs(981) <= layer0_outputs(846);
    outputs(982) <= not((layer0_outputs(1548)) or (layer0_outputs(4181)));
    outputs(983) <= (layer0_outputs(4896)) and not (layer0_outputs(4821));
    outputs(984) <= layer0_outputs(4878);
    outputs(985) <= not(layer0_outputs(3891));
    outputs(986) <= not((layer0_outputs(1777)) or (layer0_outputs(3610)));
    outputs(987) <= (layer0_outputs(4135)) xor (layer0_outputs(614));
    outputs(988) <= not((layer0_outputs(999)) or (layer0_outputs(2374)));
    outputs(989) <= (layer0_outputs(3867)) and not (layer0_outputs(2283));
    outputs(990) <= (layer0_outputs(4977)) and not (layer0_outputs(3947));
    outputs(991) <= not(layer0_outputs(2277));
    outputs(992) <= not((layer0_outputs(995)) or (layer0_outputs(3879)));
    outputs(993) <= (layer0_outputs(2584)) and not (layer0_outputs(1558));
    outputs(994) <= (layer0_outputs(3250)) and not (layer0_outputs(1761));
    outputs(995) <= not((layer0_outputs(1019)) xor (layer0_outputs(339)));
    outputs(996) <= (layer0_outputs(4486)) and not (layer0_outputs(2387));
    outputs(997) <= (layer0_outputs(2481)) and not (layer0_outputs(1505));
    outputs(998) <= (layer0_outputs(2973)) and (layer0_outputs(3992));
    outputs(999) <= (layer0_outputs(4374)) and (layer0_outputs(2393));
    outputs(1000) <= not((layer0_outputs(3671)) xor (layer0_outputs(1413)));
    outputs(1001) <= (layer0_outputs(3441)) xor (layer0_outputs(3740));
    outputs(1002) <= '0';
    outputs(1003) <= (layer0_outputs(1353)) and (layer0_outputs(617));
    outputs(1004) <= layer0_outputs(3421);
    outputs(1005) <= (layer0_outputs(3386)) and (layer0_outputs(1624));
    outputs(1006) <= (layer0_outputs(27)) and not (layer0_outputs(3756));
    outputs(1007) <= not((layer0_outputs(1259)) or (layer0_outputs(3973)));
    outputs(1008) <= (layer0_outputs(329)) and not (layer0_outputs(362));
    outputs(1009) <= (layer0_outputs(4399)) and not (layer0_outputs(2833));
    outputs(1010) <= (layer0_outputs(1869)) and (layer0_outputs(2869));
    outputs(1011) <= (layer0_outputs(656)) and (layer0_outputs(2031));
    outputs(1012) <= (layer0_outputs(3088)) and not (layer0_outputs(2939));
    outputs(1013) <= not((layer0_outputs(866)) or (layer0_outputs(955)));
    outputs(1014) <= not((layer0_outputs(738)) or (layer0_outputs(4440)));
    outputs(1015) <= (layer0_outputs(3026)) and not (layer0_outputs(4079));
    outputs(1016) <= not((layer0_outputs(284)) or (layer0_outputs(3387)));
    outputs(1017) <= layer0_outputs(4022);
    outputs(1018) <= not(layer0_outputs(2901));
    outputs(1019) <= layer0_outputs(4492);
    outputs(1020) <= not((layer0_outputs(1459)) or (layer0_outputs(3121)));
    outputs(1021) <= not((layer0_outputs(2716)) or (layer0_outputs(3078)));
    outputs(1022) <= not((layer0_outputs(3043)) or (layer0_outputs(1467)));
    outputs(1023) <= layer0_outputs(3298);
    outputs(1024) <= not(layer0_outputs(112)) or (layer0_outputs(484));
    outputs(1025) <= layer0_outputs(511);
    outputs(1026) <= layer0_outputs(274);
    outputs(1027) <= not(layer0_outputs(4252));
    outputs(1028) <= (layer0_outputs(1939)) or (layer0_outputs(3552));
    outputs(1029) <= not(layer0_outputs(2145));
    outputs(1030) <= not(layer0_outputs(4337));
    outputs(1031) <= layer0_outputs(1523);
    outputs(1032) <= layer0_outputs(3160);
    outputs(1033) <= not(layer0_outputs(4067));
    outputs(1034) <= (layer0_outputs(3387)) and (layer0_outputs(425));
    outputs(1035) <= (layer0_outputs(4838)) or (layer0_outputs(3014));
    outputs(1036) <= not((layer0_outputs(3211)) and (layer0_outputs(923)));
    outputs(1037) <= (layer0_outputs(3196)) and not (layer0_outputs(1296));
    outputs(1038) <= layer0_outputs(2257);
    outputs(1039) <= not(layer0_outputs(243));
    outputs(1040) <= not(layer0_outputs(4735)) or (layer0_outputs(2316));
    outputs(1041) <= not(layer0_outputs(4976));
    outputs(1042) <= layer0_outputs(604);
    outputs(1043) <= not(layer0_outputs(4647));
    outputs(1044) <= not(layer0_outputs(4356));
    outputs(1045) <= not(layer0_outputs(3862));
    outputs(1046) <= not(layer0_outputs(730));
    outputs(1047) <= layer0_outputs(4755);
    outputs(1048) <= not(layer0_outputs(4208));
    outputs(1049) <= layer0_outputs(2541);
    outputs(1050) <= not(layer0_outputs(2258));
    outputs(1051) <= not(layer0_outputs(2651));
    outputs(1052) <= not((layer0_outputs(3058)) xor (layer0_outputs(4317)));
    outputs(1053) <= layer0_outputs(1994);
    outputs(1054) <= layer0_outputs(2531);
    outputs(1055) <= layer0_outputs(51);
    outputs(1056) <= (layer0_outputs(4955)) and not (layer0_outputs(3010));
    outputs(1057) <= layer0_outputs(2278);
    outputs(1058) <= (layer0_outputs(3452)) and (layer0_outputs(671));
    outputs(1059) <= not((layer0_outputs(941)) xor (layer0_outputs(1156)));
    outputs(1060) <= layer0_outputs(1706);
    outputs(1061) <= layer0_outputs(3481);
    outputs(1062) <= not((layer0_outputs(2812)) xor (layer0_outputs(2201)));
    outputs(1063) <= (layer0_outputs(301)) or (layer0_outputs(1061));
    outputs(1064) <= not(layer0_outputs(2271));
    outputs(1065) <= layer0_outputs(4589);
    outputs(1066) <= not((layer0_outputs(1615)) and (layer0_outputs(4299)));
    outputs(1067) <= (layer0_outputs(4840)) xor (layer0_outputs(247));
    outputs(1068) <= layer0_outputs(1163);
    outputs(1069) <= (layer0_outputs(1484)) and not (layer0_outputs(5065));
    outputs(1070) <= not(layer0_outputs(3592)) or (layer0_outputs(3971));
    outputs(1071) <= layer0_outputs(1255);
    outputs(1072) <= layer0_outputs(279);
    outputs(1073) <= not(layer0_outputs(1543));
    outputs(1074) <= not((layer0_outputs(917)) and (layer0_outputs(3933)));
    outputs(1075) <= not((layer0_outputs(2129)) or (layer0_outputs(2985)));
    outputs(1076) <= not(layer0_outputs(4325));
    outputs(1077) <= not(layer0_outputs(4512)) or (layer0_outputs(4305));
    outputs(1078) <= layer0_outputs(1319);
    outputs(1079) <= (layer0_outputs(4706)) xor (layer0_outputs(879));
    outputs(1080) <= not(layer0_outputs(492)) or (layer0_outputs(781));
    outputs(1081) <= not((layer0_outputs(4906)) and (layer0_outputs(72)));
    outputs(1082) <= (layer0_outputs(3966)) or (layer0_outputs(2157));
    outputs(1083) <= layer0_outputs(3074);
    outputs(1084) <= not(layer0_outputs(4209));
    outputs(1085) <= not(layer0_outputs(1804));
    outputs(1086) <= layer0_outputs(4755);
    outputs(1087) <= layer0_outputs(4229);
    outputs(1088) <= not(layer0_outputs(1829)) or (layer0_outputs(1352));
    outputs(1089) <= not(layer0_outputs(2051)) or (layer0_outputs(1045));
    outputs(1090) <= layer0_outputs(1958);
    outputs(1091) <= layer0_outputs(1419);
    outputs(1092) <= not(layer0_outputs(4638)) or (layer0_outputs(3432));
    outputs(1093) <= layer0_outputs(2528);
    outputs(1094) <= (layer0_outputs(2231)) and not (layer0_outputs(413));
    outputs(1095) <= not(layer0_outputs(1412));
    outputs(1096) <= layer0_outputs(4071);
    outputs(1097) <= (layer0_outputs(1709)) xor (layer0_outputs(1941));
    outputs(1098) <= (layer0_outputs(3993)) and not (layer0_outputs(424));
    outputs(1099) <= layer0_outputs(1800);
    outputs(1100) <= not(layer0_outputs(3666));
    outputs(1101) <= not(layer0_outputs(4544)) or (layer0_outputs(2524));
    outputs(1102) <= not(layer0_outputs(2217)) or (layer0_outputs(4183));
    outputs(1103) <= not(layer0_outputs(48));
    outputs(1104) <= layer0_outputs(1029);
    outputs(1105) <= (layer0_outputs(3358)) and not (layer0_outputs(4397));
    outputs(1106) <= (layer0_outputs(1788)) or (layer0_outputs(4483));
    outputs(1107) <= not((layer0_outputs(1100)) xor (layer0_outputs(4494)));
    outputs(1108) <= layer0_outputs(1534);
    outputs(1109) <= not(layer0_outputs(818));
    outputs(1110) <= (layer0_outputs(1576)) or (layer0_outputs(1009));
    outputs(1111) <= layer0_outputs(4853);
    outputs(1112) <= (layer0_outputs(3523)) and not (layer0_outputs(3141));
    outputs(1113) <= (layer0_outputs(2859)) and (layer0_outputs(3485));
    outputs(1114) <= not((layer0_outputs(3773)) or (layer0_outputs(816)));
    outputs(1115) <= layer0_outputs(1894);
    outputs(1116) <= not(layer0_outputs(3024));
    outputs(1117) <= not((layer0_outputs(1344)) and (layer0_outputs(3677)));
    outputs(1118) <= (layer0_outputs(2881)) xor (layer0_outputs(1794));
    outputs(1119) <= layer0_outputs(209);
    outputs(1120) <= not(layer0_outputs(4276));
    outputs(1121) <= (layer0_outputs(3255)) or (layer0_outputs(2368));
    outputs(1122) <= (layer0_outputs(2392)) or (layer0_outputs(1105));
    outputs(1123) <= not(layer0_outputs(4574)) or (layer0_outputs(3757));
    outputs(1124) <= layer0_outputs(4025);
    outputs(1125) <= not((layer0_outputs(445)) and (layer0_outputs(1409)));
    outputs(1126) <= not((layer0_outputs(1168)) or (layer0_outputs(710)));
    outputs(1127) <= layer0_outputs(612);
    outputs(1128) <= layer0_outputs(154);
    outputs(1129) <= (layer0_outputs(2578)) xor (layer0_outputs(4785));
    outputs(1130) <= (layer0_outputs(3372)) and not (layer0_outputs(3251));
    outputs(1131) <= layer0_outputs(619);
    outputs(1132) <= not((layer0_outputs(4109)) xor (layer0_outputs(4206)));
    outputs(1133) <= not(layer0_outputs(2187));
    outputs(1134) <= layer0_outputs(4382);
    outputs(1135) <= (layer0_outputs(2268)) xor (layer0_outputs(1720));
    outputs(1136) <= layer0_outputs(4429);
    outputs(1137) <= not((layer0_outputs(3225)) and (layer0_outputs(2223)));
    outputs(1138) <= layer0_outputs(4040);
    outputs(1139) <= not(layer0_outputs(3826));
    outputs(1140) <= layer0_outputs(3176);
    outputs(1141) <= layer0_outputs(438);
    outputs(1142) <= not((layer0_outputs(2611)) or (layer0_outputs(700)));
    outputs(1143) <= layer0_outputs(994);
    outputs(1144) <= (layer0_outputs(1414)) xor (layer0_outputs(2083));
    outputs(1145) <= not(layer0_outputs(2486));
    outputs(1146) <= not(layer0_outputs(4622));
    outputs(1147) <= not(layer0_outputs(4849));
    outputs(1148) <= not(layer0_outputs(221));
    outputs(1149) <= layer0_outputs(5017);
    outputs(1150) <= (layer0_outputs(3820)) and (layer0_outputs(806));
    outputs(1151) <= not(layer0_outputs(3437)) or (layer0_outputs(783));
    outputs(1152) <= not((layer0_outputs(3911)) and (layer0_outputs(341)));
    outputs(1153) <= (layer0_outputs(3702)) and not (layer0_outputs(4936));
    outputs(1154) <= not(layer0_outputs(3625)) or (layer0_outputs(4542));
    outputs(1155) <= (layer0_outputs(3459)) or (layer0_outputs(4447));
    outputs(1156) <= layer0_outputs(3419);
    outputs(1157) <= not((layer0_outputs(2961)) and (layer0_outputs(3547)));
    outputs(1158) <= (layer0_outputs(1251)) and (layer0_outputs(926));
    outputs(1159) <= not(layer0_outputs(4099)) or (layer0_outputs(93));
    outputs(1160) <= not(layer0_outputs(4032)) or (layer0_outputs(3694));
    outputs(1161) <= not(layer0_outputs(3602));
    outputs(1162) <= not((layer0_outputs(3621)) xor (layer0_outputs(2284)));
    outputs(1163) <= not(layer0_outputs(3027)) or (layer0_outputs(1008));
    outputs(1164) <= not((layer0_outputs(1590)) and (layer0_outputs(469)));
    outputs(1165) <= layer0_outputs(921);
    outputs(1166) <= layer0_outputs(5031);
    outputs(1167) <= not((layer0_outputs(4617)) or (layer0_outputs(1111)));
    outputs(1168) <= (layer0_outputs(4132)) and (layer0_outputs(2629));
    outputs(1169) <= not(layer0_outputs(244));
    outputs(1170) <= not(layer0_outputs(1837));
    outputs(1171) <= not(layer0_outputs(5059));
    outputs(1172) <= not(layer0_outputs(3716));
    outputs(1173) <= layer0_outputs(2070);
    outputs(1174) <= not(layer0_outputs(2130));
    outputs(1175) <= layer0_outputs(4595);
    outputs(1176) <= layer0_outputs(1439);
    outputs(1177) <= not(layer0_outputs(2131));
    outputs(1178) <= layer0_outputs(2690);
    outputs(1179) <= (layer0_outputs(3883)) xor (layer0_outputs(3975));
    outputs(1180) <= not((layer0_outputs(2772)) xor (layer0_outputs(2570)));
    outputs(1181) <= (layer0_outputs(4634)) xor (layer0_outputs(3522));
    outputs(1182) <= not(layer0_outputs(3446)) or (layer0_outputs(1140));
    outputs(1183) <= layer0_outputs(1439);
    outputs(1184) <= not(layer0_outputs(1450));
    outputs(1185) <= (layer0_outputs(4002)) and (layer0_outputs(2805));
    outputs(1186) <= layer0_outputs(206);
    outputs(1187) <= layer0_outputs(3020);
    outputs(1188) <= not(layer0_outputs(5107)) or (layer0_outputs(3866));
    outputs(1189) <= not(layer0_outputs(1775));
    outputs(1190) <= not(layer0_outputs(532)) or (layer0_outputs(2932));
    outputs(1191) <= layer0_outputs(2390);
    outputs(1192) <= not(layer0_outputs(944));
    outputs(1193) <= not(layer0_outputs(523));
    outputs(1194) <= not(layer0_outputs(2857)) or (layer0_outputs(1257));
    outputs(1195) <= not((layer0_outputs(4753)) xor (layer0_outputs(1576)));
    outputs(1196) <= not(layer0_outputs(2263));
    outputs(1197) <= layer0_outputs(1725);
    outputs(1198) <= (layer0_outputs(2252)) and (layer0_outputs(2144));
    outputs(1199) <= (layer0_outputs(2052)) or (layer0_outputs(2838));
    outputs(1200) <= not(layer0_outputs(134));
    outputs(1201) <= (layer0_outputs(4296)) and not (layer0_outputs(2297));
    outputs(1202) <= not((layer0_outputs(4099)) and (layer0_outputs(1590)));
    outputs(1203) <= layer0_outputs(2687);
    outputs(1204) <= not(layer0_outputs(4281));
    outputs(1205) <= not(layer0_outputs(213));
    outputs(1206) <= (layer0_outputs(1538)) xor (layer0_outputs(4737));
    outputs(1207) <= not(layer0_outputs(3095));
    outputs(1208) <= layer0_outputs(3537);
    outputs(1209) <= layer0_outputs(2548);
    outputs(1210) <= not(layer0_outputs(4181)) or (layer0_outputs(285));
    outputs(1211) <= layer0_outputs(4336);
    outputs(1212) <= (layer0_outputs(2278)) and not (layer0_outputs(1412));
    outputs(1213) <= layer0_outputs(4741);
    outputs(1214) <= not(layer0_outputs(1650)) or (layer0_outputs(1137));
    outputs(1215) <= not(layer0_outputs(1836)) or (layer0_outputs(2026));
    outputs(1216) <= (layer0_outputs(375)) and (layer0_outputs(4108));
    outputs(1217) <= (layer0_outputs(3700)) or (layer0_outputs(4584));
    outputs(1218) <= layer0_outputs(385);
    outputs(1219) <= not((layer0_outputs(2521)) or (layer0_outputs(2739)));
    outputs(1220) <= not((layer0_outputs(2039)) and (layer0_outputs(3721)));
    outputs(1221) <= layer0_outputs(1404);
    outputs(1222) <= not((layer0_outputs(4604)) xor (layer0_outputs(790)));
    outputs(1223) <= layer0_outputs(3893);
    outputs(1224) <= not(layer0_outputs(1729)) or (layer0_outputs(1299));
    outputs(1225) <= layer0_outputs(3626);
    outputs(1226) <= not((layer0_outputs(668)) xor (layer0_outputs(4725)));
    outputs(1227) <= not(layer0_outputs(270)) or (layer0_outputs(4186));
    outputs(1228) <= (layer0_outputs(4342)) and not (layer0_outputs(1745));
    outputs(1229) <= layer0_outputs(4167);
    outputs(1230) <= not(layer0_outputs(1908));
    outputs(1231) <= not((layer0_outputs(273)) and (layer0_outputs(1238)));
    outputs(1232) <= not(layer0_outputs(896));
    outputs(1233) <= (layer0_outputs(771)) or (layer0_outputs(1117));
    outputs(1234) <= layer0_outputs(3816);
    outputs(1235) <= not((layer0_outputs(19)) and (layer0_outputs(3386)));
    outputs(1236) <= layer0_outputs(4933);
    outputs(1237) <= layer0_outputs(2451);
    outputs(1238) <= (layer0_outputs(2183)) and (layer0_outputs(2913));
    outputs(1239) <= not((layer0_outputs(395)) and (layer0_outputs(945)));
    outputs(1240) <= (layer0_outputs(639)) or (layer0_outputs(775));
    outputs(1241) <= (layer0_outputs(1341)) or (layer0_outputs(3951));
    outputs(1242) <= (layer0_outputs(1502)) xor (layer0_outputs(428));
    outputs(1243) <= (layer0_outputs(4452)) xor (layer0_outputs(3299));
    outputs(1244) <= (layer0_outputs(2940)) and not (layer0_outputs(4130));
    outputs(1245) <= not(layer0_outputs(3669));
    outputs(1246) <= (layer0_outputs(4938)) and (layer0_outputs(1091));
    outputs(1247) <= (layer0_outputs(3702)) and (layer0_outputs(1004));
    outputs(1248) <= layer0_outputs(1714);
    outputs(1249) <= not((layer0_outputs(1065)) or (layer0_outputs(2542)));
    outputs(1250) <= not(layer0_outputs(2878));
    outputs(1251) <= not((layer0_outputs(3732)) and (layer0_outputs(559)));
    outputs(1252) <= not(layer0_outputs(158)) or (layer0_outputs(1712));
    outputs(1253) <= not((layer0_outputs(4395)) xor (layer0_outputs(1613)));
    outputs(1254) <= layer0_outputs(1336);
    outputs(1255) <= (layer0_outputs(4336)) or (layer0_outputs(3119));
    outputs(1256) <= not(layer0_outputs(1937));
    outputs(1257) <= not(layer0_outputs(992));
    outputs(1258) <= (layer0_outputs(962)) or (layer0_outputs(792));
    outputs(1259) <= not(layer0_outputs(3565));
    outputs(1260) <= layer0_outputs(138);
    outputs(1261) <= (layer0_outputs(615)) and (layer0_outputs(4157));
    outputs(1262) <= not((layer0_outputs(983)) and (layer0_outputs(2119)));
    outputs(1263) <= (layer0_outputs(2375)) xor (layer0_outputs(1770));
    outputs(1264) <= (layer0_outputs(1193)) xor (layer0_outputs(4879));
    outputs(1265) <= (layer0_outputs(96)) xor (layer0_outputs(558));
    outputs(1266) <= layer0_outputs(29);
    outputs(1267) <= not(layer0_outputs(1619));
    outputs(1268) <= not(layer0_outputs(4829));
    outputs(1269) <= (layer0_outputs(2006)) and (layer0_outputs(2517));
    outputs(1270) <= not(layer0_outputs(4577));
    outputs(1271) <= not((layer0_outputs(4075)) or (layer0_outputs(743)));
    outputs(1272) <= not(layer0_outputs(680));
    outputs(1273) <= (layer0_outputs(1205)) and not (layer0_outputs(2915));
    outputs(1274) <= layer0_outputs(1550);
    outputs(1275) <= not(layer0_outputs(2567)) or (layer0_outputs(3218));
    outputs(1276) <= not(layer0_outputs(1057));
    outputs(1277) <= not(layer0_outputs(544));
    outputs(1278) <= not(layer0_outputs(4411));
    outputs(1279) <= not((layer0_outputs(246)) or (layer0_outputs(2379)));
    outputs(1280) <= not((layer0_outputs(630)) or (layer0_outputs(1522)));
    outputs(1281) <= layer0_outputs(3620);
    outputs(1282) <= not(layer0_outputs(3414)) or (layer0_outputs(3098));
    outputs(1283) <= (layer0_outputs(4453)) or (layer0_outputs(1530));
    outputs(1284) <= not((layer0_outputs(1991)) and (layer0_outputs(4133)));
    outputs(1285) <= not(layer0_outputs(4985));
    outputs(1286) <= not((layer0_outputs(3697)) xor (layer0_outputs(4330)));
    outputs(1287) <= layer0_outputs(4102);
    outputs(1288) <= (layer0_outputs(3801)) xor (layer0_outputs(352));
    outputs(1289) <= (layer0_outputs(1463)) and (layer0_outputs(4711));
    outputs(1290) <= not(layer0_outputs(4226));
    outputs(1291) <= (layer0_outputs(4802)) and not (layer0_outputs(3381));
    outputs(1292) <= not(layer0_outputs(3568));
    outputs(1293) <= not((layer0_outputs(3582)) or (layer0_outputs(3334)));
    outputs(1294) <= not(layer0_outputs(317)) or (layer0_outputs(2141));
    outputs(1295) <= not(layer0_outputs(4568)) or (layer0_outputs(1738));
    outputs(1296) <= not(layer0_outputs(348));
    outputs(1297) <= not((layer0_outputs(1476)) or (layer0_outputs(1056)));
    outputs(1298) <= not((layer0_outputs(3334)) or (layer0_outputs(788)));
    outputs(1299) <= not((layer0_outputs(2460)) or (layer0_outputs(1681)));
    outputs(1300) <= not((layer0_outputs(132)) and (layer0_outputs(2852)));
    outputs(1301) <= not((layer0_outputs(2796)) xor (layer0_outputs(4579)));
    outputs(1302) <= (layer0_outputs(1583)) xor (layer0_outputs(2729));
    outputs(1303) <= layer0_outputs(4169);
    outputs(1304) <= layer0_outputs(1288);
    outputs(1305) <= (layer0_outputs(4826)) and (layer0_outputs(1603));
    outputs(1306) <= not(layer0_outputs(704));
    outputs(1307) <= not((layer0_outputs(3323)) or (layer0_outputs(3712)));
    outputs(1308) <= layer0_outputs(4805);
    outputs(1309) <= layer0_outputs(1455);
    outputs(1310) <= not((layer0_outputs(4124)) xor (layer0_outputs(4299)));
    outputs(1311) <= not(layer0_outputs(2324));
    outputs(1312) <= not((layer0_outputs(2484)) xor (layer0_outputs(1277)));
    outputs(1313) <= layer0_outputs(150);
    outputs(1314) <= not(layer0_outputs(3044)) or (layer0_outputs(1950));
    outputs(1315) <= layer0_outputs(4850);
    outputs(1316) <= not(layer0_outputs(3821)) or (layer0_outputs(1982));
    outputs(1317) <= not(layer0_outputs(742));
    outputs(1318) <= not(layer0_outputs(4981));
    outputs(1319) <= not(layer0_outputs(649));
    outputs(1320) <= not(layer0_outputs(2882));
    outputs(1321) <= not(layer0_outputs(1925));
    outputs(1322) <= not(layer0_outputs(5005));
    outputs(1323) <= (layer0_outputs(5074)) and not (layer0_outputs(1888));
    outputs(1324) <= (layer0_outputs(4921)) and (layer0_outputs(1017));
    outputs(1325) <= (layer0_outputs(1325)) or (layer0_outputs(953));
    outputs(1326) <= not((layer0_outputs(2096)) or (layer0_outputs(4654)));
    outputs(1327) <= layer0_outputs(2604);
    outputs(1328) <= not(layer0_outputs(56));
    outputs(1329) <= (layer0_outputs(3894)) and not (layer0_outputs(4001));
    outputs(1330) <= not(layer0_outputs(363));
    outputs(1331) <= not(layer0_outputs(1418));
    outputs(1332) <= not((layer0_outputs(3320)) and (layer0_outputs(4661)));
    outputs(1333) <= layer0_outputs(1336);
    outputs(1334) <= not(layer0_outputs(2077));
    outputs(1335) <= not((layer0_outputs(165)) or (layer0_outputs(4110)));
    outputs(1336) <= not(layer0_outputs(313)) or (layer0_outputs(4951));
    outputs(1337) <= (layer0_outputs(3267)) or (layer0_outputs(3289));
    outputs(1338) <= not(layer0_outputs(3886));
    outputs(1339) <= layer0_outputs(306);
    outputs(1340) <= layer0_outputs(3360);
    outputs(1341) <= not((layer0_outputs(3805)) or (layer0_outputs(716)));
    outputs(1342) <= not(layer0_outputs(4535));
    outputs(1343) <= (layer0_outputs(32)) and (layer0_outputs(899));
    outputs(1344) <= layer0_outputs(4689);
    outputs(1345) <= (layer0_outputs(4357)) and not (layer0_outputs(2667));
    outputs(1346) <= not((layer0_outputs(64)) and (layer0_outputs(4812)));
    outputs(1347) <= (layer0_outputs(3119)) or (layer0_outputs(2826));
    outputs(1348) <= not((layer0_outputs(354)) xor (layer0_outputs(4669)));
    outputs(1349) <= layer0_outputs(4736);
    outputs(1350) <= not((layer0_outputs(1691)) xor (layer0_outputs(1541)));
    outputs(1351) <= (layer0_outputs(220)) and not (layer0_outputs(4454));
    outputs(1352) <= layer0_outputs(4262);
    outputs(1353) <= not(layer0_outputs(3011));
    outputs(1354) <= not(layer0_outputs(2756)) or (layer0_outputs(2156));
    outputs(1355) <= layer0_outputs(1329);
    outputs(1356) <= layer0_outputs(3738);
    outputs(1357) <= not((layer0_outputs(5117)) xor (layer0_outputs(4083)));
    outputs(1358) <= layer0_outputs(5030);
    outputs(1359) <= (layer0_outputs(760)) xor (layer0_outputs(1729));
    outputs(1360) <= not(layer0_outputs(429)) or (layer0_outputs(485));
    outputs(1361) <= (layer0_outputs(5064)) xor (layer0_outputs(3900));
    outputs(1362) <= not(layer0_outputs(4664));
    outputs(1363) <= layer0_outputs(4293);
    outputs(1364) <= not(layer0_outputs(3786));
    outputs(1365) <= layer0_outputs(2804);
    outputs(1366) <= (layer0_outputs(1090)) and not (layer0_outputs(990));
    outputs(1367) <= (layer0_outputs(5108)) or (layer0_outputs(3615));
    outputs(1368) <= not(layer0_outputs(4543));
    outputs(1369) <= layer0_outputs(4925);
    outputs(1370) <= (layer0_outputs(422)) or (layer0_outputs(4477));
    outputs(1371) <= layer0_outputs(2516);
    outputs(1372) <= (layer0_outputs(3724)) and not (layer0_outputs(5015));
    outputs(1373) <= not((layer0_outputs(259)) or (layer0_outputs(4277)));
    outputs(1374) <= not(layer0_outputs(4117)) or (layer0_outputs(2196));
    outputs(1375) <= layer0_outputs(1955);
    outputs(1376) <= not((layer0_outputs(836)) and (layer0_outputs(718)));
    outputs(1377) <= not(layer0_outputs(2205));
    outputs(1378) <= (layer0_outputs(740)) and not (layer0_outputs(2771));
    outputs(1379) <= (layer0_outputs(690)) and (layer0_outputs(4770));
    outputs(1380) <= (layer0_outputs(1618)) or (layer0_outputs(3122));
    outputs(1381) <= (layer0_outputs(4468)) or (layer0_outputs(4321));
    outputs(1382) <= not(layer0_outputs(2985));
    outputs(1383) <= not((layer0_outputs(3162)) and (layer0_outputs(4796)));
    outputs(1384) <= not((layer0_outputs(2482)) or (layer0_outputs(527)));
    outputs(1385) <= layer0_outputs(4862);
    outputs(1386) <= (layer0_outputs(2810)) and (layer0_outputs(4964));
    outputs(1387) <= not((layer0_outputs(603)) and (layer0_outputs(910)));
    outputs(1388) <= layer0_outputs(250);
    outputs(1389) <= not(layer0_outputs(680));
    outputs(1390) <= layer0_outputs(882);
    outputs(1391) <= not((layer0_outputs(2378)) or (layer0_outputs(4337)));
    outputs(1392) <= not(layer0_outputs(1152));
    outputs(1393) <= layer0_outputs(3558);
    outputs(1394) <= (layer0_outputs(2708)) and not (layer0_outputs(2120));
    outputs(1395) <= layer0_outputs(3303);
    outputs(1396) <= not(layer0_outputs(2515)) or (layer0_outputs(2377));
    outputs(1397) <= (layer0_outputs(1886)) or (layer0_outputs(468));
    outputs(1398) <= not((layer0_outputs(4157)) xor (layer0_outputs(1643)));
    outputs(1399) <= not((layer0_outputs(1151)) xor (layer0_outputs(2978)));
    outputs(1400) <= not(layer0_outputs(490));
    outputs(1401) <= not(layer0_outputs(3061));
    outputs(1402) <= (layer0_outputs(1297)) and not (layer0_outputs(900));
    outputs(1403) <= (layer0_outputs(3847)) and not (layer0_outputs(735));
    outputs(1404) <= (layer0_outputs(1680)) and not (layer0_outputs(3487));
    outputs(1405) <= not((layer0_outputs(3275)) or (layer0_outputs(3077)));
    outputs(1406) <= not((layer0_outputs(4430)) xor (layer0_outputs(4900)));
    outputs(1407) <= (layer0_outputs(4558)) and (layer0_outputs(2383));
    outputs(1408) <= layer0_outputs(3346);
    outputs(1409) <= not(layer0_outputs(4582));
    outputs(1410) <= not((layer0_outputs(4703)) or (layer0_outputs(1469)));
    outputs(1411) <= not((layer0_outputs(3965)) and (layer0_outputs(481)));
    outputs(1412) <= not((layer0_outputs(2714)) xor (layer0_outputs(298)));
    outputs(1413) <= not(layer0_outputs(1858)) or (layer0_outputs(1652));
    outputs(1414) <= not(layer0_outputs(4931)) or (layer0_outputs(754));
    outputs(1415) <= not(layer0_outputs(4136));
    outputs(1416) <= not((layer0_outputs(1710)) and (layer0_outputs(3278)));
    outputs(1417) <= (layer0_outputs(1510)) or (layer0_outputs(1646));
    outputs(1418) <= not(layer0_outputs(4180));
    outputs(1419) <= not((layer0_outputs(454)) and (layer0_outputs(436)));
    outputs(1420) <= (layer0_outputs(2088)) and not (layer0_outputs(4226));
    outputs(1421) <= not((layer0_outputs(74)) xor (layer0_outputs(4238)));
    outputs(1422) <= layer0_outputs(3481);
    outputs(1423) <= layer0_outputs(4285);
    outputs(1424) <= (layer0_outputs(4212)) and (layer0_outputs(3220));
    outputs(1425) <= not(layer0_outputs(1765));
    outputs(1426) <= layer0_outputs(1732);
    outputs(1427) <= (layer0_outputs(2088)) and not (layer0_outputs(2093));
    outputs(1428) <= not((layer0_outputs(3657)) and (layer0_outputs(782)));
    outputs(1429) <= (layer0_outputs(320)) and not (layer0_outputs(5098));
    outputs(1430) <= not(layer0_outputs(4424)) or (layer0_outputs(2680));
    outputs(1431) <= not(layer0_outputs(4393));
    outputs(1432) <= not(layer0_outputs(788));
    outputs(1433) <= not(layer0_outputs(2178));
    outputs(1434) <= not((layer0_outputs(4403)) and (layer0_outputs(3062)));
    outputs(1435) <= (layer0_outputs(5032)) xor (layer0_outputs(3375));
    outputs(1436) <= not(layer0_outputs(2182));
    outputs(1437) <= not(layer0_outputs(1962));
    outputs(1438) <= layer0_outputs(1007);
    outputs(1439) <= not(layer0_outputs(3606));
    outputs(1440) <= not(layer0_outputs(3956));
    outputs(1441) <= not(layer0_outputs(1136));
    outputs(1442) <= (layer0_outputs(4593)) and not (layer0_outputs(713));
    outputs(1443) <= layer0_outputs(3896);
    outputs(1444) <= not(layer0_outputs(2621));
    outputs(1445) <= not(layer0_outputs(2537)) or (layer0_outputs(3853));
    outputs(1446) <= not(layer0_outputs(2800));
    outputs(1447) <= not(layer0_outputs(3661));
    outputs(1448) <= not((layer0_outputs(4069)) and (layer0_outputs(1708)));
    outputs(1449) <= not(layer0_outputs(1133));
    outputs(1450) <= not(layer0_outputs(39)) or (layer0_outputs(3330));
    outputs(1451) <= not((layer0_outputs(859)) xor (layer0_outputs(1655)));
    outputs(1452) <= layer0_outputs(673);
    outputs(1453) <= not(layer0_outputs(3779)) or (layer0_outputs(2646));
    outputs(1454) <= not(layer0_outputs(2871)) or (layer0_outputs(3460));
    outputs(1455) <= (layer0_outputs(5062)) and (layer0_outputs(1985));
    outputs(1456) <= not(layer0_outputs(4867));
    outputs(1457) <= layer0_outputs(1896);
    outputs(1458) <= not(layer0_outputs(1131)) or (layer0_outputs(2552));
    outputs(1459) <= layer0_outputs(1327);
    outputs(1460) <= not(layer0_outputs(3142));
    outputs(1461) <= layer0_outputs(3161);
    outputs(1462) <= not(layer0_outputs(1821));
    outputs(1463) <= not((layer0_outputs(2596)) and (layer0_outputs(1201)));
    outputs(1464) <= not(layer0_outputs(4331)) or (layer0_outputs(1999));
    outputs(1465) <= not(layer0_outputs(3280));
    outputs(1466) <= not(layer0_outputs(2654));
    outputs(1467) <= not(layer0_outputs(2362));
    outputs(1468) <= not((layer0_outputs(4282)) xor (layer0_outputs(1311)));
    outputs(1469) <= not(layer0_outputs(4935));
    outputs(1470) <= not(layer0_outputs(1848));
    outputs(1471) <= (layer0_outputs(2939)) xor (layer0_outputs(2330));
    outputs(1472) <= layer0_outputs(387);
    outputs(1473) <= not(layer0_outputs(4118));
    outputs(1474) <= not(layer0_outputs(4493)) or (layer0_outputs(447));
    outputs(1475) <= layer0_outputs(3303);
    outputs(1476) <= layer0_outputs(2941);
    outputs(1477) <= layer0_outputs(102);
    outputs(1478) <= not(layer0_outputs(3137));
    outputs(1479) <= not(layer0_outputs(2194)) or (layer0_outputs(447));
    outputs(1480) <= not((layer0_outputs(489)) or (layer0_outputs(3883)));
    outputs(1481) <= (layer0_outputs(4850)) and not (layer0_outputs(3182));
    outputs(1482) <= not(layer0_outputs(4874));
    outputs(1483) <= layer0_outputs(4004);
    outputs(1484) <= not(layer0_outputs(4278));
    outputs(1485) <= not(layer0_outputs(1571)) or (layer0_outputs(1825));
    outputs(1486) <= not((layer0_outputs(4481)) and (layer0_outputs(4403)));
    outputs(1487) <= not((layer0_outputs(4344)) and (layer0_outputs(397)));
    outputs(1488) <= not((layer0_outputs(2859)) xor (layer0_outputs(2025)));
    outputs(1489) <= (layer0_outputs(1493)) xor (layer0_outputs(255));
    outputs(1490) <= (layer0_outputs(3788)) or (layer0_outputs(3336));
    outputs(1491) <= not(layer0_outputs(5048)) or (layer0_outputs(1679));
    outputs(1492) <= not(layer0_outputs(4190));
    outputs(1493) <= not(layer0_outputs(1253)) or (layer0_outputs(1717));
    outputs(1494) <= (layer0_outputs(496)) or (layer0_outputs(3042));
    outputs(1495) <= not(layer0_outputs(2743));
    outputs(1496) <= (layer0_outputs(2231)) and not (layer0_outputs(3311));
    outputs(1497) <= not(layer0_outputs(1193));
    outputs(1498) <= layer0_outputs(2301);
    outputs(1499) <= layer0_outputs(153);
    outputs(1500) <= (layer0_outputs(1532)) and not (layer0_outputs(4173));
    outputs(1501) <= (layer0_outputs(2733)) and (layer0_outputs(2426));
    outputs(1502) <= not(layer0_outputs(2645)) or (layer0_outputs(4004));
    outputs(1503) <= not(layer0_outputs(4891));
    outputs(1504) <= not((layer0_outputs(4709)) xor (layer0_outputs(3848)));
    outputs(1505) <= (layer0_outputs(66)) and not (layer0_outputs(4796));
    outputs(1506) <= (layer0_outputs(3599)) or (layer0_outputs(4429));
    outputs(1507) <= layer0_outputs(3739);
    outputs(1508) <= (layer0_outputs(1395)) or (layer0_outputs(3769));
    outputs(1509) <= not(layer0_outputs(3129));
    outputs(1510) <= layer0_outputs(3449);
    outputs(1511) <= not(layer0_outputs(595));
    outputs(1512) <= layer0_outputs(1555);
    outputs(1513) <= (layer0_outputs(488)) and not (layer0_outputs(1145));
    outputs(1514) <= '1';
    outputs(1515) <= layer0_outputs(2353);
    outputs(1516) <= (layer0_outputs(804)) and (layer0_outputs(5066));
    outputs(1517) <= not(layer0_outputs(758));
    outputs(1518) <= layer0_outputs(4432);
    outputs(1519) <= not(layer0_outputs(4828));
    outputs(1520) <= (layer0_outputs(1689)) and not (layer0_outputs(3843));
    outputs(1521) <= not(layer0_outputs(1038)) or (layer0_outputs(4165));
    outputs(1522) <= layer0_outputs(4296);
    outputs(1523) <= layer0_outputs(674);
    outputs(1524) <= (layer0_outputs(4343)) or (layer0_outputs(5063));
    outputs(1525) <= not((layer0_outputs(1594)) and (layer0_outputs(2607)));
    outputs(1526) <= not(layer0_outputs(3345)) or (layer0_outputs(1155));
    outputs(1527) <= layer0_outputs(4126);
    outputs(1528) <= not(layer0_outputs(4241)) or (layer0_outputs(2229));
    outputs(1529) <= not(layer0_outputs(945)) or (layer0_outputs(3363));
    outputs(1530) <= layer0_outputs(1797);
    outputs(1531) <= (layer0_outputs(4711)) and not (layer0_outputs(3859));
    outputs(1532) <= not(layer0_outputs(264));
    outputs(1533) <= not(layer0_outputs(797));
    outputs(1534) <= not((layer0_outputs(4655)) and (layer0_outputs(2139)));
    outputs(1535) <= not(layer0_outputs(4907)) or (layer0_outputs(2920));
    outputs(1536) <= not(layer0_outputs(2274)) or (layer0_outputs(1195));
    outputs(1537) <= layer0_outputs(124);
    outputs(1538) <= not((layer0_outputs(2934)) or (layer0_outputs(3349)));
    outputs(1539) <= layer0_outputs(3352);
    outputs(1540) <= layer0_outputs(2465);
    outputs(1541) <= not((layer0_outputs(3418)) or (layer0_outputs(3797)));
    outputs(1542) <= layer0_outputs(4475);
    outputs(1543) <= (layer0_outputs(4284)) and not (layer0_outputs(130));
    outputs(1544) <= not(layer0_outputs(1126));
    outputs(1545) <= (layer0_outputs(1292)) and not (layer0_outputs(3221));
    outputs(1546) <= (layer0_outputs(4330)) and not (layer0_outputs(3099));
    outputs(1547) <= (layer0_outputs(4332)) and not (layer0_outputs(3816));
    outputs(1548) <= layer0_outputs(3562);
    outputs(1549) <= not(layer0_outputs(3628));
    outputs(1550) <= (layer0_outputs(315)) and not (layer0_outputs(3120));
    outputs(1551) <= not(layer0_outputs(4592));
    outputs(1552) <= layer0_outputs(2681);
    outputs(1553) <= (layer0_outputs(2892)) and not (layer0_outputs(1974));
    outputs(1554) <= (layer0_outputs(2004)) and (layer0_outputs(4464));
    outputs(1555) <= layer0_outputs(1760);
    outputs(1556) <= (layer0_outputs(5039)) and not (layer0_outputs(4080));
    outputs(1557) <= (layer0_outputs(1410)) and not (layer0_outputs(4362));
    outputs(1558) <= not((layer0_outputs(2780)) xor (layer0_outputs(3768)));
    outputs(1559) <= not(layer0_outputs(2831)) or (layer0_outputs(2038));
    outputs(1560) <= layer0_outputs(643);
    outputs(1561) <= layer0_outputs(4764);
    outputs(1562) <= layer0_outputs(3323);
    outputs(1563) <= (layer0_outputs(4374)) and not (layer0_outputs(2288));
    outputs(1564) <= not(layer0_outputs(2331));
    outputs(1565) <= not((layer0_outputs(944)) or (layer0_outputs(1880)));
    outputs(1566) <= not((layer0_outputs(4659)) xor (layer0_outputs(789)));
    outputs(1567) <= (layer0_outputs(745)) and not (layer0_outputs(4753));
    outputs(1568) <= layer0_outputs(2943);
    outputs(1569) <= (layer0_outputs(2022)) and not (layer0_outputs(1009));
    outputs(1570) <= (layer0_outputs(4167)) and (layer0_outputs(1179));
    outputs(1571) <= (layer0_outputs(2494)) or (layer0_outputs(3385));
    outputs(1572) <= layer0_outputs(830);
    outputs(1573) <= not((layer0_outputs(545)) or (layer0_outputs(3584)));
    outputs(1574) <= layer0_outputs(4077);
    outputs(1575) <= (layer0_outputs(1921)) and not (layer0_outputs(855));
    outputs(1576) <= not(layer0_outputs(4093));
    outputs(1577) <= not(layer0_outputs(266));
    outputs(1578) <= not(layer0_outputs(2970));
    outputs(1579) <= (layer0_outputs(1943)) and (layer0_outputs(2950));
    outputs(1580) <= (layer0_outputs(1929)) xor (layer0_outputs(2627));
    outputs(1581) <= not(layer0_outputs(2475));
    outputs(1582) <= not(layer0_outputs(3246)) or (layer0_outputs(981));
    outputs(1583) <= layer0_outputs(1224);
    outputs(1584) <= (layer0_outputs(4089)) and not (layer0_outputs(4147));
    outputs(1585) <= not(layer0_outputs(4037));
    outputs(1586) <= not(layer0_outputs(2862));
    outputs(1587) <= not(layer0_outputs(4822)) or (layer0_outputs(4706));
    outputs(1588) <= layer0_outputs(4683);
    outputs(1589) <= not((layer0_outputs(4152)) or (layer0_outputs(387)));
    outputs(1590) <= not((layer0_outputs(409)) and (layer0_outputs(3688)));
    outputs(1591) <= layer0_outputs(3613);
    outputs(1592) <= not(layer0_outputs(2768));
    outputs(1593) <= (layer0_outputs(4417)) and not (layer0_outputs(1265));
    outputs(1594) <= layer0_outputs(1291);
    outputs(1595) <= layer0_outputs(259);
    outputs(1596) <= (layer0_outputs(269)) and not (layer0_outputs(2873));
    outputs(1597) <= (layer0_outputs(880)) or (layer0_outputs(2663));
    outputs(1598) <= layer0_outputs(3145);
    outputs(1599) <= (layer0_outputs(3357)) or (layer0_outputs(347));
    outputs(1600) <= layer0_outputs(1902);
    outputs(1601) <= layer0_outputs(3615);
    outputs(1602) <= layer0_outputs(4582);
    outputs(1603) <= not((layer0_outputs(3967)) or (layer0_outputs(1676)));
    outputs(1604) <= not(layer0_outputs(4266));
    outputs(1605) <= layer0_outputs(1295);
    outputs(1606) <= layer0_outputs(721);
    outputs(1607) <= not(layer0_outputs(1058));
    outputs(1608) <= (layer0_outputs(3092)) and not (layer0_outputs(4449));
    outputs(1609) <= not((layer0_outputs(3954)) xor (layer0_outputs(3858)));
    outputs(1610) <= layer0_outputs(3571);
    outputs(1611) <= not(layer0_outputs(4751));
    outputs(1612) <= not(layer0_outputs(278));
    outputs(1613) <= (layer0_outputs(382)) and not (layer0_outputs(4342));
    outputs(1614) <= (layer0_outputs(714)) xor (layer0_outputs(3369));
    outputs(1615) <= (layer0_outputs(3195)) and not (layer0_outputs(814));
    outputs(1616) <= (layer0_outputs(95)) and not (layer0_outputs(1146));
    outputs(1617) <= (layer0_outputs(4738)) or (layer0_outputs(2841));
    outputs(1618) <= (layer0_outputs(2910)) and not (layer0_outputs(3656));
    outputs(1619) <= layer0_outputs(2356);
    outputs(1620) <= (layer0_outputs(3469)) and (layer0_outputs(566));
    outputs(1621) <= not(layer0_outputs(4384)) or (layer0_outputs(1434));
    outputs(1622) <= layer0_outputs(3888);
    outputs(1623) <= layer0_outputs(594);
    outputs(1624) <= not(layer0_outputs(1687));
    outputs(1625) <= layer0_outputs(2200);
    outputs(1626) <= not((layer0_outputs(4902)) or (layer0_outputs(3711)));
    outputs(1627) <= not(layer0_outputs(104));
    outputs(1628) <= not(layer0_outputs(2678));
    outputs(1629) <= layer0_outputs(2440);
    outputs(1630) <= (layer0_outputs(4516)) and not (layer0_outputs(3227));
    outputs(1631) <= (layer0_outputs(3877)) and not (layer0_outputs(4269));
    outputs(1632) <= layer0_outputs(1110);
    outputs(1633) <= (layer0_outputs(598)) and not (layer0_outputs(3274));
    outputs(1634) <= not(layer0_outputs(4534)) or (layer0_outputs(2581));
    outputs(1635) <= (layer0_outputs(86)) or (layer0_outputs(3248));
    outputs(1636) <= layer0_outputs(1037);
    outputs(1637) <= (layer0_outputs(2415)) and (layer0_outputs(1452));
    outputs(1638) <= not((layer0_outputs(1249)) xor (layer0_outputs(3235)));
    outputs(1639) <= (layer0_outputs(1335)) xor (layer0_outputs(403));
    outputs(1640) <= layer0_outputs(681);
    outputs(1641) <= not(layer0_outputs(4486)) or (layer0_outputs(97));
    outputs(1642) <= layer0_outputs(1937);
    outputs(1643) <= not(layer0_outputs(1657));
    outputs(1644) <= not(layer0_outputs(3705));
    outputs(1645) <= (layer0_outputs(4456)) and not (layer0_outputs(593));
    outputs(1646) <= (layer0_outputs(4016)) and not (layer0_outputs(3997));
    outputs(1647) <= (layer0_outputs(4084)) xor (layer0_outputs(2692));
    outputs(1648) <= layer0_outputs(4430);
    outputs(1649) <= (layer0_outputs(4097)) and (layer0_outputs(3738));
    outputs(1650) <= (layer0_outputs(2254)) or (layer0_outputs(2761));
    outputs(1651) <= not(layer0_outputs(4263)) or (layer0_outputs(2429));
    outputs(1652) <= not(layer0_outputs(4752));
    outputs(1653) <= layer0_outputs(2127);
    outputs(1654) <= not((layer0_outputs(3025)) xor (layer0_outputs(3153)));
    outputs(1655) <= (layer0_outputs(3748)) and not (layer0_outputs(1647));
    outputs(1656) <= (layer0_outputs(4407)) and not (layer0_outputs(3314));
    outputs(1657) <= (layer0_outputs(969)) and not (layer0_outputs(3530));
    outputs(1658) <= not((layer0_outputs(4399)) xor (layer0_outputs(76)));
    outputs(1659) <= not((layer0_outputs(4231)) or (layer0_outputs(4616)));
    outputs(1660) <= not(layer0_outputs(2688));
    outputs(1661) <= (layer0_outputs(4599)) and not (layer0_outputs(4546));
    outputs(1662) <= not(layer0_outputs(704)) or (layer0_outputs(1378));
    outputs(1663) <= not(layer0_outputs(4307)) or (layer0_outputs(798));
    outputs(1664) <= not((layer0_outputs(1951)) or (layer0_outputs(350)));
    outputs(1665) <= not(layer0_outputs(309));
    outputs(1666) <= layer0_outputs(4929);
    outputs(1667) <= (layer0_outputs(3072)) and not (layer0_outputs(4350));
    outputs(1668) <= (layer0_outputs(3812)) and not (layer0_outputs(4188));
    outputs(1669) <= (layer0_outputs(1384)) and not (layer0_outputs(1357));
    outputs(1670) <= not((layer0_outputs(2412)) xor (layer0_outputs(1278)));
    outputs(1671) <= (layer0_outputs(4870)) and (layer0_outputs(105));
    outputs(1672) <= not((layer0_outputs(3938)) or (layer0_outputs(2224)));
    outputs(1673) <= layer0_outputs(336);
    outputs(1674) <= layer0_outputs(3770);
    outputs(1675) <= not(layer0_outputs(2259));
    outputs(1676) <= (layer0_outputs(2303)) and not (layer0_outputs(2375));
    outputs(1677) <= not(layer0_outputs(3663));
    outputs(1678) <= not(layer0_outputs(3263));
    outputs(1679) <= not(layer0_outputs(2153));
    outputs(1680) <= (layer0_outputs(4591)) and not (layer0_outputs(3199));
    outputs(1681) <= not(layer0_outputs(875));
    outputs(1682) <= not(layer0_outputs(1633)) or (layer0_outputs(4098));
    outputs(1683) <= not(layer0_outputs(3746));
    outputs(1684) <= not(layer0_outputs(2706));
    outputs(1685) <= not((layer0_outputs(1853)) or (layer0_outputs(1565)));
    outputs(1686) <= not((layer0_outputs(2383)) xor (layer0_outputs(3910)));
    outputs(1687) <= layer0_outputs(4475);
    outputs(1688) <= layer0_outputs(1213);
    outputs(1689) <= not((layer0_outputs(4843)) or (layer0_outputs(1724)));
    outputs(1690) <= not(layer0_outputs(2493));
    outputs(1691) <= not(layer0_outputs(1442)) or (layer0_outputs(1761));
    outputs(1692) <= (layer0_outputs(3844)) xor (layer0_outputs(1909));
    outputs(1693) <= (layer0_outputs(411)) and (layer0_outputs(337));
    outputs(1694) <= (layer0_outputs(1601)) and (layer0_outputs(316));
    outputs(1695) <= layer0_outputs(3506);
    outputs(1696) <= layer0_outputs(3516);
    outputs(1697) <= not(layer0_outputs(2792));
    outputs(1698) <= not(layer0_outputs(4719));
    outputs(1699) <= layer0_outputs(955);
    outputs(1700) <= (layer0_outputs(4868)) xor (layer0_outputs(4295));
    outputs(1701) <= not(layer0_outputs(1911));
    outputs(1702) <= not((layer0_outputs(2762)) or (layer0_outputs(157)));
    outputs(1703) <= layer0_outputs(3427);
    outputs(1704) <= layer0_outputs(248);
    outputs(1705) <= (layer0_outputs(4135)) or (layer0_outputs(3036));
    outputs(1706) <= (layer0_outputs(686)) and (layer0_outputs(1319));
    outputs(1707) <= layer0_outputs(2322);
    outputs(1708) <= (layer0_outputs(539)) and not (layer0_outputs(4836));
    outputs(1709) <= layer0_outputs(3208);
    outputs(1710) <= not((layer0_outputs(1162)) xor (layer0_outputs(991)));
    outputs(1711) <= not(layer0_outputs(2572));
    outputs(1712) <= (layer0_outputs(40)) and not (layer0_outputs(2071));
    outputs(1713) <= layer0_outputs(3456);
    outputs(1714) <= not(layer0_outputs(767));
    outputs(1715) <= (layer0_outputs(3587)) and not (layer0_outputs(4445));
    outputs(1716) <= not(layer0_outputs(2685));
    outputs(1717) <= not((layer0_outputs(2061)) and (layer0_outputs(4360)));
    outputs(1718) <= not((layer0_outputs(1198)) or (layer0_outputs(2053)));
    outputs(1719) <= (layer0_outputs(1502)) and not (layer0_outputs(4874));
    outputs(1720) <= layer0_outputs(4369);
    outputs(1721) <= (layer0_outputs(3457)) and not (layer0_outputs(1972));
    outputs(1722) <= (layer0_outputs(1296)) and (layer0_outputs(1783));
    outputs(1723) <= not(layer0_outputs(951)) or (layer0_outputs(3341));
    outputs(1724) <= layer0_outputs(4085);
    outputs(1725) <= layer0_outputs(2705);
    outputs(1726) <= not((layer0_outputs(608)) or (layer0_outputs(4256)));
    outputs(1727) <= (layer0_outputs(3803)) and not (layer0_outputs(2686));
    outputs(1728) <= not(layer0_outputs(77)) or (layer0_outputs(887));
    outputs(1729) <= not(layer0_outputs(4433));
    outputs(1730) <= not(layer0_outputs(1445)) or (layer0_outputs(973));
    outputs(1731) <= not((layer0_outputs(4761)) xor (layer0_outputs(2315)));
    outputs(1732) <= (layer0_outputs(1995)) and not (layer0_outputs(57));
    outputs(1733) <= layer0_outputs(2534);
    outputs(1734) <= (layer0_outputs(1673)) and (layer0_outputs(2577));
    outputs(1735) <= not((layer0_outputs(1524)) and (layer0_outputs(354)));
    outputs(1736) <= (layer0_outputs(2156)) or (layer0_outputs(2175));
    outputs(1737) <= not(layer0_outputs(4668)) or (layer0_outputs(147));
    outputs(1738) <= not((layer0_outputs(4313)) or (layer0_outputs(4941)));
    outputs(1739) <= not(layer0_outputs(3767)) or (layer0_outputs(1881));
    outputs(1740) <= (layer0_outputs(2989)) and not (layer0_outputs(2366));
    outputs(1741) <= not(layer0_outputs(4795));
    outputs(1742) <= (layer0_outputs(1015)) and (layer0_outputs(2897));
    outputs(1743) <= (layer0_outputs(403)) xor (layer0_outputs(3935));
    outputs(1744) <= layer0_outputs(4778);
    outputs(1745) <= not((layer0_outputs(2881)) or (layer0_outputs(1856)));
    outputs(1746) <= (layer0_outputs(4572)) and not (layer0_outputs(4926));
    outputs(1747) <= not(layer0_outputs(4614));
    outputs(1748) <= not(layer0_outputs(2926));
    outputs(1749) <= not(layer0_outputs(599));
    outputs(1750) <= not(layer0_outputs(2427));
    outputs(1751) <= (layer0_outputs(2673)) or (layer0_outputs(2867));
    outputs(1752) <= not((layer0_outputs(2543)) or (layer0_outputs(5010)));
    outputs(1753) <= layer0_outputs(4416);
    outputs(1754) <= layer0_outputs(1518);
    outputs(1755) <= layer0_outputs(2562);
    outputs(1756) <= (layer0_outputs(472)) xor (layer0_outputs(4388));
    outputs(1757) <= not(layer0_outputs(73));
    outputs(1758) <= (layer0_outputs(1942)) and not (layer0_outputs(3503));
    outputs(1759) <= not(layer0_outputs(3107));
    outputs(1760) <= (layer0_outputs(1368)) and (layer0_outputs(3953));
    outputs(1761) <= not(layer0_outputs(4422));
    outputs(1762) <= not(layer0_outputs(359));
    outputs(1763) <= not((layer0_outputs(3526)) or (layer0_outputs(3604)));
    outputs(1764) <= (layer0_outputs(3218)) xor (layer0_outputs(1254));
    outputs(1765) <= layer0_outputs(2584);
    outputs(1766) <= (layer0_outputs(2154)) xor (layer0_outputs(4694));
    outputs(1767) <= (layer0_outputs(2008)) and not (layer0_outputs(4942));
    outputs(1768) <= not(layer0_outputs(4113));
    outputs(1769) <= (layer0_outputs(2636)) and not (layer0_outputs(3373));
    outputs(1770) <= not(layer0_outputs(1578)) or (layer0_outputs(3802));
    outputs(1771) <= not(layer0_outputs(4813));
    outputs(1772) <= not(layer0_outputs(3600));
    outputs(1773) <= (layer0_outputs(3259)) and not (layer0_outputs(2253));
    outputs(1774) <= (layer0_outputs(843)) and not (layer0_outputs(4394));
    outputs(1775) <= (layer0_outputs(1053)) and not (layer0_outputs(256));
    outputs(1776) <= not(layer0_outputs(2197));
    outputs(1777) <= not(layer0_outputs(4887));
    outputs(1778) <= (layer0_outputs(3192)) or (layer0_outputs(2894));
    outputs(1779) <= (layer0_outputs(2004)) and (layer0_outputs(66));
    outputs(1780) <= not((layer0_outputs(1711)) and (layer0_outputs(1520)));
    outputs(1781) <= (layer0_outputs(2340)) and (layer0_outputs(865));
    outputs(1782) <= not((layer0_outputs(5045)) xor (layer0_outputs(5102)));
    outputs(1783) <= (layer0_outputs(4516)) and (layer0_outputs(3092));
    outputs(1784) <= not(layer0_outputs(4333));
    outputs(1785) <= (layer0_outputs(3996)) and not (layer0_outputs(2034));
    outputs(1786) <= layer0_outputs(249);
    outputs(1787) <= (layer0_outputs(2466)) and (layer0_outputs(4100));
    outputs(1788) <= (layer0_outputs(1252)) and not (layer0_outputs(42));
    outputs(1789) <= (layer0_outputs(2499)) and not (layer0_outputs(2997));
    outputs(1790) <= not((layer0_outputs(378)) or (layer0_outputs(378)));
    outputs(1791) <= (layer0_outputs(1899)) and (layer0_outputs(4637));
    outputs(1792) <= not(layer0_outputs(1129));
    outputs(1793) <= (layer0_outputs(4410)) and (layer0_outputs(2568));
    outputs(1794) <= not((layer0_outputs(2773)) or (layer0_outputs(3737)));
    outputs(1795) <= layer0_outputs(4089);
    outputs(1796) <= not((layer0_outputs(808)) xor (layer0_outputs(461)));
    outputs(1797) <= (layer0_outputs(1160)) or (layer0_outputs(3543));
    outputs(1798) <= (layer0_outputs(1850)) and not (layer0_outputs(4056));
    outputs(1799) <= not((layer0_outputs(4058)) xor (layer0_outputs(762)));
    outputs(1800) <= (layer0_outputs(4794)) and not (layer0_outputs(1116));
    outputs(1801) <= not((layer0_outputs(972)) or (layer0_outputs(2363)));
    outputs(1802) <= not((layer0_outputs(227)) and (layer0_outputs(1431)));
    outputs(1803) <= (layer0_outputs(3328)) or (layer0_outputs(2410));
    outputs(1804) <= (layer0_outputs(2512)) and not (layer0_outputs(1882));
    outputs(1805) <= (layer0_outputs(50)) and (layer0_outputs(2338));
    outputs(1806) <= not(layer0_outputs(1557));
    outputs(1807) <= not(layer0_outputs(765)) or (layer0_outputs(1999));
    outputs(1808) <= (layer0_outputs(4721)) and not (layer0_outputs(162));
    outputs(1809) <= (layer0_outputs(2351)) and (layer0_outputs(462));
    outputs(1810) <= not(layer0_outputs(2670));
    outputs(1811) <= (layer0_outputs(2294)) and not (layer0_outputs(3959));
    outputs(1812) <= (layer0_outputs(1292)) and not (layer0_outputs(688));
    outputs(1813) <= layer0_outputs(4997);
    outputs(1814) <= (layer0_outputs(4129)) and not (layer0_outputs(3880));
    outputs(1815) <= (layer0_outputs(3424)) and (layer0_outputs(3944));
    outputs(1816) <= (layer0_outputs(83)) and not (layer0_outputs(4747));
    outputs(1817) <= not(layer0_outputs(1735));
    outputs(1818) <= layer0_outputs(1479);
    outputs(1819) <= not(layer0_outputs(1880));
    outputs(1820) <= not(layer0_outputs(4346));
    outputs(1821) <= layer0_outputs(3045);
    outputs(1822) <= not(layer0_outputs(538));
    outputs(1823) <= layer0_outputs(1306);
    outputs(1824) <= not(layer0_outputs(3140));
    outputs(1825) <= not((layer0_outputs(4219)) or (layer0_outputs(3028)));
    outputs(1826) <= not(layer0_outputs(1690));
    outputs(1827) <= (layer0_outputs(3376)) xor (layer0_outputs(756));
    outputs(1828) <= (layer0_outputs(481)) and not (layer0_outputs(349));
    outputs(1829) <= not(layer0_outputs(3379));
    outputs(1830) <= not(layer0_outputs(2501));
    outputs(1831) <= not(layer0_outputs(4690));
    outputs(1832) <= layer0_outputs(3052);
    outputs(1833) <= not((layer0_outputs(4858)) or (layer0_outputs(1641)));
    outputs(1834) <= layer0_outputs(4682);
    outputs(1835) <= not(layer0_outputs(1390));
    outputs(1836) <= not(layer0_outputs(1370));
    outputs(1837) <= layer0_outputs(2801);
    outputs(1838) <= (layer0_outputs(2016)) and not (layer0_outputs(1861));
    outputs(1839) <= (layer0_outputs(3544)) and (layer0_outputs(3067));
    outputs(1840) <= not(layer0_outputs(1885)) or (layer0_outputs(3403));
    outputs(1841) <= layer0_outputs(149);
    outputs(1842) <= not(layer0_outputs(3105)) or (layer0_outputs(2048));
    outputs(1843) <= not(layer0_outputs(1178));
    outputs(1844) <= not(layer0_outputs(349));
    outputs(1845) <= not(layer0_outputs(1082));
    outputs(1846) <= not((layer0_outputs(957)) and (layer0_outputs(3842)));
    outputs(1847) <= not(layer0_outputs(3773));
    outputs(1848) <= not(layer0_outputs(242));
    outputs(1849) <= not(layer0_outputs(4833));
    outputs(1850) <= layer0_outputs(2152);
    outputs(1851) <= not((layer0_outputs(4235)) xor (layer0_outputs(3113)));
    outputs(1852) <= (layer0_outputs(345)) and (layer0_outputs(4410));
    outputs(1853) <= not((layer0_outputs(3331)) and (layer0_outputs(4716)));
    outputs(1854) <= not((layer0_outputs(4499)) xor (layer0_outputs(350)));
    outputs(1855) <= layer0_outputs(3071);
    outputs(1856) <= not(layer0_outputs(1234)) or (layer0_outputs(263));
    outputs(1857) <= not((layer0_outputs(1804)) or (layer0_outputs(2111)));
    outputs(1858) <= layer0_outputs(4327);
    outputs(1859) <= (layer0_outputs(1722)) and (layer0_outputs(2066));
    outputs(1860) <= (layer0_outputs(3354)) and not (layer0_outputs(2267));
    outputs(1861) <= (layer0_outputs(4632)) or (layer0_outputs(1377));
    outputs(1862) <= not((layer0_outputs(356)) or (layer0_outputs(940)));
    outputs(1863) <= not(layer0_outputs(677));
    outputs(1864) <= not((layer0_outputs(2834)) and (layer0_outputs(3280)));
    outputs(1865) <= not((layer0_outputs(3765)) and (layer0_outputs(4035)));
    outputs(1866) <= (layer0_outputs(1204)) xor (layer0_outputs(3684));
    outputs(1867) <= not((layer0_outputs(2706)) or (layer0_outputs(4504)));
    outputs(1868) <= not(layer0_outputs(3347));
    outputs(1869) <= not(layer0_outputs(2062));
    outputs(1870) <= layer0_outputs(4358);
    outputs(1871) <= not(layer0_outputs(2921));
    outputs(1872) <= not(layer0_outputs(4595)) or (layer0_outputs(4019));
    outputs(1873) <= not(layer0_outputs(3550));
    outputs(1874) <= (layer0_outputs(3234)) and (layer0_outputs(1363));
    outputs(1875) <= layer0_outputs(3390);
    outputs(1876) <= (layer0_outputs(4815)) and (layer0_outputs(79));
    outputs(1877) <= (layer0_outputs(4645)) and not (layer0_outputs(920));
    outputs(1878) <= (layer0_outputs(1736)) and (layer0_outputs(2637));
    outputs(1879) <= (layer0_outputs(5047)) and (layer0_outputs(3129));
    outputs(1880) <= not(layer0_outputs(1953));
    outputs(1881) <= (layer0_outputs(156)) xor (layer0_outputs(4509));
    outputs(1882) <= (layer0_outputs(4377)) xor (layer0_outputs(4373));
    outputs(1883) <= layer0_outputs(2530);
    outputs(1884) <= layer0_outputs(4357);
    outputs(1885) <= layer0_outputs(988);
    outputs(1886) <= (layer0_outputs(2634)) or (layer0_outputs(28));
    outputs(1887) <= (layer0_outputs(1478)) xor (layer0_outputs(464));
    outputs(1888) <= (layer0_outputs(100)) and not (layer0_outputs(3522));
    outputs(1889) <= not(layer0_outputs(2044)) or (layer0_outputs(3431));
    outputs(1890) <= not((layer0_outputs(1435)) or (layer0_outputs(4453)));
    outputs(1891) <= not(layer0_outputs(1380));
    outputs(1892) <= layer0_outputs(231);
    outputs(1893) <= (layer0_outputs(2138)) xor (layer0_outputs(979));
    outputs(1894) <= layer0_outputs(553);
    outputs(1895) <= (layer0_outputs(3471)) and not (layer0_outputs(243));
    outputs(1896) <= layer0_outputs(1451);
    outputs(1897) <= not(layer0_outputs(4656));
    outputs(1898) <= not(layer0_outputs(4442));
    outputs(1899) <= layer0_outputs(4683);
    outputs(1900) <= (layer0_outputs(1969)) and not (layer0_outputs(979));
    outputs(1901) <= layer0_outputs(732);
    outputs(1902) <= not((layer0_outputs(3322)) and (layer0_outputs(2328)));
    outputs(1903) <= layer0_outputs(274);
    outputs(1904) <= (layer0_outputs(116)) and not (layer0_outputs(4866));
    outputs(1905) <= not(layer0_outputs(4480));
    outputs(1906) <= layer0_outputs(1591);
    outputs(1907) <= not(layer0_outputs(2493));
    outputs(1908) <= layer0_outputs(3747);
    outputs(1909) <= not((layer0_outputs(2601)) xor (layer0_outputs(4708)));
    outputs(1910) <= layer0_outputs(575);
    outputs(1911) <= (layer0_outputs(742)) and not (layer0_outputs(4729));
    outputs(1912) <= (layer0_outputs(1054)) and not (layer0_outputs(2803));
    outputs(1913) <= layer0_outputs(2527);
    outputs(1914) <= (layer0_outputs(2877)) and (layer0_outputs(2074));
    outputs(1915) <= (layer0_outputs(1833)) and not (layer0_outputs(3557));
    outputs(1916) <= (layer0_outputs(2068)) or (layer0_outputs(4126));
    outputs(1917) <= not((layer0_outputs(3686)) or (layer0_outputs(4992)));
    outputs(1918) <= layer0_outputs(4314);
    outputs(1919) <= (layer0_outputs(2832)) and not (layer0_outputs(4876));
    outputs(1920) <= (layer0_outputs(3699)) or (layer0_outputs(200));
    outputs(1921) <= not(layer0_outputs(2500)) or (layer0_outputs(3837));
    outputs(1922) <= (layer0_outputs(1029)) and not (layer0_outputs(2021));
    outputs(1923) <= not((layer0_outputs(4597)) or (layer0_outputs(4818)));
    outputs(1924) <= not(layer0_outputs(1586));
    outputs(1925) <= not(layer0_outputs(1884));
    outputs(1926) <= not(layer0_outputs(858));
    outputs(1927) <= (layer0_outputs(4426)) and not (layer0_outputs(2591));
    outputs(1928) <= not((layer0_outputs(456)) or (layer0_outputs(4941)));
    outputs(1929) <= not(layer0_outputs(4473)) or (layer0_outputs(5042));
    outputs(1930) <= layer0_outputs(3051);
    outputs(1931) <= (layer0_outputs(2316)) and not (layer0_outputs(2129));
    outputs(1932) <= (layer0_outputs(2927)) xor (layer0_outputs(1483));
    outputs(1933) <= not(layer0_outputs(3304)) or (layer0_outputs(1720));
    outputs(1934) <= layer0_outputs(2681);
    outputs(1935) <= not(layer0_outputs(2211));
    outputs(1936) <= not(layer0_outputs(4630));
    outputs(1937) <= not(layer0_outputs(2323));
    outputs(1938) <= (layer0_outputs(2639)) and not (layer0_outputs(2650));
    outputs(1939) <= (layer0_outputs(4216)) and not (layer0_outputs(4147));
    outputs(1940) <= layer0_outputs(2295);
    outputs(1941) <= layer0_outputs(5058);
    outputs(1942) <= not(layer0_outputs(3480)) or (layer0_outputs(185));
    outputs(1943) <= layer0_outputs(2611);
    outputs(1944) <= not(layer0_outputs(1281));
    outputs(1945) <= (layer0_outputs(2470)) and not (layer0_outputs(2928));
    outputs(1946) <= not(layer0_outputs(3017)) or (layer0_outputs(4265));
    outputs(1947) <= (layer0_outputs(5069)) and (layer0_outputs(3589));
    outputs(1948) <= not(layer0_outputs(529));
    outputs(1949) <= (layer0_outputs(20)) or (layer0_outputs(884));
    outputs(1950) <= layer0_outputs(2195);
    outputs(1951) <= not(layer0_outputs(2492));
    outputs(1952) <= not(layer0_outputs(3015));
    outputs(1953) <= (layer0_outputs(210)) and (layer0_outputs(1959));
    outputs(1954) <= (layer0_outputs(94)) and (layer0_outputs(4862));
    outputs(1955) <= layer0_outputs(4434);
    outputs(1956) <= layer0_outputs(1504);
    outputs(1957) <= (layer0_outputs(4671)) xor (layer0_outputs(4040));
    outputs(1958) <= layer0_outputs(4773);
    outputs(1959) <= layer0_outputs(1867);
    outputs(1960) <= layer0_outputs(2058);
    outputs(1961) <= layer0_outputs(2230);
    outputs(1962) <= not((layer0_outputs(1124)) or (layer0_outputs(4115)));
    outputs(1963) <= (layer0_outputs(1215)) and not (layer0_outputs(2437));
    outputs(1964) <= (layer0_outputs(1212)) xor (layer0_outputs(2317));
    outputs(1965) <= not(layer0_outputs(4979));
    outputs(1966) <= not(layer0_outputs(2167)) or (layer0_outputs(4220));
    outputs(1967) <= (layer0_outputs(103)) and not (layer0_outputs(1022));
    outputs(1968) <= not((layer0_outputs(3660)) xor (layer0_outputs(932)));
    outputs(1969) <= (layer0_outputs(4275)) and not (layer0_outputs(5037));
    outputs(1970) <= (layer0_outputs(3205)) and not (layer0_outputs(2343));
    outputs(1971) <= (layer0_outputs(1491)) and not (layer0_outputs(359));
    outputs(1972) <= (layer0_outputs(3282)) and not (layer0_outputs(498));
    outputs(1973) <= (layer0_outputs(822)) and not (layer0_outputs(5116));
    outputs(1974) <= (layer0_outputs(838)) and not (layer0_outputs(399));
    outputs(1975) <= not(layer0_outputs(4967)) or (layer0_outputs(1665));
    outputs(1976) <= not(layer0_outputs(1241)) or (layer0_outputs(5118));
    outputs(1977) <= not((layer0_outputs(2454)) xor (layer0_outputs(1572)));
    outputs(1978) <= (layer0_outputs(1041)) and not (layer0_outputs(107));
    outputs(1979) <= not((layer0_outputs(4808)) xor (layer0_outputs(1621)));
    outputs(1980) <= not(layer0_outputs(1967));
    outputs(1981) <= (layer0_outputs(2098)) and not (layer0_outputs(1622));
    outputs(1982) <= layer0_outputs(4791);
    outputs(1983) <= not((layer0_outputs(1026)) or (layer0_outputs(4046)));
    outputs(1984) <= not((layer0_outputs(2235)) or (layer0_outputs(2814)));
    outputs(1985) <= (layer0_outputs(638)) or (layer0_outputs(1632));
    outputs(1986) <= not((layer0_outputs(5071)) xor (layer0_outputs(3575)));
    outputs(1987) <= not(layer0_outputs(2357)) or (layer0_outputs(4750));
    outputs(1988) <= layer0_outputs(1457);
    outputs(1989) <= (layer0_outputs(41)) and not (layer0_outputs(1046));
    outputs(1990) <= (layer0_outputs(1740)) and not (layer0_outputs(4044));
    outputs(1991) <= (layer0_outputs(1991)) and (layer0_outputs(135));
    outputs(1992) <= (layer0_outputs(4397)) or (layer0_outputs(2904));
    outputs(1993) <= (layer0_outputs(629)) and not (layer0_outputs(4845));
    outputs(1994) <= not(layer0_outputs(3413));
    outputs(1995) <= not(layer0_outputs(1159));
    outputs(1996) <= not((layer0_outputs(1705)) or (layer0_outputs(5100)));
    outputs(1997) <= not(layer0_outputs(494));
    outputs(1998) <= (layer0_outputs(420)) and (layer0_outputs(2391));
    outputs(1999) <= (layer0_outputs(4068)) and (layer0_outputs(1742));
    outputs(2000) <= layer0_outputs(365);
    outputs(2001) <= (layer0_outputs(3801)) and not (layer0_outputs(5115));
    outputs(2002) <= not((layer0_outputs(3567)) or (layer0_outputs(1962)));
    outputs(2003) <= not((layer0_outputs(3887)) or (layer0_outputs(1512)));
    outputs(2004) <= not(layer0_outputs(117)) or (layer0_outputs(3155));
    outputs(2005) <= not(layer0_outputs(3411));
    outputs(2006) <= (layer0_outputs(1242)) xor (layer0_outputs(962));
    outputs(2007) <= not(layer0_outputs(1912));
    outputs(2008) <= (layer0_outputs(4060)) or (layer0_outputs(4466));
    outputs(2009) <= (layer0_outputs(2098)) and (layer0_outputs(722));
    outputs(2010) <= not(layer0_outputs(5082)) or (layer0_outputs(4361));
    outputs(2011) <= layer0_outputs(3877);
    outputs(2012) <= not((layer0_outputs(3848)) or (layer0_outputs(2947)));
    outputs(2013) <= layer0_outputs(4441);
    outputs(2014) <= (layer0_outputs(4232)) and not (layer0_outputs(4405));
    outputs(2015) <= not(layer0_outputs(1786));
    outputs(2016) <= (layer0_outputs(2527)) and (layer0_outputs(4470));
    outputs(2017) <= not((layer0_outputs(2282)) xor (layer0_outputs(2159)));
    outputs(2018) <= not(layer0_outputs(4199)) or (layer0_outputs(3980));
    outputs(2019) <= not(layer0_outputs(4362)) or (layer0_outputs(1495));
    outputs(2020) <= (layer0_outputs(3836)) and (layer0_outputs(4848));
    outputs(2021) <= (layer0_outputs(727)) and not (layer0_outputs(3097));
    outputs(2022) <= not(layer0_outputs(723));
    outputs(2023) <= (layer0_outputs(2252)) and not (layer0_outputs(3646));
    outputs(2024) <= not((layer0_outputs(2951)) and (layer0_outputs(1816)));
    outputs(2025) <= (layer0_outputs(550)) and not (layer0_outputs(4445));
    outputs(2026) <= not((layer0_outputs(2749)) xor (layer0_outputs(324)));
    outputs(2027) <= (layer0_outputs(1114)) and (layer0_outputs(5110));
    outputs(2028) <= (layer0_outputs(225)) and (layer0_outputs(1187));
    outputs(2029) <= layer0_outputs(4464);
    outputs(2030) <= layer0_outputs(28);
    outputs(2031) <= layer0_outputs(3519);
    outputs(2032) <= not(layer0_outputs(2916));
    outputs(2033) <= (layer0_outputs(299)) xor (layer0_outputs(509));
    outputs(2034) <= not(layer0_outputs(1101)) or (layer0_outputs(4666));
    outputs(2035) <= layer0_outputs(2536);
    outputs(2036) <= not(layer0_outputs(4916));
    outputs(2037) <= not(layer0_outputs(1390)) or (layer0_outputs(1732));
    outputs(2038) <= (layer0_outputs(3858)) or (layer0_outputs(2740));
    outputs(2039) <= layer0_outputs(834);
    outputs(2040) <= (layer0_outputs(1671)) and not (layer0_outputs(3723));
    outputs(2041) <= (layer0_outputs(476)) and not (layer0_outputs(658));
    outputs(2042) <= layer0_outputs(2710);
    outputs(2043) <= (layer0_outputs(148)) and not (layer0_outputs(285));
    outputs(2044) <= (layer0_outputs(3839)) and not (layer0_outputs(280));
    outputs(2045) <= layer0_outputs(988);
    outputs(2046) <= layer0_outputs(3998);
    outputs(2047) <= (layer0_outputs(4934)) and not (layer0_outputs(4609));
    outputs(2048) <= layer0_outputs(4894);
    outputs(2049) <= not((layer0_outputs(1531)) xor (layer0_outputs(1403)));
    outputs(2050) <= (layer0_outputs(2566)) and not (layer0_outputs(1805));
    outputs(2051) <= not(layer0_outputs(1760));
    outputs(2052) <= (layer0_outputs(3732)) and not (layer0_outputs(2699));
    outputs(2053) <= layer0_outputs(1569);
    outputs(2054) <= not(layer0_outputs(2353)) or (layer0_outputs(1448));
    outputs(2055) <= not(layer0_outputs(5069));
    outputs(2056) <= (layer0_outputs(4425)) and (layer0_outputs(626));
    outputs(2057) <= layer0_outputs(2616);
    outputs(2058) <= (layer0_outputs(3383)) and not (layer0_outputs(3813));
    outputs(2059) <= (layer0_outputs(920)) and not (layer0_outputs(4601));
    outputs(2060) <= (layer0_outputs(4844)) or (layer0_outputs(4958));
    outputs(2061) <= not(layer0_outputs(2030));
    outputs(2062) <= not(layer0_outputs(4567));
    outputs(2063) <= not(layer0_outputs(4138));
    outputs(2064) <= layer0_outputs(373);
    outputs(2065) <= not((layer0_outputs(149)) or (layer0_outputs(3482)));
    outputs(2066) <= not(layer0_outputs(4628));
    outputs(2067) <= not((layer0_outputs(2176)) xor (layer0_outputs(3690)));
    outputs(2068) <= layer0_outputs(3865);
    outputs(2069) <= layer0_outputs(1385);
    outputs(2070) <= (layer0_outputs(371)) xor (layer0_outputs(2619));
    outputs(2071) <= layer0_outputs(4247);
    outputs(2072) <= layer0_outputs(4818);
    outputs(2073) <= (layer0_outputs(1745)) or (layer0_outputs(2807));
    outputs(2074) <= (layer0_outputs(2396)) and (layer0_outputs(2875));
    outputs(2075) <= not(layer0_outputs(3270)) or (layer0_outputs(4684));
    outputs(2076) <= (layer0_outputs(965)) xor (layer0_outputs(698));
    outputs(2077) <= not(layer0_outputs(528));
    outputs(2078) <= not(layer0_outputs(3497));
    outputs(2079) <= not(layer0_outputs(391));
    outputs(2080) <= (layer0_outputs(2785)) and not (layer0_outputs(4024));
    outputs(2081) <= layer0_outputs(1522);
    outputs(2082) <= (layer0_outputs(3228)) xor (layer0_outputs(736));
    outputs(2083) <= not(layer0_outputs(4996)) or (layer0_outputs(1813));
    outputs(2084) <= (layer0_outputs(4806)) and (layer0_outputs(4786));
    outputs(2085) <= not((layer0_outputs(3509)) or (layer0_outputs(2511)));
    outputs(2086) <= not(layer0_outputs(4761));
    outputs(2087) <= layer0_outputs(3649);
    outputs(2088) <= layer0_outputs(641);
    outputs(2089) <= layer0_outputs(1499);
    outputs(2090) <= layer0_outputs(3473);
    outputs(2091) <= layer0_outputs(1389);
    outputs(2092) <= (layer0_outputs(363)) and not (layer0_outputs(4173));
    outputs(2093) <= layer0_outputs(2542);
    outputs(2094) <= layer0_outputs(1644);
    outputs(2095) <= (layer0_outputs(2207)) and not (layer0_outputs(2245));
    outputs(2096) <= not((layer0_outputs(2243)) and (layer0_outputs(2592)));
    outputs(2097) <= layer0_outputs(3504);
    outputs(2098) <= not(layer0_outputs(1437));
    outputs(2099) <= (layer0_outputs(67)) and not (layer0_outputs(950));
    outputs(2100) <= not(layer0_outputs(2865)) or (layer0_outputs(358));
    outputs(2101) <= layer0_outputs(240);
    outputs(2102) <= layer0_outputs(592);
    outputs(2103) <= layer0_outputs(167);
    outputs(2104) <= not(layer0_outputs(275));
    outputs(2105) <= not(layer0_outputs(3598));
    outputs(2106) <= not(layer0_outputs(2664));
    outputs(2107) <= not(layer0_outputs(619));
    outputs(2108) <= not(layer0_outputs(5086));
    outputs(2109) <= layer0_outputs(4823);
    outputs(2110) <= layer0_outputs(3550);
    outputs(2111) <= layer0_outputs(4479);
    outputs(2112) <= not(layer0_outputs(196));
    outputs(2113) <= layer0_outputs(2760);
    outputs(2114) <= not((layer0_outputs(841)) and (layer0_outputs(1331)));
    outputs(2115) <= (layer0_outputs(1647)) and not (layer0_outputs(1198));
    outputs(2116) <= layer0_outputs(4026);
    outputs(2117) <= (layer0_outputs(568)) and (layer0_outputs(4390));
    outputs(2118) <= not(layer0_outputs(1382));
    outputs(2119) <= not(layer0_outputs(660)) or (layer0_outputs(4817));
    outputs(2120) <= not(layer0_outputs(1550));
    outputs(2121) <= (layer0_outputs(281)) and not (layer0_outputs(4074));
    outputs(2122) <= (layer0_outputs(3783)) and not (layer0_outputs(801));
    outputs(2123) <= (layer0_outputs(3254)) and (layer0_outputs(996));
    outputs(2124) <= (layer0_outputs(3044)) or (layer0_outputs(3895));
    outputs(2125) <= (layer0_outputs(4101)) and not (layer0_outputs(3400));
    outputs(2126) <= layer0_outputs(4249);
    outputs(2127) <= not(layer0_outputs(4528));
    outputs(2128) <= layer0_outputs(4479);
    outputs(2129) <= not((layer0_outputs(4569)) xor (layer0_outputs(2110)));
    outputs(2130) <= layer0_outputs(4547);
    outputs(2131) <= layer0_outputs(3902);
    outputs(2132) <= (layer0_outputs(3961)) and not (layer0_outputs(819));
    outputs(2133) <= not(layer0_outputs(3049));
    outputs(2134) <= layer0_outputs(2421);
    outputs(2135) <= not(layer0_outputs(340));
    outputs(2136) <= (layer0_outputs(1708)) and not (layer0_outputs(2242));
    outputs(2137) <= not(layer0_outputs(514));
    outputs(2138) <= layer0_outputs(3727);
    outputs(2139) <= not((layer0_outputs(1146)) xor (layer0_outputs(3658)));
    outputs(2140) <= not(layer0_outputs(3240)) or (layer0_outputs(1185));
    outputs(2141) <= layer0_outputs(2903);
    outputs(2142) <= not(layer0_outputs(3932));
    outputs(2143) <= layer0_outputs(43);
    outputs(2144) <= layer0_outputs(3236);
    outputs(2145) <= not((layer0_outputs(3381)) xor (layer0_outputs(4001)));
    outputs(2146) <= layer0_outputs(3222);
    outputs(2147) <= not(layer0_outputs(193)) or (layer0_outputs(2510));
    outputs(2148) <= layer0_outputs(2666);
    outputs(2149) <= not(layer0_outputs(2307));
    outputs(2150) <= (layer0_outputs(4553)) or (layer0_outputs(3879));
    outputs(2151) <= (layer0_outputs(2189)) and not (layer0_outputs(3616));
    outputs(2152) <= not((layer0_outputs(792)) and (layer0_outputs(4665)));
    outputs(2153) <= not(layer0_outputs(4779));
    outputs(2154) <= not(layer0_outputs(799));
    outputs(2155) <= not((layer0_outputs(4938)) or (layer0_outputs(280)));
    outputs(2156) <= (layer0_outputs(3528)) and not (layer0_outputs(1223));
    outputs(2157) <= (layer0_outputs(5051)) or (layer0_outputs(2955));
    outputs(2158) <= layer0_outputs(3823);
    outputs(2159) <= not((layer0_outputs(644)) or (layer0_outputs(3675)));
    outputs(2160) <= not(layer0_outputs(3524));
    outputs(2161) <= (layer0_outputs(4682)) and not (layer0_outputs(1718));
    outputs(2162) <= not((layer0_outputs(1978)) or (layer0_outputs(3339)));
    outputs(2163) <= not(layer0_outputs(1749));
    outputs(2164) <= not(layer0_outputs(2878)) or (layer0_outputs(2072));
    outputs(2165) <= not((layer0_outputs(3699)) or (layer0_outputs(3764)));
    outputs(2166) <= layer0_outputs(707);
    outputs(2167) <= not((layer0_outputs(4364)) xor (layer0_outputs(2830)));
    outputs(2168) <= not((layer0_outputs(1377)) or (layer0_outputs(3230)));
    outputs(2169) <= (layer0_outputs(2167)) and not (layer0_outputs(3788));
    outputs(2170) <= not((layer0_outputs(4049)) xor (layer0_outputs(3348)));
    outputs(2171) <= not(layer0_outputs(1288));
    outputs(2172) <= (layer0_outputs(4174)) and not (layer0_outputs(417));
    outputs(2173) <= layer0_outputs(3698);
    outputs(2174) <= layer0_outputs(2362);
    outputs(2175) <= layer0_outputs(2580);
    outputs(2176) <= layer0_outputs(2372);
    outputs(2177) <= not(layer0_outputs(3023));
    outputs(2178) <= not(layer0_outputs(4715));
    outputs(2179) <= (layer0_outputs(67)) and not (layer0_outputs(4462));
    outputs(2180) <= not((layer0_outputs(4841)) or (layer0_outputs(3026)));
    outputs(2181) <= (layer0_outputs(261)) and not (layer0_outputs(3827));
    outputs(2182) <= layer0_outputs(3244);
    outputs(2183) <= layer0_outputs(3554);
    outputs(2184) <= layer0_outputs(4702);
    outputs(2185) <= layer0_outputs(3661);
    outputs(2186) <= not(layer0_outputs(4221));
    outputs(2187) <= (layer0_outputs(3238)) xor (layer0_outputs(4676));
    outputs(2188) <= not((layer0_outputs(2421)) xor (layer0_outputs(1721)));
    outputs(2189) <= not(layer0_outputs(2225));
    outputs(2190) <= (layer0_outputs(2281)) and (layer0_outputs(5110));
    outputs(2191) <= layer0_outputs(25);
    outputs(2192) <= layer0_outputs(2602);
    outputs(2193) <= (layer0_outputs(3978)) and (layer0_outputs(3862));
    outputs(2194) <= layer0_outputs(2826);
    outputs(2195) <= not((layer0_outputs(1948)) or (layer0_outputs(939)));
    outputs(2196) <= (layer0_outputs(3064)) or (layer0_outputs(2208));
    outputs(2197) <= layer0_outputs(428);
    outputs(2198) <= not(layer0_outputs(1812)) or (layer0_outputs(3264));
    outputs(2199) <= layer0_outputs(4948);
    outputs(2200) <= layer0_outputs(4093);
    outputs(2201) <= layer0_outputs(2803);
    outputs(2202) <= layer0_outputs(2010);
    outputs(2203) <= not(layer0_outputs(2610));
    outputs(2204) <= not(layer0_outputs(4756)) or (layer0_outputs(430));
    outputs(2205) <= not((layer0_outputs(3852)) or (layer0_outputs(1087)));
    outputs(2206) <= not((layer0_outputs(5041)) xor (layer0_outputs(1177)));
    outputs(2207) <= not((layer0_outputs(918)) and (layer0_outputs(1109)));
    outputs(2208) <= not((layer0_outputs(4555)) or (layer0_outputs(1164)));
    outputs(2209) <= not((layer0_outputs(426)) and (layer0_outputs(224)));
    outputs(2210) <= not(layer0_outputs(3857));
    outputs(2211) <= layer0_outputs(3976);
    outputs(2212) <= layer0_outputs(3869);
    outputs(2213) <= (layer0_outputs(240)) and not (layer0_outputs(2958));
    outputs(2214) <= not(layer0_outputs(1354));
    outputs(2215) <= (layer0_outputs(63)) and not (layer0_outputs(3461));
    outputs(2216) <= layer0_outputs(1885);
    outputs(2217) <= (layer0_outputs(1216)) xor (layer0_outputs(3499));
    outputs(2218) <= not(layer0_outputs(3948)) or (layer0_outputs(3272));
    outputs(2219) <= (layer0_outputs(2115)) and not (layer0_outputs(3987));
    outputs(2220) <= not(layer0_outputs(2112));
    outputs(2221) <= not(layer0_outputs(2783)) or (layer0_outputs(2682));
    outputs(2222) <= not(layer0_outputs(4402)) or (layer0_outputs(4396));
    outputs(2223) <= not((layer0_outputs(2735)) xor (layer0_outputs(805)));
    outputs(2224) <= not(layer0_outputs(799)) or (layer0_outputs(322));
    outputs(2225) <= not(layer0_outputs(1053));
    outputs(2226) <= layer0_outputs(1782);
    outputs(2227) <= layer0_outputs(2431);
    outputs(2228) <= layer0_outputs(2622);
    outputs(2229) <= not(layer0_outputs(3841));
    outputs(2230) <= (layer0_outputs(4112)) and not (layer0_outputs(2759));
    outputs(2231) <= not(layer0_outputs(1961));
    outputs(2232) <= not(layer0_outputs(633));
    outputs(2233) <= (layer0_outputs(3931)) and (layer0_outputs(772));
    outputs(2234) <= not(layer0_outputs(1027));
    outputs(2235) <= layer0_outputs(1758);
    outputs(2236) <= not(layer0_outputs(3643));
    outputs(2237) <= (layer0_outputs(2657)) and (layer0_outputs(4318));
    outputs(2238) <= not(layer0_outputs(3517)) or (layer0_outputs(985));
    outputs(2239) <= not((layer0_outputs(3854)) or (layer0_outputs(3151)));
    outputs(2240) <= not(layer0_outputs(4772));
    outputs(2241) <= (layer0_outputs(2630)) and not (layer0_outputs(3935));
    outputs(2242) <= (layer0_outputs(3750)) or (layer0_outputs(1789));
    outputs(2243) <= not(layer0_outputs(2997));
    outputs(2244) <= not(layer0_outputs(4280)) or (layer0_outputs(1561));
    outputs(2245) <= layer0_outputs(386);
    outputs(2246) <= layer0_outputs(1790);
    outputs(2247) <= (layer0_outputs(4788)) and not (layer0_outputs(3331));
    outputs(2248) <= (layer0_outputs(5010)) and (layer0_outputs(2668));
    outputs(2249) <= not(layer0_outputs(898));
    outputs(2250) <= not(layer0_outputs(2923)) or (layer0_outputs(4728));
    outputs(2251) <= layer0_outputs(3805);
    outputs(2252) <= layer0_outputs(1625);
    outputs(2253) <= layer0_outputs(2440);
    outputs(2254) <= not(layer0_outputs(1660)) or (layer0_outputs(4664));
    outputs(2255) <= (layer0_outputs(4502)) and not (layer0_outputs(1043));
    outputs(2256) <= layer0_outputs(2154);
    outputs(2257) <= (layer0_outputs(659)) and not (layer0_outputs(3108));
    outputs(2258) <= not((layer0_outputs(3239)) and (layer0_outputs(3885)));
    outputs(2259) <= (layer0_outputs(5015)) and not (layer0_outputs(4495));
    outputs(2260) <= not(layer0_outputs(3426));
    outputs(2261) <= layer0_outputs(2472);
    outputs(2262) <= (layer0_outputs(928)) and not (layer0_outputs(5067));
    outputs(2263) <= (layer0_outputs(133)) and (layer0_outputs(4550));
    outputs(2264) <= layer0_outputs(4740);
    outputs(2265) <= (layer0_outputs(4209)) and not (layer0_outputs(3777));
    outputs(2266) <= not((layer0_outputs(875)) xor (layer0_outputs(3016)));
    outputs(2267) <= (layer0_outputs(3611)) and not (layer0_outputs(4322));
    outputs(2268) <= not(layer0_outputs(3674)) or (layer0_outputs(412));
    outputs(2269) <= not(layer0_outputs(453));
    outputs(2270) <= (layer0_outputs(3454)) and (layer0_outputs(1888));
    outputs(2271) <= (layer0_outputs(4612)) xor (layer0_outputs(1387));
    outputs(2272) <= (layer0_outputs(4626)) and not (layer0_outputs(980));
    outputs(2273) <= not((layer0_outputs(1043)) or (layer0_outputs(1749)));
    outputs(2274) <= not(layer0_outputs(2917));
    outputs(2275) <= layer0_outputs(506);
    outputs(2276) <= (layer0_outputs(1511)) and (layer0_outputs(3030));
    outputs(2277) <= not(layer0_outputs(2799));
    outputs(2278) <= (layer0_outputs(4307)) and not (layer0_outputs(4267));
    outputs(2279) <= (layer0_outputs(2428)) and not (layer0_outputs(4678));
    outputs(2280) <= (layer0_outputs(5073)) and not (layer0_outputs(632));
    outputs(2281) <= (layer0_outputs(3476)) and not (layer0_outputs(770));
    outputs(2282) <= not(layer0_outputs(2086));
    outputs(2283) <= layer0_outputs(1221);
    outputs(2284) <= not(layer0_outputs(1460));
    outputs(2285) <= not(layer0_outputs(1839));
    outputs(2286) <= not(layer0_outputs(4669));
    outputs(2287) <= (layer0_outputs(2096)) or (layer0_outputs(2514));
    outputs(2288) <= not(layer0_outputs(1703));
    outputs(2289) <= not(layer0_outputs(417));
    outputs(2290) <= (layer0_outputs(2509)) and (layer0_outputs(2896));
    outputs(2291) <= layer0_outputs(2622);
    outputs(2292) <= (layer0_outputs(3656)) and not (layer0_outputs(2104));
    outputs(2293) <= (layer0_outputs(560)) and not (layer0_outputs(3754));
    outputs(2294) <= (layer0_outputs(1821)) and (layer0_outputs(368));
    outputs(2295) <= not((layer0_outputs(3647)) or (layer0_outputs(3798)));
    outputs(2296) <= layer0_outputs(3634);
    outputs(2297) <= not(layer0_outputs(460));
    outputs(2298) <= not(layer0_outputs(2128)) or (layer0_outputs(2795));
    outputs(2299) <= layer0_outputs(1584);
    outputs(2300) <= (layer0_outputs(2010)) and not (layer0_outputs(2262));
    outputs(2301) <= (layer0_outputs(2755)) and not (layer0_outputs(438));
    outputs(2302) <= layer0_outputs(3175);
    outputs(2303) <= not((layer0_outputs(5092)) xor (layer0_outputs(3646)));
    outputs(2304) <= (layer0_outputs(4799)) or (layer0_outputs(2297));
    outputs(2305) <= not(layer0_outputs(3409));
    outputs(2306) <= not((layer0_outputs(497)) xor (layer0_outputs(4940)));
    outputs(2307) <= (layer0_outputs(4245)) and (layer0_outputs(592));
    outputs(2308) <= not((layer0_outputs(3209)) or (layer0_outputs(1895)));
    outputs(2309) <= (layer0_outputs(763)) and (layer0_outputs(4249));
    outputs(2310) <= layer0_outputs(3904);
    outputs(2311) <= layer0_outputs(879);
    outputs(2312) <= layer0_outputs(104);
    outputs(2313) <= (layer0_outputs(160)) or (layer0_outputs(3473));
    outputs(2314) <= not(layer0_outputs(2105));
    outputs(2315) <= (layer0_outputs(2715)) and (layer0_outputs(4737));
    outputs(2316) <= (layer0_outputs(948)) and not (layer0_outputs(3726));
    outputs(2317) <= layer0_outputs(1754);
    outputs(2318) <= not(layer0_outputs(3691));
    outputs(2319) <= (layer0_outputs(3181)) and (layer0_outputs(1050));
    outputs(2320) <= (layer0_outputs(2827)) and not (layer0_outputs(4));
    outputs(2321) <= (layer0_outputs(692)) xor (layer0_outputs(822));
    outputs(2322) <= not((layer0_outputs(2172)) xor (layer0_outputs(355)));
    outputs(2323) <= not((layer0_outputs(201)) and (layer0_outputs(2468)));
    outputs(2324) <= not(layer0_outputs(2109));
    outputs(2325) <= not(layer0_outputs(660));
    outputs(2326) <= (layer0_outputs(1392)) and not (layer0_outputs(301));
    outputs(2327) <= not(layer0_outputs(1567));
    outputs(2328) <= not(layer0_outputs(778));
    outputs(2329) <= (layer0_outputs(4300)) and (layer0_outputs(3408));
    outputs(2330) <= not(layer0_outputs(1384));
    outputs(2331) <= not((layer0_outputs(4499)) or (layer0_outputs(2338)));
    outputs(2332) <= not((layer0_outputs(647)) or (layer0_outputs(4222)));
    outputs(2333) <= (layer0_outputs(3048)) and (layer0_outputs(3994));
    outputs(2334) <= not((layer0_outputs(2839)) or (layer0_outputs(3163)));
    outputs(2335) <= layer0_outputs(750);
    outputs(2336) <= not(layer0_outputs(4298));
    outputs(2337) <= layer0_outputs(862);
    outputs(2338) <= (layer0_outputs(1083)) and not (layer0_outputs(636));
    outputs(2339) <= layer0_outputs(914);
    outputs(2340) <= (layer0_outputs(1873)) and not (layer0_outputs(2005));
    outputs(2341) <= not(layer0_outputs(3948));
    outputs(2342) <= not((layer0_outputs(2665)) or (layer0_outputs(1694)));
    outputs(2343) <= layer0_outputs(1116);
    outputs(2344) <= not((layer0_outputs(1640)) or (layer0_outputs(3400)));
    outputs(2345) <= layer0_outputs(1341);
    outputs(2346) <= (layer0_outputs(4473)) and not (layer0_outputs(4841));
    outputs(2347) <= (layer0_outputs(1381)) and not (layer0_outputs(1272));
    outputs(2348) <= layer0_outputs(159);
    outputs(2349) <= layer0_outputs(322);
    outputs(2350) <= layer0_outputs(4515);
    outputs(2351) <= (layer0_outputs(4396)) or (layer0_outputs(1099));
    outputs(2352) <= not((layer0_outputs(4946)) or (layer0_outputs(1161)));
    outputs(2353) <= (layer0_outputs(321)) xor (layer0_outputs(4120));
    outputs(2354) <= layer0_outputs(3897);
    outputs(2355) <= (layer0_outputs(1947)) and not (layer0_outputs(4413));
    outputs(2356) <= (layer0_outputs(3063)) or (layer0_outputs(3241));
    outputs(2357) <= layer0_outputs(4185);
    outputs(2358) <= (layer0_outputs(19)) and (layer0_outputs(3812));
    outputs(2359) <= not(layer0_outputs(2059));
    outputs(2360) <= not(layer0_outputs(1875));
    outputs(2361) <= layer0_outputs(1766);
    outputs(2362) <= layer0_outputs(1780);
    outputs(2363) <= layer0_outputs(1699);
    outputs(2364) <= layer0_outputs(1369);
    outputs(2365) <= (layer0_outputs(1766)) xor (layer0_outputs(1267));
    outputs(2366) <= not((layer0_outputs(4446)) or (layer0_outputs(499)));
    outputs(2367) <= not((layer0_outputs(1978)) and (layer0_outputs(876)));
    outputs(2368) <= not(layer0_outputs(1361));
    outputs(2369) <= layer0_outputs(4489);
    outputs(2370) <= layer0_outputs(745);
    outputs(2371) <= (layer0_outputs(3143)) and (layer0_outputs(2593));
    outputs(2372) <= not((layer0_outputs(3633)) or (layer0_outputs(4168)));
    outputs(2373) <= (layer0_outputs(4985)) and (layer0_outputs(173));
    outputs(2374) <= not((layer0_outputs(3612)) or (layer0_outputs(1379)));
    outputs(2375) <= layer0_outputs(4393);
    outputs(2376) <= not(layer0_outputs(2114)) or (layer0_outputs(1705));
    outputs(2377) <= not(layer0_outputs(4833));
    outputs(2378) <= (layer0_outputs(4269)) and not (layer0_outputs(2037));
    outputs(2379) <= not(layer0_outputs(4270)) or (layer0_outputs(1039));
    outputs(2380) <= (layer0_outputs(4326)) xor (layer0_outputs(3019));
    outputs(2381) <= layer0_outputs(2337);
    outputs(2382) <= (layer0_outputs(2048)) xor (layer0_outputs(1434));
    outputs(2383) <= (layer0_outputs(4936)) and not (layer0_outputs(3014));
    outputs(2384) <= (layer0_outputs(1515)) and not (layer0_outputs(4901));
    outputs(2385) <= not((layer0_outputs(4161)) xor (layer0_outputs(5046)));
    outputs(2386) <= layer0_outputs(3210);
    outputs(2387) <= (layer0_outputs(1608)) and not (layer0_outputs(3443));
    outputs(2388) <= (layer0_outputs(2644)) and (layer0_outputs(4554));
    outputs(2389) <= not((layer0_outputs(5050)) or (layer0_outputs(4419)));
    outputs(2390) <= layer0_outputs(5051);
    outputs(2391) <= not(layer0_outputs(591));
    outputs(2392) <= not(layer0_outputs(1471));
    outputs(2393) <= layer0_outputs(4793);
    outputs(2394) <= (layer0_outputs(2234)) and not (layer0_outputs(2471));
    outputs(2395) <= not(layer0_outputs(1311)) or (layer0_outputs(1918));
    outputs(2396) <= layer0_outputs(4541);
    outputs(2397) <= not((layer0_outputs(1148)) or (layer0_outputs(2467)));
    outputs(2398) <= (layer0_outputs(4272)) and not (layer0_outputs(839));
    outputs(2399) <= not((layer0_outputs(4763)) and (layer0_outputs(648)));
    outputs(2400) <= (layer0_outputs(195)) and not (layer0_outputs(2134));
    outputs(2401) <= not(layer0_outputs(3108));
    outputs(2402) <= not((layer0_outputs(3128)) or (layer0_outputs(2577)));
    outputs(2403) <= (layer0_outputs(2498)) and not (layer0_outputs(3616));
    outputs(2404) <= not((layer0_outputs(3514)) or (layer0_outputs(500)));
    outputs(2405) <= not((layer0_outputs(3059)) or (layer0_outputs(3153)));
    outputs(2406) <= (layer0_outputs(4328)) xor (layer0_outputs(4973));
    outputs(2407) <= (layer0_outputs(1695)) and (layer0_outputs(3478));
    outputs(2408) <= layer0_outputs(3568);
    outputs(2409) <= (layer0_outputs(2938)) and not (layer0_outputs(146));
    outputs(2410) <= not((layer0_outputs(470)) or (layer0_outputs(620)));
    outputs(2411) <= (layer0_outputs(4560)) xor (layer0_outputs(1905));
    outputs(2412) <= not(layer0_outputs(1752));
    outputs(2413) <= not(layer0_outputs(252));
    outputs(2414) <= layer0_outputs(4733);
    outputs(2415) <= not((layer0_outputs(1062)) and (layer0_outputs(1287)));
    outputs(2416) <= layer0_outputs(1560);
    outputs(2417) <= not((layer0_outputs(302)) or (layer0_outputs(1788)));
    outputs(2418) <= not(layer0_outputs(4491));
    outputs(2419) <= not(layer0_outputs(1961)) or (layer0_outputs(4095));
    outputs(2420) <= not((layer0_outputs(1638)) xor (layer0_outputs(2786)));
    outputs(2421) <= layer0_outputs(613);
    outputs(2422) <= (layer0_outputs(4170)) and not (layer0_outputs(1120));
    outputs(2423) <= (layer0_outputs(2202)) and not (layer0_outputs(4448));
    outputs(2424) <= not(layer0_outputs(1949)) or (layer0_outputs(3027));
    outputs(2425) <= not(layer0_outputs(1451));
    outputs(2426) <= not((layer0_outputs(3196)) xor (layer0_outputs(2860)));
    outputs(2427) <= layer0_outputs(1607);
    outputs(2428) <= layer0_outputs(1954);
    outputs(2429) <= layer0_outputs(2121);
    outputs(2430) <= layer0_outputs(187);
    outputs(2431) <= layer0_outputs(1247);
    outputs(2432) <= layer0_outputs(1877);
    outputs(2433) <= not(layer0_outputs(3975));
    outputs(2434) <= not((layer0_outputs(1061)) and (layer0_outputs(674)));
    outputs(2435) <= not((layer0_outputs(3237)) xor (layer0_outputs(868)));
    outputs(2436) <= layer0_outputs(116);
    outputs(2437) <= layer0_outputs(1581);
    outputs(2438) <= not(layer0_outputs(1601)) or (layer0_outputs(229));
    outputs(2439) <= layer0_outputs(938);
    outputs(2440) <= not((layer0_outputs(3913)) or (layer0_outputs(4508)));
    outputs(2441) <= (layer0_outputs(3592)) and not (layer0_outputs(622));
    outputs(2442) <= (layer0_outputs(688)) and (layer0_outputs(2778));
    outputs(2443) <= not((layer0_outputs(1684)) or (layer0_outputs(2432)));
    outputs(2444) <= not((layer0_outputs(828)) or (layer0_outputs(1712)));
    outputs(2445) <= (layer0_outputs(1841)) and not (layer0_outputs(100));
    outputs(2446) <= not((layer0_outputs(1023)) and (layer0_outputs(3434)));
    outputs(2447) <= (layer0_outputs(3149)) xor (layer0_outputs(3845));
    outputs(2448) <= not(layer0_outputs(2441));
    outputs(2449) <= not(layer0_outputs(1382));
    outputs(2450) <= layer0_outputs(2847);
    outputs(2451) <= not(layer0_outputs(2957));
    outputs(2452) <= not(layer0_outputs(2942)) or (layer0_outputs(3629));
    outputs(2453) <= not(layer0_outputs(1985));
    outputs(2454) <= layer0_outputs(997);
    outputs(2455) <= not(layer0_outputs(4757)) or (layer0_outputs(787));
    outputs(2456) <= not(layer0_outputs(4614));
    outputs(2457) <= not(layer0_outputs(1033));
    outputs(2458) <= layer0_outputs(4743);
    outputs(2459) <= not((layer0_outputs(4477)) xor (layer0_outputs(3795)));
    outputs(2460) <= (layer0_outputs(2264)) and not (layer0_outputs(916));
    outputs(2461) <= not(layer0_outputs(1580)) or (layer0_outputs(3810));
    outputs(2462) <= layer0_outputs(5088);
    outputs(2463) <= (layer0_outputs(2313)) and not (layer0_outputs(4013));
    outputs(2464) <= not((layer0_outputs(21)) and (layer0_outputs(4061)));
    outputs(2465) <= not(layer0_outputs(2235)) or (layer0_outputs(2712));
    outputs(2466) <= (layer0_outputs(997)) or (layer0_outputs(909));
    outputs(2467) <= not(layer0_outputs(1229));
    outputs(2468) <= (layer0_outputs(1039)) and not (layer0_outputs(4476));
    outputs(2469) <= (layer0_outputs(4442)) and not (layer0_outputs(4871));
    outputs(2470) <= (layer0_outputs(2994)) and (layer0_outputs(2899));
    outputs(2471) <= not((layer0_outputs(4315)) or (layer0_outputs(2070)));
    outputs(2472) <= not(layer0_outputs(4137)) or (layer0_outputs(442));
    outputs(2473) <= (layer0_outputs(1135)) xor (layer0_outputs(4642));
    outputs(2474) <= not((layer0_outputs(2802)) or (layer0_outputs(82)));
    outputs(2475) <= not(layer0_outputs(2897)) or (layer0_outputs(4028));
    outputs(2476) <= (layer0_outputs(3185)) and not (layer0_outputs(3428));
    outputs(2477) <= (layer0_outputs(2232)) and not (layer0_outputs(4142));
    outputs(2478) <= not((layer0_outputs(181)) and (layer0_outputs(2322)));
    outputs(2479) <= not((layer0_outputs(960)) or (layer0_outputs(4096)));
    outputs(2480) <= not(layer0_outputs(1941));
    outputs(2481) <= layer0_outputs(4141);
    outputs(2482) <= not(layer0_outputs(3861));
    outputs(2483) <= not(layer0_outputs(1171));
    outputs(2484) <= (layer0_outputs(5053)) and not (layer0_outputs(4897));
    outputs(2485) <= (layer0_outputs(506)) and (layer0_outputs(2189));
    outputs(2486) <= not(layer0_outputs(3043));
    outputs(2487) <= not((layer0_outputs(1275)) or (layer0_outputs(3675)));
    outputs(2488) <= not((layer0_outputs(5081)) xor (layer0_outputs(1211)));
    outputs(2489) <= not(layer0_outputs(4540));
    outputs(2490) <= not((layer0_outputs(3182)) and (layer0_outputs(445)));
    outputs(2491) <= not(layer0_outputs(1482));
    outputs(2492) <= not(layer0_outputs(4472));
    outputs(2493) <= layer0_outputs(2781);
    outputs(2494) <= not(layer0_outputs(3617));
    outputs(2495) <= not((layer0_outputs(4518)) and (layer0_outputs(2744)));
    outputs(2496) <= layer0_outputs(3157);
    outputs(2497) <= (layer0_outputs(2131)) and not (layer0_outputs(3852));
    outputs(2498) <= layer0_outputs(1284);
    outputs(2499) <= not((layer0_outputs(4341)) or (layer0_outputs(3080)));
    outputs(2500) <= (layer0_outputs(3963)) and not (layer0_outputs(3249));
    outputs(2501) <= (layer0_outputs(4954)) and not (layer0_outputs(4641));
    outputs(2502) <= not((layer0_outputs(2485)) xor (layer0_outputs(2893)));
    outputs(2503) <= layer0_outputs(3403);
    outputs(2504) <= not(layer0_outputs(96));
    outputs(2505) <= (layer0_outputs(4899)) and not (layer0_outputs(255));
    outputs(2506) <= (layer0_outputs(3070)) and not (layer0_outputs(2448));
    outputs(2507) <= not(layer0_outputs(4401));
    outputs(2508) <= not(layer0_outputs(3943));
    outputs(2509) <= (layer0_outputs(195)) and (layer0_outputs(1200));
    outputs(2510) <= not((layer0_outputs(3086)) or (layer0_outputs(3985)));
    outputs(2511) <= not(layer0_outputs(856));
    outputs(2512) <= layer0_outputs(3914);
    outputs(2513) <= not((layer0_outputs(3864)) xor (layer0_outputs(3062)));
    outputs(2514) <= (layer0_outputs(4825)) and (layer0_outputs(1501));
    outputs(2515) <= not(layer0_outputs(1271));
    outputs(2516) <= layer0_outputs(4839);
    outputs(2517) <= not((layer0_outputs(582)) and (layer0_outputs(488)));
    outputs(2518) <= not(layer0_outputs(4524));
    outputs(2519) <= layer0_outputs(833);
    outputs(2520) <= layer0_outputs(1701);
    outputs(2521) <= (layer0_outputs(4261)) and not (layer0_outputs(1340));
    outputs(2522) <= not(layer0_outputs(2815));
    outputs(2523) <= not(layer0_outputs(664));
    outputs(2524) <= not((layer0_outputs(2127)) or (layer0_outputs(1495)));
    outputs(2525) <= not(layer0_outputs(1670)) or (layer0_outputs(211));
    outputs(2526) <= not((layer0_outputs(2769)) or (layer0_outputs(1479)));
    outputs(2527) <= (layer0_outputs(2558)) xor (layer0_outputs(1282));
    outputs(2528) <= not(layer0_outputs(1063));
    outputs(2529) <= (layer0_outputs(173)) and not (layer0_outputs(2293));
    outputs(2530) <= layer0_outputs(2975);
    outputs(2531) <= not(layer0_outputs(3969));
    outputs(2532) <= not(layer0_outputs(4522));
    outputs(2533) <= (layer0_outputs(465)) and not (layer0_outputs(1202));
    outputs(2534) <= not(layer0_outputs(491));
    outputs(2535) <= layer0_outputs(4353);
    outputs(2536) <= (layer0_outputs(4220)) xor (layer0_outputs(1722));
    outputs(2537) <= layer0_outputs(3445);
    outputs(2538) <= (layer0_outputs(478)) or (layer0_outputs(1125));
    outputs(2539) <= (layer0_outputs(646)) or (layer0_outputs(4515));
    outputs(2540) <= (layer0_outputs(5016)) and (layer0_outputs(2615));
    outputs(2541) <= layer0_outputs(3495);
    outputs(2542) <= layer0_outputs(119);
    outputs(2543) <= (layer0_outputs(4550)) or (layer0_outputs(4624));
    outputs(2544) <= not((layer0_outputs(4198)) xor (layer0_outputs(1308)));
    outputs(2545) <= not(layer0_outputs(2816)) or (layer0_outputs(2239));
    outputs(2546) <= not((layer0_outputs(1653)) or (layer0_outputs(1612)));
    outputs(2547) <= (layer0_outputs(2549)) and not (layer0_outputs(3353));
    outputs(2548) <= not(layer0_outputs(874)) or (layer0_outputs(2718));
    outputs(2549) <= layer0_outputs(547);
    outputs(2550) <= layer0_outputs(4055);
    outputs(2551) <= layer0_outputs(3890);
    outputs(2552) <= not(layer0_outputs(1990));
    outputs(2553) <= layer0_outputs(1370);
    outputs(2554) <= (layer0_outputs(1408)) and not (layer0_outputs(1348));
    outputs(2555) <= layer0_outputs(3398);
    outputs(2556) <= not((layer0_outputs(4551)) or (layer0_outputs(3341)));
    outputs(2557) <= (layer0_outputs(1013)) or (layer0_outputs(4834));
    outputs(2558) <= (layer0_outputs(724)) xor (layer0_outputs(1582));
    outputs(2559) <= not(layer0_outputs(110)) or (layer0_outputs(2296));
    outputs(2560) <= not(layer0_outputs(1794)) or (layer0_outputs(1924));
    outputs(2561) <= not(layer0_outputs(5024));
    outputs(2562) <= layer0_outputs(3729);
    outputs(2563) <= not((layer0_outputs(2931)) xor (layer0_outputs(1697)));
    outputs(2564) <= (layer0_outputs(3052)) and (layer0_outputs(1723));
    outputs(2565) <= not(layer0_outputs(3853));
    outputs(2566) <= layer0_outputs(1087);
    outputs(2567) <= not((layer0_outputs(1963)) xor (layer0_outputs(1757)));
    outputs(2568) <= layer0_outputs(2328);
    outputs(2569) <= layer0_outputs(2524);
    outputs(2570) <= (layer0_outputs(4705)) and not (layer0_outputs(4439));
    outputs(2571) <= not(layer0_outputs(4662));
    outputs(2572) <= (layer0_outputs(554)) and not (layer0_outputs(257));
    outputs(2573) <= not(layer0_outputs(2123));
    outputs(2574) <= (layer0_outputs(2144)) xor (layer0_outputs(4889));
    outputs(2575) <= not((layer0_outputs(3766)) xor (layer0_outputs(1175)));
    outputs(2576) <= not(layer0_outputs(1807));
    outputs(2577) <= (layer0_outputs(650)) xor (layer0_outputs(2399));
    outputs(2578) <= (layer0_outputs(4633)) or (layer0_outputs(4730));
    outputs(2579) <= not(layer0_outputs(4436));
    outputs(2580) <= (layer0_outputs(2794)) and not (layer0_outputs(3290));
    outputs(2581) <= layer0_outputs(2251);
    outputs(2582) <= not(layer0_outputs(2836)) or (layer0_outputs(146));
    outputs(2583) <= not(layer0_outputs(618)) or (layer0_outputs(4654));
    outputs(2584) <= not(layer0_outputs(1889));
    outputs(2585) <= (layer0_outputs(4240)) or (layer0_outputs(2382));
    outputs(2586) <= not(layer0_outputs(3329));
    outputs(2587) <= layer0_outputs(2228);
    outputs(2588) <= (layer0_outputs(784)) and not (layer0_outputs(743));
    outputs(2589) <= not(layer0_outputs(366));
    outputs(2590) <= not((layer0_outputs(4982)) or (layer0_outputs(4131)));
    outputs(2591) <= (layer0_outputs(4203)) xor (layer0_outputs(856));
    outputs(2592) <= (layer0_outputs(1458)) and not (layer0_outputs(2649));
    outputs(2593) <= not(layer0_outputs(5021));
    outputs(2594) <= layer0_outputs(2641);
    outputs(2595) <= not((layer0_outputs(1843)) and (layer0_outputs(4919)));
    outputs(2596) <= not((layer0_outputs(2388)) or (layer0_outputs(1875)));
    outputs(2597) <= layer0_outputs(4350);
    outputs(2598) <= not((layer0_outputs(1730)) xor (layer0_outputs(1082)));
    outputs(2599) <= not(layer0_outputs(4659));
    outputs(2600) <= not(layer0_outputs(214));
    outputs(2601) <= not((layer0_outputs(4670)) xor (layer0_outputs(1366)));
    outputs(2602) <= (layer0_outputs(270)) and not (layer0_outputs(3677));
    outputs(2603) <= (layer0_outputs(393)) and (layer0_outputs(3057));
    outputs(2604) <= not((layer0_outputs(5094)) xor (layer0_outputs(254)));
    outputs(2605) <= (layer0_outputs(453)) and (layer0_outputs(2165));
    outputs(2606) <= not((layer0_outputs(1209)) xor (layer0_outputs(4895)));
    outputs(2607) <= not((layer0_outputs(3382)) xor (layer0_outputs(3451)));
    outputs(2608) <= not(layer0_outputs(729));
    outputs(2609) <= layer0_outputs(4949);
    outputs(2610) <= layer0_outputs(1752);
    outputs(2611) <= not(layer0_outputs(755));
    outputs(2612) <= layer0_outputs(4343);
    outputs(2613) <= layer0_outputs(4687);
    outputs(2614) <= not((layer0_outputs(824)) or (layer0_outputs(1980)));
    outputs(2615) <= (layer0_outputs(3394)) xor (layer0_outputs(4389));
    outputs(2616) <= not(layer0_outputs(3489));
    outputs(2617) <= not(layer0_outputs(311));
    outputs(2618) <= not((layer0_outputs(2333)) xor (layer0_outputs(99)));
    outputs(2619) <= layer0_outputs(3388);
    outputs(2620) <= not((layer0_outputs(1628)) and (layer0_outputs(3556)));
    outputs(2621) <= (layer0_outputs(4378)) and not (layer0_outputs(2974));
    outputs(2622) <= (layer0_outputs(3431)) xor (layer0_outputs(3257));
    outputs(2623) <= not(layer0_outputs(1137));
    outputs(2624) <= layer0_outputs(4788);
    outputs(2625) <= not(layer0_outputs(1351));
    outputs(2626) <= layer0_outputs(4766);
    outputs(2627) <= layer0_outputs(1810);
    outputs(2628) <= (layer0_outputs(2906)) and not (layer0_outputs(1883));
    outputs(2629) <= (layer0_outputs(3179)) and not (layer0_outputs(2825));
    outputs(2630) <= (layer0_outputs(78)) xor (layer0_outputs(3846));
    outputs(2631) <= (layer0_outputs(3241)) and not (layer0_outputs(1604));
    outputs(2632) <= layer0_outputs(1148);
    outputs(2633) <= (layer0_outputs(4349)) or (layer0_outputs(1672));
    outputs(2634) <= not((layer0_outputs(1339)) and (layer0_outputs(4586)));
    outputs(2635) <= not((layer0_outputs(294)) xor (layer0_outputs(4602)));
    outputs(2636) <= (layer0_outputs(1397)) and (layer0_outputs(1027));
    outputs(2637) <= (layer0_outputs(297)) and (layer0_outputs(4428));
    outputs(2638) <= (layer0_outputs(198)) xor (layer0_outputs(2084));
    outputs(2639) <= not(layer0_outputs(3295));
    outputs(2640) <= not(layer0_outputs(2302));
    outputs(2641) <= (layer0_outputs(3055)) and not (layer0_outputs(5112));
    outputs(2642) <= layer0_outputs(1402);
    outputs(2643) <= (layer0_outputs(2943)) and (layer0_outputs(2407));
    outputs(2644) <= not(layer0_outputs(4900));
    outputs(2645) <= (layer0_outputs(2423)) and not (layer0_outputs(2065));
    outputs(2646) <= not(layer0_outputs(4365));
    outputs(2647) <= (layer0_outputs(3785)) or (layer0_outputs(1460));
    outputs(2648) <= (layer0_outputs(1772)) and not (layer0_outputs(929));
    outputs(2649) <= (layer0_outputs(2570)) xor (layer0_outputs(2461));
    outputs(2650) <= not((layer0_outputs(1199)) xor (layer0_outputs(2193)));
    outputs(2651) <= not((layer0_outputs(2614)) xor (layer0_outputs(3035)));
    outputs(2652) <= not(layer0_outputs(1919)) or (layer0_outputs(2550));
    outputs(2653) <= not((layer0_outputs(3013)) xor (layer0_outputs(2766)));
    outputs(2654) <= not(layer0_outputs(3704));
    outputs(2655) <= not((layer0_outputs(812)) xor (layer0_outputs(3237)));
    outputs(2656) <= not(layer0_outputs(4644)) or (layer0_outputs(144));
    outputs(2657) <= not((layer0_outputs(3955)) xor (layer0_outputs(2896)));
    outputs(2658) <= (layer0_outputs(3327)) xor (layer0_outputs(4932));
    outputs(2659) <= not((layer0_outputs(975)) and (layer0_outputs(4943)));
    outputs(2660) <= layer0_outputs(4853);
    outputs(2661) <= layer0_outputs(2080);
    outputs(2662) <= not((layer0_outputs(3492)) or (layer0_outputs(2207)));
    outputs(2663) <= not(layer0_outputs(3926)) or (layer0_outputs(4322));
    outputs(2664) <= not((layer0_outputs(53)) xor (layer0_outputs(3892)));
    outputs(2665) <= layer0_outputs(2521);
    outputs(2666) <= not((layer0_outputs(3091)) xor (layer0_outputs(2550)));
    outputs(2667) <= not(layer0_outputs(3045)) or (layer0_outputs(207));
    outputs(2668) <= not(layer0_outputs(1048));
    outputs(2669) <= not(layer0_outputs(4314));
    outputs(2670) <= (layer0_outputs(2922)) and (layer0_outputs(2758));
    outputs(2671) <= (layer0_outputs(293)) xor (layer0_outputs(4366));
    outputs(2672) <= not(layer0_outputs(2473)) or (layer0_outputs(4836));
    outputs(2673) <= (layer0_outputs(3776)) and (layer0_outputs(292));
    outputs(2674) <= not(layer0_outputs(2815));
    outputs(2675) <= (layer0_outputs(3521)) xor (layer0_outputs(3501));
    outputs(2676) <= (layer0_outputs(2468)) and not (layer0_outputs(4627));
    outputs(2677) <= not(layer0_outputs(177));
    outputs(2678) <= layer0_outputs(3261);
    outputs(2679) <= layer0_outputs(3189);
    outputs(2680) <= not((layer0_outputs(1648)) and (layer0_outputs(1814)));
    outputs(2681) <= not(layer0_outputs(2559));
    outputs(2682) <= layer0_outputs(2012);
    outputs(2683) <= layer0_outputs(4831);
    outputs(2684) <= (layer0_outputs(3091)) xor (layer0_outputs(4500));
    outputs(2685) <= layer0_outputs(2270);
    outputs(2686) <= (layer0_outputs(1383)) xor (layer0_outputs(2945));
    outputs(2687) <= not(layer0_outputs(4122));
    outputs(2688) <= not((layer0_outputs(3133)) xor (layer0_outputs(2905)));
    outputs(2689) <= (layer0_outputs(943)) xor (layer0_outputs(1641));
    outputs(2690) <= not((layer0_outputs(3203)) or (layer0_outputs(4217)));
    outputs(2691) <= (layer0_outputs(892)) and (layer0_outputs(857));
    outputs(2692) <= layer0_outputs(4023);
    outputs(2693) <= layer0_outputs(561);
    outputs(2694) <= not(layer0_outputs(1687));
    outputs(2695) <= layer0_outputs(2843);
    outputs(2696) <= (layer0_outputs(1663)) and not (layer0_outputs(2659));
    outputs(2697) <= not((layer0_outputs(3617)) xor (layer0_outputs(1393)));
    outputs(2698) <= (layer0_outputs(2915)) and (layer0_outputs(530));
    outputs(2699) <= not(layer0_outputs(4188));
    outputs(2700) <= (layer0_outputs(1863)) and (layer0_outputs(2643));
    outputs(2701) <= not(layer0_outputs(463));
    outputs(2702) <= (layer0_outputs(3187)) and (layer0_outputs(3051));
    outputs(2703) <= (layer0_outputs(4064)) and not (layer0_outputs(3876));
    outputs(2704) <= not(layer0_outputs(1577));
    outputs(2705) <= not(layer0_outputs(4482));
    outputs(2706) <= not(layer0_outputs(4341));
    outputs(2707) <= (layer0_outputs(5009)) xor (layer0_outputs(4966));
    outputs(2708) <= not((layer0_outputs(1834)) and (layer0_outputs(5077)));
    outputs(2709) <= (layer0_outputs(3422)) or (layer0_outputs(2150));
    outputs(2710) <= not(layer0_outputs(3004));
    outputs(2711) <= not((layer0_outputs(2980)) xor (layer0_outputs(3813)));
    outputs(2712) <= (layer0_outputs(603)) and (layer0_outputs(3111));
    outputs(2713) <= layer0_outputs(125);
    outputs(2714) <= not((layer0_outputs(1263)) xor (layer0_outputs(828)));
    outputs(2715) <= layer0_outputs(3071);
    outputs(2716) <= (layer0_outputs(3013)) xor (layer0_outputs(4692));
    outputs(2717) <= layer0_outputs(690);
    outputs(2718) <= (layer0_outputs(2965)) and not (layer0_outputs(4237));
    outputs(2719) <= not(layer0_outputs(4263));
    outputs(2720) <= not(layer0_outputs(1052));
    outputs(2721) <= (layer0_outputs(5)) xor (layer0_outputs(1162));
    outputs(2722) <= (layer0_outputs(4670)) xor (layer0_outputs(4620));
    outputs(2723) <= not(layer0_outputs(4045));
    outputs(2724) <= (layer0_outputs(2215)) and not (layer0_outputs(3073));
    outputs(2725) <= (layer0_outputs(1602)) or (layer0_outputs(4267));
    outputs(2726) <= (layer0_outputs(3860)) and (layer0_outputs(368));
    outputs(2727) <= not(layer0_outputs(2825));
    outputs(2728) <= not((layer0_outputs(4573)) or (layer0_outputs(4803)));
    outputs(2729) <= not(layer0_outputs(2807));
    outputs(2730) <= (layer0_outputs(2742)) and not (layer0_outputs(3324));
    outputs(2731) <= (layer0_outputs(4538)) and (layer0_outputs(520));
    outputs(2732) <= (layer0_outputs(1387)) and (layer0_outputs(1753));
    outputs(2733) <= (layer0_outputs(687)) and not (layer0_outputs(2565));
    outputs(2734) <= layer0_outputs(4107);
    outputs(2735) <= not(layer0_outputs(1407));
    outputs(2736) <= (layer0_outputs(3781)) and (layer0_outputs(2456));
    outputs(2737) <= not(layer0_outputs(4171));
    outputs(2738) <= not((layer0_outputs(3439)) or (layer0_outputs(2159)));
    outputs(2739) <= layer0_outputs(1784);
    outputs(2740) <= layer0_outputs(715);
    outputs(2741) <= layer0_outputs(2621);
    outputs(2742) <= (layer0_outputs(3685)) and (layer0_outputs(4965));
    outputs(2743) <= layer0_outputs(3139);
    outputs(2744) <= not(layer0_outputs(3979));
    outputs(2745) <= not((layer0_outputs(2854)) and (layer0_outputs(904)));
    outputs(2746) <= not(layer0_outputs(705)) or (layer0_outputs(129));
    outputs(2747) <= not(layer0_outputs(4536));
    outputs(2748) <= layer0_outputs(4658);
    outputs(2749) <= not((layer0_outputs(3150)) and (layer0_outputs(741)));
    outputs(2750) <= not(layer0_outputs(627));
    outputs(2751) <= layer0_outputs(1122);
    outputs(2752) <= (layer0_outputs(2574)) and not (layer0_outputs(583));
    outputs(2753) <= layer0_outputs(3057);
    outputs(2754) <= layer0_outputs(4653);
    outputs(2755) <= not(layer0_outputs(1060));
    outputs(2756) <= (layer0_outputs(1650)) xor (layer0_outputs(1897));
    outputs(2757) <= layer0_outputs(3986);
    outputs(2758) <= (layer0_outputs(253)) and not (layer0_outputs(1415));
    outputs(2759) <= not(layer0_outputs(5080));
    outputs(2760) <= not(layer0_outputs(3613));
    outputs(2761) <= (layer0_outputs(2725)) xor (layer0_outputs(759));
    outputs(2762) <= (layer0_outputs(3638)) and not (layer0_outputs(4439));
    outputs(2763) <= layer0_outputs(1946);
    outputs(2764) <= (layer0_outputs(3337)) and not (layer0_outputs(4876));
    outputs(2765) <= not(layer0_outputs(926));
    outputs(2766) <= not((layer0_outputs(584)) or (layer0_outputs(3128)));
    outputs(2767) <= not((layer0_outputs(3223)) and (layer0_outputs(610)));
    outputs(2768) <= not(layer0_outputs(2246));
    outputs(2769) <= not(layer0_outputs(2365));
    outputs(2770) <= (layer0_outputs(1220)) and not (layer0_outputs(2206));
    outputs(2771) <= layer0_outputs(297);
    outputs(2772) <= not(layer0_outputs(3594));
    outputs(2773) <= not((layer0_outputs(2244)) xor (layer0_outputs(513)));
    outputs(2774) <= not((layer0_outputs(2757)) or (layer0_outputs(4021)));
    outputs(2775) <= not(layer0_outputs(2367)) or (layer0_outputs(1904));
    outputs(2776) <= layer0_outputs(310);
    outputs(2777) <= not(layer0_outputs(1933));
    outputs(2778) <= (layer0_outputs(3977)) xor (layer0_outputs(3996));
    outputs(2779) <= not((layer0_outputs(4826)) and (layer0_outputs(679)));
    outputs(2780) <= not(layer0_outputs(3075));
    outputs(2781) <= (layer0_outputs(527)) and not (layer0_outputs(4034));
    outputs(2782) <= (layer0_outputs(4225)) xor (layer0_outputs(3751));
    outputs(2783) <= not((layer0_outputs(2488)) xor (layer0_outputs(739)));
    outputs(2784) <= layer0_outputs(968);
    outputs(2785) <= (layer0_outputs(1809)) and not (layer0_outputs(4244));
    outputs(2786) <= layer0_outputs(1389);
    outputs(2787) <= not(layer0_outputs(1324));
    outputs(2788) <= (layer0_outputs(1465)) and not (layer0_outputs(2269));
    outputs(2789) <= not(layer0_outputs(435));
    outputs(2790) <= layer0_outputs(3266);
    outputs(2791) <= not(layer0_outputs(203)) or (layer0_outputs(4498));
    outputs(2792) <= not(layer0_outputs(3719));
    outputs(2793) <= not((layer0_outputs(4623)) and (layer0_outputs(425)));
    outputs(2794) <= not((layer0_outputs(4465)) xor (layer0_outputs(3856)));
    outputs(2795) <= not(layer0_outputs(3467)) or (layer0_outputs(889));
    outputs(2796) <= not((layer0_outputs(3121)) xor (layer0_outputs(1755)));
    outputs(2797) <= not(layer0_outputs(3086));
    outputs(2798) <= not((layer0_outputs(4864)) xor (layer0_outputs(4090)));
    outputs(2799) <= (layer0_outputs(4498)) xor (layer0_outputs(4733));
    outputs(2800) <= (layer0_outputs(1067)) and not (layer0_outputs(4387));
    outputs(2801) <= not((layer0_outputs(98)) xor (layer0_outputs(9)));
    outputs(2802) <= layer0_outputs(3809);
    outputs(2803) <= (layer0_outputs(3185)) xor (layer0_outputs(2487));
    outputs(2804) <= (layer0_outputs(2279)) and (layer0_outputs(446));
    outputs(2805) <= not(layer0_outputs(2056));
    outputs(2806) <= not(layer0_outputs(3374));
    outputs(2807) <= not((layer0_outputs(4643)) xor (layer0_outputs(4043)));
    outputs(2808) <= not(layer0_outputs(2463));
    outputs(2809) <= (layer0_outputs(2520)) or (layer0_outputs(456));
    outputs(2810) <= (layer0_outputs(4011)) xor (layer0_outputs(178));
    outputs(2811) <= (layer0_outputs(4532)) xor (layer0_outputs(1635));
    outputs(2812) <= (layer0_outputs(3934)) or (layer0_outputs(4162));
    outputs(2813) <= not(layer0_outputs(2173)) or (layer0_outputs(5052));
    outputs(2814) <= not((layer0_outputs(543)) xor (layer0_outputs(1315)));
    outputs(2815) <= layer0_outputs(1396);
    outputs(2816) <= layer0_outputs(2177);
    outputs(2817) <= layer0_outputs(4289);
    outputs(2818) <= not(layer0_outputs(4196));
    outputs(2819) <= not(layer0_outputs(1263)) or (layer0_outputs(3964));
    outputs(2820) <= not(layer0_outputs(178));
    outputs(2821) <= (layer0_outputs(3204)) or (layer0_outputs(3414));
    outputs(2822) <= not((layer0_outputs(1223)) xor (layer0_outputs(568)));
    outputs(2823) <= (layer0_outputs(2217)) and not (layer0_outputs(52));
    outputs(2824) <= layer0_outputs(4210);
    outputs(2825) <= layer0_outputs(1425);
    outputs(2826) <= not((layer0_outputs(2332)) xor (layer0_outputs(4323)));
    outputs(2827) <= not((layer0_outputs(1365)) xor (layer0_outputs(2404)));
    outputs(2828) <= not(layer0_outputs(222));
    outputs(2829) <= layer0_outputs(593);
    outputs(2830) <= layer0_outputs(338);
    outputs(2831) <= (layer0_outputs(115)) and not (layer0_outputs(4053));
    outputs(2832) <= not((layer0_outputs(858)) xor (layer0_outputs(1917)));
    outputs(2833) <= (layer0_outputs(1527)) or (layer0_outputs(4294));
    outputs(2834) <= layer0_outputs(1178);
    outputs(2835) <= not(layer0_outputs(2902)) or (layer0_outputs(2618));
    outputs(2836) <= (layer0_outputs(4324)) and not (layer0_outputs(4775));
    outputs(2837) <= layer0_outputs(3767);
    outputs(2838) <= layer0_outputs(4581);
    outputs(2839) <= (layer0_outputs(2961)) xor (layer0_outputs(1907));
    outputs(2840) <= layer0_outputs(2183);
    outputs(2841) <= not((layer0_outputs(720)) or (layer0_outputs(3479)));
    outputs(2842) <= (layer0_outputs(2220)) or (layer0_outputs(5090));
    outputs(2843) <= not(layer0_outputs(5001));
    outputs(2844) <= not(layer0_outputs(2136));
    outputs(2845) <= (layer0_outputs(2198)) and (layer0_outputs(2490));
    outputs(2846) <= (layer0_outputs(2787)) xor (layer0_outputs(4967));
    outputs(2847) <= (layer0_outputs(2003)) and (layer0_outputs(3892));
    outputs(2848) <= not(layer0_outputs(2647));
    outputs(2849) <= not(layer0_outputs(4907));
    outputs(2850) <= (layer0_outputs(1747)) and (layer0_outputs(2624));
    outputs(2851) <= layer0_outputs(190);
    outputs(2852) <= not(layer0_outputs(2264)) or (layer0_outputs(3468));
    outputs(2853) <= layer0_outputs(5025);
    outputs(2854) <= layer0_outputs(1737);
    outputs(2855) <= not(layer0_outputs(1682));
    outputs(2856) <= not((layer0_outputs(1805)) and (layer0_outputs(2771)));
    outputs(2857) <= not(layer0_outputs(1304));
    outputs(2858) <= not(layer0_outputs(3093)) or (layer0_outputs(1921));
    outputs(2859) <= not(layer0_outputs(4110));
    outputs(2860) <= not((layer0_outputs(1440)) or (layer0_outputs(1423)));
    outputs(2861) <= not(layer0_outputs(3730));
    outputs(2862) <= not(layer0_outputs(4698));
    outputs(2863) <= not(layer0_outputs(2394));
    outputs(2864) <= not((layer0_outputs(3459)) and (layer0_outputs(4339)));
    outputs(2865) <= not(layer0_outputs(3493)) or (layer0_outputs(3308));
    outputs(2866) <= not((layer0_outputs(4146)) xor (layer0_outputs(3713)));
    outputs(2867) <= not(layer0_outputs(1285));
    outputs(2868) <= not(layer0_outputs(3455));
    outputs(2869) <= not((layer0_outputs(35)) xor (layer0_outputs(391)));
    outputs(2870) <= not(layer0_outputs(2365));
    outputs(2871) <= layer0_outputs(1523);
    outputs(2872) <= not(layer0_outputs(1305));
    outputs(2873) <= not(layer0_outputs(3824));
    outputs(2874) <= (layer0_outputs(3297)) and (layer0_outputs(5109));
    outputs(2875) <= not((layer0_outputs(850)) and (layer0_outputs(2828)));
    outputs(2876) <= layer0_outputs(3055);
    outputs(2877) <= (layer0_outputs(2668)) xor (layer0_outputs(3233));
    outputs(2878) <= not((layer0_outputs(984)) xor (layer0_outputs(2579)));
    outputs(2879) <= not((layer0_outputs(3713)) xor (layer0_outputs(7)));
    outputs(2880) <= layer0_outputs(1847);
    outputs(2881) <= layer0_outputs(1862);
    outputs(2882) <= not(layer0_outputs(969));
    outputs(2883) <= (layer0_outputs(2447)) or (layer0_outputs(1726));
    outputs(2884) <= (layer0_outputs(1675)) and (layer0_outputs(642));
    outputs(2885) <= (layer0_outputs(719)) or (layer0_outputs(3968));
    outputs(2886) <= layer0_outputs(2425);
    outputs(2887) <= not(layer0_outputs(3192)) or (layer0_outputs(1072));
    outputs(2888) <= not((layer0_outputs(982)) xor (layer0_outputs(5072)));
    outputs(2889) <= not(layer0_outputs(1424)) or (layer0_outputs(4118));
    outputs(2890) <= (layer0_outputs(5075)) xor (layer0_outputs(1074));
    outputs(2891) <= (layer0_outputs(2750)) and (layer0_outputs(3519));
    outputs(2892) <= not((layer0_outputs(2289)) xor (layer0_outputs(4104)));
    outputs(2893) <= not(layer0_outputs(4630)) or (layer0_outputs(4624));
    outputs(2894) <= not((layer0_outputs(1103)) xor (layer0_outputs(4461)));
    outputs(2895) <= not((layer0_outputs(4784)) xor (layer0_outputs(2301)));
    outputs(2896) <= not(layer0_outputs(2464));
    outputs(2897) <= not(layer0_outputs(1380));
    outputs(2898) <= not((layer0_outputs(1021)) or (layer0_outputs(10)));
    outputs(2899) <= not((layer0_outputs(2829)) xor (layer0_outputs(4090)));
    outputs(2900) <= not((layer0_outputs(365)) xor (layer0_outputs(2956)));
    outputs(2901) <= (layer0_outputs(810)) xor (layer0_outputs(307));
    outputs(2902) <= layer0_outputs(3743);
    outputs(2903) <= (layer0_outputs(2790)) and (layer0_outputs(3426));
    outputs(2904) <= layer0_outputs(4673);
    outputs(2905) <= not(layer0_outputs(3962));
    outputs(2906) <= layer0_outputs(2064);
    outputs(2907) <= layer0_outputs(2742);
    outputs(2908) <= (layer0_outputs(2979)) or (layer0_outputs(2963));
    outputs(2909) <= not(layer0_outputs(2646));
    outputs(2910) <= not((layer0_outputs(4003)) xor (layer0_outputs(783)));
    outputs(2911) <= (layer0_outputs(4888)) and (layer0_outputs(4041));
    outputs(2912) <= (layer0_outputs(3502)) and not (layer0_outputs(3662));
    outputs(2913) <= (layer0_outputs(163)) or (layer0_outputs(1470));
    outputs(2914) <= layer0_outputs(1150);
    outputs(2915) <= layer0_outputs(3706);
    outputs(2916) <= (layer0_outputs(477)) xor (layer0_outputs(2989));
    outputs(2917) <= not(layer0_outputs(3377)) or (layer0_outputs(2138));
    outputs(2918) <= not(layer0_outputs(2571));
    outputs(2919) <= (layer0_outputs(2489)) xor (layer0_outputs(668));
    outputs(2920) <= not(layer0_outputs(1400));
    outputs(2921) <= (layer0_outputs(3760)) xor (layer0_outputs(4904));
    outputs(2922) <= layer0_outputs(1236);
    outputs(2923) <= not((layer0_outputs(2327)) or (layer0_outputs(3420)));
    outputs(2924) <= (layer0_outputs(3219)) xor (layer0_outputs(2917));
    outputs(2925) <= not(layer0_outputs(4129));
    outputs(2926) <= not(layer0_outputs(4373));
    outputs(2927) <= (layer0_outputs(2441)) or (layer0_outputs(282));
    outputs(2928) <= layer0_outputs(129);
    outputs(2929) <= (layer0_outputs(2617)) xor (layer0_outputs(3553));
    outputs(2930) <= not((layer0_outputs(906)) and (layer0_outputs(1879)));
    outputs(2931) <= not(layer0_outputs(4880));
    outputs(2932) <= (layer0_outputs(1700)) and (layer0_outputs(1673));
    outputs(2933) <= not((layer0_outputs(3479)) or (layer0_outputs(2341)));
    outputs(2934) <= (layer0_outputs(5049)) and (layer0_outputs(3600));
    outputs(2935) <= layer0_outputs(3136);
    outputs(2936) <= (layer0_outputs(4132)) xor (layer0_outputs(2320));
    outputs(2937) <= not(layer0_outputs(3730));
    outputs(2938) <= (layer0_outputs(2998)) and not (layer0_outputs(3279));
    outputs(2939) <= not(layer0_outputs(1207));
    outputs(2940) <= not((layer0_outputs(933)) xor (layer0_outputs(1176)));
    outputs(2941) <= layer0_outputs(1249);
    outputs(2942) <= layer0_outputs(602);
    outputs(2943) <= not((layer0_outputs(2879)) xor (layer0_outputs(4485)));
    outputs(2944) <= (layer0_outputs(3867)) and not (layer0_outputs(2458));
    outputs(2945) <= (layer0_outputs(4306)) and (layer0_outputs(4751));
    outputs(2946) <= layer0_outputs(2560);
    outputs(2947) <= not(layer0_outputs(2060)) or (layer0_outputs(4338));
    outputs(2948) <= not((layer0_outputs(1247)) and (layer0_outputs(3850)));
    outputs(2949) <= (layer0_outputs(1527)) or (layer0_outputs(1227));
    outputs(2950) <= (layer0_outputs(4885)) and not (layer0_outputs(1305));
    outputs(2951) <= layer0_outputs(938);
    outputs(2952) <= not(layer0_outputs(5040));
    outputs(2953) <= not((layer0_outputs(2185)) or (layer0_outputs(2578)));
    outputs(2954) <= (layer0_outputs(2)) xor (layer0_outputs(3451));
    outputs(2955) <= not((layer0_outputs(2831)) xor (layer0_outputs(333)));
    outputs(2956) <= layer0_outputs(2024);
    outputs(2957) <= not(layer0_outputs(3244));
    outputs(2958) <= (layer0_outputs(2456)) and not (layer0_outputs(1391));
    outputs(2959) <= not((layer0_outputs(448)) xor (layer0_outputs(3759)));
    outputs(2960) <= not(layer0_outputs(3210)) or (layer0_outputs(2835));
    outputs(2961) <= not((layer0_outputs(1578)) and (layer0_outputs(2066)));
    outputs(2962) <= (layer0_outputs(1881)) xor (layer0_outputs(2987));
    outputs(2963) <= not((layer0_outputs(1366)) and (layer0_outputs(1907)));
    outputs(2964) <= (layer0_outputs(4041)) and not (layer0_outputs(2659));
    outputs(2965) <= (layer0_outputs(549)) or (layer0_outputs(4039));
    outputs(2966) <= (layer0_outputs(4386)) and (layer0_outputs(3379));
    outputs(2967) <= layer0_outputs(2724);
    outputs(2968) <= not(layer0_outputs(653));
    outputs(2969) <= layer0_outputs(1675);
    outputs(2970) <= layer0_outputs(3743);
    outputs(2971) <= not((layer0_outputs(3289)) or (layer0_outputs(3573)));
    outputs(2972) <= layer0_outputs(2923);
    outputs(2973) <= not(layer0_outputs(277));
    outputs(2974) <= (layer0_outputs(1763)) xor (layer0_outputs(820));
    outputs(2975) <= not(layer0_outputs(2761));
    outputs(2976) <= not(layer0_outputs(3486)) or (layer0_outputs(3851));
    outputs(2977) <= (layer0_outputs(1605)) or (layer0_outputs(1698));
    outputs(2978) <= not((layer0_outputs(4301)) xor (layer0_outputs(2914)));
    outputs(2979) <= not(layer0_outputs(345));
    outputs(2980) <= layer0_outputs(4636);
    outputs(2981) <= (layer0_outputs(4235)) or (layer0_outputs(4246));
    outputs(2982) <= not((layer0_outputs(1280)) or (layer0_outputs(4166)));
    outputs(2983) <= not(layer0_outputs(407));
    outputs(2984) <= layer0_outputs(2233);
    outputs(2985) <= (layer0_outputs(525)) xor (layer0_outputs(1149));
    outputs(2986) <= (layer0_outputs(3822)) and not (layer0_outputs(262));
    outputs(2987) <= (layer0_outputs(780)) xor (layer0_outputs(5084));
    outputs(2988) <= (layer0_outputs(144)) and (layer0_outputs(3190));
    outputs(2989) <= (layer0_outputs(5046)) xor (layer0_outputs(1113));
    outputs(2990) <= not((layer0_outputs(2289)) xor (layer0_outputs(757)));
    outputs(2991) <= not(layer0_outputs(3995));
    outputs(2992) <= not((layer0_outputs(2255)) or (layer0_outputs(2538)));
    outputs(2993) <= layer0_outputs(936);
    outputs(2994) <= (layer0_outputs(3614)) and not (layer0_outputs(3463));
    outputs(2995) <= layer0_outputs(1491);
    outputs(2996) <= layer0_outputs(1121);
    outputs(2997) <= not((layer0_outputs(101)) and (layer0_outputs(708)));
    outputs(2998) <= not(layer0_outputs(392));
    outputs(2999) <= not(layer0_outputs(2017)) or (layer0_outputs(1586));
    outputs(3000) <= not(layer0_outputs(4194));
    outputs(3001) <= (layer0_outputs(2325)) or (layer0_outputs(3020));
    outputs(3002) <= (layer0_outputs(1936)) and (layer0_outputs(3293));
    outputs(3003) <= layer0_outputs(1782);
    outputs(3004) <= layer0_outputs(2852);
    outputs(3005) <= layer0_outputs(1938);
    outputs(3006) <= (layer0_outputs(4583)) and (layer0_outputs(821));
    outputs(3007) <= not(layer0_outputs(3510));
    outputs(3008) <= not(layer0_outputs(1485));
    outputs(3009) <= not((layer0_outputs(2228)) xor (layer0_outputs(4697)));
    outputs(3010) <= (layer0_outputs(1992)) and not (layer0_outputs(1690));
    outputs(3011) <= (layer0_outputs(1762)) xor (layer0_outputs(5019));
    outputs(3012) <= not((layer0_outputs(4361)) or (layer0_outputs(529)));
    outputs(3013) <= (layer0_outputs(2357)) and not (layer0_outputs(758));
    outputs(3014) <= not((layer0_outputs(443)) xor (layer0_outputs(2863)));
    outputs(3015) <= (layer0_outputs(3815)) xor (layer0_outputs(59));
    outputs(3016) <= (layer0_outputs(232)) xor (layer0_outputs(1142));
    outputs(3017) <= not(layer0_outputs(444));
    outputs(3018) <= (layer0_outputs(1069)) xor (layer0_outputs(1680));
    outputs(3019) <= not(layer0_outputs(4130)) or (layer0_outputs(3795));
    outputs(3020) <= not(layer0_outputs(2707));
    outputs(3021) <= not((layer0_outputs(1758)) or (layer0_outputs(1626)));
    outputs(3022) <= layer0_outputs(1287);
    outputs(3023) <= not(layer0_outputs(4559)) or (layer0_outputs(4657));
    outputs(3024) <= not(layer0_outputs(1514)) or (layer0_outputs(4547));
    outputs(3025) <= (layer0_outputs(4631)) xor (layer0_outputs(987));
    outputs(3026) <= layer0_outputs(849);
    outputs(3027) <= not(layer0_outputs(3203));
    outputs(3028) <= layer0_outputs(4344);
    outputs(3029) <= (layer0_outputs(4264)) and (layer0_outputs(582));
    outputs(3030) <= not((layer0_outputs(410)) xor (layer0_outputs(3925)));
    outputs(3031) <= (layer0_outputs(4048)) or (layer0_outputs(3640));
    outputs(3032) <= not(layer0_outputs(820));
    outputs(3033) <= layer0_outputs(4278);
    outputs(3034) <= not(layer0_outputs(2971));
    outputs(3035) <= layer0_outputs(1915);
    outputs(3036) <= (layer0_outputs(4902)) xor (layer0_outputs(3603));
    outputs(3037) <= not(layer0_outputs(4768));
    outputs(3038) <= not((layer0_outputs(1980)) or (layer0_outputs(844)));
    outputs(3039) <= (layer0_outputs(4522)) and not (layer0_outputs(2381));
    outputs(3040) <= not(layer0_outputs(4138));
    outputs(3041) <= layer0_outputs(1219);
    outputs(3042) <= (layer0_outputs(2835)) and (layer0_outputs(226));
    outputs(3043) <= not((layer0_outputs(623)) xor (layer0_outputs(1822)));
    outputs(3044) <= (layer0_outputs(1817)) and (layer0_outputs(3521));
    outputs(3045) <= not(layer0_outputs(2347));
    outputs(3046) <= (layer0_outputs(4017)) and not (layer0_outputs(3639));
    outputs(3047) <= not(layer0_outputs(4723));
    outputs(3048) <= not((layer0_outputs(251)) xor (layer0_outputs(3865)));
    outputs(3049) <= (layer0_outputs(3141)) and not (layer0_outputs(4727));
    outputs(3050) <= not(layer0_outputs(3637));
    outputs(3051) <= not((layer0_outputs(1836)) and (layer0_outputs(837)));
    outputs(3052) <= layer0_outputs(386);
    outputs(3053) <= layer0_outputs(796);
    outputs(3054) <= not((layer0_outputs(4178)) xor (layer0_outputs(531)));
    outputs(3055) <= (layer0_outputs(658)) and (layer0_outputs(2702));
    outputs(3056) <= not(layer0_outputs(4055)) or (layer0_outputs(4154));
    outputs(3057) <= layer0_outputs(2309);
    outputs(3058) <= layer0_outputs(2309);
    outputs(3059) <= not(layer0_outputs(4381));
    outputs(3060) <= not((layer0_outputs(699)) and (layer0_outputs(2630)));
    outputs(3061) <= not(layer0_outputs(1731));
    outputs(3062) <= not(layer0_outputs(2107));
    outputs(3063) <= not((layer0_outputs(164)) or (layer0_outputs(4358)));
    outputs(3064) <= not((layer0_outputs(3072)) or (layer0_outputs(186)));
    outputs(3065) <= not((layer0_outputs(1313)) or (layer0_outputs(1682)));
    outputs(3066) <= (layer0_outputs(1979)) xor (layer0_outputs(1354));
    outputs(3067) <= layer0_outputs(3186);
    outputs(3068) <= not(layer0_outputs(4404));
    outputs(3069) <= (layer0_outputs(1449)) and not (layer0_outputs(706));
    outputs(3070) <= (layer0_outputs(2262)) or (layer0_outputs(989));
    outputs(3071) <= not(layer0_outputs(4282));
    outputs(3072) <= layer0_outputs(1079);
    outputs(3073) <= layer0_outputs(83);
    outputs(3074) <= not(layer0_outputs(4461));
    outputs(3075) <= layer0_outputs(3370);
    outputs(3076) <= not(layer0_outputs(3870));
    outputs(3077) <= (layer0_outputs(1011)) and (layer0_outputs(633));
    outputs(3078) <= layer0_outputs(3421);
    outputs(3079) <= (layer0_outputs(4993)) and (layer0_outputs(4541));
    outputs(3080) <= not((layer0_outputs(1768)) or (layer0_outputs(963)));
    outputs(3081) <= (layer0_outputs(4561)) and not (layer0_outputs(4195));
    outputs(3082) <= not(layer0_outputs(1850));
    outputs(3083) <= layer0_outputs(3977);
    outputs(3084) <= (layer0_outputs(4444)) or (layer0_outputs(722));
    outputs(3085) <= layer0_outputs(4202);
    outputs(3086) <= layer0_outputs(1243);
    outputs(3087) <= layer0_outputs(4072);
    outputs(3088) <= not(layer0_outputs(577));
    outputs(3089) <= not(layer0_outputs(1717));
    outputs(3090) <= (layer0_outputs(714)) and not (layer0_outputs(3389));
    outputs(3091) <= not((layer0_outputs(2655)) or (layer0_outputs(3313)));
    outputs(3092) <= not((layer0_outputs(343)) xor (layer0_outputs(389)));
    outputs(3093) <= (layer0_outputs(3999)) and not (layer0_outputs(1948));
    outputs(3094) <= not(layer0_outputs(4046));
    outputs(3095) <= not(layer0_outputs(3609));
    outputs(3096) <= not(layer0_outputs(1151));
    outputs(3097) <= (layer0_outputs(3265)) and not (layer0_outputs(4746));
    outputs(3098) <= (layer0_outputs(2147)) and not (layer0_outputs(4644));
    outputs(3099) <= layer0_outputs(4691);
    outputs(3100) <= not(layer0_outputs(2962));
    outputs(3101) <= not(layer0_outputs(3520));
    outputs(3102) <= not(layer0_outputs(2876)) or (layer0_outputs(579));
    outputs(3103) <= not(layer0_outputs(4622));
    outputs(3104) <= layer0_outputs(4290);
    outputs(3105) <= layer0_outputs(5034);
    outputs(3106) <= (layer0_outputs(71)) and (layer0_outputs(1952));
    outputs(3107) <= not(layer0_outputs(4197)) or (layer0_outputs(1115));
    outputs(3108) <= not((layer0_outputs(1330)) xor (layer0_outputs(3596)));
    outputs(3109) <= (layer0_outputs(851)) or (layer0_outputs(3577));
    outputs(3110) <= layer0_outputs(4044);
    outputs(3111) <= not(layer0_outputs(2367));
    outputs(3112) <= not(layer0_outputs(4859));
    outputs(3113) <= not((layer0_outputs(1887)) or (layer0_outputs(1543)));
    outputs(3114) <= not(layer0_outputs(3463));
    outputs(3115) <= not(layer0_outputs(2920));
    outputs(3116) <= layer0_outputs(3029);
    outputs(3117) <= not((layer0_outputs(3563)) or (layer0_outputs(2928)));
    outputs(3118) <= not(layer0_outputs(1972));
    outputs(3119) <= (layer0_outputs(2186)) and not (layer0_outputs(4744));
    outputs(3120) <= (layer0_outputs(2603)) and (layer0_outputs(2147));
    outputs(3121) <= (layer0_outputs(4521)) and not (layer0_outputs(4873));
    outputs(3122) <= (layer0_outputs(1642)) and not (layer0_outputs(589));
    outputs(3123) <= not(layer0_outputs(897));
    outputs(3124) <= (layer0_outputs(1317)) and not (layer0_outputs(750));
    outputs(3125) <= not(layer0_outputs(3409));
    outputs(3126) <= not(layer0_outputs(1883));
    outputs(3127) <= (layer0_outputs(4718)) and not (layer0_outputs(1240));
    outputs(3128) <= not(layer0_outputs(3255));
    outputs(3129) <= layer0_outputs(4366);
    outputs(3130) <= not(layer0_outputs(222));
    outputs(3131) <= layer0_outputs(1756);
    outputs(3132) <= (layer0_outputs(76)) and not (layer0_outputs(2890));
    outputs(3133) <= not(layer0_outputs(2623));
    outputs(3134) <= (layer0_outputs(3138)) xor (layer0_outputs(3972));
    outputs(3135) <= layer0_outputs(4583);
    outputs(3136) <= layer0_outputs(3791);
    outputs(3137) <= (layer0_outputs(3194)) and (layer0_outputs(4619));
    outputs(3138) <= (layer0_outputs(693)) and (layer0_outputs(1290));
    outputs(3139) <= (layer0_outputs(2689)) xor (layer0_outputs(3957));
    outputs(3140) <= not(layer0_outputs(231)) or (layer0_outputs(4285));
    outputs(3141) <= not((layer0_outputs(2968)) or (layer0_outputs(3342)));
    outputs(3142) <= not(layer0_outputs(5078));
    outputs(3143) <= layer0_outputs(4452);
    outputs(3144) <= not((layer0_outputs(1015)) xor (layer0_outputs(4293)));
    outputs(3145) <= not((layer0_outputs(1848)) and (layer0_outputs(316)));
    outputs(3146) <= (layer0_outputs(3246)) and (layer0_outputs(4015));
    outputs(3147) <= layer0_outputs(4769);
    outputs(3148) <= (layer0_outputs(1651)) and not (layer0_outputs(4496));
    outputs(3149) <= layer0_outputs(5070);
    outputs(3150) <= not(layer0_outputs(946)) or (layer0_outputs(2929));
    outputs(3151) <= not(layer0_outputs(1001));
    outputs(3152) <= (layer0_outputs(976)) and not (layer0_outputs(5078));
    outputs(3153) <= layer0_outputs(3008);
    outputs(3154) <= not(layer0_outputs(159));
    outputs(3155) <= not((layer0_outputs(1615)) xor (layer0_outputs(525)));
    outputs(3156) <= layer0_outputs(1483);
    outputs(3157) <= not(layer0_outputs(214));
    outputs(3158) <= layer0_outputs(4487);
    outputs(3159) <= not(layer0_outputs(3290));
    outputs(3160) <= (layer0_outputs(4813)) and not (layer0_outputs(2428));
    outputs(3161) <= (layer0_outputs(831)) and not (layer0_outputs(260));
    outputs(3162) <= layer0_outputs(1410);
    outputs(3163) <= (layer0_outputs(1545)) and not (layer0_outputs(443));
    outputs(3164) <= not(layer0_outputs(5029)) or (layer0_outputs(1696));
    outputs(3165) <= (layer0_outputs(2115)) and not (layer0_outputs(2658));
    outputs(3166) <= layer0_outputs(3678);
    outputs(3167) <= layer0_outputs(1933);
    outputs(3168) <= layer0_outputs(2018);
    outputs(3169) <= (layer0_outputs(4832)) and not (layer0_outputs(3564));
    outputs(3170) <= (layer0_outputs(520)) and (layer0_outputs(2111));
    outputs(3171) <= layer0_outputs(972);
    outputs(3172) <= not(layer0_outputs(4954));
    outputs(3173) <= layer0_outputs(720);
    outputs(3174) <= (layer0_outputs(4423)) and not (layer0_outputs(3904));
    outputs(3175) <= layer0_outputs(3195);
    outputs(3176) <= not(layer0_outputs(2373)) or (layer0_outputs(1168));
    outputs(3177) <= not(layer0_outputs(621));
    outputs(3178) <= (layer0_outputs(2522)) and not (layer0_outputs(1214));
    outputs(3179) <= layer0_outputs(2121);
    outputs(3180) <= (layer0_outputs(4869)) and not (layer0_outputs(1379));
    outputs(3181) <= not((layer0_outputs(1018)) or (layer0_outputs(5091)));
    outputs(3182) <= layer0_outputs(3302);
    outputs(3183) <= (layer0_outputs(567)) and (layer0_outputs(3169));
    outputs(3184) <= layer0_outputs(4326);
    outputs(3185) <= (layer0_outputs(1591)) and not (layer0_outputs(3881));
    outputs(3186) <= (layer0_outputs(4949)) and not (layer0_outputs(1312));
    outputs(3187) <= (layer0_outputs(1531)) xor (layer0_outputs(3042));
    outputs(3188) <= (layer0_outputs(1109)) and not (layer0_outputs(2675));
    outputs(3189) <= layer0_outputs(1826);
    outputs(3190) <= (layer0_outputs(1620)) and not (layer0_outputs(731));
    outputs(3191) <= not((layer0_outputs(3978)) or (layer0_outputs(3158)));
    outputs(3192) <= (layer0_outputs(1158)) and (layer0_outputs(4381));
    outputs(3193) <= (layer0_outputs(3737)) or (layer0_outputs(3159));
    outputs(3194) <= not(layer0_outputs(4717));
    outputs(3195) <= not(layer0_outputs(1436));
    outputs(3196) <= (layer0_outputs(3603)) or (layer0_outputs(5017));
    outputs(3197) <= layer0_outputs(802);
    outputs(3198) <= layer0_outputs(925);
    outputs(3199) <= not(layer0_outputs(4230));
    outputs(3200) <= (layer0_outputs(2560)) and (layer0_outputs(4885));
    outputs(3201) <= not((layer0_outputs(1157)) and (layer0_outputs(3105)));
    outputs(3202) <= not((layer0_outputs(930)) xor (layer0_outputs(4268)));
    outputs(3203) <= (layer0_outputs(3416)) xor (layer0_outputs(1554));
    outputs(3204) <= not((layer0_outputs(805)) or (layer0_outputs(1904)));
    outputs(3205) <= (layer0_outputs(1529)) and (layer0_outputs(3884));
    outputs(3206) <= layer0_outputs(188);
    outputs(3207) <= not((layer0_outputs(1068)) or (layer0_outputs(3087)));
    outputs(3208) <= not((layer0_outputs(4544)) or (layer0_outputs(1927)));
    outputs(3209) <= (layer0_outputs(625)) and (layer0_outputs(2336));
    outputs(3210) <= (layer0_outputs(37)) and not (layer0_outputs(3226));
    outputs(3211) <= not(layer0_outputs(4153));
    outputs(3212) <= (layer0_outputs(4087)) or (layer0_outputs(1122));
    outputs(3213) <= layer0_outputs(3683);
    outputs(3214) <= not(layer0_outputs(3505));
    outputs(3215) <= (layer0_outputs(4251)) and (layer0_outputs(4734));
    outputs(3216) <= (layer0_outputs(4368)) and not (layer0_outputs(4039));
    outputs(3217) <= (layer0_outputs(4898)) xor (layer0_outputs(171));
    outputs(3218) <= (layer0_outputs(3492)) and (layer0_outputs(122));
    outputs(3219) <= (layer0_outputs(472)) and (layer0_outputs(4704));
    outputs(3220) <= layer0_outputs(1477);
    outputs(3221) <= not(layer0_outputs(1186));
    outputs(3222) <= (layer0_outputs(60)) and not (layer0_outputs(4722));
    outputs(3223) <= (layer0_outputs(2698)) and not (layer0_outputs(4484));
    outputs(3224) <= layer0_outputs(4308);
    outputs(3225) <= (layer0_outputs(2163)) and (layer0_outputs(3839));
    outputs(3226) <= layer0_outputs(3938);
    outputs(3227) <= not((layer0_outputs(323)) or (layer0_outputs(3626)));
    outputs(3228) <= (layer0_outputs(2469)) xor (layer0_outputs(3761));
    outputs(3229) <= (layer0_outputs(2310)) and not (layer0_outputs(3802));
    outputs(3230) <= (layer0_outputs(4172)) and not (layer0_outputs(1789));
    outputs(3231) <= not((layer0_outputs(1347)) xor (layer0_outputs(1147)));
    outputs(3232) <= (layer0_outputs(3132)) and not (layer0_outputs(2495));
    outputs(3233) <= not((layer0_outputs(1692)) xor (layer0_outputs(600)));
    outputs(3234) <= layer0_outputs(1096);
    outputs(3235) <= layer0_outputs(2466);
    outputs(3236) <= (layer0_outputs(3474)) and (layer0_outputs(208));
    outputs(3237) <= not(layer0_outputs(4248)) or (layer0_outputs(4971));
    outputs(3238) <= not(layer0_outputs(1279));
    outputs(3239) <= not(layer0_outputs(2747));
    outputs(3240) <= not(layer0_outputs(258));
    outputs(3241) <= layer0_outputs(196);
    outputs(3242) <= layer0_outputs(976);
    outputs(3243) <= not((layer0_outputs(1508)) and (layer0_outputs(1506)));
    outputs(3244) <= (layer0_outputs(791)) and (layer0_outputs(1374));
    outputs(3245) <= not(layer0_outputs(3103));
    outputs(3246) <= (layer0_outputs(5067)) xor (layer0_outputs(3696));
    outputs(3247) <= layer0_outputs(3926);
    outputs(3248) <= not((layer0_outputs(2890)) or (layer0_outputs(1216)));
    outputs(3249) <= not((layer0_outputs(1036)) or (layer0_outputs(3563)));
    outputs(3250) <= layer0_outputs(1454);
    outputs(3251) <= not(layer0_outputs(958));
    outputs(3252) <= not(layer0_outputs(898));
    outputs(3253) <= layer0_outputs(1900);
    outputs(3254) <= (layer0_outputs(2085)) or (layer0_outputs(1289));
    outputs(3255) <= not(layer0_outputs(2424));
    outputs(3256) <= layer0_outputs(2462);
    outputs(3257) <= (layer0_outputs(1784)) xor (layer0_outputs(2452));
    outputs(3258) <= not(layer0_outputs(1050));
    outputs(3259) <= layer0_outputs(1658);
    outputs(3260) <= not(layer0_outputs(2526));
    outputs(3261) <= not(layer0_outputs(2882)) or (layer0_outputs(4171));
    outputs(3262) <= not(layer0_outputs(4163)) or (layer0_outputs(2426));
    outputs(3263) <= (layer0_outputs(2477)) or (layer0_outputs(1012));
    outputs(3264) <= not(layer0_outputs(886)) or (layer0_outputs(4335));
    outputs(3265) <= not((layer0_outputs(3395)) xor (layer0_outputs(903)));
    outputs(3266) <= not((layer0_outputs(2846)) or (layer0_outputs(3083)));
    outputs(3267) <= (layer0_outputs(3577)) and not (layer0_outputs(4369));
    outputs(3268) <= not(layer0_outputs(2731));
    outputs(3269) <= (layer0_outputs(3097)) or (layer0_outputs(1327));
    outputs(3270) <= layer0_outputs(3015);
    outputs(3271) <= layer0_outputs(4953);
    outputs(3272) <= not(layer0_outputs(3686)) or (layer0_outputs(3283));
    outputs(3273) <= not((layer0_outputs(1441)) or (layer0_outputs(1360)));
    outputs(3274) <= not(layer0_outputs(5029));
    outputs(3275) <= not(layer0_outputs(1824));
    outputs(3276) <= layer0_outputs(2692);
    outputs(3277) <= not((layer0_outputs(3457)) xor (layer0_outputs(4905)));
    outputs(3278) <= (layer0_outputs(3372)) and not (layer0_outputs(3855));
    outputs(3279) <= not(layer0_outputs(3230));
    outputs(3280) <= not(layer0_outputs(3742));
    outputs(3281) <= not(layer0_outputs(1191));
    outputs(3282) <= layer0_outputs(3622);
    outputs(3283) <= not(layer0_outputs(4016));
    outputs(3284) <= not(layer0_outputs(2545));
    outputs(3285) <= not(layer0_outputs(1695));
    outputs(3286) <= layer0_outputs(2113);
    outputs(3287) <= not((layer0_outputs(465)) or (layer0_outputs(4610)));
    outputs(3288) <= layer0_outputs(3493);
    outputs(3289) <= (layer0_outputs(4754)) or (layer0_outputs(3901));
    outputs(3290) <= layer0_outputs(1361);
    outputs(3291) <= not(layer0_outputs(3930));
    outputs(3292) <= (layer0_outputs(2288)) and (layer0_outputs(5076));
    outputs(3293) <= not(layer0_outputs(854));
    outputs(3294) <= not((layer0_outputs(2036)) or (layer0_outputs(1194)));
    outputs(3295) <= not(layer0_outputs(1599));
    outputs(3296) <= not(layer0_outputs(3698));
    outputs(3297) <= not(layer0_outputs(3962)) or (layer0_outputs(1621));
    outputs(3298) <= (layer0_outputs(2755)) and not (layer0_outputs(3731));
    outputs(3299) <= not(layer0_outputs(1630));
    outputs(3300) <= not((layer0_outputs(1445)) or (layer0_outputs(2893)));
    outputs(3301) <= (layer0_outputs(1607)) and not (layer0_outputs(2823));
    outputs(3302) <= (layer0_outputs(724)) and not (layer0_outputs(3271));
    outputs(3303) <= (layer0_outputs(2728)) and not (layer0_outputs(4940));
    outputs(3304) <= (layer0_outputs(5103)) and not (layer0_outputs(1496));
    outputs(3305) <= not(layer0_outputs(3494)) or (layer0_outputs(1349));
    outputs(3306) <= layer0_outputs(1225);
    outputs(3307) <= layer0_outputs(335);
    outputs(3308) <= not((layer0_outputs(1422)) and (layer0_outputs(3498)));
    outputs(3309) <= layer0_outputs(3081);
    outputs(3310) <= (layer0_outputs(3081)) and (layer0_outputs(1667));
    outputs(3311) <= not((layer0_outputs(1494)) or (layer0_outputs(2393)));
    outputs(3312) <= not(layer0_outputs(2885));
    outputs(3313) <= not(layer0_outputs(1792));
    outputs(3314) <= not(layer0_outputs(1791));
    outputs(3315) <= (layer0_outputs(2683)) xor (layer0_outputs(3559));
    outputs(3316) <= layer0_outputs(3651);
    outputs(3317) <= not((layer0_outputs(3582)) or (layer0_outputs(2160)));
    outputs(3318) <= (layer0_outputs(3907)) and (layer0_outputs(2907));
    outputs(3319) <= not(layer0_outputs(4460)) or (layer0_outputs(3002));
    outputs(3320) <= (layer0_outputs(1060)) xor (layer0_outputs(4987));
    outputs(3321) <= (layer0_outputs(4024)) and (layer0_outputs(4086));
    outputs(3322) <= (layer0_outputs(933)) and not (layer0_outputs(1528));
    outputs(3323) <= not((layer0_outputs(40)) xor (layer0_outputs(3478)));
    outputs(3324) <= not(layer0_outputs(1628)) or (layer0_outputs(1893));
    outputs(3325) <= (layer0_outputs(4685)) and (layer0_outputs(4619));
    outputs(3326) <= (layer0_outputs(2056)) and not (layer0_outputs(1486));
    outputs(3327) <= (layer0_outputs(3458)) and not (layer0_outputs(954));
    outputs(3328) <= (layer0_outputs(3559)) and not (layer0_outputs(4400));
    outputs(3329) <= (layer0_outputs(3595)) and not (layer0_outputs(2371));
    outputs(3330) <= not((layer0_outputs(347)) xor (layer0_outputs(2952)));
    outputs(3331) <= (layer0_outputs(556)) and not (layer0_outputs(1897));
    outputs(3332) <= (layer0_outputs(2364)) and not (layer0_outputs(1406));
    outputs(3333) <= (layer0_outputs(4008)) and not (layer0_outputs(3634));
    outputs(3334) <= layer0_outputs(1802);
    outputs(3335) <= (layer0_outputs(3546)) and not (layer0_outputs(1332));
    outputs(3336) <= not(layer0_outputs(467));
    outputs(3337) <= not(layer0_outputs(1353)) or (layer0_outputs(1970));
    outputs(3338) <= not((layer0_outputs(415)) xor (layer0_outputs(4052)));
    outputs(3339) <= layer0_outputs(4294);
    outputs(3340) <= not((layer0_outputs(1118)) xor (layer0_outputs(4313)));
    outputs(3341) <= (layer0_outputs(3570)) and not (layer0_outputs(4005));
    outputs(3342) <= (layer0_outputs(2990)) and not (layer0_outputs(4134));
    outputs(3343) <= layer0_outputs(4304);
    outputs(3344) <= layer0_outputs(2349);
    outputs(3345) <= layer0_outputs(4033);
    outputs(3346) <= layer0_outputs(2506);
    outputs(3347) <= (layer0_outputs(3058)) and not (layer0_outputs(3583));
    outputs(3348) <= not(layer0_outputs(2863));
    outputs(3349) <= not(layer0_outputs(49));
    outputs(3350) <= not(layer0_outputs(2095));
    outputs(3351) <= not(layer0_outputs(4182));
    outputs(3352) <= not(layer0_outputs(2443)) or (layer0_outputs(2329));
    outputs(3353) <= (layer0_outputs(3721)) and not (layer0_outputs(2704));
    outputs(3354) <= (layer0_outputs(1433)) and (layer0_outputs(1025));
    outputs(3355) <= layer0_outputs(3539);
    outputs(3356) <= layer0_outputs(4121);
    outputs(3357) <= (layer0_outputs(3810)) and not (layer0_outputs(2069));
    outputs(3358) <= layer0_outputs(2188);
    outputs(3359) <= (layer0_outputs(4291)) and (layer0_outputs(309));
    outputs(3360) <= not((layer0_outputs(3854)) or (layer0_outputs(3833)));
    outputs(3361) <= layer0_outputs(4632);
    outputs(3362) <= layer0_outputs(3429);
    outputs(3363) <= layer0_outputs(4668);
    outputs(3364) <= not((layer0_outputs(2957)) and (layer0_outputs(62)));
    outputs(3365) <= not(layer0_outputs(3349));
    outputs(3366) <= not(layer0_outputs(731));
    outputs(3367) <= layer0_outputs(4511);
    outputs(3368) <= not((layer0_outputs(3301)) or (layer0_outputs(2766)));
    outputs(3369) <= not((layer0_outputs(1051)) xor (layer0_outputs(2602)));
    outputs(3370) <= (layer0_outputs(1242)) and (layer0_outputs(2569));
    outputs(3371) <= not(layer0_outputs(4828));
    outputs(3372) <= layer0_outputs(3650);
    outputs(3373) <= not(layer0_outputs(3932));
    outputs(3374) <= not(layer0_outputs(545));
    outputs(3375) <= (layer0_outputs(5106)) xor (layer0_outputs(1812));
    outputs(3376) <= (layer0_outputs(2588)) and (layer0_outputs(39));
    outputs(3377) <= (layer0_outputs(2068)) xor (layer0_outputs(3929));
    outputs(3378) <= layer0_outputs(701);
    outputs(3379) <= (layer0_outputs(3869)) xor (layer0_outputs(905));
    outputs(3380) <= not(layer0_outputs(4301));
    outputs(3381) <= (layer0_outputs(2723)) and not (layer0_outputs(2774));
    outputs(3382) <= not(layer0_outputs(62)) or (layer0_outputs(3385));
    outputs(3383) <= not((layer0_outputs(1372)) or (layer0_outputs(1355)));
    outputs(3384) <= (layer0_outputs(3611)) and not (layer0_outputs(887));
    outputs(3385) <= not(layer0_outputs(4591)) or (layer0_outputs(2065));
    outputs(3386) <= (layer0_outputs(3485)) and not (layer0_outputs(3061));
    outputs(3387) <= (layer0_outputs(4047)) and (layer0_outputs(4050));
    outputs(3388) <= not((layer0_outputs(4204)) and (layer0_outputs(847)));
    outputs(3389) <= layer0_outputs(331);
    outputs(3390) <= not(layer0_outputs(1874));
    outputs(3391) <= (layer0_outputs(2953)) and not (layer0_outputs(1160));
    outputs(3392) <= (layer0_outputs(418)) and not (layer0_outputs(853));
    outputs(3393) <= layer0_outputs(2206);
    outputs(3394) <= (layer0_outputs(4290)) xor (layer0_outputs(5112));
    outputs(3395) <= not(layer0_outputs(1236));
    outputs(3396) <= not(layer0_outputs(70));
    outputs(3397) <= (layer0_outputs(974)) xor (layer0_outputs(215));
    outputs(3398) <= not(layer0_outputs(3910));
    outputs(3399) <= not(layer0_outputs(3838));
    outputs(3400) <= not(layer0_outputs(913));
    outputs(3401) <= layer0_outputs(3114);
    outputs(3402) <= not((layer0_outputs(3117)) xor (layer0_outputs(624)));
    outputs(3403) <= (layer0_outputs(5068)) and not (layer0_outputs(3912));
    outputs(3404) <= layer0_outputs(5055);
    outputs(3405) <= layer0_outputs(4677);
    outputs(3406) <= layer0_outputs(763);
    outputs(3407) <= not(layer0_outputs(4648));
    outputs(3408) <= not(layer0_outputs(1417));
    outputs(3409) <= layer0_outputs(2389);
    outputs(3410) <= (layer0_outputs(1073)) and (layer0_outputs(3365));
    outputs(3411) <= (layer0_outputs(4963)) and not (layer0_outputs(1208));
    outputs(3412) <= layer0_outputs(52);
    outputs(3413) <= not(layer0_outputs(3438));
    outputs(3414) <= not((layer0_outputs(2693)) or (layer0_outputs(4085)));
    outputs(3415) <= not(layer0_outputs(832)) or (layer0_outputs(1800));
    outputs(3416) <= (layer0_outputs(191)) and not (layer0_outputs(2846));
    outputs(3417) <= (layer0_outputs(825)) xor (layer0_outputs(3435));
    outputs(3418) <= (layer0_outputs(2960)) and (layer0_outputs(4956));
    outputs(3419) <= (layer0_outputs(2343)) and not (layer0_outputs(3306));
    outputs(3420) <= not(layer0_outputs(3759));
    outputs(3421) <= (layer0_outputs(4237)) and not (layer0_outputs(1859));
    outputs(3422) <= not((layer0_outputs(2536)) or (layer0_outputs(118)));
    outputs(3423) <= not((layer0_outputs(4892)) or (layer0_outputs(1103)));
    outputs(3424) <= (layer0_outputs(114)) and not (layer0_outputs(2142));
    outputs(3425) <= layer0_outputs(4713);
    outputs(3426) <= not(layer0_outputs(2416));
    outputs(3427) <= (layer0_outputs(3047)) or (layer0_outputs(1408));
    outputs(3428) <= not(layer0_outputs(1908));
    outputs(3429) <= not(layer0_outputs(1388));
    outputs(3430) <= (layer0_outputs(3720)) and (layer0_outputs(1339));
    outputs(3431) <= (layer0_outputs(4152)) and not (layer0_outputs(1131));
    outputs(3432) <= not(layer0_outputs(1924));
    outputs(3433) <= not(layer0_outputs(3540));
    outputs(3434) <= (layer0_outputs(1031)) and (layer0_outputs(718));
    outputs(3435) <= (layer0_outputs(1678)) xor (layer0_outputs(2520));
    outputs(3436) <= not(layer0_outputs(4214));
    outputs(3437) <= (layer0_outputs(730)) or (layer0_outputs(3543));
    outputs(3438) <= not(layer0_outputs(4598));
    outputs(3439) <= (layer0_outputs(2081)) or (layer0_outputs(5071));
    outputs(3440) <= not(layer0_outputs(3495));
    outputs(3441) <= layer0_outputs(2918);
    outputs(3442) <= layer0_outputs(1241);
    outputs(3443) <= layer0_outputs(4769);
    outputs(3444) <= not(layer0_outputs(2808));
    outputs(3445) <= not(layer0_outputs(3088));
    outputs(3446) <= (layer0_outputs(1598)) or (layer0_outputs(2218));
    outputs(3447) <= not(layer0_outputs(97));
    outputs(3448) <= (layer0_outputs(2049)) and not (layer0_outputs(140));
    outputs(3449) <= not(layer0_outputs(3727));
    outputs(3450) <= layer0_outputs(4088);
    outputs(3451) <= not(layer0_outputs(372));
    outputs(3452) <= (layer0_outputs(1579)) and (layer0_outputs(3305));
    outputs(3453) <= not((layer0_outputs(3591)) xor (layer0_outputs(3338)));
    outputs(3454) <= (layer0_outputs(766)) xor (layer0_outputs(2151));
    outputs(3455) <= not((layer0_outputs(1828)) or (layer0_outputs(3005)));
    outputs(3456) <= layer0_outputs(851);
    outputs(3457) <= not((layer0_outputs(137)) xor (layer0_outputs(2053)));
    outputs(3458) <= not(layer0_outputs(3000));
    outputs(3459) <= not(layer0_outputs(2059));
    outputs(3460) <= (layer0_outputs(2580)) xor (layer0_outputs(4320));
    outputs(3461) <= (layer0_outputs(4712)) and not (layer0_outputs(4328));
    outputs(3462) <= layer0_outputs(1226);
    outputs(3463) <= (layer0_outputs(4113)) or (layer0_outputs(3968));
    outputs(3464) <= not(layer0_outputs(2335));
    outputs(3465) <= (layer0_outputs(2259)) and not (layer0_outputs(1840));
    outputs(3466) <= layer0_outputs(2974);
    outputs(3467) <= layer0_outputs(3325);
    outputs(3468) <= not(layer0_outputs(1350));
    outputs(3469) <= (layer0_outputs(1320)) xor (layer0_outputs(3547));
    outputs(3470) <= not(layer0_outputs(1923));
    outputs(3471) <= (layer0_outputs(1290)) xor (layer0_outputs(3664));
    outputs(3472) <= not(layer0_outputs(539));
    outputs(3473) <= not(layer0_outputs(912));
    outputs(3474) <= not(layer0_outputs(3806));
    outputs(3475) <= (layer0_outputs(12)) and (layer0_outputs(3944));
    outputs(3476) <= layer0_outputs(4611);
    outputs(3477) <= not((layer0_outputs(3276)) and (layer0_outputs(124)));
    outputs(3478) <= not(layer0_outputs(501));
    outputs(3479) <= layer0_outputs(327);
    outputs(3480) <= not(layer0_outputs(3695));
    outputs(3481) <= layer0_outputs(421);
    outputs(3482) <= (layer0_outputs(629)) and not (layer0_outputs(1617));
    outputs(3483) <= (layer0_outputs(774)) and not (layer0_outputs(3472));
    outputs(3484) <= (layer0_outputs(1637)) and (layer0_outputs(2973));
    outputs(3485) <= not(layer0_outputs(854));
    outputs(3486) <= not(layer0_outputs(3628)) or (layer0_outputs(3916));
    outputs(3487) <= layer0_outputs(1016);
    outputs(3488) <= (layer0_outputs(4562)) and not (layer0_outputs(2450));
    outputs(3489) <= not(layer0_outputs(1394));
    outputs(3490) <= not(layer0_outputs(3116));
    outputs(3491) <= (layer0_outputs(4109)) and not (layer0_outputs(4571));
    outputs(3492) <= not(layer0_outputs(1260));
    outputs(3493) <= (layer0_outputs(4420)) and not (layer0_outputs(2406));
    outputs(3494) <= not((layer0_outputs(721)) or (layer0_outputs(3164)));
    outputs(3495) <= not(layer0_outputs(1797));
    outputs(3496) <= not((layer0_outputs(2355)) xor (layer0_outputs(4292)));
    outputs(3497) <= not((layer0_outputs(823)) and (layer0_outputs(2705)));
    outputs(3498) <= not(layer0_outputs(3937));
    outputs(3499) <= layer0_outputs(4288);
    outputs(3500) <= not(layer0_outputs(3454)) or (layer0_outputs(2776));
    outputs(3501) <= layer0_outputs(778);
    outputs(3502) <= not((layer0_outputs(2478)) and (layer0_outputs(2319)));
    outputs(3503) <= layer0_outputs(2819);
    outputs(3504) <= layer0_outputs(3428);
    outputs(3505) <= not(layer0_outputs(4742));
    outputs(3506) <= layer0_outputs(524);
    outputs(3507) <= layer0_outputs(4986);
    outputs(3508) <= layer0_outputs(1868);
    outputs(3509) <= not(layer0_outputs(1858)) or (layer0_outputs(4160));
    outputs(3510) <= (layer0_outputs(1986)) or (layer0_outputs(1852));
    outputs(3511) <= not(layer0_outputs(1930)) or (layer0_outputs(1843));
    outputs(3512) <= layer0_outputs(286);
    outputs(3513) <= not(layer0_outputs(1743)) or (layer0_outputs(1863));
    outputs(3514) <= not(layer0_outputs(3496));
    outputs(3515) <= not((layer0_outputs(3033)) or (layer0_outputs(1170)));
    outputs(3516) <= layer0_outputs(2272);
    outputs(3517) <= (layer0_outputs(4311)) and not (layer0_outputs(1152));
    outputs(3518) <= not(layer0_outputs(1613));
    outputs(3519) <= not(layer0_outputs(4814));
    outputs(3520) <= (layer0_outputs(2241)) or (layer0_outputs(1481));
    outputs(3521) <= (layer0_outputs(4655)) and not (layer0_outputs(1164));
    outputs(3522) <= (layer0_outputs(3760)) and not (layer0_outputs(3464));
    outputs(3523) <= not(layer0_outputs(351));
    outputs(3524) <= not(layer0_outputs(2684)) or (layer0_outputs(3585));
    outputs(3525) <= not((layer0_outputs(1215)) and (layer0_outputs(413)));
    outputs(3526) <= not((layer0_outputs(2724)) or (layer0_outputs(794)));
    outputs(3527) <= not((layer0_outputs(2830)) or (layer0_outputs(2023)));
    outputs(3528) <= not(layer0_outputs(4409));
    outputs(3529) <= layer0_outputs(1099);
    outputs(3530) <= not(layer0_outputs(4520));
    outputs(3531) <= (layer0_outputs(228)) and not (layer0_outputs(422));
    outputs(3532) <= (layer0_outputs(1125)) xor (layer0_outputs(4474));
    outputs(3533) <= (layer0_outputs(2936)) and not (layer0_outputs(2718));
    outputs(3534) <= (layer0_outputs(654)) and not (layer0_outputs(230));
    outputs(3535) <= (layer0_outputs(2872)) and not (layer0_outputs(3012));
    outputs(3536) <= (layer0_outputs(2057)) and not (layer0_outputs(3919));
    outputs(3537) <= (layer0_outputs(4407)) xor (layer0_outputs(4579));
    outputs(3538) <= layer0_outputs(2117);
    outputs(3539) <= not(layer0_outputs(4758));
    outputs(3540) <= layer0_outputs(768);
    outputs(3541) <= (layer0_outputs(748)) xor (layer0_outputs(949));
    outputs(3542) <= (layer0_outputs(4259)) or (layer0_outputs(2305));
    outputs(3543) <= (layer0_outputs(2656)) and not (layer0_outputs(1609));
    outputs(3544) <= not((layer0_outputs(3217)) xor (layer0_outputs(2153)));
    outputs(3545) <= layer0_outputs(3183);
    outputs(3546) <= (layer0_outputs(2557)) and not (layer0_outputs(4648));
    outputs(3547) <= not(layer0_outputs(2984));
    outputs(3548) <= layer0_outputs(1891);
    outputs(3549) <= layer0_outputs(4740);
    outputs(3550) <= (layer0_outputs(4904)) and (layer0_outputs(3383));
    outputs(3551) <= not(layer0_outputs(3462));
    outputs(3552) <= layer0_outputs(4310);
    outputs(3553) <= not((layer0_outputs(2688)) or (layer0_outputs(4651)));
    outputs(3554) <= not(layer0_outputs(1165));
    outputs(3555) <= not((layer0_outputs(248)) or (layer0_outputs(4554)));
    outputs(3556) <= (layer0_outputs(2097)) and not (layer0_outputs(258));
    outputs(3557) <= not(layer0_outputs(1427)) or (layer0_outputs(3411));
    outputs(3558) <= (layer0_outputs(4613)) and not (layer0_outputs(676));
    outputs(3559) <= (layer0_outputs(1126)) and not (layer0_outputs(2419));
    outputs(3560) <= not(layer0_outputs(873));
    outputs(3561) <= layer0_outputs(98);
    outputs(3562) <= not(layer0_outputs(1314));
    outputs(3563) <= not(layer0_outputs(2658));
    outputs(3564) <= not(layer0_outputs(356));
    outputs(3565) <= (layer0_outputs(69)) and not (layer0_outputs(3744));
    outputs(3566) <= (layer0_outputs(3791)) and not (layer0_outputs(1604));
    outputs(3567) <= not(layer0_outputs(202));
    outputs(3568) <= (layer0_outputs(915)) and not (layer0_outputs(2952));
    outputs(3569) <= (layer0_outputs(4243)) and (layer0_outputs(2459));
    outputs(3570) <= not(layer0_outputs(558));
    outputs(3571) <= not(layer0_outputs(3984)) or (layer0_outputs(448));
    outputs(3572) <= not(layer0_outputs(3540));
    outputs(3573) <= layer0_outputs(1965);
    outputs(3574) <= not(layer0_outputs(166));
    outputs(3575) <= layer0_outputs(2931);
    outputs(3576) <= layer0_outputs(1143);
    outputs(3577) <= layer0_outputs(4086);
    outputs(3578) <= (layer0_outputs(712)) and not (layer0_outputs(1337));
    outputs(3579) <= layer0_outputs(192);
    outputs(3580) <= (layer0_outputs(3796)) and not (layer0_outputs(2339));
    outputs(3581) <= not((layer0_outputs(1819)) or (layer0_outputs(4543)));
    outputs(3582) <= not(layer0_outputs(4371));
    outputs(3583) <= not(layer0_outputs(2976));
    outputs(3584) <= (layer0_outputs(587)) and (layer0_outputs(3225));
    outputs(3585) <= layer0_outputs(3660);
    outputs(3586) <= not(layer0_outputs(4137));
    outputs(3587) <= layer0_outputs(4517);
    outputs(3588) <= (layer0_outputs(1246)) and not (layer0_outputs(1870));
    outputs(3589) <= not((layer0_outputs(1419)) xor (layer0_outputs(332)));
    outputs(3590) <= not(layer0_outputs(3665));
    outputs(3591) <= not((layer0_outputs(925)) or (layer0_outputs(3796)));
    outputs(3592) <= (layer0_outputs(3937)) or (layer0_outputs(1371));
    outputs(3593) <= not(layer0_outputs(4242));
    outputs(3594) <= not(layer0_outputs(3095));
    outputs(3595) <= not((layer0_outputs(2895)) or (layer0_outputs(2990)));
    outputs(3596) <= not(layer0_outputs(115));
    outputs(3597) <= layer0_outputs(897);
    outputs(3598) <= not((layer0_outputs(4455)) or (layer0_outputs(3855)));
    outputs(3599) <= layer0_outputs(1453);
    outputs(3600) <= not(layer0_outputs(1964));
    outputs(3601) <= layer0_outputs(952);
    outputs(3602) <= not(layer0_outputs(4978));
    outputs(3603) <= (layer0_outputs(1820)) and not (layer0_outputs(4618));
    outputs(3604) <= layer0_outputs(2052);
    outputs(3605) <= (layer0_outputs(3115)) or (layer0_outputs(2605));
    outputs(3606) <= not(layer0_outputs(1134));
    outputs(3607) <= (layer0_outputs(2158)) and not (layer0_outputs(75));
    outputs(3608) <= (layer0_outputs(4292)) and not (layer0_outputs(4730));
    outputs(3609) <= not(layer0_outputs(1431));
    outputs(3610) <= (layer0_outputs(1427)) and not (layer0_outputs(3715));
    outputs(3611) <= not(layer0_outputs(4081));
    outputs(3612) <= layer0_outputs(3291);
    outputs(3613) <= not(layer0_outputs(4692));
    outputs(3614) <= layer0_outputs(2227);
    outputs(3615) <= (layer0_outputs(2196)) and not (layer0_outputs(4059));
    outputs(3616) <= layer0_outputs(1362);
    outputs(3617) <= (layer0_outputs(3209)) and not (layer0_outputs(3461));
    outputs(3618) <= (layer0_outputs(2248)) and not (layer0_outputs(2505));
    outputs(3619) <= not((layer0_outputs(2255)) xor (layer0_outputs(1653)));
    outputs(3620) <= not((layer0_outputs(2491)) or (layer0_outputs(4437)));
    outputs(3621) <= layer0_outputs(4933);
    outputs(3622) <= layer0_outputs(2369);
    outputs(3623) <= not(layer0_outputs(4660));
    outputs(3624) <= not((layer0_outputs(3555)) and (layer0_outputs(1746)));
    outputs(3625) <= not((layer0_outputs(1476)) or (layer0_outputs(3516)));
    outputs(3626) <= layer0_outputs(697);
    outputs(3627) <= not((layer0_outputs(2855)) xor (layer0_outputs(3388)));
    outputs(3628) <= not(layer0_outputs(4525)) or (layer0_outputs(4094));
    outputs(3629) <= layer0_outputs(1954);
    outputs(3630) <= layer0_outputs(239);
    outputs(3631) <= not(layer0_outputs(370));
    outputs(3632) <= (layer0_outputs(4032)) and not (layer0_outputs(2628));
    outputs(3633) <= not(layer0_outputs(2205));
    outputs(3634) <= not(layer0_outputs(1997));
    outputs(3635) <= not(layer0_outputs(1458));
    outputs(3636) <= not((layer0_outputs(3778)) or (layer0_outputs(375)));
    outputs(3637) <= (layer0_outputs(1248)) xor (layer0_outputs(1430));
    outputs(3638) <= (layer0_outputs(4042)) and not (layer0_outputs(564));
    outputs(3639) <= not(layer0_outputs(2191));
    outputs(3640) <= not(layer0_outputs(5100));
    outputs(3641) <= not((layer0_outputs(2799)) xor (layer0_outputs(2033)));
    outputs(3642) <= not((layer0_outputs(3507)) or (layer0_outputs(1028)));
    outputs(3643) <= (layer0_outputs(4404)) or (layer0_outputs(2083));
    outputs(3644) <= not(layer0_outputs(4463)) or (layer0_outputs(1260));
    outputs(3645) <= layer0_outputs(683);
    outputs(3646) <= (layer0_outputs(2040)) and (layer0_outputs(4563));
    outputs(3647) <= not(layer0_outputs(4986));
    outputs(3648) <= not(layer0_outputs(2200));
    outputs(3649) <= not(layer0_outputs(1559));
    outputs(3650) <= not(layer0_outputs(290)) or (layer0_outputs(3560));
    outputs(3651) <= not((layer0_outputs(4605)) or (layer0_outputs(2845)));
    outputs(3652) <= (layer0_outputs(4810)) and not (layer0_outputs(1506));
    outputs(3653) <= not(layer0_outputs(2145));
    outputs(3654) <= not(layer0_outputs(3757));
    outputs(3655) <= not((layer0_outputs(4899)) or (layer0_outputs(540)));
    outputs(3656) <= layer0_outputs(1574);
    outputs(3657) <= (layer0_outputs(807)) and (layer0_outputs(2727));
    outputs(3658) <= not(layer0_outputs(2462));
    outputs(3659) <= (layer0_outputs(1928)) and not (layer0_outputs(2758));
    outputs(3660) <= not(layer0_outputs(4107));
    outputs(3661) <= layer0_outputs(3012);
    outputs(3662) <= layer0_outputs(3419);
    outputs(3663) <= (layer0_outputs(4960)) xor (layer0_outputs(4324));
    outputs(3664) <= not(layer0_outputs(228)) or (layer0_outputs(223));
    outputs(3665) <= layer0_outputs(2809);
    outputs(3666) <= layer0_outputs(3874);
    outputs(3667) <= (layer0_outputs(326)) and not (layer0_outputs(3966));
    outputs(3668) <= (layer0_outputs(2029)) and not (layer0_outputs(1102));
    outputs(3669) <= (layer0_outputs(1153)) and not (layer0_outputs(1556));
    outputs(3670) <= not((layer0_outputs(3729)) xor (layer0_outputs(3434)));
    outputs(3671) <= not(layer0_outputs(3650));
    outputs(3672) <= not(layer0_outputs(1767)) or (layer0_outputs(499));
    outputs(3673) <= layer0_outputs(3639);
    outputs(3674) <= (layer0_outputs(1733)) and not (layer0_outputs(217));
    outputs(3675) <= not(layer0_outputs(867));
    outputs(3676) <= (layer0_outputs(3068)) xor (layer0_outputs(161));
    outputs(3677) <= layer0_outputs(2384);
    outputs(3678) <= not((layer0_outputs(2204)) or (layer0_outputs(4799)));
    outputs(3679) <= (layer0_outputs(881)) or (layer0_outputs(3054));
    outputs(3680) <= (layer0_outputs(340)) and not (layer0_outputs(344));
    outputs(3681) <= layer0_outputs(4593);
    outputs(3682) <= layer0_outputs(4199);
    outputs(3683) <= not((layer0_outputs(68)) or (layer0_outputs(1326)));
    outputs(3684) <= not(layer0_outputs(60)) or (layer0_outputs(650));
    outputs(3685) <= (layer0_outputs(1969)) and not (layer0_outputs(352));
    outputs(3686) <= (layer0_outputs(2461)) or (layer0_outputs(1391));
    outputs(3687) <= not(layer0_outputs(1209));
    outputs(3688) <= layer0_outputs(1453);
    outputs(3689) <= not(layer0_outputs(5054));
    outputs(3690) <= not(layer0_outputs(1940));
    outputs(3691) <= (layer0_outputs(2779)) xor (layer0_outputs(967));
    outputs(3692) <= (layer0_outputs(184)) and not (layer0_outputs(3310));
    outputs(3693) <= (layer0_outputs(3312)) and not (layer0_outputs(4305));
    outputs(3694) <= not(layer0_outputs(3793));
    outputs(3695) <= not(layer0_outputs(860));
    outputs(3696) <= (layer0_outputs(994)) and (layer0_outputs(70));
    outputs(3697) <= not(layer0_outputs(1734));
    outputs(3698) <= not((layer0_outputs(92)) or (layer0_outputs(4070)));
    outputs(3699) <= not(layer0_outputs(4100)) or (layer0_outputs(1212));
    outputs(3700) <= not(layer0_outputs(4254));
    outputs(3701) <= layer0_outputs(276);
    outputs(3702) <= not(layer0_outputs(504));
    outputs(3703) <= not(layer0_outputs(2334));
    outputs(3704) <= not(layer0_outputs(1993));
    outputs(3705) <= not(layer0_outputs(4053));
    outputs(3706) <= layer0_outputs(2436);
    outputs(3707) <= (layer0_outputs(3399)) and (layer0_outputs(3529));
    outputs(3708) <= (layer0_outputs(1957)) and not (layer0_outputs(1174));
    outputs(3709) <= (layer0_outputs(4523)) and (layer0_outputs(2158));
    outputs(3710) <= (layer0_outputs(2838)) and not (layer0_outputs(2993));
    outputs(3711) <= not(layer0_outputs(4572));
    outputs(3712) <= not(layer0_outputs(1228));
    outputs(3713) <= not(layer0_outputs(2652)) or (layer0_outputs(964));
    outputs(3714) <= (layer0_outputs(4519)) and (layer0_outputs(2661));
    outputs(3715) <= layer0_outputs(1066);
    outputs(3716) <= not(layer0_outputs(34));
    outputs(3717) <= layer0_outputs(1791);
    outputs(3718) <= not((layer0_outputs(3701)) or (layer0_outputs(253)));
    outputs(3719) <= not(layer0_outputs(2308));
    outputs(3720) <= (layer0_outputs(4281)) and not (layer0_outputs(2967));
    outputs(3721) <= not(layer0_outputs(3404));
    outputs(3722) <= (layer0_outputs(3000)) and (layer0_outputs(1906));
    outputs(3723) <= layer0_outputs(3542);
    outputs(3724) <= (layer0_outputs(2788)) and not (layer0_outputs(4029));
    outputs(3725) <= (layer0_outputs(3060)) xor (layer0_outputs(4480));
    outputs(3726) <= not(layer0_outputs(956));
    outputs(3727) <= layer0_outputs(1239);
    outputs(3728) <= (layer0_outputs(4801)) and not (layer0_outputs(430));
    outputs(3729) <= (layer0_outputs(2079)) and not (layer0_outputs(5030));
    outputs(3730) <= (layer0_outputs(2532)) and not (layer0_outputs(4072));
    outputs(3731) <= (layer0_outputs(2526)) and not (layer0_outputs(4542));
    outputs(3732) <= not(layer0_outputs(535));
    outputs(3733) <= not(layer0_outputs(3248));
    outputs(3734) <= not(layer0_outputs(421));
    outputs(3735) <= not((layer0_outputs(1855)) or (layer0_outputs(265)));
    outputs(3736) <= (layer0_outputs(4354)) or (layer0_outputs(546));
    outputs(3737) <= (layer0_outputs(3223)) and not (layer0_outputs(5101));
    outputs(3738) <= not((layer0_outputs(2738)) or (layer0_outputs(3008)));
    outputs(3739) <= (layer0_outputs(4252)) or (layer0_outputs(2617));
    outputs(3740) <= not(layer0_outputs(2506));
    outputs(3741) <= (layer0_outputs(180)) and not (layer0_outputs(1396));
    outputs(3742) <= not(layer0_outputs(1094)) or (layer0_outputs(1661));
    outputs(3743) <= not((layer0_outputs(4427)) or (layer0_outputs(4731)));
    outputs(3744) <= layer0_outputs(2380);
    outputs(3745) <= layer0_outputs(2025);
    outputs(3746) <= layer0_outputs(2894);
    outputs(3747) <= not(layer0_outputs(4531));
    outputs(3748) <= (layer0_outputs(3807)) and not (layer0_outputs(3672));
    outputs(3749) <= not(layer0_outputs(4088));
    outputs(3750) <= layer0_outputs(1803);
    outputs(3751) <= not(layer0_outputs(1633));
    outputs(3752) <= (layer0_outputs(4555)) and (layer0_outputs(2089));
    outputs(3753) <= (layer0_outputs(3749)) and not (layer0_outputs(2055));
    outputs(3754) <= not((layer0_outputs(3171)) or (layer0_outputs(5090)));
    outputs(3755) <= (layer0_outputs(4164)) and (layer0_outputs(4127));
    outputs(3756) <= not(layer0_outputs(3169));
    outputs(3757) <= layer0_outputs(151);
    outputs(3758) <= (layer0_outputs(3317)) xor (layer0_outputs(3));
    outputs(3759) <= (layer0_outputs(3364)) and not (layer0_outputs(1741));
    outputs(3760) <= not(layer0_outputs(1402));
    outputs(3761) <= (layer0_outputs(1121)) xor (layer0_outputs(1801));
    outputs(3762) <= layer0_outputs(2800);
    outputs(3763) <= (layer0_outputs(3155)) and (layer0_outputs(461));
    outputs(3764) <= layer0_outputs(113);
    outputs(3765) <= layer0_outputs(895);
    outputs(3766) <= (layer0_outputs(1893)) and not (layer0_outputs(4201));
    outputs(3767) <= (layer0_outputs(5055)) xor (layer0_outputs(986));
    outputs(3768) <= not((layer0_outputs(5061)) or (layer0_outputs(215)));
    outputs(3769) <= layer0_outputs(1318);
    outputs(3770) <= not((layer0_outputs(510)) or (layer0_outputs(2483)));
    outputs(3771) <= not((layer0_outputs(956)) or (layer0_outputs(167)));
    outputs(3772) <= layer0_outputs(930);
    outputs(3773) <= (layer0_outputs(2087)) and (layer0_outputs(4638));
    outputs(3774) <= not(layer0_outputs(2988)) or (layer0_outputs(2038));
    outputs(3775) <= (layer0_outputs(2452)) and not (layer0_outputs(4741));
    outputs(3776) <= (layer0_outputs(4189)) xor (layer0_outputs(4125));
    outputs(3777) <= (layer0_outputs(3814)) and not (layer0_outputs(1289));
    outputs(3778) <= (layer0_outputs(266)) and not (layer0_outputs(4977));
    outputs(3779) <= (layer0_outputs(2566)) and not (layer0_outputs(635));
    outputs(3780) <= layer0_outputs(1733);
    outputs(3781) <= (layer0_outputs(4184)) xor (layer0_outputs(4571));
    outputs(3782) <= not(layer0_outputs(4789)) or (layer0_outputs(1422));
    outputs(3783) <= not(layer0_outputs(4608));
    outputs(3784) <= layer0_outputs(392);
    outputs(3785) <= layer0_outputs(678);
    outputs(3786) <= (layer0_outputs(3176)) and (layer0_outputs(4414));
    outputs(3787) <= (layer0_outputs(543)) and not (layer0_outputs(2492));
    outputs(3788) <= not((layer0_outputs(4144)) and (layer0_outputs(4435)));
    outputs(3789) <= layer0_outputs(1874);
    outputs(3790) <= layer0_outputs(2401);
    outputs(3791) <= not(layer0_outputs(42)) or (layer0_outputs(2075));
    outputs(3792) <= layer0_outputs(435);
    outputs(3793) <= not((layer0_outputs(424)) or (layer0_outputs(3243)));
    outputs(3794) <= (layer0_outputs(3536)) and not (layer0_outputs(503));
    outputs(3795) <= not(layer0_outputs(3945));
    outputs(3796) <= not(layer0_outputs(423));
    outputs(3797) <= layer0_outputs(1813);
    outputs(3798) <= layer0_outputs(2093);
    outputs(3799) <= (layer0_outputs(977)) xor (layer0_outputs(3294));
    outputs(3800) <= not((layer0_outputs(109)) and (layer0_outputs(1011)));
    outputs(3801) <= not(layer0_outputs(2503));
    outputs(3802) <= (layer0_outputs(2164)) and not (layer0_outputs(992));
    outputs(3803) <= (layer0_outputs(4812)) and not (layer0_outputs(1277));
    outputs(3804) <= (layer0_outputs(216)) and (layer0_outputs(1301));
    outputs(3805) <= (layer0_outputs(2401)) and not (layer0_outputs(4259));
    outputs(3806) <= (layer0_outputs(4776)) and not (layer0_outputs(4070));
    outputs(3807) <= not(layer0_outputs(1898));
    outputs(3808) <= (layer0_outputs(2750)) and not (layer0_outputs(3733));
    outputs(3809) <= (layer0_outputs(3295)) or (layer0_outputs(2317));
    outputs(3810) <= not((layer0_outputs(3986)) or (layer0_outputs(1181)));
    outputs(3811) <= (layer0_outputs(3533)) or (layer0_outputs(4010));
    outputs(3812) <= not(layer0_outputs(2007));
    outputs(3813) <= (layer0_outputs(2433)) and (layer0_outputs(3270));
    outputs(3814) <= not(layer0_outputs(2457));
    outputs(3815) <= (layer0_outputs(4991)) and not (layer0_outputs(3665));
    outputs(3816) <= not(layer0_outputs(4158));
    outputs(3817) <= layer0_outputs(4643);
    outputs(3818) <= (layer0_outputs(1936)) and (layer0_outputs(3405));
    outputs(3819) <= not(layer0_outputs(5097));
    outputs(3820) <= (layer0_outputs(4411)) and (layer0_outputs(3754));
    outputs(3821) <= not((layer0_outputs(2143)) or (layer0_outputs(4026)));
    outputs(3822) <= not((layer0_outputs(4553)) or (layer0_outputs(4106)));
    outputs(3823) <= not((layer0_outputs(2995)) or (layer0_outputs(1174)));
    outputs(3824) <= (layer0_outputs(2279)) or (layer0_outputs(2891));
    outputs(3825) <= not((layer0_outputs(869)) or (layer0_outputs(3003)));
    outputs(3826) <= (layer0_outputs(5095)) or (layer0_outputs(323));
    outputs(3827) <= not((layer0_outputs(313)) and (layer0_outputs(1739)));
    outputs(3828) <= layer0_outputs(1819);
    outputs(3829) <= not(layer0_outputs(302));
    outputs(3830) <= (layer0_outputs(1177)) or (layer0_outputs(4536));
    outputs(3831) <= (layer0_outputs(1526)) and (layer0_outputs(1192));
    outputs(3832) <= not((layer0_outputs(4715)) xor (layer0_outputs(3638)));
    outputs(3833) <= not(layer0_outputs(3269)) or (layer0_outputs(1112));
    outputs(3834) <= not((layer0_outputs(1046)) or (layer0_outputs(1317)));
    outputs(3835) <= not(layer0_outputs(1737)) or (layer0_outputs(3065));
    outputs(3836) <= not(layer0_outputs(661));
    outputs(3837) <= (layer0_outputs(94)) and not (layer0_outputs(3508));
    outputs(3838) <= layer0_outputs(3818);
    outputs(3839) <= (layer0_outputs(640)) and (layer0_outputs(809));
    outputs(3840) <= layer0_outputs(1057);
    outputs(3841) <= layer0_outputs(4877);
    outputs(3842) <= not((layer0_outputs(597)) or (layer0_outputs(4739)));
    outputs(3843) <= layer0_outputs(108);
    outputs(3844) <= not((layer0_outputs(597)) or (layer0_outputs(3351)));
    outputs(3845) <= not(layer0_outputs(4092));
    outputs(3846) <= layer0_outputs(233);
    outputs(3847) <= (layer0_outputs(1666)) xor (layer0_outputs(886));
    outputs(3848) <= not((layer0_outputs(1147)) or (layer0_outputs(3285)));
    outputs(3849) <= layer0_outputs(3056);
    outputs(3850) <= (layer0_outputs(4005)) and not (layer0_outputs(1561));
    outputs(3851) <= not(layer0_outputs(3453));
    outputs(3852) <= layer0_outputs(2839);
    outputs(3853) <= (layer0_outputs(4460)) and not (layer0_outputs(2457));
    outputs(3854) <= (layer0_outputs(1274)) and (layer0_outputs(517));
    outputs(3855) <= not(layer0_outputs(2813)) or (layer0_outputs(4496));
    outputs(3856) <= not(layer0_outputs(4851));
    outputs(3857) <= not((layer0_outputs(2548)) or (layer0_outputs(1532)));
    outputs(3858) <= not(layer0_outputs(3173));
    outputs(3859) <= layer0_outputs(581);
    outputs(3860) <= (layer0_outputs(2026)) and not (layer0_outputs(4993));
    outputs(3861) <= (layer0_outputs(4168)) and (layer0_outputs(3147));
    outputs(3862) <= not(layer0_outputs(4143));
    outputs(3863) <= not(layer0_outputs(1181));
    outputs(3864) <= (layer0_outputs(4526)) or (layer0_outputs(2719));
    outputs(3865) <= not(layer0_outputs(4909));
    outputs(3866) <= not((layer0_outputs(4549)) or (layer0_outputs(752)));
    outputs(3867) <= (layer0_outputs(1367)) and (layer0_outputs(2672));
    outputs(3868) <= (layer0_outputs(3985)) or (layer0_outputs(2730));
    outputs(3869) <= not(layer0_outputs(4513));
    outputs(3870) <= not(layer0_outputs(2402));
    outputs(3871) <= (layer0_outputs(3146)) and not (layer0_outputs(1822));
    outputs(3872) <= not((layer0_outputs(4924)) xor (layer0_outputs(5114)));
    outputs(3873) <= not((layer0_outputs(4320)) xor (layer0_outputs(2300)));
    outputs(3874) <= not(layer0_outputs(318));
    outputs(3875) <= not(layer0_outputs(2508));
    outputs(3876) <= (layer0_outputs(1208)) and (layer0_outputs(3150));
    outputs(3877) <= not(layer0_outputs(3427));
    outputs(3878) <= not((layer0_outputs(4177)) and (layer0_outputs(891)));
    outputs(3879) <= layer0_outputs(4675);
    outputs(3880) <= (layer0_outputs(4821)) and not (layer0_outputs(106));
    outputs(3881) <= not(layer0_outputs(4082));
    outputs(3882) <= (layer0_outputs(4983)) and not (layer0_outputs(3911));
    outputs(3883) <= not(layer0_outputs(712));
    outputs(3884) <= (layer0_outputs(1052)) and (layer0_outputs(1346));
    outputs(3885) <= (layer0_outputs(3717)) and not (layer0_outputs(2028));
    outputs(3886) <= not(layer0_outputs(2503));
    outputs(3887) <= (layer0_outputs(3201)) and not (layer0_outputs(734));
    outputs(3888) <= (layer0_outputs(4645)) and (layer0_outputs(871));
    outputs(3889) <= not(layer0_outputs(2350));
    outputs(3890) <= layer0_outputs(1070);
    outputs(3891) <= (layer0_outputs(4216)) and (layer0_outputs(2190));
    outputs(3892) <= (layer0_outputs(4991)) and not (layer0_outputs(3332));
    outputs(3893) <= (layer0_outputs(1759)) xor (layer0_outputs(1114));
    outputs(3894) <= (layer0_outputs(1)) xor (layer0_outputs(768));
    outputs(3895) <= not((layer0_outputs(3148)) or (layer0_outputs(3832)));
    outputs(3896) <= not(layer0_outputs(2449)) or (layer0_outputs(4974));
    outputs(3897) <= layer0_outputs(4574);
    outputs(3898) <= not(layer0_outputs(4155)) or (layer0_outputs(2125));
    outputs(3899) <= layer0_outputs(4802);
    outputs(3900) <= layer0_outputs(3915);
    outputs(3901) <= layer0_outputs(4400);
    outputs(3902) <= (layer0_outputs(4526)) or (layer0_outputs(931));
    outputs(3903) <= not((layer0_outputs(574)) and (layer0_outputs(2249)));
    outputs(3904) <= not(layer0_outputs(5057));
    outputs(3905) <= (layer0_outputs(3484)) and not (layer0_outputs(3830));
    outputs(3906) <= layer0_outputs(4623);
    outputs(3907) <= (layer0_outputs(3783)) and (layer0_outputs(4935));
    outputs(3908) <= (layer0_outputs(471)) and not (layer0_outputs(1988));
    outputs(3909) <= (layer0_outputs(843)) and not (layer0_outputs(901));
    outputs(3910) <= (layer0_outputs(2998)) and not (layer0_outputs(2689));
    outputs(3911) <= (layer0_outputs(645)) and not (layer0_outputs(537));
    outputs(3912) <= layer0_outputs(4686);
    outputs(3913) <= (layer0_outputs(3789)) and (layer0_outputs(5026));
    outputs(3914) <= (layer0_outputs(2478)) and not (layer0_outputs(1672));
    outputs(3915) <= (layer0_outputs(3396)) and (layer0_outputs(4912));
    outputs(3916) <= not((layer0_outputs(4463)) and (layer0_outputs(2011)));
    outputs(3917) <= not(layer0_outputs(737));
    outputs(3918) <= (layer0_outputs(748)) and not (layer0_outputs(511));
    outputs(3919) <= layer0_outputs(3359);
    outputs(3920) <= layer0_outputs(4119);
    outputs(3921) <= not((layer0_outputs(942)) xor (layer0_outputs(44)));
    outputs(3922) <= (layer0_outputs(4896)) and (layer0_outputs(2439));
    outputs(3923) <= (layer0_outputs(3205)) and not (layer0_outputs(2575));
    outputs(3924) <= not(layer0_outputs(2241));
    outputs(3925) <= (layer0_outputs(968)) and not (layer0_outputs(2364));
    outputs(3926) <= not(layer0_outputs(2429));
    outputs(3927) <= (layer0_outputs(4008)) and not (layer0_outputs(1213));
    outputs(3928) <= (layer0_outputs(850)) xor (layer0_outputs(1847));
    outputs(3929) <= not(layer0_outputs(2505));
    outputs(3930) <= layer0_outputs(2515);
    outputs(3931) <= not(layer0_outputs(623)) or (layer0_outputs(1528));
    outputs(3932) <= (layer0_outputs(2703)) and not (layer0_outputs(3991));
    outputs(3933) <= (layer0_outputs(3886)) and (layer0_outputs(4060));
    outputs(3934) <= (layer0_outputs(4273)) and not (layer0_outputs(4852));
    outputs(3935) <= (layer0_outputs(1778)) and not (layer0_outputs(1461));
    outputs(3936) <= (layer0_outputs(618)) and not (layer0_outputs(737));
    outputs(3937) <= not((layer0_outputs(4673)) or (layer0_outputs(1036)));
    outputs(3938) <= (layer0_outputs(234)) xor (layer0_outputs(3202));
    outputs(3939) <= layer0_outputs(4919);
    outputs(3940) <= not(layer0_outputs(4773));
    outputs(3941) <= layer0_outputs(4844);
    outputs(3942) <= not(layer0_outputs(1129));
    outputs(3943) <= not(layer0_outputs(4058));
    outputs(3944) <= (layer0_outputs(2763)) and not (layer0_outputs(4162));
    outputs(3945) <= layer0_outputs(2642);
    outputs(3946) <= layer0_outputs(954);
    outputs(3947) <= (layer0_outputs(1186)) and not (layer0_outputs(4006));
    outputs(3948) <= not(layer0_outputs(1659));
    outputs(3949) <= not(layer0_outputs(370));
    outputs(3950) <= (layer0_outputs(2722)) xor (layer0_outputs(2414));
    outputs(3951) <= layer0_outputs(3115);
    outputs(3952) <= not((layer0_outputs(2152)) or (layer0_outputs(3374)));
    outputs(3953) <= layer0_outputs(3447);
    outputs(3954) <= (layer0_outputs(3337)) and (layer0_outputs(624));
    outputs(3955) <= not(layer0_outputs(2020));
    outputs(3956) <= not((layer0_outputs(2379)) or (layer0_outputs(117)));
    outputs(3957) <= (layer0_outputs(606)) and not (layer0_outputs(3003));
    outputs(3958) <= (layer0_outputs(3528)) and (layer0_outputs(1548));
    outputs(3959) <= (layer0_outputs(397)) and (layer0_outputs(3017));
    outputs(3960) <= (layer0_outputs(2002)) xor (layer0_outputs(659));
    outputs(3961) <= not((layer0_outputs(3907)) xor (layer0_outputs(2808)));
    outputs(3962) <= not(layer0_outputs(4806)) or (layer0_outputs(4824));
    outputs(3963) <= (layer0_outputs(4450)) and (layer0_outputs(741));
    outputs(3964) <= not(layer0_outputs(3982));
    outputs(3965) <= (layer0_outputs(1765)) and (layer0_outputs(4507));
    outputs(3966) <= (layer0_outputs(1189)) and not (layer0_outputs(2555));
    outputs(3967) <= not((layer0_outputs(1929)) or (layer0_outputs(1157)));
    outputs(3968) <= not((layer0_outputs(1489)) and (layer0_outputs(2833)));
    outputs(3969) <= (layer0_outputs(1333)) and not (layer0_outputs(3588));
    outputs(3970) <= not((layer0_outputs(4057)) xor (layer0_outputs(1952)));
    outputs(3971) <= not((layer0_outputs(2856)) or (layer0_outputs(1549)));
    outputs(3972) <= not((layer0_outputs(1990)) and (layer0_outputs(1994)));
    outputs(3973) <= not((layer0_outputs(4037)) and (layer0_outputs(705)));
    outputs(3974) <= (layer0_outputs(3494)) and not (layer0_outputs(3768));
    outputs(3975) <= (layer0_outputs(5023)) and not (layer0_outputs(1726));
    outputs(3976) <= (layer0_outputs(2582)) and (layer0_outputs(4194));
    outputs(3977) <= layer0_outputs(4105);
    outputs(3978) <= not((layer0_outputs(528)) or (layer0_outputs(4048)));
    outputs(3979) <= (layer0_outputs(5021)) and not (layer0_outputs(5061));
    outputs(3980) <= not(layer0_outputs(3720));
    outputs(3981) <= (layer0_outputs(4348)) and (layer0_outputs(2073));
    outputs(3982) <= not(layer0_outputs(601));
    outputs(3983) <= (layer0_outputs(80)) xor (layer0_outputs(1669));
    outputs(3984) <= layer0_outputs(1221);
    outputs(3985) <= not((layer0_outputs(1047)) and (layer0_outputs(4585)));
    outputs(3986) <= (layer0_outputs(3)) xor (layer0_outputs(2430));
    outputs(3987) <= not(layer0_outputs(1466)) or (layer0_outputs(2050));
    outputs(3988) <= layer0_outputs(3448);
    outputs(3989) <= (layer0_outputs(3025)) and (layer0_outputs(3585));
    outputs(3990) <= not(layer0_outputs(1017)) or (layer0_outputs(2454));
    outputs(3991) <= (layer0_outputs(3110)) and (layer0_outputs(369));
    outputs(3992) <= (layer0_outputs(3124)) and not (layer0_outputs(1566));
    outputs(3993) <= not(layer0_outputs(3671));
    outputs(3994) <= (layer0_outputs(3313)) xor (layer0_outputs(4924));
    outputs(3995) <= not(layer0_outputs(1884));
    outputs(3996) <= (layer0_outputs(4017)) and not (layer0_outputs(2910));
    outputs(3997) <= layer0_outputs(3035);
    outputs(3998) <= not((layer0_outputs(1352)) xor (layer0_outputs(5036)));
    outputs(3999) <= (layer0_outputs(4038)) and not (layer0_outputs(4495));
    outputs(4000) <= not((layer0_outputs(3772)) and (layer0_outputs(4635)));
    outputs(4001) <= (layer0_outputs(1405)) and not (layer0_outputs(3758));
    outputs(4002) <= not(layer0_outputs(1309)) or (layer0_outputs(3198));
    outputs(4003) <= not(layer0_outputs(23));
    outputs(4004) <= (layer0_outputs(4651)) or (layer0_outputs(1574));
    outputs(4005) <= layer0_outputs(3464);
    outputs(4006) <= (layer0_outputs(2439)) and (layer0_outputs(1097));
    outputs(4007) <= not(layer0_outputs(2146));
    outputs(4008) <= layer0_outputs(1261);
    outputs(4009) <= layer0_outputs(1404);
    outputs(4010) <= not((layer0_outputs(3283)) or (layer0_outputs(552)));
    outputs(4011) <= not((layer0_outputs(1997)) or (layer0_outputs(1430)));
    outputs(4012) <= layer0_outputs(4105);
    outputs(4013) <= layer0_outputs(644);
    outputs(4014) <= not((layer0_outputs(2678)) or (layer0_outputs(3598)));
    outputs(4015) <= (layer0_outputs(4816)) and (layer0_outputs(3147));
    outputs(4016) <= layer0_outputs(3152);
    outputs(4017) <= not(layer0_outputs(2133));
    outputs(4018) <= (layer0_outputs(1544)) and (layer0_outputs(711));
    outputs(4019) <= not(layer0_outputs(4353));
    outputs(4020) <= (layer0_outputs(1906)) and not (layer0_outputs(3575));
    outputs(4021) <= not((layer0_outputs(2954)) xor (layer0_outputs(1727)));
    outputs(4022) <= layer0_outputs(3974);
    outputs(4023) <= layer0_outputs(2245);
    outputs(4024) <= layer0_outputs(3239);
    outputs(4025) <= not((layer0_outputs(4809)) or (layer0_outputs(3310)));
    outputs(4026) <= not((layer0_outputs(4856)) xor (layer0_outputs(912)));
    outputs(4027) <= not(layer0_outputs(23));
    outputs(4028) <= (layer0_outputs(273)) and not (layer0_outputs(3599));
    outputs(4029) <= layer0_outputs(4918);
    outputs(4030) <= (layer0_outputs(2639)) or (layer0_outputs(1348));
    outputs(4031) <= layer0_outputs(922);
    outputs(4032) <= not(layer0_outputs(4205)) or (layer0_outputs(4260));
    outputs(4033) <= layer0_outputs(1210);
    outputs(4034) <= layer0_outputs(1269);
    outputs(4035) <= (layer0_outputs(4073)) and not (layer0_outputs(4165));
    outputs(4036) <= not((layer0_outputs(4175)) and (layer0_outputs(2148)));
    outputs(4037) <= layer0_outputs(1945);
    outputs(4038) <= not(layer0_outputs(4405));
    outputs(4039) <= not(layer0_outputs(2966));
    outputs(4040) <= not(layer0_outputs(4793));
    outputs(4041) <= not((layer0_outputs(4754)) and (layer0_outputs(1511)));
    outputs(4042) <= (layer0_outputs(4956)) and not (layer0_outputs(3212));
    outputs(4043) <= not((layer0_outputs(2948)) and (layer0_outputs(4426)));
    outputs(4044) <= not((layer0_outputs(3756)) or (layer0_outputs(440)));
    outputs(4045) <= not(layer0_outputs(2820));
    outputs(4046) <= layer0_outputs(4996);
    outputs(4047) <= not(layer0_outputs(5083));
    outputs(4048) <= not(layer0_outputs(4437));
    outputs(4049) <= layer0_outputs(4948);
    outputs(4050) <= (layer0_outputs(2265)) and not (layer0_outputs(2594));
    outputs(4051) <= layer0_outputs(4700);
    outputs(4052) <= not((layer0_outputs(2348)) xor (layer0_outputs(2099)));
    outputs(4053) <= not(layer0_outputs(4203));
    outputs(4054) <= not(layer0_outputs(2044)) or (layer0_outputs(4139));
    outputs(4055) <= not((layer0_outputs(900)) or (layer0_outputs(1939)));
    outputs(4056) <= (layer0_outputs(2563)) and not (layer0_outputs(3871));
    outputs(4057) <= layer0_outputs(3815);
    outputs(4058) <= not((layer0_outputs(3920)) or (layer0_outputs(3220)));
    outputs(4059) <= not(layer0_outputs(2664));
    outputs(4060) <= not(layer0_outputs(3154));
    outputs(4061) <= layer0_outputs(3350);
    outputs(4062) <= (layer0_outputs(3497)) or (layer0_outputs(3949));
    outputs(4063) <= (layer0_outputs(1831)) and not (layer0_outputs(3096));
    outputs(4064) <= layer0_outputs(3467);
    outputs(4065) <= layer0_outputs(325);
    outputs(4066) <= layer0_outputs(1456);
    outputs(4067) <= (layer0_outputs(4383)) and not (layer0_outputs(1480));
    outputs(4068) <= (layer0_outputs(3390)) and not (layer0_outputs(1910));
    outputs(4069) <= not(layer0_outputs(3118));
    outputs(4070) <= layer0_outputs(4964);
    outputs(4071) <= layer0_outputs(4973);
    outputs(4072) <= (layer0_outputs(1284)) and (layer0_outputs(2824));
    outputs(4073) <= layer0_outputs(4140);
    outputs(4074) <= not((layer0_outputs(251)) xor (layer0_outputs(4556)));
    outputs(4075) <= (layer0_outputs(4881)) and (layer0_outputs(2532));
    outputs(4076) <= (layer0_outputs(2132)) and not (layer0_outputs(4219));
    outputs(4077) <= not(layer0_outputs(1493));
    outputs(4078) <= not((layer0_outputs(75)) or (layer0_outputs(79)));
    outputs(4079) <= not((layer0_outputs(2061)) or (layer0_outputs(869)));
    outputs(4080) <= (layer0_outputs(1614)) and not (layer0_outputs(4601));
    outputs(4081) <= (layer0_outputs(4227)) and (layer0_outputs(2657));
    outputs(4082) <= layer0_outputs(2314);
    outputs(4083) <= (layer0_outputs(637)) and not (layer0_outputs(4448));
    outputs(4084) <= layer0_outputs(2169);
    outputs(4085) <= (layer0_outputs(4367)) and not (layer0_outputs(995));
    outputs(4086) <= (layer0_outputs(1496)) and (layer0_outputs(2806));
    outputs(4087) <= layer0_outputs(3327);
    outputs(4088) <= not((layer0_outputs(2192)) or (layer0_outputs(3274)));
    outputs(4089) <= not(layer0_outputs(2287)) or (layer0_outputs(3041));
    outputs(4090) <= not(layer0_outputs(749));
    outputs(4091) <= layer0_outputs(77);
    outputs(4092) <= (layer0_outputs(2109)) and (layer0_outputs(1323));
    outputs(4093) <= not(layer0_outputs(2222));
    outputs(4094) <= (layer0_outputs(3531)) and (layer0_outputs(2729));
    outputs(4095) <= not(layer0_outputs(68));
    outputs(4096) <= not(layer0_outputs(1432));
    outputs(4097) <= (layer0_outputs(811)) and not (layer0_outputs(2690));
    outputs(4098) <= (layer0_outputs(2007)) and (layer0_outputs(4681));
    outputs(4099) <= layer0_outputs(1521);
    outputs(4100) <= layer0_outputs(3170);
    outputs(4101) <= not(layer0_outputs(204));
    outputs(4102) <= not(layer0_outputs(1136));
    outputs(4103) <= layer0_outputs(4577);
    outputs(4104) <= not(layer0_outputs(1016));
    outputs(4105) <= layer0_outputs(1489);
    outputs(4106) <= (layer0_outputs(510)) and not (layer0_outputs(4969));
    outputs(4107) <= layer0_outputs(536);
    outputs(4108) <= (layer0_outputs(176)) and (layer0_outputs(3717));
    outputs(4109) <= layer0_outputs(4739);
    outputs(4110) <= layer0_outputs(3583);
    outputs(4111) <= not(layer0_outputs(1989)) or (layer0_outputs(3227));
    outputs(4112) <= not(layer0_outputs(2547));
    outputs(4113) <= layer0_outputs(264);
    outputs(4114) <= not(layer0_outputs(4192)) or (layer0_outputs(4244));
    outputs(4115) <= layer0_outputs(3474);
    outputs(4116) <= not((layer0_outputs(4871)) and (layer0_outputs(1964)));
    outputs(4117) <= not((layer0_outputs(2898)) or (layer0_outputs(2699)));
    outputs(4118) <= not(layer0_outputs(3288));
    outputs(4119) <= not((layer0_outputs(1777)) xor (layer0_outputs(1845)));
    outputs(4120) <= (layer0_outputs(1595)) and (layer0_outputs(1557));
    outputs(4121) <= not(layer0_outputs(841));
    outputs(4122) <= (layer0_outputs(319)) or (layer0_outputs(3217));
    outputs(4123) <= not(layer0_outputs(3351)) or (layer0_outputs(2472));
    outputs(4124) <= not((layer0_outputs(136)) and (layer0_outputs(4607)));
    outputs(4125) <= not(layer0_outputs(2444)) or (layer0_outputs(2950));
    outputs(4126) <= not(layer0_outputs(4076)) or (layer0_outputs(2123));
    outputs(4127) <= not(layer0_outputs(1096)) or (layer0_outputs(3034));
    outputs(4128) <= not(layer0_outputs(1763));
    outputs(4129) <= not(layer0_outputs(4533));
    outputs(4130) <= not(layer0_outputs(406)) or (layer0_outputs(2079));
    outputs(4131) <= layer0_outputs(1744);
    outputs(4132) <= (layer0_outputs(1228)) xor (layer0_outputs(1256));
    outputs(4133) <= (layer0_outputs(521)) and not (layer0_outputs(188));
    outputs(4134) <= not((layer0_outputs(3405)) xor (layer0_outputs(4251)));
    outputs(4135) <= (layer0_outputs(665)) xor (layer0_outputs(2308));
    outputs(4136) <= layer0_outputs(541);
    outputs(4137) <= not(layer0_outputs(4148));
    outputs(4138) <= (layer0_outputs(3619)) and not (layer0_outputs(761));
    outputs(4139) <= not(layer0_outputs(4629));
    outputs(4140) <= (layer0_outputs(3906)) and not (layer0_outputs(3849));
    outputs(4141) <= layer0_outputs(1751);
    outputs(4142) <= not((layer0_outputs(2984)) xor (layer0_outputs(4062)));
    outputs(4143) <= not(layer0_outputs(773)) or (layer0_outputs(2370));
    outputs(4144) <= not((layer0_outputs(3347)) xor (layer0_outputs(605)));
    outputs(4145) <= layer0_outputs(1214);
    outputs(4146) <= (layer0_outputs(304)) and not (layer0_outputs(2798));
    outputs(4147) <= layer0_outputs(4356);
    outputs(4148) <= not(layer0_outputs(171));
    outputs(4149) <= not(layer0_outputs(357));
    outputs(4150) <= not(layer0_outputs(342)) or (layer0_outputs(2740));
    outputs(4151) <= not(layer0_outputs(1355));
    outputs(4152) <= not((layer0_outputs(1088)) xor (layer0_outputs(1762)));
    outputs(4153) <= (layer0_outputs(1235)) xor (layer0_outputs(2027));
    outputs(4154) <= not((layer0_outputs(353)) and (layer0_outputs(809)));
    outputs(4155) <= (layer0_outputs(2168)) and not (layer0_outputs(1104));
    outputs(4156) <= (layer0_outputs(1328)) and (layer0_outputs(2476));
    outputs(4157) <= not(layer0_outputs(2942));
    outputs(4158) <= layer0_outputs(3546);
    outputs(4159) <= (layer0_outputs(180)) xor (layer0_outputs(4066));
    outputs(4160) <= not(layer0_outputs(4057));
    outputs(4161) <= not(layer0_outputs(3807));
    outputs(4162) <= not(layer0_outputs(360)) or (layer0_outputs(3098));
    outputs(4163) <= layer0_outputs(1079);
    outputs(4164) <= not(layer0_outputs(3123));
    outputs(4165) <= not(layer0_outputs(1320));
    outputs(4166) <= layer0_outputs(2391);
    outputs(4167) <= not((layer0_outputs(2661)) and (layer0_outputs(2340)));
    outputs(4168) <= (layer0_outputs(1218)) and (layer0_outputs(3089));
    outputs(4169) <= layer0_outputs(2358);
    outputs(4170) <= (layer0_outputs(1900)) xor (layer0_outputs(3642));
    outputs(4171) <= (layer0_outputs(2105)) and not (layer0_outputs(774));
    outputs(4172) <= not(layer0_outputs(65));
    outputs(4173) <= layer0_outputs(1481);
    outputs(4174) <= (layer0_outputs(3201)) or (layer0_outputs(4641));
    outputs(4175) <= layer0_outputs(2594);
    outputs(4176) <= not((layer0_outputs(4784)) xor (layer0_outputs(1616)));
    outputs(4177) <= not(layer0_outputs(896));
    outputs(4178) <= not(layer0_outputs(3122)) or (layer0_outputs(1895));
    outputs(4179) <= not(layer0_outputs(3402)) or (layer0_outputs(3871));
    outputs(4180) <= (layer0_outputs(1424)) and (layer0_outputs(5065));
    outputs(4181) <= not((layer0_outputs(1282)) xor (layer0_outputs(427)));
    outputs(4182) <= (layer0_outputs(4149)) and not (layer0_outputs(2402));
    outputs(4183) <= not(layer0_outputs(137));
    outputs(4184) <= not((layer0_outputs(1645)) or (layer0_outputs(139)));
    outputs(4185) <= layer0_outputs(2965);
    outputs(4186) <= layer0_outputs(1702);
    outputs(4187) <= layer0_outputs(3679);
    outputs(4188) <= not(layer0_outputs(3366));
    outputs(4189) <= not(layer0_outputs(4562)) or (layer0_outputs(2665));
    outputs(4190) <= not(layer0_outputs(937));
    outputs(4191) <= layer0_outputs(779);
    outputs(4192) <= (layer0_outputs(1605)) or (layer0_outputs(3723));
    outputs(4193) <= not(layer0_outputs(3622));
    outputs(4194) <= layer0_outputs(2161);
    outputs(4195) <= not(layer0_outputs(4955));
    outputs(4196) <= (layer0_outputs(2864)) or (layer0_outputs(2363));
    outputs(4197) <= (layer0_outputs(2424)) xor (layer0_outputs(2430));
    outputs(4198) <= not(layer0_outputs(3273));
    outputs(4199) <= not((layer0_outputs(4890)) xor (layer0_outputs(1982)));
    outputs(4200) <= (layer0_outputs(3685)) and not (layer0_outputs(1659));
    outputs(4201) <= layer0_outputs(4217);
    outputs(4202) <= not(layer0_outputs(3918));
    outputs(4203) <= not(layer0_outputs(267)) or (layer0_outputs(314));
    outputs(4204) <= layer0_outputs(4432);
    outputs(4205) <= not(layer0_outputs(1237));
    outputs(4206) <= not((layer0_outputs(1509)) xor (layer0_outputs(1799)));
    outputs(4207) <= layer0_outputs(3083);
    outputs(4208) <= not((layer0_outputs(20)) xor (layer0_outputs(4805)));
    outputs(4209) <= (layer0_outputs(667)) and not (layer0_outputs(798));
    outputs(4210) <= layer0_outputs(2596);
    outputs(4211) <= not((layer0_outputs(235)) or (layer0_outputs(4014)));
    outputs(4212) <= (layer0_outputs(4175)) xor (layer0_outputs(4656));
    outputs(4213) <= not(layer0_outputs(4745)) or (layer0_outputs(191));
    outputs(4214) <= layer0_outputs(310);
    outputs(4215) <= not(layer0_outputs(1006));
    outputs(4216) <= not(layer0_outputs(1303)) or (layer0_outputs(4743));
    outputs(4217) <= not((layer0_outputs(412)) and (layer0_outputs(2545)));
    outputs(4218) <= not(layer0_outputs(1492));
    outputs(4219) <= not((layer0_outputs(1335)) xor (layer0_outputs(418)));
    outputs(4220) <= not(layer0_outputs(4412));
    outputs(4221) <= not((layer0_outputs(2802)) or (layer0_outputs(4695)));
    outputs(4222) <= not((layer0_outputs(1200)) xor (layer0_outputs(3734)));
    outputs(4223) <= (layer0_outputs(2298)) and (layer0_outputs(4401));
    outputs(4224) <= layer0_outputs(903);
    outputs(4225) <= not((layer0_outputs(2320)) xor (layer0_outputs(331)));
    outputs(4226) <= not(layer0_outputs(2442));
    outputs(4227) <= not((layer0_outputs(3549)) and (layer0_outputs(3373)));
    outputs(4228) <= (layer0_outputs(702)) xor (layer0_outputs(449));
    outputs(4229) <= not(layer0_outputs(3942));
    outputs(4230) <= not((layer0_outputs(3551)) or (layer0_outputs(1095)));
    outputs(4231) <= (layer0_outputs(1392)) and not (layer0_outputs(1106));
    outputs(4232) <= (layer0_outputs(664)) and not (layer0_outputs(4819));
    outputs(4233) <= not(layer0_outputs(2921));
    outputs(4234) <= layer0_outputs(4663);
    outputs(4235) <= layer0_outputs(3527);
    outputs(4236) <= not((layer0_outputs(4580)) or (layer0_outputs(2444)));
    outputs(4237) <= not((layer0_outputs(2967)) xor (layer0_outputs(1540)));
    outputs(4238) <= not(layer0_outputs(2164));
    outputs(4239) <= (layer0_outputs(3885)) xor (layer0_outputs(1257));
    outputs(4240) <= not(layer0_outputs(3101));
    outputs(4241) <= (layer0_outputs(2811)) xor (layer0_outputs(4861));
    outputs(4242) <= layer0_outputs(671);
    outputs(4243) <= (layer0_outputs(4262)) xor (layer0_outputs(2209));
    outputs(4244) <= not(layer0_outputs(2116)) or (layer0_outputs(376));
    outputs(4245) <= layer0_outputs(2866);
    outputs(4246) <= layer0_outputs(2948);
    outputs(4247) <= (layer0_outputs(902)) xor (layer0_outputs(405));
    outputs(4248) <= not((layer0_outputs(2132)) xor (layer0_outputs(380)));
    outputs(4249) <= not(layer0_outputs(3384));
    outputs(4250) <= not(layer0_outputs(1283)) or (layer0_outputs(5042));
    outputs(4251) <= not(layer0_outputs(3016));
    outputs(4252) <= not(layer0_outputs(2579));
    outputs(4253) <= layer0_outputs(5054);
    outputs(4254) <= not((layer0_outputs(630)) xor (layer0_outputs(3955)));
    outputs(4255) <= (layer0_outputs(1161)) or (layer0_outputs(3792));
    outputs(4256) <= layer0_outputs(4271);
    outputs(4257) <= (layer0_outputs(3346)) and not (layer0_outputs(3936));
    outputs(4258) <= not(layer0_outputs(431));
    outputs(4259) <= layer0_outputs(4845);
    outputs(4260) <= (layer0_outputs(4317)) and (layer0_outputs(795));
    outputs(4261) <= layer0_outputs(295);
    outputs(4262) <= layer0_outputs(2085);
    outputs(4263) <= not(layer0_outputs(3988));
    outputs(4264) <= layer0_outputs(2911);
    outputs(4265) <= not((layer0_outputs(3144)) or (layer0_outputs(4376)));
    outputs(4266) <= layer0_outputs(1115);
    outputs(4267) <= not((layer0_outputs(1375)) xor (layer0_outputs(2844)));
    outputs(4268) <= not(layer0_outputs(2649));
    outputs(4269) <= (layer0_outputs(1995)) and not (layer0_outputs(367));
    outputs(4270) <= (layer0_outputs(2270)) xor (layer0_outputs(4846));
    outputs(4271) <= layer0_outputs(4087);
    outputs(4272) <= not(layer0_outputs(3994));
    outputs(4273) <= layer0_outputs(2494);
    outputs(4274) <= (layer0_outputs(3391)) or (layer0_outputs(1038));
    outputs(4275) <= not(layer0_outputs(1582));
    outputs(4276) <= not((layer0_outputs(3054)) or (layer0_outputs(2251)));
    outputs(4277) <= not(layer0_outputs(917));
    outputs(4278) <= layer0_outputs(2005);
    outputs(4279) <= not(layer0_outputs(3766)) or (layer0_outputs(1163));
    outputs(4280) <= not((layer0_outputs(2273)) xor (layer0_outputs(3505)));
    outputs(4281) <= layer0_outputs(4887);
    outputs(4282) <= (layer0_outputs(3272)) or (layer0_outputs(163));
    outputs(4283) <= not(layer0_outputs(1830));
    outputs(4284) <= not(layer0_outputs(4872));
    outputs(4285) <= layer0_outputs(503);
    outputs(4286) <= not((layer0_outputs(729)) or (layer0_outputs(4415)));
    outputs(4287) <= not((layer0_outputs(4990)) or (layer0_outputs(557)));
    outputs(4288) <= not(layer0_outputs(4865));
    outputs(4289) <= layer0_outputs(2953);
    outputs(4290) <= not(layer0_outputs(3151));
    outputs(4291) <= not(layer0_outputs(3159));
    outputs(4292) <= not((layer0_outputs(5068)) and (layer0_outputs(1464)));
    outputs(4293) <= not((layer0_outputs(164)) xor (layer0_outputs(3064)));
    outputs(4294) <= (layer0_outputs(1781)) or (layer0_outputs(1310));
    outputs(4295) <= not(layer0_outputs(4575));
    outputs(4296) <= not((layer0_outputs(1866)) or (layer0_outputs(3279)));
    outputs(4297) <= not((layer0_outputs(4148)) xor (layer0_outputs(5)));
    outputs(4298) <= not((layer0_outputs(3593)) and (layer0_outputs(4386)));
    outputs(4299) <= layer0_outputs(1446);
    outputs(4300) <= layer0_outputs(4451);
    outputs(4301) <= (layer0_outputs(110)) and (layer0_outputs(1844));
    outputs(4302) <= not(layer0_outputs(3645)) or (layer0_outputs(2071));
    outputs(4303) <= not(layer0_outputs(3123));
    outputs(4304) <= not(layer0_outputs(2377));
    outputs(4305) <= layer0_outputs(2250);
    outputs(4306) <= layer0_outputs(4288);
    outputs(4307) <= layer0_outputs(4061);
    outputs(4308) <= layer0_outputs(2504);
    outputs(4309) <= not(layer0_outputs(3458)) or (layer0_outputs(3066));
    outputs(4310) <= not((layer0_outputs(1623)) or (layer0_outputs(4684)));
    outputs(4311) <= (layer0_outputs(4377)) or (layer0_outputs(1993));
    outputs(4312) <= not(layer0_outputs(4872)) or (layer0_outputs(2773));
    outputs(4313) <= not((layer0_outputs(2820)) xor (layer0_outputs(1425)));
    outputs(4314) <= layer0_outputs(3669);
    outputs(4315) <= not(layer0_outputs(3984)) or (layer0_outputs(3007));
    outputs(4316) <= (layer0_outputs(657)) xor (layer0_outputs(2049));
    outputs(4317) <= not(layer0_outputs(3328));
    outputs(4318) <= not(layer0_outputs(817)) or (layer0_outputs(3846));
    outputs(4319) <= not(layer0_outputs(4859));
    outputs(4320) <= not(layer0_outputs(3317));
    outputs(4321) <= layer0_outputs(241);
    outputs(4322) <= '1';
    outputs(4323) <= layer0_outputs(2955);
    outputs(4324) <= (layer0_outputs(3566)) xor (layer0_outputs(1037));
    outputs(4325) <= (layer0_outputs(3676)) xor (layer0_outputs(1832));
    outputs(4326) <= (layer0_outputs(3640)) or (layer0_outputs(2962));
    outputs(4327) <= not((layer0_outputs(2860)) xor (layer0_outputs(434)));
    outputs(4328) <= (layer0_outputs(2176)) and not (layer0_outputs(635));
    outputs(4329) <= (layer0_outputs(2874)) and not (layer0_outputs(4634));
    outputs(4330) <= not((layer0_outputs(1699)) or (layer0_outputs(1575)));
    outputs(4331) <= not(layer0_outputs(3593));
    outputs(4332) <= layer0_outputs(1139);
    outputs(4333) <= not((layer0_outputs(3511)) and (layer0_outputs(3242)));
    outputs(4334) <= (layer0_outputs(1393)) xor (layer0_outputs(4992));
    outputs(4335) <= layer0_outputs(573);
    outputs(4336) <= (layer0_outputs(1723)) and not (layer0_outputs(4835));
    outputs(4337) <= layer0_outputs(4650);
    outputs(4338) <= not(layer0_outputs(3692));
    outputs(4339) <= not(layer0_outputs(4253)) or (layer0_outputs(2137));
    outputs(4340) <= not(layer0_outputs(4193)) or (layer0_outputs(2516));
    outputs(4341) <= (layer0_outputs(3838)) and not (layer0_outputs(170));
    outputs(4342) <= not((layer0_outputs(3800)) xor (layer0_outputs(4334)));
    outputs(4343) <= (layer0_outputs(3362)) or (layer0_outputs(3395));
    outputs(4344) <= layer0_outputs(1864);
    outputs(4345) <= not(layer0_outputs(3590)) or (layer0_outputs(2559));
    outputs(4346) <= not(layer0_outputs(426));
    outputs(4347) <= layer0_outputs(3432);
    outputs(4348) <= (layer0_outputs(3232)) xor (layer0_outputs(3407));
    outputs(4349) <= (layer0_outputs(4260)) or (layer0_outputs(2911));
    outputs(4350) <= (layer0_outputs(482)) and not (layer0_outputs(1094));
    outputs(4351) <= not(layer0_outputs(5074)) or (layer0_outputs(3127));
    outputs(4352) <= not((layer0_outputs(4747)) and (layer0_outputs(927)));
    outputs(4353) <= not(layer0_outputs(4418));
    outputs(4354) <= layer0_outputs(2663);
    outputs(4355) <= layer0_outputs(1092);
    outputs(4356) <= not(layer0_outputs(2660));
    outputs(4357) <= layer0_outputs(5073);
    outputs(4358) <= not((layer0_outputs(893)) and (layer0_outputs(2772)));
    outputs(4359) <= (layer0_outputs(4178)) xor (layer0_outputs(3232));
    outputs(4360) <= (layer0_outputs(999)) or (layer0_outputs(4768));
    outputs(4361) <= layer0_outputs(4119);
    outputs(4362) <= not((layer0_outputs(4759)) or (layer0_outputs(5012)));
    outputs(4363) <= not(layer0_outputs(111));
    outputs(4364) <= not(layer0_outputs(4839));
    outputs(4365) <= layer0_outputs(1089);
    outputs(4366) <= not(layer0_outputs(4602)) or (layer0_outputs(1344));
    outputs(4367) <= not(layer0_outputs(2670));
    outputs(4368) <= not(layer0_outputs(3148));
    outputs(4369) <= not(layer0_outputs(1266));
    outputs(4370) <= not(layer0_outputs(3586)) or (layer0_outputs(3782));
    outputs(4371) <= not((layer0_outputs(2446)) xor (layer0_outputs(4014)));
    outputs(4372) <= not((layer0_outputs(1896)) xor (layer0_outputs(1187)));
    outputs(4373) <= not((layer0_outputs(973)) xor (layer0_outputs(1525)));
    outputs(4374) <= (layer0_outputs(1546)) and not (layer0_outputs(4545));
    outputs(4375) <= layer0_outputs(777);
    outputs(4376) <= (layer0_outputs(1342)) or (layer0_outputs(4676));
    outputs(4377) <= (layer0_outputs(230)) xor (layer0_outputs(2609));
    outputs(4378) <= (layer0_outputs(2272)) xor (layer0_outputs(3142));
    outputs(4379) <= not((layer0_outputs(4206)) xor (layer0_outputs(2598)));
    outputs(4380) <= (layer0_outputs(4509)) or (layer0_outputs(2135));
    outputs(4381) <= not(layer0_outputs(3612));
    outputs(4382) <= not((layer0_outputs(1536)) xor (layer0_outputs(1189)));
    outputs(4383) <= (layer0_outputs(2679)) and (layer0_outputs(4215));
    outputs(4384) <= not(layer0_outputs(3216)) or (layer0_outputs(5085));
    outputs(4385) <= (layer0_outputs(596)) xor (layer0_outputs(555));
    outputs(4386) <= not((layer0_outputs(2606)) and (layer0_outputs(1878)));
    outputs(4387) <= (layer0_outputs(491)) or (layer0_outputs(1059));
    outputs(4388) <= layer0_outputs(3263);
    outputs(4389) <= (layer0_outputs(4030)) and not (layer0_outputs(1865));
    outputs(4390) <= not((layer0_outputs(1285)) xor (layer0_outputs(1987)));
    outputs(4391) <= layer0_outputs(1047);
    outputs(4392) <= (layer0_outputs(21)) and not (layer0_outputs(5013));
    outputs(4393) <= not(layer0_outputs(3672));
    outputs(4394) <= not((layer0_outputs(1367)) and (layer0_outputs(2817)));
    outputs(4395) <= layer0_outputs(867);
    outputs(4396) <= (layer0_outputs(1067)) and not (layer0_outputs(4421));
    outputs(4397) <= layer0_outputs(379);
    outputs(4398) <= (layer0_outputs(2504)) and not (layer0_outputs(2879));
    outputs(4399) <= not((layer0_outputs(151)) xor (layer0_outputs(4297)));
    outputs(4400) <= layer0_outputs(71);
    outputs(4401) <= layer0_outputs(1551);
    outputs(4402) <= not(layer0_outputs(1140));
    outputs(4403) <= not(layer0_outputs(3484));
    outputs(4404) <= not(layer0_outputs(1802));
    outputs(4405) <= not(layer0_outputs(427));
    outputs(4406) <= layer0_outputs(1133);
    outputs(4407) <= not((layer0_outputs(3696)) and (layer0_outputs(1184)));
    outputs(4408) <= not((layer0_outputs(3030)) and (layer0_outputs(4719)));
    outputs(4409) <= layer0_outputs(1639);
    outputs(4410) <= not((layer0_outputs(776)) xor (layer0_outputs(2275)));
    outputs(4411) <= not((layer0_outputs(1172)) xor (layer0_outputs(1474)));
    outputs(4412) <= (layer0_outputs(835)) and (layer0_outputs(655));
    outputs(4413) <= (layer0_outputs(1707)) xor (layer0_outputs(5089));
    outputs(4414) <= not((layer0_outputs(3954)) and (layer0_outputs(18)));
    outputs(4415) <= (layer0_outputs(454)) and (layer0_outputs(3820));
    outputs(4416) <= not((layer0_outputs(2346)) xor (layer0_outputs(1851)));
    outputs(4417) <= not(layer0_outputs(4537));
    outputs(4418) <= not((layer0_outputs(4408)) xor (layer0_outputs(2126)));
    outputs(4419) <= (layer0_outputs(3188)) xor (layer0_outputs(2937));
    outputs(4420) <= not(layer0_outputs(4183));
    outputs(4421) <= layer0_outputs(3909);
    outputs(4422) <= not((layer0_outputs(2774)) and (layer0_outputs(4576)));
    outputs(4423) <= not(layer0_outputs(2119)) or (layer0_outputs(2266));
    outputs(4424) <= not((layer0_outputs(1144)) xor (layer0_outputs(1892)));
    outputs(4425) <= not((layer0_outputs(1513)) or (layer0_outputs(4184)));
    outputs(4426) <= layer0_outputs(221);
    outputs(4427) <= not((layer0_outputs(1307)) xor (layer0_outputs(4915)));
    outputs(4428) <= not(layer0_outputs(2792));
    outputs(4429) <= not(layer0_outputs(2788));
    outputs(4430) <= (layer0_outputs(2438)) or (layer0_outputs(3247));
    outputs(4431) <= not((layer0_outputs(1811)) xor (layer0_outputs(1683)));
    outputs(4432) <= (layer0_outputs(3774)) xor (layer0_outputs(4316));
    outputs(4433) <= not(layer0_outputs(874));
    outputs(4434) <= not(layer0_outputs(3983)) or (layer0_outputs(1406));
    outputs(4435) <= layer0_outputs(2509);
    outputs(4436) <= (layer0_outputs(3125)) or (layer0_outputs(1542));
    outputs(4437) <= not(layer0_outputs(1902));
    outputs(4438) <= layer0_outputs(4521);
    outputs(4439) <= (layer0_outputs(2824)) xor (layer0_outputs(981));
    outputs(4440) <= not((layer0_outputs(1854)) and (layer0_outputs(965)));
    outputs(4441) <= not((layer0_outputs(3539)) xor (layer0_outputs(1757)));
    outputs(4442) <= not(layer0_outputs(1376));
    outputs(4443) <= (layer0_outputs(1537)) and (layer0_outputs(3607));
    outputs(4444) <= not(layer0_outputs(4707));
    outputs(4445) <= (layer0_outputs(1030)) xor (layer0_outputs(682));
    outputs(4446) <= layer0_outputs(4957);
    outputs(4447) <= not(layer0_outputs(2475)) or (layer0_outputs(2487));
    outputs(4448) <= layer0_outputs(3179);
    outputs(4449) <= (layer0_outputs(3371)) xor (layer0_outputs(4392));
    outputs(4450) <= not((layer0_outputs(577)) xor (layer0_outputs(3552)));
    outputs(4451) <= not((layer0_outputs(2753)) and (layer0_outputs(3594)));
    outputs(4452) <= not(layer0_outputs(3070));
    outputs(4453) <= (layer0_outputs(5091)) xor (layer0_outputs(3641));
    outputs(4454) <= not(layer0_outputs(58));
    outputs(4455) <= layer0_outputs(2479);
    outputs(4456) <= (layer0_outputs(2373)) and (layer0_outputs(1086));
    outputs(4457) <= not((layer0_outputs(5079)) xor (layer0_outputs(4975)));
    outputs(4458) <= layer0_outputs(4201);
    outputs(4459) <= layer0_outputs(3470);
    outputs(4460) <= not(layer0_outputs(4633));
    outputs(4461) <= (layer0_outputs(1867)) xor (layer0_outputs(5060));
    outputs(4462) <= not(layer0_outputs(2711)) or (layer0_outputs(327));
    outputs(4463) <= not(layer0_outputs(572)) or (layer0_outputs(2084));
    outputs(4464) <= not((layer0_outputs(2969)) xor (layer0_outputs(940)));
    outputs(4465) <= layer0_outputs(3728);
    outputs(4466) <= layer0_outputs(1343);
    outputs(4467) <= layer0_outputs(4212);
    outputs(4468) <= not((layer0_outputs(1587)) and (layer0_outputs(877)));
    outputs(4469) <= not(layer0_outputs(5082)) or (layer0_outputs(5000));
    outputs(4470) <= (layer0_outputs(3654)) and not (layer0_outputs(3368));
    outputs(4471) <= not(layer0_outputs(394));
    outputs(4472) <= (layer0_outputs(3641)) xor (layer0_outputs(2118));
    outputs(4473) <= not(layer0_outputs(4686));
    outputs(4474) <= not(layer0_outputs(4096));
    outputs(4475) <= not(layer0_outputs(3063));
    outputs(4476) <= (layer0_outputs(485)) and not (layer0_outputs(2620));
    outputs(4477) <= layer0_outputs(3753);
    outputs(4478) <= not(layer0_outputs(1764));
    outputs(4479) <= (layer0_outputs(1920)) and not (layer0_outputs(88));
    outputs(4480) <= layer0_outputs(3406);
    outputs(4481) <= not(layer0_outputs(2868));
    outputs(4482) <= not(layer0_outputs(1827)) or (layer0_outputs(2283));
    outputs(4483) <= (layer0_outputs(3919)) or (layer0_outputs(3007));
    outputs(4484) <= (layer0_outputs(4408)) or (layer0_outputs(676));
    outputs(4485) <= layer0_outputs(4360);
    outputs(4486) <= not(layer0_outputs(3029)) or (layer0_outputs(4567));
    outputs(4487) <= (layer0_outputs(1973)) and (layer0_outputs(3709));
    outputs(4488) <= not(layer0_outputs(3068)) or (layer0_outputs(4081));
    outputs(4489) <= not((layer0_outputs(1632)) xor (layer0_outputs(2975)));
    outputs(4490) <= not(layer0_outputs(1307));
    outputs(4491) <= not((layer0_outputs(1173)) and (layer0_outputs(696)));
    outputs(4492) <= not((layer0_outputs(1062)) xor (layer0_outputs(4064)));
    outputs(4493) <= not(layer0_outputs(4540)) or (layer0_outputs(1610));
    outputs(4494) <= not((layer0_outputs(5097)) xor (layer0_outputs(1911)));
    outputs(4495) <= not(layer0_outputs(35)) or (layer0_outputs(4459));
    outputs(4496) <= not((layer0_outputs(921)) xor (layer0_outputs(33)));
    outputs(4497) <= (layer0_outputs(871)) xor (layer0_outputs(2011));
    outputs(4498) <= layer0_outputs(2981);
    outputs(4499) <= not(layer0_outputs(5102));
    outputs(4500) <= not(layer0_outputs(4636));
    outputs(4501) <= layer0_outputs(2151);
    outputs(4502) <= (layer0_outputs(4804)) or (layer0_outputs(673));
    outputs(4503) <= not(layer0_outputs(3902));
    outputs(4504) <= layer0_outputs(4351);
    outputs(4505) <= not(layer0_outputs(4415));
    outputs(4506) <= not((layer0_outputs(3549)) xor (layer0_outputs(3335)));
    outputs(4507) <= (layer0_outputs(1967)) and (layer0_outputs(515));
    outputs(4508) <= (layer0_outputs(1689)) and not (layer0_outputs(2339));
    outputs(4509) <= not(layer0_outputs(4198));
    outputs(4510) <= not((layer0_outputs(4418)) or (layer0_outputs(3591)));
    outputs(4511) <= not((layer0_outputs(2959)) and (layer0_outputs(314)));
    outputs(4512) <= layer0_outputs(3186);
    outputs(4513) <= (layer0_outputs(1702)) and not (layer0_outputs(889));
    outputs(4514) <= (layer0_outputs(3916)) xor (layer0_outputs(1684));
    outputs(4515) <= not(layer0_outputs(4937)) or (layer0_outputs(4398));
    outputs(4516) <= layer0_outputs(118);
    outputs(4517) <= layer0_outputs(1595);
    outputs(4518) <= not(layer0_outputs(3262));
    outputs(4519) <= (layer0_outputs(3199)) and not (layer0_outputs(78));
    outputs(4520) <= not(layer0_outputs(2342));
    outputs(4521) <= layer0_outputs(3980);
    outputs(4522) <= not(layer0_outputs(3752));
    outputs(4523) <= (layer0_outputs(3060)) and not (layer0_outputs(200));
    outputs(4524) <= not(layer0_outputs(2405));
    outputs(4525) <= not((layer0_outputs(1835)) xor (layer0_outputs(993)));
    outputs(4526) <= not(layer0_outputs(1019)) or (layer0_outputs(911));
    outputs(4527) <= layer0_outputs(2382);
    outputs(4528) <= layer0_outputs(966);
    outputs(4529) <= not((layer0_outputs(4639)) or (layer0_outputs(594)));
    outputs(4530) <= (layer0_outputs(4488)) and (layer0_outputs(505));
    outputs(4531) <= (layer0_outputs(194)) and not (layer0_outputs(81));
    outputs(4532) <= layer0_outputs(4994);
    outputs(4533) <= (layer0_outputs(4243)) xor (layer0_outputs(2590));
    outputs(4534) <= not(layer0_outputs(3533));
    outputs(4535) <= (layer0_outputs(717)) and not (layer0_outputs(1138));
    outputs(4536) <= (layer0_outputs(924)) and (layer0_outputs(396));
    outputs(4537) <= not((layer0_outputs(1190)) xor (layer0_outputs(2543)));
    outputs(4538) <= not(layer0_outputs(2418));
    outputs(4539) <= not(layer0_outputs(1032));
    outputs(4540) <= not(layer0_outputs(2107)) or (layer0_outputs(1724));
    outputs(4541) <= not(layer0_outputs(172)) or (layer0_outputs(4854));
    outputs(4542) <= layer0_outputs(3154);
    outputs(4543) <= layer0_outputs(1414);
    outputs(4544) <= not(layer0_outputs(4240));
    outputs(4545) <= (layer0_outputs(2000)) xor (layer0_outputs(4422));
    outputs(4546) <= not(layer0_outputs(2239)) or (layer0_outputs(2793));
    outputs(4547) <= not((layer0_outputs(3113)) xor (layer0_outputs(3338)));
    outputs(4548) <= not(layer0_outputs(4667)) or (layer0_outputs(563));
    outputs(4549) <= not(layer0_outputs(859));
    outputs(4550) <= not(layer0_outputs(1711));
    outputs(4551) <= (layer0_outputs(1010)) or (layer0_outputs(4476));
    outputs(4552) <= not((layer0_outputs(1872)) and (layer0_outputs(353)));
    outputs(4553) <= (layer0_outputs(3573)) and (layer0_outputs(580));
    outputs(4554) <= not(layer0_outputs(17)) or (layer0_outputs(3778));
    outputs(4555) <= (layer0_outputs(4355)) xor (layer0_outputs(2662));
    outputs(4556) <= not(layer0_outputs(2783));
    outputs(4557) <= not((layer0_outputs(4279)) or (layer0_outputs(91)));
    outputs(4558) <= layer0_outputs(3566);
    outputs(4559) <= not((layer0_outputs(591)) or (layer0_outputs(3899)));
    outputs(4560) <= not((layer0_outputs(2716)) or (layer0_outputs(2642)));
    outputs(4561) <= layer0_outputs(4449);
    outputs(4562) <= layer0_outputs(1454);
    outputs(4563) <= not(layer0_outputs(3021)) or (layer0_outputs(3362));
    outputs(4564) <= (layer0_outputs(2529)) and (layer0_outputs(1529));
    outputs(4565) <= not(layer0_outputs(1971)) or (layer0_outputs(4984));
    outputs(4566) <= not(layer0_outputs(3508));
    outputs(4567) <= not(layer0_outputs(4678));
    outputs(4568) <= (layer0_outputs(89)) xor (layer0_outputs(5063));
    outputs(4569) <= (layer0_outputs(2564)) or (layer0_outputs(1066));
    outputs(4570) <= not((layer0_outputs(608)) xor (layer0_outputs(1669)));
    outputs(4571) <= not(layer0_outputs(3116));
    outputs(4572) <= (layer0_outputs(4539)) and not (layer0_outputs(1919));
    outputs(4573) <= not(layer0_outputs(11)) or (layer0_outputs(1507));
    outputs(4574) <= not((layer0_outputs(440)) and (layer0_outputs(5027)));
    outputs(4575) <= (layer0_outputs(5081)) and not (layer0_outputs(1824));
    outputs(4576) <= not(layer0_outputs(1810)) or (layer0_outputs(4007));
    outputs(4577) <= not((layer0_outputs(4587)) and (layer0_outputs(4823)));
    outputs(4578) <= layer0_outputs(746);
    outputs(4579) <= not((layer0_outputs(5002)) or (layer0_outputs(5038)));
    outputs(4580) <= not((layer0_outputs(408)) and (layer0_outputs(3266)));
    outputs(4581) <= not(layer0_outputs(3172));
    outputs(4582) <= not(layer0_outputs(1210));
    outputs(4583) <= not(layer0_outputs(4858));
    outputs(4584) <= not((layer0_outputs(57)) xor (layer0_outputs(4481)));
    outputs(4585) <= (layer0_outputs(2117)) xor (layer0_outputs(3226));
    outputs(4586) <= not(layer0_outputs(1956)) or (layer0_outputs(4742));
    outputs(4587) <= not(layer0_outputs(4457));
    outputs(4588) <= not((layer0_outputs(2488)) xor (layer0_outputs(1872)));
    outputs(4589) <= not(layer0_outputs(357));
    outputs(4590) <= not((layer0_outputs(271)) xor (layer0_outputs(4814)));
    outputs(4591) <= not(layer0_outputs(174));
    outputs(4592) <= not((layer0_outputs(3167)) or (layer0_outputs(3921)));
    outputs(4593) <= layer0_outputs(3769);
    outputs(4594) <= layer0_outputs(2734);
    outputs(4595) <= not(layer0_outputs(2992));
    outputs(4596) <= not((layer0_outputs(2752)) xor (layer0_outputs(2767)));
    outputs(4597) <= not((layer0_outputs(121)) xor (layer0_outputs(530)));
    outputs(4598) <= layer0_outputs(3728);
    outputs(4599) <= not((layer0_outputs(4303)) and (layer0_outputs(2458)));
    outputs(4600) <= not(layer0_outputs(982));
    outputs(4601) <= (layer0_outputs(4510)) and (layer0_outputs(1755));
    outputs(4602) <= (layer0_outputs(3398)) or (layer0_outputs(4394));
    outputs(4603) <= (layer0_outputs(2700)) and (layer0_outputs(4398));
    outputs(4604) <= layer0_outputs(2168);
    outputs(4605) <= not(layer0_outputs(5040));
    outputs(4606) <= not(layer0_outputs(888));
    outputs(4607) <= (layer0_outputs(4124)) or (layer0_outputs(423));
    outputs(4608) <= layer0_outputs(4866);
    outputs(4609) <= not((layer0_outputs(3194)) and (layer0_outputs(1631)));
    outputs(4610) <= layer0_outputs(2669);
    outputs(4611) <= not((layer0_outputs(2013)) or (layer0_outputs(1401)));
    outputs(4612) <= not((layer0_outputs(524)) and (layer0_outputs(1399)));
    outputs(4613) <= layer0_outputs(2063);
    outputs(4614) <= (layer0_outputs(518)) and not (layer0_outputs(2789));
    outputs(4615) <= (layer0_outputs(2345)) and not (layer0_outputs(4469));
    outputs(4616) <= not(layer0_outputs(2796)) or (layer0_outputs(2996));
    outputs(4617) <= layer0_outputs(4416);
    outputs(4618) <= not(layer0_outputs(4));
    outputs(4619) <= layer0_outputs(959);
    outputs(4620) <= not(layer0_outputs(245));
    outputs(4621) <= not(layer0_outputs(5085));
    outputs(4622) <= layer0_outputs(1312);
    outputs(4623) <= (layer0_outputs(154)) and not (layer0_outputs(3780));
    outputs(4624) <= (layer0_outputs(91)) and not (layer0_outputs(4471));
    outputs(4625) <= not(layer0_outputs(3970)) or (layer0_outputs(4942));
    outputs(4626) <= (layer0_outputs(2291)) xor (layer0_outputs(2230));
    outputs(4627) <= layer0_outputs(637);
    outputs(4628) <= layer0_outputs(260);
    outputs(4629) <= layer0_outputs(162);
    outputs(4630) <= layer0_outputs(4196);
    outputs(4631) <= not(layer0_outputs(2978));
    outputs(4632) <= not(layer0_outputs(890)) or (layer0_outputs(2797));
    outputs(4633) <= not((layer0_outputs(2031)) and (layer0_outputs(1166)));
    outputs(4634) <= (layer0_outputs(3891)) and (layer0_outputs(3765));
    outputs(4635) <= (layer0_outputs(4995)) and not (layer0_outputs(752));
    outputs(4636) <= (layer0_outputs(2498)) and (layer0_outputs(3574));
    outputs(4637) <= (layer0_outputs(1876)) and not (layer0_outputs(3189));
    outputs(4638) <= layer0_outputs(3939);
    outputs(4639) <= (layer0_outputs(388)) and (layer0_outputs(4287));
    outputs(4640) <= not((layer0_outputs(2687)) or (layer0_outputs(1374)));
    outputs(4641) <= not(layer0_outputs(2276));
    outputs(4642) <= (layer0_outputs(4725)) and not (layer0_outputs(3618));
    outputs(4643) <= layer0_outputs(1394);
    outputs(4644) <= (layer0_outputs(3475)) and (layer0_outputs(1005));
    outputs(4645) <= not(layer0_outputs(4777));
    outputs(4646) <= layer0_outputs(2946);
    outputs(4647) <= layer0_outputs(3178);
    outputs(4648) <= layer0_outputs(2313);
    outputs(4649) <= not(layer0_outputs(2848));
    outputs(4650) <= (layer0_outputs(1983)) and not (layer0_outputs(1592));
    outputs(4651) <= not((layer0_outputs(4852)) xor (layer0_outputs(450)));
    outputs(4652) <= not(layer0_outputs(84));
    outputs(4653) <= layer0_outputs(401);
    outputs(4654) <= (layer0_outputs(4153)) and not (layer0_outputs(1894));
    outputs(4655) <= (layer0_outputs(5008)) and not (layer0_outputs(1901));
    outputs(4656) <= not((layer0_outputs(1472)) or (layer0_outputs(2221)));
    outputs(4657) <= (layer0_outputs(3321)) and not (layer0_outputs(2572));
    outputs(4658) <= not((layer0_outputs(3171)) or (layer0_outputs(1386)));
    outputs(4659) <= (layer0_outputs(3089)) and not (layer0_outputs(616));
    outputs(4660) <= (layer0_outputs(4010)) and not (layer0_outputs(2392));
    outputs(4661) <= not((layer0_outputs(1646)) or (layer0_outputs(2769)));
    outputs(4662) <= not((layer0_outputs(4710)) or (layer0_outputs(1741)));
    outputs(4663) <= layer0_outputs(4459);
    outputs(4664) <= (layer0_outputs(2895)) and (layer0_outputs(4097));
    outputs(4665) <= not((layer0_outputs(2710)) or (layer0_outputs(4798)));
    outputs(4666) <= not((layer0_outputs(3305)) or (layer0_outputs(1233)));
    outputs(4667) <= not((layer0_outputs(1325)) xor (layer0_outputs(838)));
    outputs(4668) <= (layer0_outputs(1524)) and not (layer0_outputs(1751));
    outputs(4669) <= not(layer0_outputs(1655));
    outputs(4670) <= (layer0_outputs(3536)) xor (layer0_outputs(2091));
    outputs(4671) <= (layer0_outputs(2108)) and not (layer0_outputs(1432));
    outputs(4672) <= not((layer0_outputs(3234)) or (layer0_outputs(4501)));
    outputs(4673) <= not(layer0_outputs(452));
    outputs(4674) <= layer0_outputs(4960);
    outputs(4675) <= not(layer0_outputs(3090));
    outputs(4676) <= not((layer0_outputs(2418)) xor (layer0_outputs(4421)));
    outputs(4677) <= not(layer0_outputs(4283));
    outputs(4678) <= not(layer0_outputs(420)) or (layer0_outputs(4424));
    outputs(4679) <= (layer0_outputs(2713)) xor (layer0_outputs(578));
    outputs(4680) <= layer0_outputs(3417);
    outputs(4681) <= layer0_outputs(2616);
    outputs(4682) <= not(layer0_outputs(2157));
    outputs(4683) <= not(layer0_outputs(1654)) or (layer0_outputs(182));
    outputs(4684) <= not(layer0_outputs(3127)) or (layer0_outputs(3039));
    outputs(4685) <= layer0_outputs(941);
    outputs(4686) <= not(layer0_outputs(3532));
    outputs(4687) <= not(layer0_outputs(4345));
    outputs(4688) <= not(layer0_outputs(3297)) or (layer0_outputs(1998));
    outputs(4689) <= not((layer0_outputs(4980)) or (layer0_outputs(616)));
    outputs(4690) <= (layer0_outputs(4075)) and not (layer0_outputs(168));
    outputs(4691) <= layer0_outputs(2553);
    outputs(4692) <= (layer0_outputs(2979)) and not (layer0_outputs(1167));
    outputs(4693) <= layer0_outputs(2103);
    outputs(4694) <= not((layer0_outputs(3595)) or (layer0_outputs(640)));
    outputs(4695) <= not((layer0_outputs(583)) or (layer0_outputs(4054)));
    outputs(4696) <= not((layer0_outputs(4271)) and (layer0_outputs(1490)));
    outputs(4697) <= (layer0_outputs(2946)) and not (layer0_outputs(1603));
    outputs(4698) <= layer0_outputs(2822);
    outputs(4699) <= not((layer0_outputs(106)) or (layer0_outputs(3309)));
    outputs(4700) <= (layer0_outputs(815)) or (layer0_outputs(785));
    outputs(4701) <= layer0_outputs(516);
    outputs(4702) <= (layer0_outputs(3875)) and not (layer0_outputs(3288));
    outputs(4703) <= not(layer0_outputs(4065));
    outputs(4704) <= not((layer0_outputs(570)) or (layer0_outputs(744)));
    outputs(4705) <= not((layer0_outputs(1007)) or (layer0_outputs(2323)));
    outputs(4706) <= not(layer0_outputs(4131)) or (layer0_outputs(3576));
    outputs(4707) <= not(layer0_outputs(2192));
    outputs(4708) <= not(layer0_outputs(3560));
    outputs(4709) <= not((layer0_outputs(607)) or (layer0_outputs(2933)));
    outputs(4710) <= (layer0_outputs(3369)) and (layer0_outputs(4650));
    outputs(4711) <= layer0_outputs(1842);
    outputs(4712) <= layer0_outputs(4728);
    outputs(4713) <= layer0_outputs(713);
    outputs(4714) <= not((layer0_outputs(148)) xor (layer0_outputs(3422)));
    outputs(4715) <= (layer0_outputs(2034)) and not (layer0_outputs(3367));
    outputs(4716) <= (layer0_outputs(3228)) or (layer0_outputs(4652));
    outputs(4717) <= layer0_outputs(4558);
    outputs(4718) <= not((layer0_outputs(3293)) or (layer0_outputs(2219)));
    outputs(4719) <= not(layer0_outputs(4713));
    outputs(4720) <= (layer0_outputs(2464)) xor (layer0_outputs(317));
    outputs(4721) <= (layer0_outputs(1536)) and not (layer0_outputs(4718));
    outputs(4722) <= (layer0_outputs(475)) and (layer0_outputs(2925));
    outputs(4723) <= (layer0_outputs(2601)) and not (layer0_outputs(2858));
    outputs(4724) <= not((layer0_outputs(4564)) xor (layer0_outputs(2813)));
    outputs(4725) <= not((layer0_outputs(3597)) or (layer0_outputs(384)));
    outputs(4726) <= (layer0_outputs(4607)) and (layer0_outputs(1049));
    outputs(4727) <= (layer0_outputs(2741)) and not (layer0_outputs(2791));
    outputs(4728) <= not(layer0_outputs(2784)) or (layer0_outputs(753));
    outputs(4729) <= layer0_outputs(677);
    outputs(4730) <= (layer0_outputs(840)) xor (layer0_outputs(1513));
    outputs(4731) <= not((layer0_outputs(759)) or (layer0_outputs(2355)));
    outputs(4732) <= not((layer0_outputs(2739)) xor (layer0_outputs(2708)));
    outputs(4733) <= layer0_outputs(395);
    outputs(4734) <= layer0_outputs(1796);
    outputs(4735) <= not(layer0_outputs(2919));
    outputs(4736) <= layer0_outputs(1877);
    outputs(4737) <= not(layer0_outputs(1229));
    outputs(4738) <= not(layer0_outputs(4820));
    outputs(4739) <= not(layer0_outputs(2581)) or (layer0_outputs(855));
    outputs(4740) <= (layer0_outputs(4557)) xor (layer0_outputs(823));
    outputs(4741) <= not(layer0_outputs(2567)) or (layer0_outputs(1362));
    outputs(4742) <= not(layer0_outputs(320));
    outputs(4743) <= layer0_outputs(3439);
    outputs(4744) <= (layer0_outputs(2177)) and not (layer0_outputs(2583));
    outputs(4745) <= not(layer0_outputs(1662));
    outputs(4746) <= layer0_outputs(864);
    outputs(4747) <= not((layer0_outputs(1071)) or (layer0_outputs(4191)));
    outputs(4748) <= not(layer0_outputs(3716));
    outputs(4749) <= not((layer0_outputs(3969)) or (layer0_outputs(2075)));
    outputs(4750) <= layer0_outputs(2058);
    outputs(4751) <= layer0_outputs(3333);
    outputs(4752) <= layer0_outputs(3031);
    outputs(4753) <= not(layer0_outputs(4431));
    outputs(4754) <= not((layer0_outputs(1128)) xor (layer0_outputs(4389)));
    outputs(4755) <= not(layer0_outputs(3253));
    outputs(4756) <= (layer0_outputs(2691)) and not (layer0_outputs(2422));
    outputs(4757) <= not((layer0_outputs(4011)) xor (layer0_outputs(562)));
    outputs(4758) <= not(layer0_outputs(2352));
    outputs(4759) <= not((layer0_outputs(3993)) xor (layer0_outputs(3523)));
    outputs(4760) <= layer0_outputs(4570);
    outputs(4761) <= layer0_outputs(2397);
    outputs(4762) <= not(layer0_outputs(5022)) or (layer0_outputs(649));
    outputs(4763) <= (layer0_outputs(1141)) and not (layer0_outputs(1637));
    outputs(4764) <= (layer0_outputs(610)) xor (layer0_outputs(1728));
    outputs(4765) <= not(layer0_outputs(1926));
    outputs(4766) <= not((layer0_outputs(3868)) xor (layer0_outputs(971)));
    outputs(4767) <= (layer0_outputs(4390)) and not (layer0_outputs(1423));
    outputs(4768) <= (layer0_outputs(2345)) or (layer0_outputs(4694));
    outputs(4769) <= layer0_outputs(2888);
    outputs(4770) <= not(layer0_outputs(1105));
    outputs(4771) <= not((layer0_outputs(3572)) or (layer0_outputs(3339)));
    outputs(4772) <= not(layer0_outputs(970));
    outputs(4773) <= not(layer0_outputs(2851));
    outputs(4774) <= not((layer0_outputs(4379)) xor (layer0_outputs(2546)));
    outputs(4775) <= layer0_outputs(2082);
    outputs(4776) <= layer0_outputs(2745);
    outputs(4777) <= (layer0_outputs(328)) xor (layer0_outputs(815));
    outputs(4778) <= not(layer0_outputs(4311));
    outputs(4779) <= layer0_outputs(1544);
    outputs(4780) <= not(layer0_outputs(1718));
    outputs(4781) <= (layer0_outputs(1570)) and not (layer0_outputs(4677));
    outputs(4782) <= not((layer0_outputs(468)) or (layer0_outputs(4392)));
    outputs(4783) <= layer0_outputs(2886);
    outputs(4784) <= not(layer0_outputs(4920));
    outputs(4785) <= (layer0_outputs(3960)) and not (layer0_outputs(5118));
    outputs(4786) <= not(layer0_outputs(3831));
    outputs(4787) <= (layer0_outputs(5019)) and not (layer0_outputs(1270));
    outputs(4788) <= (layer0_outputs(18)) and (layer0_outputs(4665));
    outputs(4789) <= layer0_outputs(661);
    outputs(4790) <= (layer0_outputs(4490)) and not (layer0_outputs(3922));
    outputs(4791) <= not(layer0_outputs(1677));
    outputs(4792) <= layer0_outputs(181);
    outputs(4793) <= not(layer0_outputs(471));
    outputs(4794) <= not(layer0_outputs(296));
    outputs(4795) <= layer0_outputs(2683);
    outputs(4796) <= not(layer0_outputs(3249));
    outputs(4797) <= (layer0_outputs(3666)) and (layer0_outputs(3988));
    outputs(4798) <= not((layer0_outputs(55)) xor (layer0_outputs(3262)));
    outputs(4799) <= layer0_outputs(469);
    outputs(4800) <= (layer0_outputs(330)) and not (layer0_outputs(366));
    outputs(4801) <= layer0_outputs(1664);
    outputs(4802) <= not((layer0_outputs(24)) xor (layer0_outputs(2087)));
    outputs(4803) <= not(layer0_outputs(3504)) or (layer0_outputs(3082));
    outputs(4804) <= layer0_outputs(1000);
    outputs(4805) <= not(layer0_outputs(2988));
    outputs(4806) <= (layer0_outputs(991)) and not (layer0_outputs(578));
    outputs(4807) <= (layer0_outputs(4842)) and (layer0_outputs(1359));
    outputs(4808) <= layer0_outputs(3527);
    outputs(4809) <= layer0_outputs(4827);
    outputs(4810) <= (layer0_outputs(3576)) and not (layer0_outputs(4565));
    outputs(4811) <= not(layer0_outputs(2398));
    outputs(4812) <= (layer0_outputs(952)) and not (layer0_outputs(123));
    outputs(4813) <= not((layer0_outputs(691)) and (layer0_outputs(4635)));
    outputs(4814) <= (layer0_outputs(1968)) and not (layer0_outputs(4795));
    outputs(4815) <= layer0_outputs(1315);
    outputs(4816) <= not(layer0_outputs(344));
    outputs(4817) <= (layer0_outputs(2431)) and (layer0_outputs(2763));
    outputs(4818) <= (layer0_outputs(4797)) and not (layer0_outputs(3156));
    outputs(4819) <= not((layer0_outputs(1357)) xor (layer0_outputs(687)));
    outputs(4820) <= (layer0_outputs(3087)) and not (layer0_outputs(2537));
    outputs(4821) <= not(layer0_outputs(1429));
    outputs(4822) <= not(layer0_outputs(2875));
    outputs(4823) <= not(layer0_outputs(1364)) or (layer0_outputs(383));
    outputs(4824) <= layer0_outputs(457);
    outputs(4825) <= (layer0_outputs(1593)) and not (layer0_outputs(5099));
    outputs(4826) <= layer0_outputs(3670);
    outputs(4827) <= (layer0_outputs(2880)) xor (layer0_outputs(496));
    outputs(4828) <= not(layer0_outputs(88));
    outputs(4829) <= not((layer0_outputs(1852)) and (layer0_outputs(3221)));
    outputs(4830) <= (layer0_outputs(2982)) xor (layer0_outputs(1243));
    outputs(4831) <= not((layer0_outputs(556)) and (layer0_outputs(2214)));
    outputs(4832) <= (layer0_outputs(1485)) and not (layer0_outputs(3040));
    outputs(4833) <= (layer0_outputs(1467)) and not (layer0_outputs(2210));
    outputs(4834) <= (layer0_outputs(834)) and not (layer0_outputs(4472));
    outputs(4835) <= layer0_outputs(2314);
    outputs(4836) <= not(layer0_outputs(150));
    outputs(4837) <= not(layer0_outputs(2865));
    outputs(4838) <= not(layer0_outputs(2455));
    outputs(4839) <= not((layer0_outputs(1662)) or (layer0_outputs(1889)));
    outputs(4840) <= (layer0_outputs(651)) and not (layer0_outputs(4059));
    outputs(4841) <= (layer0_outputs(3009)) and (layer0_outputs(1022));
    outputs(4842) <= layer0_outputs(237);
    outputs(4843) <= not((layer0_outputs(2376)) or (layer0_outputs(1558)));
    outputs(4844) <= layer0_outputs(2434);
    outputs(4845) <= (layer0_outputs(4906)) and (layer0_outputs(1979));
    outputs(4846) <= not(layer0_outputs(109));
    outputs(4847) <= layer0_outputs(1110);
    outputs(4848) <= not((layer0_outputs(648)) and (layer0_outputs(4695)));
    outputs(4849) <= layer0_outputs(3762);
    outputs(4850) <= layer0_outputs(2913);
    outputs(4851) <= layer0_outputs(3145);
    outputs(4852) <= (layer0_outputs(4270)) xor (layer0_outputs(134));
    outputs(4853) <= layer0_outputs(1668);
    outputs(4854) <= (layer0_outputs(1873)) and not (layer0_outputs(3038));
    outputs(4855) <= not(layer0_outputs(2991));
    outputs(4856) <= (layer0_outputs(1450)) and not (layer0_outputs(205));
    outputs(4857) <= not(layer0_outputs(3069));
    outputs(4858) <= (layer0_outputs(4214)) and not (layer0_outputs(1826));
    outputs(4859) <= not((layer0_outputs(1316)) and (layer0_outputs(114)));
    outputs(4860) <= not(layer0_outputs(2907)) or (layer0_outputs(4646));
    outputs(4861) <= not(layer0_outputs(3771)) or (layer0_outputs(1927));
    outputs(4862) <= not(layer0_outputs(1167));
    outputs(4863) <= (layer0_outputs(4255)) and not (layer0_outputs(4298));
    outputs(4864) <= layer0_outputs(3596);
    outputs(4865) <= (layer0_outputs(512)) and (layer0_outputs(1245));
    outputs(4866) <= not(layer0_outputs(4830));
    outputs(4867) <= not(layer0_outputs(2057));
    outputs(4868) <= not(layer0_outputs(3687));
    outputs(4869) <= (layer0_outputs(2332)) xor (layer0_outputs(2295));
    outputs(4870) <= not(layer0_outputs(3923));
    outputs(4871) <= not((layer0_outputs(4145)) xor (layer0_outputs(1035)));
    outputs(4872) <= not(layer0_outputs(3136)) or (layer0_outputs(2335));
    outputs(4873) <= (layer0_outputs(4500)) and (layer0_outputs(949));
    outputs(4874) <= (layer0_outputs(3198)) or (layer0_outputs(1664));
    outputs(4875) <= (layer0_outputs(2556)) and not (layer0_outputs(3987));
    outputs(4876) <= (layer0_outputs(166)) and not (layer0_outputs(4265));
    outputs(4877) <= not(layer0_outputs(1775));
    outputs(4878) <= not((layer0_outputs(1913)) xor (layer0_outputs(1546)));
    outputs(4879) <= (layer0_outputs(3864)) and not (layer0_outputs(1054));
    outputs(4880) <= not((layer0_outputs(2855)) or (layer0_outputs(4224)));
    outputs(4881) <= not(layer0_outputs(5066)) or (layer0_outputs(4531));
    outputs(4882) <= (layer0_outputs(3392)) and (layer0_outputs(1468));
    outputs(4883) <= not(layer0_outputs(947));
    outputs(4884) <= (layer0_outputs(2656)) and not (layer0_outputs(2638));
    outputs(4885) <= not(layer0_outputs(1226));
    outputs(4886) <= not((layer0_outputs(1150)) and (layer0_outputs(4116)));
    outputs(4887) <= not(layer0_outputs(2078)) or (layer0_outputs(252));
    outputs(4888) <= not(layer0_outputs(402));
    outputs(4889) <= (layer0_outputs(3233)) and not (layer0_outputs(3623));
    outputs(4890) <= not(layer0_outputs(4078));
    outputs(4891) <= (layer0_outputs(2318)) and (layer0_outputs(3695));
    outputs(4892) <= (layer0_outputs(910)) and (layer0_outputs(411));
    outputs(4893) <= not(layer0_outputs(1308));
    outputs(4894) <= (layer0_outputs(2732)) and not (layer0_outputs(4965));
    outputs(4895) <= (layer0_outputs(2250)) and not (layer0_outputs(3874));
    outputs(4896) <= not(layer0_outputs(3828));
    outputs(4897) <= layer0_outputs(2036);
    outputs(4898) <= layer0_outputs(2089);
    outputs(4899) <= layer0_outputs(4156);
    outputs(4900) <= not(layer0_outputs(708)) or (layer0_outputs(1443));
    outputs(4901) <= not((layer0_outputs(3120)) or (layer0_outputs(2290)));
    outputs(4902) <= not(layer0_outputs(3630)) or (layer0_outputs(3784));
    outputs(4903) <= (layer0_outputs(2073)) and not (layer0_outputs(1104));
    outputs(4904) <= (layer0_outputs(695)) and (layer0_outputs(2682));
    outputs(4905) <= not(layer0_outputs(2818));
    outputs(4906) <= not(layer0_outputs(3834));
    outputs(4907) <= (layer0_outputs(3407)) and not (layer0_outputs(1642));
    outputs(4908) <= (layer0_outputs(872)) and (layer0_outputs(3747));
    outputs(4909) <= not(layer0_outputs(177));
    outputs(4910) <= not(layer0_outputs(2330));
    outputs(4911) <= (layer0_outputs(2847)) and (layer0_outputs(490));
    outputs(4912) <= layer0_outputs(3079);
    outputs(4913) <= (layer0_outputs(2654)) and not (layer0_outputs(953));
    outputs(4914) <= (layer0_outputs(400)) and not (layer0_outputs(2606));
    outputs(4915) <= not(layer0_outputs(1299));
    outputs(4916) <= not(layer0_outputs(296));
    outputs(4917) <= (layer0_outputs(2582)) and not (layer0_outputs(1084));
    outputs(4918) <= (layer0_outputs(3556)) and not (layer0_outputs(145));
    outputs(4919) <= (layer0_outputs(2994)) and not (layer0_outputs(3630));
    outputs(4920) <= not((layer0_outputs(1069)) or (layer0_outputs(4736)));
    outputs(4921) <= not((layer0_outputs(1049)) xor (layer0_outputs(4756)));
    outputs(4922) <= (layer0_outputs(15)) and (layer0_outputs(74));
    outputs(4923) <= (layer0_outputs(2286)) and not (layer0_outputs(1457));
    outputs(4924) <= layer0_outputs(5024);
    outputs(4925) <= layer0_outputs(2120);
    outputs(4926) <= layer0_outputs(1072);
    outputs(4927) <= layer0_outputs(4253);
    outputs(4928) <= (layer0_outputs(2185)) xor (layer0_outputs(5096));
    outputs(4929) <= (layer0_outputs(5119)) and (layer0_outputs(1338));
    outputs(4930) <= layer0_outputs(4771);
    outputs(4931) <= not(layer0_outputs(3307));
    outputs(4932) <= not(layer0_outputs(504));
    outputs(4933) <= (layer0_outputs(3207)) xor (layer0_outputs(3197));
    outputs(4934) <= (layer0_outputs(2908)) and not (layer0_outputs(908));
    outputs(4935) <= layer0_outputs(864);
    outputs(4936) <= (layer0_outputs(4893)) and not (layer0_outputs(2165));
    outputs(4937) <= layer0_outputs(1400);
    outputs(4938) <= (layer0_outputs(2823)) or (layer0_outputs(1245));
    outputs(4939) <= not((layer0_outputs(600)) xor (layer0_outputs(4615)));
    outputs(4940) <= layer0_outputs(361);
    outputs(4941) <= not(layer0_outputs(3779));
    outputs(4942) <= (layer0_outputs(2619)) and not (layer0_outputs(1823));
    outputs(4943) <= (layer0_outputs(588)) xor (layer0_outputs(2963));
    outputs(4944) <= not(layer0_outputs(58));
    outputs(4945) <= (layer0_outputs(627)) and (layer0_outputs(2161));
    outputs(4946) <= layer0_outputs(3619);
    outputs(4947) <= not((layer0_outputs(133)) xor (layer0_outputs(2104)));
    outputs(4948) <= layer0_outputs(4359);
    outputs(4949) <= not((layer0_outputs(2047)) xor (layer0_outputs(4968)));
    outputs(4950) <= (layer0_outputs(1665)) xor (layer0_outputs(4916));
    outputs(4951) <= layer0_outputs(1790);
    outputs(4952) <= not((layer0_outputs(3849)) or (layer0_outputs(2866)));
    outputs(4953) <= not((layer0_outputs(1127)) or (layer0_outputs(3059)));
    outputs(4954) <= not(layer0_outputs(398));
    outputs(4955) <= layer0_outputs(2644);
    outputs(4956) <= layer0_outputs(1465);
    outputs(4957) <= (layer0_outputs(1398)) and (layer0_outputs(2886));
    outputs(4958) <= not((layer0_outputs(287)) xor (layer0_outputs(16)));
    outputs(4959) <= layer0_outputs(478);
    outputs(4960) <= (layer0_outputs(183)) and (layer0_outputs(3018));
    outputs(4961) <= not((layer0_outputs(1563)) or (layer0_outputs(1730)));
    outputs(4962) <= (layer0_outputs(1251)) and not (layer0_outputs(3748));
    outputs(4963) <= not(layer0_outputs(1580));
    outputs(4964) <= (layer0_outputs(433)) or (layer0_outputs(2082));
    outputs(4965) <= not((layer0_outputs(3581)) xor (layer0_outputs(4409)));
    outputs(4966) <= not((layer0_outputs(1091)) or (layer0_outputs(3735)));
    outputs(4967) <= (layer0_outputs(3749)) and not (layer0_outputs(1770));
    outputs(4968) <= layer0_outputs(189);
    outputs(4969) <= not(layer0_outputs(2112));
    outputs(4970) <= (layer0_outputs(87)) and (layer0_outputs(3541));
    outputs(4971) <= (layer0_outputs(2060)) and (layer0_outputs(2046));
    outputs(4972) <= not((layer0_outputs(4458)) or (layer0_outputs(862)));
    outputs(4973) <= layer0_outputs(519);
    outputs(4974) <= not((layer0_outputs(1916)) or (layer0_outputs(2013)));
    outputs(4975) <= layer0_outputs(431);
    outputs(4976) <= (layer0_outputs(2263)) and (layer0_outputs(3537));
    outputs(4977) <= (layer0_outputs(3322)) xor (layer0_outputs(4438));
    outputs(4978) <= layer0_outputs(2341);
    outputs(4979) <= not(layer0_outputs(4658));
    outputs(4980) <= not(layer0_outputs(1622));
    outputs(4981) <= not((layer0_outputs(4027)) or (layer0_outputs(3618)));
    outputs(4982) <= layer0_outputs(1111);
    outputs(4983) <= layer0_outputs(3610);
    outputs(4984) <= layer0_outputs(1426);
    outputs(4985) <= (layer0_outputs(31)) and (layer0_outputs(642));
    outputs(4986) <= not(layer0_outputs(4625));
    outputs(4987) <= (layer0_outputs(3416)) and (layer0_outputs(4114));
    outputs(4988) <= (layer0_outputs(911)) xor (layer0_outputs(3967));
    outputs(4989) <= layer0_outputs(281);
    outputs(4990) <= layer0_outputs(3036);
    outputs(4991) <= layer0_outputs(3350);
    outputs(4992) <= (layer0_outputs(2585)) and not (layer0_outputs(4501));
    outputs(4993) <= layer0_outputs(3718);
    outputs(4994) <= (layer0_outputs(41)) xor (layer0_outputs(5056));
    outputs(4995) <= layer0_outputs(3719);
    outputs(4996) <= not(layer0_outputs(288));
    outputs(4997) <= not(layer0_outputs(2)) or (layer0_outputs(2982));
    outputs(4998) <= layer0_outputs(811);
    outputs(4999) <= (layer0_outputs(2837)) and not (layer0_outputs(3655));
    outputs(5000) <= layer0_outputs(3632);
    outputs(5001) <= not(layer0_outputs(45));
    outputs(5002) <= not(layer0_outputs(4525));
    outputs(5003) <= not(layer0_outputs(3325));
    outputs(5004) <= not(layer0_outputs(3370));
    outputs(5005) <= layer0_outputs(2986);
    outputs(5006) <= not(layer0_outputs(4457));
    outputs(5007) <= (layer0_outputs(3833)) and (layer0_outputs(4534));
    outputs(5008) <= (layer0_outputs(4256)) and (layer0_outputs(4156));
    outputs(5009) <= not((layer0_outputs(2853)) or (layer0_outputs(2150)));
    outputs(5010) <= (layer0_outputs(3445)) and (layer0_outputs(3075));
    outputs(5011) <= not(layer0_outputs(1701));
    outputs(5012) <= not((layer0_outputs(1227)) xor (layer0_outputs(3294)));
    outputs(5013) <= not((layer0_outputs(4561)) or (layer0_outputs(1772)));
    outputs(5014) <= not(layer0_outputs(905)) or (layer0_outputs(1203));
    outputs(5015) <= not(layer0_outputs(3681));
    outputs(5016) <= (layer0_outputs(2032)) xor (layer0_outputs(390));
    outputs(5017) <= (layer0_outputs(2040)) and not (layer0_outputs(647));
    outputs(5018) <= not(layer0_outputs(4870)) or (layer0_outputs(2008));
    outputs(5019) <= not(layer0_outputs(1206));
    outputs(5020) <= (layer0_outputs(3296)) xor (layer0_outputs(598));
    outputs(5021) <= layer0_outputs(4325);
    outputs(5022) <= not(layer0_outputs(2163));
    outputs(5023) <= not(layer0_outputs(4351));
    outputs(5024) <= not(layer0_outputs(4832));
    outputs(5025) <= (layer0_outputs(4807)) and (layer0_outputs(4748));
    outputs(5026) <= not(layer0_outputs(1469));
    outputs(5027) <= (layer0_outputs(3741)) and not (layer0_outputs(1592));
    outputs(5028) <= not((layer0_outputs(2954)) xor (layer0_outputs(786)));
    outputs(5029) <= layer0_outputs(5052);
    outputs(5030) <= not(layer0_outputs(3857));
    outputs(5031) <= layer0_outputs(3882);
    outputs(5032) <= not((layer0_outputs(4144)) or (layer0_outputs(4352)));
    outputs(5033) <= (layer0_outputs(3637)) and not (layer0_outputs(1738));
    outputs(5034) <= not(layer0_outputs(3453));
    outputs(5035) <= not(layer0_outputs(4639));
    outputs(5036) <= not(layer0_outputs(2425));
    outputs(5037) <= not(layer0_outputs(3423));
    outputs(5038) <= (layer0_outputs(3440)) and not (layer0_outputs(2697));
    outputs(5039) <= not((layer0_outputs(901)) xor (layer0_outputs(559)));
    outputs(5040) <= (layer0_outputs(4837)) and (layer0_outputs(1503));
    outputs(5041) <= not((layer0_outputs(2591)) or (layer0_outputs(1934)));
    outputs(5042) <= not((layer0_outputs(2819)) or (layer0_outputs(3156)));
    outputs(5043) <= (layer0_outputs(581)) and not (layer0_outputs(4927));
    outputs(5044) <= not(layer0_outputs(3555));
    outputs(5045) <= (layer0_outputs(4860)) and (layer0_outputs(3006));
    outputs(5046) <= not((layer0_outputs(1444)) xor (layer0_outputs(290)));
    outputs(5047) <= not(layer0_outputs(1438));
    outputs(5048) <= layer0_outputs(3112);
    outputs(5049) <= (layer0_outputs(2626)) xor (layer0_outputs(4817));
    outputs(5050) <= not((layer0_outputs(3763)) or (layer0_outputs(2149)));
    outputs(5051) <= (layer0_outputs(120)) and (layer0_outputs(2756));
    outputs(5052) <= (layer0_outputs(4208)) and not (layer0_outputs(726));
    outputs(5053) <= (layer0_outputs(5003)) and (layer0_outputs(2336));
    outputs(5054) <= layer0_outputs(958);
    outputs(5055) <= not(layer0_outputs(522));
    outputs(5056) <= (layer0_outputs(1776)) and not (layer0_outputs(3970));
    outputs(5057) <= not((layer0_outputs(2551)) or (layer0_outputs(2864)));
    outputs(5058) <= not(layer0_outputs(1264));
    outputs(5059) <= (layer0_outputs(143)) and (layer0_outputs(2326));
    outputs(5060) <= (layer0_outputs(432)) or (layer0_outputs(3032));
    outputs(5061) <= layer0_outputs(913);
    outputs(5062) <= not((layer0_outputs(3124)) or (layer0_outputs(2216)));
    outputs(5063) <= not((layer0_outputs(2039)) xor (layer0_outputs(3897)));
    outputs(5064) <= layer0_outputs(4610);
    outputs(5065) <= (layer0_outputs(4319)) xor (layer0_outputs(2754));
    outputs(5066) <= (layer0_outputs(2585)) and not (layer0_outputs(4015));
    outputs(5067) <= layer0_outputs(1955);
    outputs(5068) <= (layer0_outputs(1182)) and not (layer0_outputs(2945));
    outputs(5069) <= not((layer0_outputs(1144)) and (layer0_outputs(1399)));
    outputs(5070) <= not((layer0_outputs(4631)) xor (layer0_outputs(3488)));
    outputs(5071) <= not((layer0_outputs(3001)) or (layer0_outputs(3627)));
    outputs(5072) <= layer0_outputs(5038);
    outputs(5073) <= not((layer0_outputs(620)) or (layer0_outputs(2390)));
    outputs(5074) <= layer0_outputs(3863);
    outputs(5075) <= not(layer0_outputs(1739));
    outputs(5076) <= not(layer0_outputs(2199));
    outputs(5077) <= not((layer0_outputs(1716)) xor (layer0_outputs(2037)));
    outputs(5078) <= not(layer0_outputs(2889));
    outputs(5079) <= not(layer0_outputs(2041));
    outputs(5080) <= layer0_outputs(526);
    outputs(5081) <= not(layer0_outputs(1986));
    outputs(5082) <= layer0_outputs(1648);
    outputs(5083) <= (layer0_outputs(3084)) and (layer0_outputs(4149));
    outputs(5084) <= (layer0_outputs(2563)) and (layer0_outputs(26));
    outputs(5085) <= not((layer0_outputs(3469)) or (layer0_outputs(919)));
    outputs(5086) <= layer0_outputs(3835);
    outputs(5087) <= not(layer0_outputs(2993));
    outputs(5088) <= not((layer0_outputs(2076)) and (layer0_outputs(3465)));
    outputs(5089) <= (layer0_outputs(4594)) and not (layer0_outputs(5080));
    outputs(5090) <= layer0_outputs(1818);
    outputs(5091) <= layer0_outputs(4801);
    outputs(5092) <= (layer0_outputs(4084)) and not (layer0_outputs(358));
    outputs(5093) <= layer0_outputs(560);
    outputs(5094) <= layer0_outputs(3870);
    outputs(5095) <= (layer0_outputs(3216)) and not (layer0_outputs(2569));
    outputs(5096) <= (layer0_outputs(526)) and not (layer0_outputs(4744));
    outputs(5097) <= (layer0_outputs(3094)) and (layer0_outputs(3301));
    outputs(5098) <= not((layer0_outputs(2926)) xor (layer0_outputs(1838)));
    outputs(5099) <= (layer0_outputs(2213)) and not (layer0_outputs(3140));
    outputs(5100) <= not((layer0_outputs(2557)) or (layer0_outputs(5095)));
    outputs(5101) <= (layer0_outputs(2139)) and not (layer0_outputs(2590));
    outputs(5102) <= (layer0_outputs(1232)) and not (layer0_outputs(3828));
    outputs(5103) <= not(layer0_outputs(1703));
    outputs(5104) <= not(layer0_outputs(2469));
    outputs(5105) <= layer0_outputs(4056);
    outputs(5106) <= (layer0_outputs(628)) and (layer0_outputs(3753));
    outputs(5107) <= not((layer0_outputs(2253)) or (layer0_outputs(2361)));
    outputs(5108) <= not(layer0_outputs(4371));
    outputs(5109) <= (layer0_outputs(4140)) and not (layer0_outputs(333));
    outputs(5110) <= layer0_outputs(4383);
    outputs(5111) <= (layer0_outputs(4808)) and not (layer0_outputs(1006));
    outputs(5112) <= layer0_outputs(2691);
    outputs(5113) <= (layer0_outputs(1183)) and not (layer0_outputs(848));
    outputs(5114) <= not(layer0_outputs(1914));
    outputs(5115) <= not(layer0_outputs(2141));
    outputs(5116) <= (layer0_outputs(351)) and (layer0_outputs(4803));
    outputs(5117) <= not((layer0_outputs(2275)) or (layer0_outputs(3286)));
    outputs(5118) <= layer0_outputs(2265);
    outputs(5119) <= layer0_outputs(2996);

end Behavioral;
